.subckt sky130_fd_sc_hs__inv_1 A VGND VNB VPB VPWR Y
X0 Y.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1 Y.t1 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
R0 A.n0 A.t0 240.197
R1 A.n0 A.t1 181.407
R2 A A.n0 133.847
R3 VPWR VPWR.t0 263.572
R4 Y.n3 Y 589.85
R5 Y.n3 Y.n0 585
R6 Y.n4 Y.n3 585
R7 Y.n2 Y.t1 279.738
R8 Y.t1 Y.n1 279.738
R9 Y.n3 Y.t0 26.3844
R10 Y Y.n4 12.9944
R11 Y.n1 Y 12.6066
R12 Y Y.n0 11.249
R13 Y Y.n2 9.50353
R14 Y.n2 Y 4.84898
R15 Y Y.n0 3.10353
R16 Y.n1 Y 1.74595
R17 Y.n4 Y 1.35808
R18 VPB VPB.t0 472.447
R19 VGND VGND.t0 160.762
R20 VNB VNB.t0 2159.58
C0 VPB VPWR 0.067823f
C1 Y VPWR 0.124588f
C2 A VPWR 0.062459f
C3 VPWR VGND 0.026947f
C4 Y VPB 0.014642f
C5 A VPB 0.075723f
C6 VPB VGND 0.0075f
C7 Y A 0.073611f
C8 Y VGND 0.10291f
C9 A VGND 0.061935f
C10 VGND VNB 0.269359f
C11 Y VNB 0.11805f
C12 VPWR VNB 0.218384f
C13 A VNB 0.244142f
C14 VPB VNB 0.406224f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t2 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VPWR.t1 A.t1 Y.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t0 A.t2 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t0 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
R0 A.n0 A.t1 308.481
R1 A.n2 A.t3 256.765
R2 A.n0 A.t2 200.03
R3 A.n1 A.t0 187.478
R4 A A.n2 155.067
R5 A.n1 A.n0 86.7605
R6 A.n2 A.n1 9.038
R7 VGND.n0 VGND.t0 178.792
R8 VGND.n0 VGND.t1 178.577
R9 VGND VGND.n0 0.515549
R10 Y.n1 Y 590.615
R11 Y.n1 Y.n0 585
R12 Y.n2 Y.n1 585
R13 Y.n4 Y.n3 185
R14 Y.n5 Y.n4 185
R15 Y.n1 Y.t3 26.3844
R16 Y.n1 Y.t0 26.3844
R17 Y.n4 Y.t1 22.7032
R18 Y.n4 Y.t2 22.7032
R19 Y.n2 Y 15.0461
R20 Y.n0 Y 13.0251
R21 Y.n5 Y 12.6066
R22 Y.n3 Y 9.99348
R23 Y.n3 Y 4.84898
R24 Y.n0 Y 3.59348
R25 Y Y.n5 1.74595
R26 Y Y.n2 1.57243
R27 VNB VNB.t1 1177.95
R28 VNB.t1 VNB.t0 993.177
R29 VPWR.n0 VPWR.t1 266.2
R30 VPWR.n0 VPWR.t0 255.296
R31 VPWR VPWR.n0 0.552461
R32 VPB VPB.t0 252.823
R33 VPB.t0 VPB.t1 229.839
C0 VPB A 0.077592f
C1 VGND A 0.061731f
C2 Y A 0.113885f
C3 VPWR A 0.075328f
C4 VPB VGND 0.005232f
C5 VPB Y 0.006413f
C6 Y VGND 0.164244f
C7 VPWR VPB 0.063146f
C8 VPWR VGND 0.037599f
C9 VPWR Y 0.211648f
C10 VGND VNB 0.303237f
C11 Y VNB 0.041457f
C12 VPWR VNB 0.267578f
C13 A VNB 0.305477f
C14 VPB VNB 0.406224f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y
X0 Y.t5 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t1 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2 Y.t7 A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3 VPWR.t2 A.t3 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t1 A.t4 Y.t6 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5 Y.t3 A.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t0 A.t6 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t0 A.t7 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n0 A.t3 226.809
R1 A.n3 A.t5 226.809
R2 A.n9 A.t7 226.809
R3 A.n4 A.t0 226.809
R4 A.n4 A.t1 198.204
R5 A.n0 A.t6 198.204
R6 A.n10 A.t4 196.013
R7 A.n2 A.t2 196.013
R8 A A.n1 153.191
R9 A.n12 A.n11 152
R10 A.n8 A.n7 152
R11 A.n6 A.n5 152
R12 A.n8 A.n5 49.6611
R13 A.n11 A.n10 43.8187
R14 A.n1 A.n0 37.246
R15 A.n2 A.n1 23.3702
R16 A.n11 A.n3 21.1793
R17 A.n6 A 13.6935
R18 A.n5 A.n4 10.955
R19 A.n7 A 9.52608
R20 A A.n12 8.93073
R21 A.n12 A 5.35864
R22 A.n3 A.n2 5.11262
R23 A.n9 A.n8 5.11262
R24 A.n7 A 4.76329
R25 A.n10 A.n9 0.730803
R26 A A.n6 0.595849
R27 VPWR.n3 VPWR.t2 355.3
R28 VPWR.n2 VPWR.n1 331.5
R29 VPWR.n7 VPWR.t3 257.433
R30 VPWR.n3 VPWR.n2 40.4499
R31 VPWR.n6 VPWR.n5 36.1417
R32 VPWR.n1 VPWR.t1 26.3844
R33 VPWR.n1 VPWR.t0 26.3844
R34 VPWR.n7 VPWR.n6 24.0946
R35 VPWR.n5 VPWR.n4 9.3005
R36 VPWR.n6 VPWR.n0 9.3005
R37 VPWR.n8 VPWR.n7 9.3005
R38 VPWR.n4 VPWR.n3 2.0675
R39 VPWR.n5 VPWR.n2 1.12991
R40 VPWR.n4 VPWR.n0 0.122949
R41 VPWR.n8 VPWR.n0 0.122949
R42 VPWR VPWR.n8 0.0617245
R43 Y.n2 Y.n0 248.405
R44 Y.n2 Y.n1 205.487
R45 Y.n5 Y.n4 166.697
R46 Y.n5 Y.n3 103.65
R47 Y Y.n2 62.1018
R48 Y Y.n5 33.1299
R49 Y.n4 Y.t1 29.1897
R50 Y.n0 Y.t2 26.3844
R51 Y.n0 Y.t5 26.3844
R52 Y.n1 Y.t4 26.3844
R53 Y.n1 Y.t3 26.3844
R54 Y.n4 Y.t6 22.7032
R55 Y.n3 Y.t0 22.7032
R56 Y.n3 Y.t7 22.7032
R57 VPB VPB.t3 275.807
R58 VPB.t1 VPB.t2 229.839
R59 VPB.t0 VPB.t1 229.839
R60 VPB.t3 VPB.t0 229.839
R61 VGND.n1 VGND.t0 275.735
R62 VGND.n3 VGND.n2 208.079
R63 VGND.n5 VGND.t3 159.561
R64 VGND.n2 VGND.t2 30.8113
R65 VGND.n4 VGND.n3 24.4711
R66 VGND.n2 VGND.t1 22.7032
R67 VGND.n5 VGND.n4 20.7064
R68 VGND.n6 VGND.n5 9.3005
R69 VGND.n4 VGND.n0 9.3005
R70 VGND.n3 VGND.n1 6.55879
R71 VGND.n1 VGND.n0 0.675741
R72 VGND.n6 VGND.n0 0.122949
R73 VGND VGND.n6 0.0617245
R74 VNB VNB.t3 1212.6
R75 VNB.t1 VNB.t2 1108.66
R76 VNB.t3 VNB.t1 1085.56
R77 VNB.t2 VNB.t0 993.177
C0 A Y 0.373135f
C1 VPWR VPB 0.086151f
C2 VPWR VGND 0.043024f
C3 VPB Y 0.01352f
C4 A VPB 0.143465f
C5 VGND Y 0.312664f
C6 VGND A 0.103868f
C7 VPWR Y 0.382254f
C8 VGND VPB 0.005607f
C9 VPWR A 0.092902f
C10 VGND VNB 0.384929f
C11 Y VNB 0.084683f
C12 VPWR VNB 0.329316f
C13 A VNB 0.476918f
C14 VPB VNB 0.620496f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_8 A VGND VNB VPB VPWR Y
X0 Y.t12 A.t0 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t6 A.t1 Y.t11 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t15 A.t2 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 Y.t10 A.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t14 A.t4 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 VPWR.t2 A.t5 Y.t9 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t8 A.t6 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7 VGND.t5 A.t7 Y.t13 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VGND.t4 A.t8 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t0 A.t9 Y.t7 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t3 A.t10 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 Y.t2 A.t11 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X12 Y.t1 A.t12 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t4 A.t13 Y.t6 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y.t5 A.t14 VPWR.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X15 VGND.t0 A.t15 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n1 A.t13 230.459
R1 A.n15 A.t0 227.31
R2 A.n2 A.t14 226.809
R3 A.n4 A.t1 226.809
R4 A.n6 A.t3 226.809
R5 A.n9 A.t5 226.809
R6 A.n12 A.t6 226.809
R7 A.n13 A.t9 225.838
R8 A.n20 A.t12 196.013
R9 A.n10 A.t8 196.013
R10 A.n7 A.t4 196.013
R11 A.n5 A.t15 196.013
R12 A.n3 A.t11 196.013
R13 A.n1 A.t7 196.013
R14 A.n8 A.n0 162.121
R15 A.n11 A.n0 152
R16 A.n22 A.n21 152
R17 A.n19 A.n18 152
R18 A.n17 A.n16 152
R19 A.n14 A.t10 147.814
R20 A.n15 A.t2 147.814
R21 A.n4 A.n3 72.3005
R22 A.n2 A.n1 62.0763
R23 A.n6 A.n5 54.7732
R24 A.n20 A.n19 44.549
R25 A.n12 A.n11 42.3581
R26 A.n8 A.n7 31.4035
R27 A.n9 A.n8 26.2914
R28 A.n16 A.n14 21.5901
R29 A.n16 A.n15 21.5901
R30 A.n10 A.n9 15.3369
R31 A.n19 A.n13 12.3079
R32 A.n5 A.n4 10.955
R33 A.n18 A.n17 10.1214
R34 A.n22 A 8.63306
R35 A.n7 A.n6 8.03383
R36 A.n11 A.n10 8.03383
R37 A.n21 A.n12 7.30353
R38 A A.n22 5.65631
R39 A.n21 A.n20 5.11262
R40 A A.n0 4.46562
R41 A.n17 A 2.67957
R42 A.n18 A 1.48887
R43 A.n14 A.n13 1.43996
R44 A.n3 A.n2 0.730803
R45 VPWR.n4 VPWR.n3 323.406
R46 VPWR.n13 VPWR.n2 315.928
R47 VPWR.n5 VPWR.t4 265.531
R48 VPWR.n15 VPWR.t7 259.171
R49 VPWR.n7 VPWR.n6 223.696
R50 VPWR.n2 VPWR.t1 35.1791
R51 VPWR.n6 VPWR.t3 35.1791
R52 VPWR.n12 VPWR.n4 27.4829
R53 VPWR.n15 VPWR.n14 26.7299
R54 VPWR.n2 VPWR.t0 26.3844
R55 VPWR.n3 VPWR.t5 26.3844
R56 VPWR.n3 VPWR.t2 26.3844
R57 VPWR.n6 VPWR.t6 26.3844
R58 VPWR.n8 VPWR.n4 25.977
R59 VPWR.n13 VPWR.n12 25.224
R60 VPWR.n14 VPWR.n13 22.2123
R61 VPWR.n8 VPWR.n7 16.9417
R62 VPWR.n9 VPWR.n8 9.3005
R63 VPWR.n10 VPWR.n4 9.3005
R64 VPWR.n12 VPWR.n11 9.3005
R65 VPWR.n13 VPWR.n1 9.3005
R66 VPWR.n14 VPWR.n0 9.3005
R67 VPWR.n16 VPWR.n15 9.3005
R68 VPWR.n7 VPWR.n5 6.98721
R69 VPWR.n9 VPWR.n5 0.596295
R70 VPWR.n10 VPWR.n9 0.122949
R71 VPWR.n11 VPWR.n10 0.122949
R72 VPWR.n11 VPWR.n1 0.122949
R73 VPWR.n1 VPWR.n0 0.122949
R74 VPWR.n16 VPWR.n0 0.122949
R75 VPWR VPWR.n16 0.0617245
R76 Y.n5 Y.n3 261.483
R77 Y.n14 Y.n0 217.879
R78 Y.n6 Y.n2 207.349
R79 Y.n5 Y.n4 205.487
R80 Y.n10 Y.n9 162.933
R81 Y.n11 Y.n10 123.76
R82 Y.n13 Y.n1 106.343
R83 Y.n10 Y.n8 103.65
R84 Y.n11 Y.n7 95.3729
R85 Y.n6 Y.n5 55.3417
R86 Y.n12 Y.n6 41.453
R87 Y.n12 Y.n11 33.0223
R88 Y.n2 Y.t11 26.3844
R89 Y.n2 Y.t10 26.3844
R90 Y.n3 Y.t7 26.3844
R91 Y.n3 Y.t12 26.3844
R92 Y.n4 Y.t9 26.3844
R93 Y.n4 Y.t8 26.3844
R94 Y.n0 Y.t6 26.3844
R95 Y.n0 Y.t5 26.3844
R96 Y.n7 Y.t0 22.7032
R97 Y.n7 Y.t14 22.7032
R98 Y.n9 Y.t3 22.7032
R99 Y.n9 Y.t15 22.7032
R100 Y.n8 Y.t4 22.7032
R101 Y.n8 Y.t1 22.7032
R102 Y.n1 Y.t13 22.7032
R103 Y.n1 Y.t2 22.7032
R104 Y.n13 Y.n12 21.3338
R105 Y Y.n14 12.4005
R106 Y.n14 Y.n13 1.33383
R107 VPB VPB.t7 257.93
R108 VPB.t6 VPB.t0 255.376
R109 VPB.t2 VPB.t3 255.376
R110 VPB.t0 VPB.t1 229.839
R111 VPB.t5 VPB.t6 229.839
R112 VPB.t4 VPB.t5 229.839
R113 VPB.t3 VPB.t4 229.839
R114 VPB.t7 VPB.t2 229.839
R115 VGND.n9 VGND.n8 211.183
R116 VGND.n13 VGND.n2 211.183
R117 VGND.n15 VGND.t7 171.77
R118 VGND.n4 VGND.t5 160.25
R119 VGND.n6 VGND.n5 115.245
R120 VGND.n9 VGND.n7 34.6358
R121 VGND.n5 VGND.t2 34.0546
R122 VGND.n5 VGND.t0 34.0546
R123 VGND.n8 VGND.t6 34.0546
R124 VGND.n13 VGND.n1 27.1064
R125 VGND.n15 VGND.n14 25.6005
R126 VGND.n8 VGND.t4 22.7032
R127 VGND.n2 VGND.t1 22.7032
R128 VGND.n2 VGND.t3 22.7032
R129 VGND.n14 VGND.n13 20.3299
R130 VGND.n7 VGND.n6 15.8123
R131 VGND.n9 VGND.n1 12.8005
R132 VGND.n16 VGND.n15 9.3005
R133 VGND.n7 VGND.n3 9.3005
R134 VGND.n10 VGND.n9 9.3005
R135 VGND.n11 VGND.n1 9.3005
R136 VGND.n13 VGND.n12 9.3005
R137 VGND.n14 VGND.n0 9.3005
R138 VGND.n6 VGND.n4 6.93285
R139 VGND.n4 VGND.n3 0.677147
R140 VGND.n10 VGND.n3 0.122949
R141 VGND.n11 VGND.n10 0.122949
R142 VGND.n12 VGND.n11 0.122949
R143 VGND.n12 VGND.n0 0.122949
R144 VGND.n16 VGND.n0 0.122949
R145 VGND VGND.n16 0.0617245
R146 VNB.t0 VNB.t2 1316.54
R147 VNB VNB.t7 1177.95
R148 VNB.t4 VNB.t6 1154.86
R149 VNB.t2 VNB.t5 993.177
R150 VNB.t6 VNB.t0 993.177
R151 VNB.t1 VNB.t4 993.177
R152 VNB.t3 VNB.t1 993.177
R153 VNB.t7 VNB.t3 993.177
C0 VPB Y 0.020569f
C1 VGND Y 0.66808f
C2 A VPWR 0.174992f
C3 A VPB 0.29059f
C4 A VGND 0.141994f
C5 VPB VPWR 0.138167f
C6 A Y 0.664082f
C7 VPWR VGND 0.085813f
C8 VPB VGND 0.007616f
C9 VPWR Y 0.856977f
C10 VGND VNB 0.59851f
C11 Y VNB 0.083993f
C12 VPWR VNB 0.502892f
C13 A VNB 0.881288f
C14 VPB VNB 1.04904f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y
X0 Y.t31 A.t0 VPWR.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1 Y.t30 A.t1 VPWR.t4 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t3 A.t2 Y.t29 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t28 A.t3 VPWR.t2 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X4 Y.t2 A.t4 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 VGND.t14 A.t5 Y.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 Y.t27 A.t6 VPWR.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.1792 ps=1.44 w=1.12 l=0.15
X7 VGND.t13 A.t7 Y.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t0 A.t8 Y.t26 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.1848 ps=1.45 w=1.12 l=0.15
X9 VPWR.t11 A.t9 Y.t25 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t24 A.t10 VPWR.t10 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X11 Y.t5 A.t11 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X12 VGND.t11 A.t12 Y.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VGND.t10 A.t13 Y.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t9 A.t14 Y.t23 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Y.t15 A.t15 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 Y.t22 A.t16 VPWR.t8 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 VGND.t8 A.t17 Y.t14 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VPWR.t7 A.t18 Y.t21 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t13 A.t19 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X20 VPWR.t6 A.t20 Y.t20 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X21 Y.t19 A.t21 VPWR.t13 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X22 VPWR.t12 A.t22 Y.t18 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X23 VGND.t6 A.t23 Y.t11 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 Y.t17 A.t24 VPWR.t15 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X25 VGND.t5 A.t25 Y.t10 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 Y.t9 A.t26 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 VGND.t3 A.t27 Y.t8 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 Y.t7 A.t28 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X29 VPWR.t14 A.t29 Y.t16 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X30 Y.t6 A.t30 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X31 Y.t12 A.t31 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1628 ps=1.18 w=0.74 l=0.15
R0 A.n4 A.t2 235.571
R1 A.n36 A.t1 235.571
R2 A.n5 A.t3 226.809
R3 A.n9 A.t22 226.809
R4 A.n7 A.t24 226.809
R5 A.n13 A.t8 226.809
R6 A.n15 A.t6 226.809
R7 A.n18 A.t14 226.809
R8 A.n20 A.t16 226.809
R9 A.n23 A.t18 226.809
R10 A.n1 A.t21 226.809
R11 A.n28 A.t29 226.809
R12 A.n30 A.t0 226.809
R13 A.n33 A.t9 226.809
R14 A.n35 A.t10 226.809
R15 A.n37 A.t20 226.809
R16 A.n1 A.t28 196.013
R17 A.n28 A.t5 196.013
R18 A.n36 A.t11 196.013
R19 A.n38 A.t25 196.013
R20 A.n34 A.t15 196.013
R21 A.n32 A.t7 196.013
R22 A.n29 A.t30 196.013
R23 A.n22 A.t17 196.013
R24 A.n21 A.t26 196.013
R25 A.n19 A.t13 196.013
R26 A.n16 A.t4 196.013
R27 A.n14 A.t27 196.013
R28 A.n3 A.t19 196.013
R29 A.n8 A.t12 196.013
R30 A.n6 A.t31 196.013
R31 A.n4 A.t23 196.013
R32 A.n27 A.n26 168.282
R33 A.n25 A.n24 168.157
R34 A.n31 A.n0 167.922
R35 A.n11 A.n10 167.841
R36 A.n40 A.n39 167.494
R37 A.n17 A.n2 167.395
R38 A.n12 A.n11 167.031
R39 A.n22 A.n1 62.8066
R40 A.n29 A.n28 62.8066
R41 A.n34 A.n33 59.8853
R42 A.n15 A.n14 58.4247
R43 A.n5 A.n4 56.9641
R44 A.n20 A.n19 56.9641
R45 A.n37 A.n36 56.9641
R46 A.n8 A.n7 54.0429
R47 A.n13 A.n12 40.1672
R48 A.n10 A.n9 39.4369
R49 A.n28 A.n27 37.246
R50 A.n27 A.n1 35.7853
R51 A.n32 A.n31 35.7853
R52 A.n10 A.n6 35.055
R53 A.n31 A.n30 34.3247
R54 A.n39 A.n38 34.3247
R55 A.n18 A.n17 33.5944
R56 A.n39 A.n35 32.8641
R57 A.n24 A.n23 32.1338
R58 A.n12 A.n3 31.4035
R59 A.n17 A.n16 30.6732
R60 A.n24 A.n21 27.752
R61 A.n9 A.n8 11.6853
R62 A.n14 A.n13 11.6853
R63 A.n7 A.n3 8.76414
R64 A.n19 A.n18 8.76414
R65 A.n6 A.n5 5.84292
R66 A.n21 A.n20 5.84292
R67 A.n35 A.n34 5.84292
R68 A.n38 A.n37 5.84292
R69 A.n16 A.n15 4.38232
R70 A.n23 A.n22 2.92171
R71 A.n30 A.n29 2.92171
R72 A.n33 A.n32 2.92171
R73 A.n11 A.n2 0.541261
R74 A.n26 A.n0 0.51137
R75 A.n40 A.n0 0.51137
R76 A.n26 A.n25 0.497783
R77 A.n25 A.n2 0.495065
R78 A A.n40 0.0793043
R79 VPWR.n35 VPWR.t4 259.171
R80 VPWR.n13 VPWR.t3 258.68
R81 VPWR.n8 VPWR.n7 233.734
R82 VPWR.n4 VPWR.n3 231.429
R83 VPWR.n27 VPWR.n6 231.429
R84 VPWR.n21 VPWR.n10 226.987
R85 VPWR.n33 VPWR.n2 226.439
R86 VPWR.n12 VPWR.n11 222.651
R87 VPWR.n15 VPWR.n14 222.651
R88 VPWR.n2 VPWR.t10 35.1791
R89 VPWR.n3 VPWR.t5 35.1791
R90 VPWR.n6 VPWR.t13 35.1791
R91 VPWR.n11 VPWR.t15 35.1791
R92 VPWR.n11 VPWR.t0 35.1791
R93 VPWR.n14 VPWR.t2 35.1791
R94 VPWR.n14 VPWR.t12 35.1791
R95 VPWR.n21 VPWR.n20 32.0005
R96 VPWR.n22 VPWR.n8 30.8711
R97 VPWR.n10 VPWR.t1 29.9023
R98 VPWR.n16 VPWR.n12 28.9887
R99 VPWR.n32 VPWR.n4 27.4829
R100 VPWR.n35 VPWR.n34 26.7299
R101 VPWR.n28 VPWR.n27 26.7299
R102 VPWR.n27 VPWR.n26 26.7299
R103 VPWR.n2 VPWR.t6 26.3844
R104 VPWR.n3 VPWR.t11 26.3844
R105 VPWR.n6 VPWR.t14 26.3844
R106 VPWR.n7 VPWR.t8 26.3844
R107 VPWR.n7 VPWR.t7 26.3844
R108 VPWR.n10 VPWR.t9 26.3844
R109 VPWR.n28 VPWR.n4 25.977
R110 VPWR.n34 VPWR.n33 25.224
R111 VPWR.n33 VPWR.n32 25.224
R112 VPWR.n26 VPWR.n8 23.7181
R113 VPWR.n16 VPWR.n15 21.4593
R114 VPWR.n22 VPWR.n21 18.824
R115 VPWR.n20 VPWR.n12 18.4476
R116 VPWR.n17 VPWR.n16 9.3005
R117 VPWR.n18 VPWR.n12 9.3005
R118 VPWR.n20 VPWR.n19 9.3005
R119 VPWR.n21 VPWR.n9 9.3005
R120 VPWR.n23 VPWR.n22 9.3005
R121 VPWR.n24 VPWR.n8 9.3005
R122 VPWR.n26 VPWR.n25 9.3005
R123 VPWR.n27 VPWR.n5 9.3005
R124 VPWR.n29 VPWR.n28 9.3005
R125 VPWR.n30 VPWR.n4 9.3005
R126 VPWR.n32 VPWR.n31 9.3005
R127 VPWR.n33 VPWR.n1 9.3005
R128 VPWR.n34 VPWR.n0 9.3005
R129 VPWR.n36 VPWR.n35 9.3005
R130 VPWR.n15 VPWR.n13 6.77577
R131 VPWR.n17 VPWR.n13 0.617781
R132 VPWR.n18 VPWR.n17 0.122949
R133 VPWR.n19 VPWR.n18 0.122949
R134 VPWR.n19 VPWR.n9 0.122949
R135 VPWR.n23 VPWR.n9 0.122949
R136 VPWR.n24 VPWR.n23 0.122949
R137 VPWR.n25 VPWR.n24 0.122949
R138 VPWR.n25 VPWR.n5 0.122949
R139 VPWR.n29 VPWR.n5 0.122949
R140 VPWR.n30 VPWR.n29 0.122949
R141 VPWR.n31 VPWR.n30 0.122949
R142 VPWR.n31 VPWR.n1 0.122949
R143 VPWR.n1 VPWR.n0 0.122949
R144 VPWR.n36 VPWR.n0 0.122949
R145 VPWR VPWR.n36 0.0617245
R146 Y.n2 Y.n1 203.748
R147 Y.n13 Y.n12 203.454
R148 Y.n17 Y.n16 203.315
R149 Y.n25 Y.n24 203.056
R150 Y.n9 Y.n8 202.802
R151 Y.n29 Y.n27 202.684
R152 Y.n21 Y.n20 202.457
R153 Y.n5 Y.n4 202.457
R154 Y.n13 Y.n11 150.185
R155 Y.n25 Y.n23 143.799
R156 Y.n2 Y.n0 143.638
R157 Y.n17 Y.n15 142.806
R158 Y.n9 Y.n7 140.738
R159 Y.n21 Y.n19 140.192
R160 Y.n29 Y.n28 140.054
R161 Y.n5 Y.n3 138.594
R162 Y.n8 Y.t27 31.6612
R163 Y.n27 Y.t20 26.3844
R164 Y.n27 Y.t30 26.3844
R165 Y.n24 Y.t25 26.3844
R166 Y.n24 Y.t24 26.3844
R167 Y.n20 Y.t16 26.3844
R168 Y.n20 Y.t31 26.3844
R169 Y.n16 Y.t21 26.3844
R170 Y.n16 Y.t19 26.3844
R171 Y.n12 Y.t23 26.3844
R172 Y.n12 Y.t22 26.3844
R173 Y.n8 Y.t26 26.3844
R174 Y.n4 Y.t18 26.3844
R175 Y.n4 Y.t17 26.3844
R176 Y.n1 Y.t29 26.3844
R177 Y.n1 Y.t28 26.3844
R178 Y.n28 Y.t10 22.7032
R179 Y.n28 Y.t5 22.7032
R180 Y.n23 Y.t0 22.7032
R181 Y.n23 Y.t15 22.7032
R182 Y.n19 Y.t1 22.7032
R183 Y.n19 Y.t6 22.7032
R184 Y.n15 Y.t14 22.7032
R185 Y.n15 Y.t7 22.7032
R186 Y.n11 Y.t3 22.7032
R187 Y.n11 Y.t9 22.7032
R188 Y.n7 Y.t8 22.7032
R189 Y.n7 Y.t2 22.7032
R190 Y.n3 Y.t4 22.7032
R191 Y.n3 Y.t13 22.7032
R192 Y.n0 Y.t11 22.7032
R193 Y.n0 Y.t12 22.7032
R194 Y.n6 Y.n2 10.6406
R195 Y.n14 Y.n13 10.0685
R196 Y.n18 Y.n17 10.055
R197 Y.n10 Y.n9 10.0053
R198 Y.n30 Y.n29 9.99393
R199 Y.n22 Y.n21 9.97218
R200 Y.n6 Y.n5 9.97218
R201 Y.n26 Y.n25 9.43563
R202 Y.n10 Y.n6 0.543978
R203 Y.n14 Y.n10 0.516804
R204 Y.n22 Y.n18 0.516804
R205 Y.n26 Y.n22 0.516804
R206 Y.n30 Y.n26 0.516804
R207 Y.n18 Y.n14 0.48963
R208 Y Y.n30 0.0793043
R209 VPB.t2 VPB.t12 280.914
R210 VPB.t10 VPB.t1 280.914
R211 VPB VPB.t14 257.93
R212 VPB.t0 VPB.t3 255.376
R213 VPB.t9 VPB.t15 255.376
R214 VPB.t4 VPB.t8 255.376
R215 VPB.t11 VPB.t10 245.161
R216 VPB.t7 VPB.t11 240.054
R217 VPB.t12 VPB.t13 229.839
R218 VPB.t1 VPB.t2 229.839
R219 VPB.t6 VPB.t7 229.839
R220 VPB.t5 VPB.t6 229.839
R221 VPB.t3 VPB.t5 229.839
R222 VPB.t15 VPB.t0 229.839
R223 VPB.t8 VPB.t9 229.839
R224 VPB.t14 VPB.t4 229.839
R225 VGND.n9 VGND.t6 174.359
R226 VGND.n36 VGND.t12 174.131
R227 VGND.n20 VGND.n19 123.653
R228 VGND.n23 VGND.n22 123.079
R229 VGND.n34 VGND.n2 123.079
R230 VGND.n27 VGND.n5 121.957
R231 VGND.n30 VGND.n29 120.915
R232 VGND.n14 VGND.n13 117.856
R233 VGND.n11 VGND.n10 116.374
R234 VGND.n18 VGND.n7 36.1417
R235 VGND.n10 VGND.t0 35.6762
R236 VGND.n10 VGND.t11 35.6762
R237 VGND.n14 VGND.n12 34.2593
R238 VGND.n13 VGND.t7 34.0546
R239 VGND.n13 VGND.t3 34.0546
R240 VGND.n29 VGND.t1 34.0546
R241 VGND.n2 VGND.t5 34.0546
R242 VGND.n23 VGND.n21 30.8711
R243 VGND.n5 VGND.t14 30.8113
R244 VGND.n35 VGND.n34 29.7417
R245 VGND.n19 VGND.t15 28.3789
R246 VGND.n19 VGND.t10 28.3789
R247 VGND.n27 VGND.n4 26.7299
R248 VGND.n30 VGND.n1 25.977
R249 VGND.n5 VGND.t2 25.9464
R250 VGND.n28 VGND.n27 25.224
R251 VGND.n30 VGND.n28 25.224
R252 VGND.n34 VGND.n1 22.9652
R253 VGND.n22 VGND.t4 22.7032
R254 VGND.n22 VGND.t8 22.7032
R255 VGND.n29 VGND.t13 22.7032
R256 VGND.n2 VGND.t9 22.7032
R257 VGND.n23 VGND.n4 21.8358
R258 VGND.n36 VGND.n35 20.7064
R259 VGND.n12 VGND.n11 16.9417
R260 VGND.n21 VGND.n20 15.4358
R261 VGND.n14 VGND.n7 13.9299
R262 VGND.n37 VGND.n36 9.3005
R263 VGND.n12 VGND.n8 9.3005
R264 VGND.n15 VGND.n14 9.3005
R265 VGND.n16 VGND.n7 9.3005
R266 VGND.n18 VGND.n17 9.3005
R267 VGND.n21 VGND.n6 9.3005
R268 VGND.n24 VGND.n23 9.3005
R269 VGND.n25 VGND.n4 9.3005
R270 VGND.n27 VGND.n26 9.3005
R271 VGND.n28 VGND.n3 9.3005
R272 VGND.n31 VGND.n30 9.3005
R273 VGND.n32 VGND.n1 9.3005
R274 VGND.n34 VGND.n33 9.3005
R275 VGND.n35 VGND.n0 9.3005
R276 VGND.n11 VGND.n9 6.96039
R277 VGND.n20 VGND.n18 1.12991
R278 VGND.n9 VGND.n8 0.594857
R279 VGND.n15 VGND.n8 0.122949
R280 VGND.n16 VGND.n15 0.122949
R281 VGND.n17 VGND.n16 0.122949
R282 VGND.n17 VGND.n6 0.122949
R283 VGND.n24 VGND.n6 0.122949
R284 VGND.n25 VGND.n24 0.122949
R285 VGND.n26 VGND.n25 0.122949
R286 VGND.n26 VGND.n3 0.122949
R287 VGND.n31 VGND.n3 0.122949
R288 VGND.n32 VGND.n31 0.122949
R289 VGND.n33 VGND.n32 0.122949
R290 VGND.n33 VGND.n0 0.122949
R291 VGND.n37 VGND.n0 0.122949
R292 VGND VGND.n37 0.0617245
R293 VNB.t11 VNB.t0 1362.73
R294 VNB.t3 VNB.t7 1316.54
R295 VNB VNB.t12 1304.99
R296 VNB.t10 VNB.t15 1154.86
R297 VNB.t14 VNB.t2 1154.86
R298 VNB.t13 VNB.t1 1154.86
R299 VNB.t5 VNB.t9 1154.86
R300 VNB.t0 VNB.t6 993.177
R301 VNB.t7 VNB.t11 993.177
R302 VNB.t15 VNB.t3 993.177
R303 VNB.t4 VNB.t10 993.177
R304 VNB.t8 VNB.t4 993.177
R305 VNB.t2 VNB.t8 993.177
R306 VNB.t1 VNB.t14 993.177
R307 VNB.t9 VNB.t13 993.177
R308 VNB.t12 VNB.t5 993.177
C0 Y VPB 0.045372f
C1 VGND VPWR 0.064897f
C2 VPWR A 0.529164f
C3 VPWR Y 2.08315f
C4 VGND A 0.686864f
C5 VPWR VPB 0.231595f
C6 VGND Y 1.31768f
C7 VGND VPB 0.008245f
C8 A Y 2.0772f
C9 A VPB 0.601473f
C10 VGND VNB 1.02743f
C11 Y VNB 0.09351f
C12 VPWR VNB 0.825774f
C13 A VNB 1.727695f
C14 VPB VNB 1.90613f
C15 Y.t11 VNB 0.017533f
C16 Y.t12 VNB 0.017533f
C17 Y.n0 VNB 0.077558f
C18 Y.t29 VNB 0.028432f
C19 Y.t28 VNB 0.028432f
C20 Y.n1 VNB 0.061755f
C21 Y.n2 VNB 0.211114f
C22 Y.t4 VNB 0.017533f
C23 Y.t13 VNB 0.017533f
C24 Y.n3 VNB 0.075471f
C25 Y.t18 VNB 0.028432f
C26 Y.t17 VNB 0.028432f
C27 Y.n4 VNB 0.061808f
C28 Y.n5 VNB 0.238955f
C29 Y.n6 VNB 0.138977f
C30 Y.t8 VNB 0.017533f
C31 Y.t2 VNB 0.017533f
C32 Y.n7 VNB 0.074431f
C33 Y.t26 VNB 0.028432f
C34 Y.t27 VNB 0.034118f
C35 Y.n8 VNB 0.067479f
C36 Y.n9 VNB 0.225797f
C37 Y.n10 VNB 0.082839f
C38 Y.t3 VNB 0.017533f
C39 Y.t9 VNB 0.017533f
C40 Y.n11 VNB 0.071679f
C41 Y.t23 VNB 0.028432f
C42 Y.t22 VNB 0.028432f
C43 Y.n12 VNB 0.061767f
C44 Y.n13 VNB 0.190901f
C45 Y.n14 VNB 0.078899f
C46 Y.t14 VNB 0.017533f
C47 Y.t7 VNB 0.017533f
C48 Y.n15 VNB 0.074045f
C49 Y.t21 VNB 0.028432f
C50 Y.t19 VNB 0.028432f
C51 Y.n16 VNB 0.061772f
C52 Y.n17 VNB 0.2118f
C53 Y.n18 VNB 0.078908f
C54 Y.t1 VNB 0.017533f
C55 Y.t6 VNB 0.017533f
C56 Y.n19 VNB 0.074551f
C57 Y.t16 VNB 0.028432f
C58 Y.t31 VNB 0.028432f
C59 Y.n20 VNB 0.061808f
C60 Y.n21 VNB 0.2316f
C61 Y.n22 VNB 0.080921f
C62 Y.t0 VNB 0.017533f
C63 Y.t15 VNB 0.017533f
C64 Y.n23 VNB 0.073941f
C65 Y.t25 VNB 0.028432f
C66 Y.t24 VNB 0.028432f
C67 Y.n24 VNB 0.06188f
C68 Y.n25 VNB 0.226892f
C69 Y.n26 VNB 0.075404f
C70 Y.t20 VNB 0.028432f
C71 Y.t30 VNB 0.028432f
C72 Y.n27 VNB 0.061918f
C73 Y.t10 VNB 0.017533f
C74 Y.t5 VNB 0.017533f
C75 Y.n28 VNB 0.075754f
C76 Y.n29 VNB 0.232942f
C77 Y.n30 VNB 0.049674f
C78 VPWR.n0 VNB 0.040808f
C79 VPWR.t4 VNB 0.060735f
C80 VPWR.n1 VNB 0.040808f
C81 VPWR.t10 VNB 0.019433f
C82 VPWR.t6 VNB 0.014574f
C83 VPWR.n2 VNB 0.041719f
C84 VPWR.t5 VNB 0.019433f
C85 VPWR.t11 VNB 0.014574f
C86 VPWR.n3 VNB 0.041545f
C87 VPWR.n4 VNB 0.066913f
C88 VPWR.n5 VNB 0.040808f
C89 VPWR.t13 VNB 0.019433f
C90 VPWR.t14 VNB 0.014574f
C91 VPWR.n6 VNB 0.041545f
C92 VPWR.t8 VNB 0.014574f
C93 VPWR.t7 VNB 0.014574f
C94 VPWR.n7 VNB 0.036609f
C95 VPWR.n8 VNB 0.063369f
C96 VPWR.n9 VNB 0.040808f
C97 VPWR.t1 VNB 0.016518f
C98 VPWR.t9 VNB 0.014574f
C99 VPWR.n10 VNB 0.038784f
C100 VPWR.t15 VNB 0.019433f
C101 VPWR.t0 VNB 0.019433f
C102 VPWR.n11 VNB 0.046714f
C103 VPWR.n12 VNB 0.085896f
C104 VPWR.t3 VNB 0.063115f
C105 VPWR.n13 VNB 0.117088f
C106 VPWR.t2 VNB 0.019433f
C107 VPWR.t12 VNB 0.019433f
C108 VPWR.n14 VNB 0.046714f
C109 VPWR.n15 VNB 0.087431f
C110 VPWR.n16 VNB 0.009881f
C111 VPWR.n17 VNB 0.135007f
C112 VPWR.n18 VNB 0.040808f
C113 VPWR.n19 VNB 0.040808f
C114 VPWR.n20 VNB 0.009881f
C115 VPWR.n21 VNB 0.075195f
C116 VPWR.n22 VNB 0.009734f
C117 VPWR.n23 VNB 0.040808f
C118 VPWR.n24 VNB 0.040808f
C119 VPWR.n25 VNB 0.040808f
C120 VPWR.n26 VNB 0.009881f
C121 VPWR.n27 VNB 0.066913f
C122 VPWR.n28 VNB 0.010323f
C123 VPWR.n29 VNB 0.040808f
C124 VPWR.n30 VNB 0.040808f
C125 VPWR.n31 VNB 0.040808f
C126 VPWR.n32 VNB 0.010323f
C127 VPWR.n33 VNB 0.076386f
C128 VPWR.n34 VNB 0.010176f
C129 VPWR.n35 VNB 0.06762f
C130 VPWR.n36 VNB 0.030606f
C131 A.n0 VNB 0.072399f
C132 A.t10 VNB 0.025933f
C133 A.t15 VNB 0.018017f
C134 A.t9 VNB 0.025933f
C135 A.t7 VNB 0.018017f
C136 A.t0 VNB 0.025933f
C137 A.t30 VNB 0.018017f
C138 A.t29 VNB 0.025933f
C139 A.t5 VNB 0.018017f
C140 A.t21 VNB 0.025933f
C141 A.t28 VNB 0.018017f
C142 A.n1 VNB 0.047273f
C143 A.n2 VNB 0.075212f
C144 A.t26 VNB 0.018017f
C145 A.t16 VNB 0.025933f
C146 A.t13 VNB 0.018017f
C147 A.t14 VNB 0.025933f
C148 A.t4 VNB 0.018017f
C149 A.t6 VNB 0.025933f
C150 A.t27 VNB 0.018017f
C151 A.t8 VNB 0.025933f
C152 A.t19 VNB 0.018017f
C153 A.n3 VNB 0.020083f
C154 A.t31 VNB 0.018017f
C155 A.t3 VNB 0.025933f
C156 A.t23 VNB 0.018017f
C157 A.t2 VNB 0.026728f
C158 A.n4 VNB 0.047024f
C159 A.n5 VNB 0.028282f
C160 A.n6 VNB 0.020264f
C161 A.t22 VNB 0.025933f
C162 A.t12 VNB 0.018017f
C163 A.t24 VNB 0.025933f
C164 A.n7 VNB 0.028282f
C165 A.n8 VNB 0.026446f
C166 A.n9 VNB 0.025372f
C167 A.n10 VNB 0.020992f
C168 A.n11 VNB 0.13885f
C169 A.n12 VNB 0.020153f
C170 A.n13 VNB 0.025554f
C171 A.n14 VNB 0.027537f
C172 A.n15 VNB 0.028282f
C173 A.n16 VNB 0.01881f
C174 A.n17 VNB 0.018227f
C175 A.n18 VNB 0.023191f
C176 A.n19 VNB 0.026446f
C177 A.n20 VNB 0.028282f
C178 A.n21 VNB 0.018446f
C179 A.t18 VNB 0.025933f
C180 A.t17 VNB 0.018017f
C181 A.n22 VNB 0.026446f
C182 A.n23 VNB 0.021372f
C183 A.n24 VNB 0.016946f
C184 A.n25 VNB 0.070133f
C185 A.n26 VNB 0.070458f
C186 A.n27 VNB 0.020192f
C187 A.n28 VNB 0.047637f
C188 A.n29 VNB 0.026446f
C189 A.n30 VNB 0.021918f
C190 A.n31 VNB 0.019546f
C191 A.n32 VNB 0.019719f
C192 A.n33 VNB 0.028282f
C193 A.n34 VNB 0.026446f
C194 A.n35 VNB 0.022282f
C195 A.t25 VNB 0.018017f
C196 A.t20 VNB 0.025933f
C197 A.t11 VNB 0.018017f
C198 A.t1 VNB 0.026728f
C199 A.n36 VNB 0.047024f
C200 A.n37 VNB 0.028282f
C201 A.n38 VNB 0.020083f
C202 A.n39 VNB 0.018927f
C203 A.n40 VNB 0.053993f
.ends
