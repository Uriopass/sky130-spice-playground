* NGSPICE file created from sky130_fd_sc_hs__inv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_1 A VGND VNB VPB VPWR Y
X0 Y.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1 Y.t1 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
R0 A.n0 A.t0 240.197
R1 A.n0 A.t1 181.407
R2 A A.n0 133.847
R3 VPWR VPWR.t0 263.572
R4 Y.n3 Y 589.85
R5 Y.n3 Y.n0 585
R6 Y.n4 Y.n3 585
R7 Y.n2 Y.t1 279.738
R8 Y.t1 Y.n1 279.738
R9 Y.n3 Y.t0 26.3844
R10 Y Y.n4 12.9944
R11 Y.n1 Y 12.6066
R12 Y Y.n0 11.249
R13 Y Y.n2 9.50353
R14 Y.n2 Y 4.84898
R15 Y Y.n0 3.10353
R16 Y.n1 Y 1.74595
R17 Y.n4 Y 1.35808
R18 VPB VPB.t0 472.447
R19 VGND VGND.t0 160.762
R20 VNB VNB.t0 2159.58
C0 VPB VPWR 0.067823f
C1 Y VPWR 0.124588f
C2 A VPWR 0.062459f
C3 VPWR VGND 0.026947f
C4 Y VPB 0.014642f
C5 A VPB 0.075723f
C6 VPB VGND 0.0075f
C7 Y A 0.073611f
C8 Y VGND 0.10291f
C9 A VGND 0.061935f
C10 VGND VNB 0.269359f
C11 Y VNB 0.11805f
C12 VPWR VNB 0.218384f
C13 A VNB 0.244142f
C14 VPB VNB 0.406224f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t2 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VPWR.t1 A.t1 Y.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t0 A.t2 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t0 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
R0 A.n0 A.t1 308.481
R1 A.n2 A.t3 256.765
R2 A.n0 A.t2 200.03
R3 A.n1 A.t0 187.478
R4 A A.n2 155.067
R5 A.n1 A.n0 86.7605
R6 A.n2 A.n1 9.038
R7 VGND.n0 VGND.t0 178.792
R8 VGND.n0 VGND.t1 178.577
R9 VGND VGND.n0 0.515549
R10 Y.n1 Y 590.615
R11 Y.n1 Y.n0 585
R12 Y.n2 Y.n1 585
R13 Y.n4 Y.n3 185
R14 Y.n5 Y.n4 185
R15 Y.n1 Y.t3 26.3844
R16 Y.n1 Y.t0 26.3844
R17 Y.n4 Y.t1 22.7032
R18 Y.n4 Y.t2 22.7032
R19 Y.n2 Y 15.0461
R20 Y.n0 Y 13.0251
R21 Y.n5 Y 12.6066
R22 Y.n3 Y 9.99348
R23 Y.n3 Y 4.84898
R24 Y.n0 Y 3.59348
R25 Y Y.n5 1.74595
R26 Y Y.n2 1.57243
R27 VNB VNB.t1 1177.95
R28 VNB.t1 VNB.t0 993.177
R29 VPWR.n0 VPWR.t1 266.2
R30 VPWR.n0 VPWR.t0 255.296
R31 VPWR VPWR.n0 0.552461
R32 VPB VPB.t0 252.823
R33 VPB.t0 VPB.t1 229.839
C0 VPB A 0.077592f
C1 VGND A 0.061731f
C2 Y A 0.113885f
C3 VPWR A 0.075328f
C4 VPB VGND 0.005232f
C5 VPB Y 0.006413f
C6 Y VGND 0.164244f
C7 VPWR VPB 0.063146f
C8 VPWR VGND 0.037599f
C9 VPWR Y 0.211648f
C10 VGND VNB 0.303237f
C11 Y VNB 0.041457f
C12 VPWR VNB 0.267578f
C13 A VNB 0.305477f
C14 VPB VNB 0.406224f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y
X0 Y.t5 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t1 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2 Y.t7 A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3 VPWR.t2 A.t3 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t1 A.t4 Y.t6 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5 Y.t3 A.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t0 A.t6 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t0 A.t7 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n0 A.t3 226.809
R1 A.n3 A.t5 226.809
R2 A.n9 A.t7 226.809
R3 A.n4 A.t0 226.809
R4 A.n4 A.t1 198.204
R5 A.n0 A.t6 198.204
R6 A.n10 A.t4 196.013
R7 A.n2 A.t2 196.013
R8 A A.n1 153.191
R9 A.n12 A.n11 152
R10 A.n8 A.n7 152
R11 A.n6 A.n5 152
R12 A.n8 A.n5 49.6611
R13 A.n11 A.n10 43.8187
R14 A.n1 A.n0 37.246
R15 A.n2 A.n1 23.3702
R16 A.n11 A.n3 21.1793
R17 A.n6 A 13.6935
R18 A.n5 A.n4 10.955
R19 A.n7 A 9.52608
R20 A A.n12 8.93073
R21 A.n12 A 5.35864
R22 A.n3 A.n2 5.11262
R23 A.n9 A.n8 5.11262
R24 A.n7 A 4.76329
R25 A.n10 A.n9 0.730803
R26 A A.n6 0.595849
R27 VPWR.n3 VPWR.t2 355.3
R28 VPWR.n2 VPWR.n1 331.5
R29 VPWR.n7 VPWR.t3 257.433
R30 VPWR.n3 VPWR.n2 40.4499
R31 VPWR.n6 VPWR.n5 36.1417
R32 VPWR.n1 VPWR.t1 26.3844
R33 VPWR.n1 VPWR.t0 26.3844
R34 VPWR.n7 VPWR.n6 24.0946
R35 VPWR.n5 VPWR.n4 9.3005
R36 VPWR.n6 VPWR.n0 9.3005
R37 VPWR.n8 VPWR.n7 9.3005
R38 VPWR.n4 VPWR.n3 2.0675
R39 VPWR.n5 VPWR.n2 1.12991
R40 VPWR.n4 VPWR.n0 0.122949
R41 VPWR.n8 VPWR.n0 0.122949
R42 VPWR VPWR.n8 0.0617245
R43 Y.n2 Y.n0 248.405
R44 Y.n2 Y.n1 205.487
R45 Y.n5 Y.n4 166.697
R46 Y.n5 Y.n3 103.65
R47 Y Y.n2 62.1018
R48 Y Y.n5 33.1299
R49 Y.n4 Y.t1 29.1897
R50 Y.n0 Y.t2 26.3844
R51 Y.n0 Y.t5 26.3844
R52 Y.n1 Y.t4 26.3844
R53 Y.n1 Y.t3 26.3844
R54 Y.n4 Y.t6 22.7032
R55 Y.n3 Y.t0 22.7032
R56 Y.n3 Y.t7 22.7032
R57 VPB VPB.t3 275.807
R58 VPB.t1 VPB.t2 229.839
R59 VPB.t0 VPB.t1 229.839
R60 VPB.t3 VPB.t0 229.839
R61 VGND.n1 VGND.t0 275.735
R62 VGND.n3 VGND.n2 208.079
R63 VGND.n5 VGND.t3 159.561
R64 VGND.n2 VGND.t2 30.8113
R65 VGND.n4 VGND.n3 24.4711
R66 VGND.n2 VGND.t1 22.7032
R67 VGND.n5 VGND.n4 20.7064
R68 VGND.n6 VGND.n5 9.3005
R69 VGND.n4 VGND.n0 9.3005
R70 VGND.n3 VGND.n1 6.55879
R71 VGND.n1 VGND.n0 0.675741
R72 VGND.n6 VGND.n0 0.122949
R73 VGND VGND.n6 0.0617245
R74 VNB VNB.t3 1212.6
R75 VNB.t1 VNB.t2 1108.66
R76 VNB.t3 VNB.t1 1085.56
R77 VNB.t2 VNB.t0 993.177
C0 A Y 0.373135f
C1 VPWR VPB 0.086151f
C2 VPWR VGND 0.043024f
C3 VPB Y 0.01352f
C4 A VPB 0.143465f
C5 VGND Y 0.312664f
C6 VGND A 0.103868f
C7 VPWR Y 0.382254f
C8 VGND VPB 0.005607f
C9 VPWR A 0.092902f
C10 VGND VNB 0.384929f
C11 Y VNB 0.084683f
C12 VPWR VNB 0.329316f
C13 A VNB 0.476918f
C14 VPB VNB 0.620496f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_8 A VGND VNB VPB VPWR Y
X0 Y.t12 A.t0 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t6 A.t1 Y.t11 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t15 A.t2 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 Y.t10 A.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t14 A.t4 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 VPWR.t2 A.t5 Y.t9 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t8 A.t6 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7 VGND.t5 A.t7 Y.t13 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VGND.t4 A.t8 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t0 A.t9 Y.t7 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t3 A.t10 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 Y.t2 A.t11 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X12 Y.t1 A.t12 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t4 A.t13 Y.t6 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y.t5 A.t14 VPWR.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X15 VGND.t0 A.t15 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n1 A.t13 230.459
R1 A.n15 A.t0 227.31
R2 A.n2 A.t14 226.809
R3 A.n4 A.t1 226.809
R4 A.n6 A.t3 226.809
R5 A.n9 A.t5 226.809
R6 A.n12 A.t6 226.809
R7 A.n13 A.t9 225.838
R8 A.n20 A.t12 196.013
R9 A.n10 A.t8 196.013
R10 A.n7 A.t4 196.013
R11 A.n5 A.t15 196.013
R12 A.n3 A.t11 196.013
R13 A.n1 A.t7 196.013
R14 A.n8 A.n0 162.121
R15 A.n11 A.n0 152
R16 A.n22 A.n21 152
R17 A.n19 A.n18 152
R18 A.n17 A.n16 152
R19 A.n14 A.t10 147.814
R20 A.n15 A.t2 147.814
R21 A.n4 A.n3 72.3005
R22 A.n2 A.n1 62.0763
R23 A.n6 A.n5 54.7732
R24 A.n20 A.n19 44.549
R25 A.n12 A.n11 42.3581
R26 A.n8 A.n7 31.4035
R27 A.n9 A.n8 26.2914
R28 A.n16 A.n14 21.5901
R29 A.n16 A.n15 21.5901
R30 A.n10 A.n9 15.3369
R31 A.n19 A.n13 12.3079
R32 A.n5 A.n4 10.955
R33 A.n18 A.n17 10.1214
R34 A.n22 A 8.63306
R35 A.n7 A.n6 8.03383
R36 A.n11 A.n10 8.03383
R37 A.n21 A.n12 7.30353
R38 A A.n22 5.65631
R39 A.n21 A.n20 5.11262
R40 A A.n0 4.46562
R41 A.n17 A 2.67957
R42 A.n18 A 1.48887
R43 A.n14 A.n13 1.43996
R44 A.n3 A.n2 0.730803
R45 VPWR.n4 VPWR.n3 323.406
R46 VPWR.n13 VPWR.n2 315.928
R47 VPWR.n5 VPWR.t4 265.531
R48 VPWR.n15 VPWR.t7 259.171
R49 VPWR.n7 VPWR.n6 223.696
R50 VPWR.n2 VPWR.t1 35.1791
R51 VPWR.n6 VPWR.t3 35.1791
R52 VPWR.n12 VPWR.n4 27.4829
R53 VPWR.n15 VPWR.n14 26.7299
R54 VPWR.n2 VPWR.t0 26.3844
R55 VPWR.n3 VPWR.t5 26.3844
R56 VPWR.n3 VPWR.t2 26.3844
R57 VPWR.n6 VPWR.t6 26.3844
R58 VPWR.n8 VPWR.n4 25.977
R59 VPWR.n13 VPWR.n12 25.224
R60 VPWR.n14 VPWR.n13 22.2123
R61 VPWR.n8 VPWR.n7 16.9417
R62 VPWR.n9 VPWR.n8 9.3005
R63 VPWR.n10 VPWR.n4 9.3005
R64 VPWR.n12 VPWR.n11 9.3005
R65 VPWR.n13 VPWR.n1 9.3005
R66 VPWR.n14 VPWR.n0 9.3005
R67 VPWR.n16 VPWR.n15 9.3005
R68 VPWR.n7 VPWR.n5 6.98721
R69 VPWR.n9 VPWR.n5 0.596295
R70 VPWR.n10 VPWR.n9 0.122949
R71 VPWR.n11 VPWR.n10 0.122949
R72 VPWR.n11 VPWR.n1 0.122949
R73 VPWR.n1 VPWR.n0 0.122949
R74 VPWR.n16 VPWR.n0 0.122949
R75 VPWR VPWR.n16 0.0617245
R76 Y.n5 Y.n3 261.483
R77 Y.n14 Y.n0 217.879
R78 Y.n6 Y.n2 207.349
R79 Y.n5 Y.n4 205.487
R80 Y.n10 Y.n9 162.933
R81 Y.n11 Y.n10 123.76
R82 Y.n13 Y.n1 106.343
R83 Y.n10 Y.n8 103.65
R84 Y.n11 Y.n7 95.3729
R85 Y.n6 Y.n5 55.3417
R86 Y.n12 Y.n6 41.453
R87 Y.n12 Y.n11 33.0223
R88 Y.n2 Y.t11 26.3844
R89 Y.n2 Y.t10 26.3844
R90 Y.n3 Y.t7 26.3844
R91 Y.n3 Y.t12 26.3844
R92 Y.n4 Y.t9 26.3844
R93 Y.n4 Y.t8 26.3844
R94 Y.n0 Y.t6 26.3844
R95 Y.n0 Y.t5 26.3844
R96 Y.n7 Y.t0 22.7032
R97 Y.n7 Y.t14 22.7032
R98 Y.n9 Y.t3 22.7032
R99 Y.n9 Y.t15 22.7032
R100 Y.n8 Y.t4 22.7032
R101 Y.n8 Y.t1 22.7032
R102 Y.n1 Y.t13 22.7032
R103 Y.n1 Y.t2 22.7032
R104 Y.n13 Y.n12 21.3338
R105 Y Y.n14 12.4005
R106 Y.n14 Y.n13 1.33383
R107 VPB VPB.t7 257.93
R108 VPB.t6 VPB.t0 255.376
R109 VPB.t2 VPB.t3 255.376
R110 VPB.t0 VPB.t1 229.839
R111 VPB.t5 VPB.t6 229.839
R112 VPB.t4 VPB.t5 229.839
R113 VPB.t3 VPB.t4 229.839
R114 VPB.t7 VPB.t2 229.839
R115 VGND.n9 VGND.n8 211.183
R116 VGND.n13 VGND.n2 211.183
R117 VGND.n15 VGND.t7 171.77
R118 VGND.n4 VGND.t5 160.25
R119 VGND.n6 VGND.n5 115.245
R120 VGND.n9 VGND.n7 34.6358
R121 VGND.n5 VGND.t2 34.0546
R122 VGND.n5 VGND.t0 34.0546
R123 VGND.n8 VGND.t6 34.0546
R124 VGND.n13 VGND.n1 27.1064
R125 VGND.n15 VGND.n14 25.6005
R126 VGND.n8 VGND.t4 22.7032
R127 VGND.n2 VGND.t1 22.7032
R128 VGND.n2 VGND.t3 22.7032
R129 VGND.n14 VGND.n13 20.3299
R130 VGND.n7 VGND.n6 15.8123
R131 VGND.n9 VGND.n1 12.8005
R132 VGND.n16 VGND.n15 9.3005
R133 VGND.n7 VGND.n3 9.3005
R134 VGND.n10 VGND.n9 9.3005
R135 VGND.n11 VGND.n1 9.3005
R136 VGND.n13 VGND.n12 9.3005
R137 VGND.n14 VGND.n0 9.3005
R138 VGND.n6 VGND.n4 6.93285
R139 VGND.n4 VGND.n3 0.677147
R140 VGND.n10 VGND.n3 0.122949
R141 VGND.n11 VGND.n10 0.122949
R142 VGND.n12 VGND.n11 0.122949
R143 VGND.n12 VGND.n0 0.122949
R144 VGND.n16 VGND.n0 0.122949
R145 VGND VGND.n16 0.0617245
R146 VNB.t0 VNB.t2 1316.54
R147 VNB VNB.t7 1177.95
R148 VNB.t4 VNB.t6 1154.86
R149 VNB.t2 VNB.t5 993.177
R150 VNB.t6 VNB.t0 993.177
R151 VNB.t1 VNB.t4 993.177
R152 VNB.t3 VNB.t1 993.177
R153 VNB.t7 VNB.t3 993.177
C0 VPB Y 0.020569f
C1 VGND Y 0.66808f
C2 A VPWR 0.174992f
C3 A VPB 0.29059f
C4 A VGND 0.141994f
C5 VPB VPWR 0.138167f
C6 A Y 0.664082f
C7 VPWR VGND 0.085813f
C8 VPB VGND 0.007616f
C9 VPWR Y 0.856977f
C10 VGND VNB 0.59851f
C11 Y VNB 0.083993f
C12 VPWR VNB 0.502892f
C13 A VNB 0.881288f
C14 VPB VNB 1.04904f
.ends


* NGSPICE file created from sky130_fd_sc_hs__inv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y
X0 Y.t31 A.t0 VPWR.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1 Y.t30 A.t1 VPWR.t4 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t3 A.t2 Y.t29 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t28 A.t3 VPWR.t2 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X4 Y.t2 A.t4 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 VGND.t14 A.t5 Y.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 Y.t27 A.t6 VPWR.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.1792 ps=1.44 w=1.12 l=0.15
X7 VGND.t13 A.t7 Y.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t0 A.t8 Y.t26 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.1848 ps=1.45 w=1.12 l=0.15
X9 VPWR.t11 A.t9 Y.t25 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t24 A.t10 VPWR.t10 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X11 Y.t5 A.t11 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X12 VGND.t11 A.t12 Y.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VGND.t10 A.t13 Y.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t9 A.t14 Y.t23 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Y.t15 A.t15 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 Y.t22 A.t16 VPWR.t8 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 VGND.t8 A.t17 Y.t14 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VPWR.t7 A.t18 Y.t21 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t13 A.t19 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X20 VPWR.t6 A.t20 Y.t20 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X21 Y.t19 A.t21 VPWR.t13 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X22 VPWR.t12 A.t22 Y.t18 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X23 VGND.t6 A.t23 Y.t11 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 Y.t17 A.t24 VPWR.t15 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X25 VGND.t5 A.t25 Y.t10 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 Y.t9 A.t26 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 VGND.t3 A.t27 Y.t8 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 Y.t7 A.t28 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X29 VPWR.t14 A.t29 Y.t16 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X30 Y.t6 A.t30 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X31 Y.t12 A.t31 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1628 ps=1.18 w=0.74 l=0.15
R0 A.n4 A.t2 235.571
R1 A.n36 A.t1 235.571
R2 A.n5 A.t3 226.809
R3 A.n9 A.t22 226.809
R4 A.n7 A.t24 226.809
R5 A.n13 A.t8 226.809
R6 A.n15 A.t6 226.809
R7 A.n18 A.t14 226.809
R8 A.n20 A.t16 226.809
R9 A.n23 A.t18 226.809
R10 A.n1 A.t21 226.809
R11 A.n28 A.t29 226.809
R12 A.n30 A.t0 226.809
R13 A.n33 A.t9 226.809
R14 A.n35 A.t10 226.809
R15 A.n37 A.t20 226.809
R16 A.n1 A.t28 196.013
R17 A.n28 A.t5 196.013
R18 A.n36 A.t11 196.013
R19 A.n38 A.t25 196.013
R20 A.n34 A.t15 196.013
R21 A.n32 A.t7 196.013
R22 A.n29 A.t30 196.013
R23 A.n22 A.t17 196.013
R24 A.n21 A.t26 196.013
R25 A.n19 A.t13 196.013
R26 A.n16 A.t4 196.013
R27 A.n14 A.t27 196.013
R28 A.n3 A.t19 196.013
R29 A.n8 A.t12 196.013
R30 A.n6 A.t31 196.013
R31 A.n4 A.t23 196.013
R32 A.n27 A.n26 168.282
R33 A.n25 A.n24 168.157
R34 A.n31 A.n0 167.922
R35 A.n11 A.n10 167.841
R36 A.n40 A.n39 167.494
R37 A.n17 A.n2 167.395
R38 A.n12 A.n11 167.031
R39 A.n22 A.n1 62.8066
R40 A.n29 A.n28 62.8066
R41 A.n34 A.n33 59.8853
R42 A.n15 A.n14 58.4247
R43 A.n5 A.n4 56.9641
R44 A.n20 A.n19 56.9641
R45 A.n37 A.n36 56.9641
R46 A.n8 A.n7 54.0429
R47 A.n13 A.n12 40.1672
R48 A.n10 A.n9 39.4369
R49 A.n28 A.n27 37.246
R50 A.n27 A.n1 35.7853
R51 A.n32 A.n31 35.7853
R52 A.n10 A.n6 35.055
R53 A.n31 A.n30 34.3247
R54 A.n39 A.n38 34.3247
R55 A.n18 A.n17 33.5944
R56 A.n39 A.n35 32.8641
R57 A.n24 A.n23 32.1338
R58 A.n12 A.n3 31.4035
R59 A.n17 A.n16 30.6732
R60 A.n24 A.n21 27.752
R61 A.n9 A.n8 11.6853
R62 A.n14 A.n13 11.6853
R63 A.n7 A.n3 8.76414
R64 A.n19 A.n18 8.76414
R65 A.n6 A.n5 5.84292
R66 A.n21 A.n20 5.84292
R67 A.n35 A.n34 5.84292
R68 A.n38 A.n37 5.84292
R69 A.n16 A.n15 4.38232
R70 A.n23 A.n22 2.92171
R71 A.n30 A.n29 2.92171
R72 A.n33 A.n32 2.92171
R73 A.n11 A.n2 0.541261
R74 A.n26 A.n0 0.51137
R75 A.n40 A.n0 0.51137
R76 A.n26 A.n25 0.497783
R77 A.n25 A.n2 0.495065
R78 A A.n40 0.0793043
R79 VPWR.n35 VPWR.t4 259.171
R80 VPWR.n13 VPWR.t3 258.68
R81 VPWR.n8 VPWR.n7 233.734
R82 VPWR.n4 VPWR.n3 231.429
R83 VPWR.n27 VPWR.n6 231.429
R84 VPWR.n21 VPWR.n10 226.987
R85 VPWR.n33 VPWR.n2 226.439
R86 VPWR.n12 VPWR.n11 222.651
R87 VPWR.n15 VPWR.n14 222.651
R88 VPWR.n2 VPWR.t10 35.1791
R89 VPWR.n3 VPWR.t5 35.1791
R90 VPWR.n6 VPWR.t13 35.1791
R91 VPWR.n11 VPWR.t15 35.1791
R92 VPWR.n11 VPWR.t0 35.1791
R93 VPWR.n14 VPWR.t2 35.1791
R94 VPWR.n14 VPWR.t12 35.1791
R95 VPWR.n21 VPWR.n20 32.0005
R96 VPWR.n22 VPWR.n8 30.8711
R97 VPWR.n10 VPWR.t1 29.9023
R98 VPWR.n16 VPWR.n12 28.9887
R99 VPWR.n32 VPWR.n4 27.4829
R100 VPWR.n35 VPWR.n34 26.7299
R101 VPWR.n28 VPWR.n27 26.7299
R102 VPWR.n27 VPWR.n26 26.7299
R103 VPWR.n2 VPWR.t6 26.3844
R104 VPWR.n3 VPWR.t11 26.3844
R105 VPWR.n6 VPWR.t14 26.3844
R106 VPWR.n7 VPWR.t8 26.3844
R107 VPWR.n7 VPWR.t7 26.3844
R108 VPWR.n10 VPWR.t9 26.3844
R109 VPWR.n28 VPWR.n4 25.977
R110 VPWR.n34 VPWR.n33 25.224
R111 VPWR.n33 VPWR.n32 25.224
R112 VPWR.n26 VPWR.n8 23.7181
R113 VPWR.n16 VPWR.n15 21.4593
R114 VPWR.n22 VPWR.n21 18.824
R115 VPWR.n20 VPWR.n12 18.4476
R116 VPWR.n17 VPWR.n16 9.3005
R117 VPWR.n18 VPWR.n12 9.3005
R118 VPWR.n20 VPWR.n19 9.3005
R119 VPWR.n21 VPWR.n9 9.3005
R120 VPWR.n23 VPWR.n22 9.3005
R121 VPWR.n24 VPWR.n8 9.3005
R122 VPWR.n26 VPWR.n25 9.3005
R123 VPWR.n27 VPWR.n5 9.3005
R124 VPWR.n29 VPWR.n28 9.3005
R125 VPWR.n30 VPWR.n4 9.3005
R126 VPWR.n32 VPWR.n31 9.3005
R127 VPWR.n33 VPWR.n1 9.3005
R128 VPWR.n34 VPWR.n0 9.3005
R129 VPWR.n36 VPWR.n35 9.3005
R130 VPWR.n15 VPWR.n13 6.77577
R131 VPWR.n17 VPWR.n13 0.617781
R132 VPWR.n18 VPWR.n17 0.122949
R133 VPWR.n19 VPWR.n18 0.122949
R134 VPWR.n19 VPWR.n9 0.122949
R135 VPWR.n23 VPWR.n9 0.122949
R136 VPWR.n24 VPWR.n23 0.122949
R137 VPWR.n25 VPWR.n24 0.122949
R138 VPWR.n25 VPWR.n5 0.122949
R139 VPWR.n29 VPWR.n5 0.122949
R140 VPWR.n30 VPWR.n29 0.122949
R141 VPWR.n31 VPWR.n30 0.122949
R142 VPWR.n31 VPWR.n1 0.122949
R143 VPWR.n1 VPWR.n0 0.122949
R144 VPWR.n36 VPWR.n0 0.122949
R145 VPWR VPWR.n36 0.0617245
R146 Y.n2 Y.n1 203.748
R147 Y.n13 Y.n12 203.454
R148 Y.n17 Y.n16 203.315
R149 Y.n25 Y.n24 203.056
R150 Y.n9 Y.n8 202.802
R151 Y.n29 Y.n27 202.684
R152 Y.n21 Y.n20 202.457
R153 Y.n5 Y.n4 202.457
R154 Y.n13 Y.n11 150.185
R155 Y.n25 Y.n23 143.799
R156 Y.n2 Y.n0 143.638
R157 Y.n17 Y.n15 142.806
R158 Y.n9 Y.n7 140.738
R159 Y.n21 Y.n19 140.192
R160 Y.n29 Y.n28 140.054
R161 Y.n5 Y.n3 138.594
R162 Y.n8 Y.t27 31.6612
R163 Y.n27 Y.t20 26.3844
R164 Y.n27 Y.t30 26.3844
R165 Y.n24 Y.t25 26.3844
R166 Y.n24 Y.t24 26.3844
R167 Y.n20 Y.t16 26.3844
R168 Y.n20 Y.t31 26.3844
R169 Y.n16 Y.t21 26.3844
R170 Y.n16 Y.t19 26.3844
R171 Y.n12 Y.t23 26.3844
R172 Y.n12 Y.t22 26.3844
R173 Y.n8 Y.t26 26.3844
R174 Y.n4 Y.t18 26.3844
R175 Y.n4 Y.t17 26.3844
R176 Y.n1 Y.t29 26.3844
R177 Y.n1 Y.t28 26.3844
R178 Y.n28 Y.t10 22.7032
R179 Y.n28 Y.t5 22.7032
R180 Y.n23 Y.t0 22.7032
R181 Y.n23 Y.t15 22.7032
R182 Y.n19 Y.t1 22.7032
R183 Y.n19 Y.t6 22.7032
R184 Y.n15 Y.t14 22.7032
R185 Y.n15 Y.t7 22.7032
R186 Y.n11 Y.t3 22.7032
R187 Y.n11 Y.t9 22.7032
R188 Y.n7 Y.t8 22.7032
R189 Y.n7 Y.t2 22.7032
R190 Y.n3 Y.t4 22.7032
R191 Y.n3 Y.t13 22.7032
R192 Y.n0 Y.t11 22.7032
R193 Y.n0 Y.t12 22.7032
R194 Y.n6 Y.n2 10.6406
R195 Y.n14 Y.n13 10.0685
R196 Y.n18 Y.n17 10.055
R197 Y.n10 Y.n9 10.0053
R198 Y.n30 Y.n29 9.99393
R199 Y.n22 Y.n21 9.97218
R200 Y.n6 Y.n5 9.97218
R201 Y.n26 Y.n25 9.43563
R202 Y.n10 Y.n6 0.543978
R203 Y.n14 Y.n10 0.516804
R204 Y.n22 Y.n18 0.516804
R205 Y.n26 Y.n22 0.516804
R206 Y.n30 Y.n26 0.516804
R207 Y.n18 Y.n14 0.48963
R208 Y Y.n30 0.0793043
R209 VPB.t2 VPB.t12 280.914
R210 VPB.t10 VPB.t1 280.914
R211 VPB VPB.t14 257.93
R212 VPB.t0 VPB.t3 255.376
R213 VPB.t9 VPB.t15 255.376
R214 VPB.t4 VPB.t8 255.376
R215 VPB.t11 VPB.t10 245.161
R216 VPB.t7 VPB.t11 240.054
R217 VPB.t12 VPB.t13 229.839
R218 VPB.t1 VPB.t2 229.839
R219 VPB.t6 VPB.t7 229.839
R220 VPB.t5 VPB.t6 229.839
R221 VPB.t3 VPB.t5 229.839
R222 VPB.t15 VPB.t0 229.839
R223 VPB.t8 VPB.t9 229.839
R224 VPB.t14 VPB.t4 229.839
R225 VGND.n9 VGND.t6 174.359
R226 VGND.n36 VGND.t12 174.131
R227 VGND.n20 VGND.n19 123.653
R228 VGND.n23 VGND.n22 123.079
R229 VGND.n34 VGND.n2 123.079
R230 VGND.n27 VGND.n5 121.957
R231 VGND.n30 VGND.n29 120.915
R232 VGND.n14 VGND.n13 117.856
R233 VGND.n11 VGND.n10 116.374
R234 VGND.n18 VGND.n7 36.1417
R235 VGND.n10 VGND.t0 35.6762
R236 VGND.n10 VGND.t11 35.6762
R237 VGND.n14 VGND.n12 34.2593
R238 VGND.n13 VGND.t7 34.0546
R239 VGND.n13 VGND.t3 34.0546
R240 VGND.n29 VGND.t1 34.0546
R241 VGND.n2 VGND.t5 34.0546
R242 VGND.n23 VGND.n21 30.8711
R243 VGND.n5 VGND.t14 30.8113
R244 VGND.n35 VGND.n34 29.7417
R245 VGND.n19 VGND.t15 28.3789
R246 VGND.n19 VGND.t10 28.3789
R247 VGND.n27 VGND.n4 26.7299
R248 VGND.n30 VGND.n1 25.977
R249 VGND.n5 VGND.t2 25.9464
R250 VGND.n28 VGND.n27 25.224
R251 VGND.n30 VGND.n28 25.224
R252 VGND.n34 VGND.n1 22.9652
R253 VGND.n22 VGND.t4 22.7032
R254 VGND.n22 VGND.t8 22.7032
R255 VGND.n29 VGND.t13 22.7032
R256 VGND.n2 VGND.t9 22.7032
R257 VGND.n23 VGND.n4 21.8358
R258 VGND.n36 VGND.n35 20.7064
R259 VGND.n12 VGND.n11 16.9417
R260 VGND.n21 VGND.n20 15.4358
R261 VGND.n14 VGND.n7 13.9299
R262 VGND.n37 VGND.n36 9.3005
R263 VGND.n12 VGND.n8 9.3005
R264 VGND.n15 VGND.n14 9.3005
R265 VGND.n16 VGND.n7 9.3005
R266 VGND.n18 VGND.n17 9.3005
R267 VGND.n21 VGND.n6 9.3005
R268 VGND.n24 VGND.n23 9.3005
R269 VGND.n25 VGND.n4 9.3005
R270 VGND.n27 VGND.n26 9.3005
R271 VGND.n28 VGND.n3 9.3005
R272 VGND.n31 VGND.n30 9.3005
R273 VGND.n32 VGND.n1 9.3005
R274 VGND.n34 VGND.n33 9.3005
R275 VGND.n35 VGND.n0 9.3005
R276 VGND.n11 VGND.n9 6.96039
R277 VGND.n20 VGND.n18 1.12991
R278 VGND.n9 VGND.n8 0.594857
R279 VGND.n15 VGND.n8 0.122949
R280 VGND.n16 VGND.n15 0.122949
R281 VGND.n17 VGND.n16 0.122949
R282 VGND.n17 VGND.n6 0.122949
R283 VGND.n24 VGND.n6 0.122949
R284 VGND.n25 VGND.n24 0.122949
R285 VGND.n26 VGND.n25 0.122949
R286 VGND.n26 VGND.n3 0.122949
R287 VGND.n31 VGND.n3 0.122949
R288 VGND.n32 VGND.n31 0.122949
R289 VGND.n33 VGND.n32 0.122949
R290 VGND.n33 VGND.n0 0.122949
R291 VGND.n37 VGND.n0 0.122949
R292 VGND VGND.n37 0.0617245
R293 VNB.t11 VNB.t0 1362.73
R294 VNB.t3 VNB.t7 1316.54
R295 VNB VNB.t12 1304.99
R296 VNB.t10 VNB.t15 1154.86
R297 VNB.t14 VNB.t2 1154.86
R298 VNB.t13 VNB.t1 1154.86
R299 VNB.t5 VNB.t9 1154.86
R300 VNB.t0 VNB.t6 993.177
R301 VNB.t7 VNB.t11 993.177
R302 VNB.t15 VNB.t3 993.177
R303 VNB.t4 VNB.t10 993.177
R304 VNB.t8 VNB.t4 993.177
R305 VNB.t2 VNB.t8 993.177
R306 VNB.t1 VNB.t14 993.177
R307 VNB.t9 VNB.t13 993.177
R308 VNB.t12 VNB.t5 993.177
C0 Y VPB 0.045372f
C1 VGND VPWR 0.064897f
C2 VPWR A 0.529164f
C3 VPWR Y 2.08315f
C4 VGND A 0.686864f
C5 VPWR VPB 0.231595f
C6 VGND Y 1.31768f
C7 VGND VPB 0.008245f
C8 A Y 2.0772f
C9 A VPB 0.601473f
C10 VGND VNB 1.02743f
C11 Y VNB 0.09351f
C12 VPWR VNB 0.825774f
C13 A VNB 1.727695f
C14 VPB VNB 1.90613f
C15 Y.t11 VNB 0.017533f
C16 Y.t12 VNB 0.017533f
C17 Y.n0 VNB 0.077558f
C18 Y.t29 VNB 0.028432f
C19 Y.t28 VNB 0.028432f
C20 Y.n1 VNB 0.061755f
C21 Y.n2 VNB 0.211114f
C22 Y.t4 VNB 0.017533f
C23 Y.t13 VNB 0.017533f
C24 Y.n3 VNB 0.075471f
C25 Y.t18 VNB 0.028432f
C26 Y.t17 VNB 0.028432f
C27 Y.n4 VNB 0.061808f
C28 Y.n5 VNB 0.238955f
C29 Y.n6 VNB 0.138977f
C30 Y.t8 VNB 0.017533f
C31 Y.t2 VNB 0.017533f
C32 Y.n7 VNB 0.074431f
C33 Y.t26 VNB 0.028432f
C34 Y.t27 VNB 0.034118f
C35 Y.n8 VNB 0.067479f
C36 Y.n9 VNB 0.225797f
C37 Y.n10 VNB 0.082839f
C38 Y.t3 VNB 0.017533f
C39 Y.t9 VNB 0.017533f
C40 Y.n11 VNB 0.071679f
C41 Y.t23 VNB 0.028432f
C42 Y.t22 VNB 0.028432f
C43 Y.n12 VNB 0.061767f
C44 Y.n13 VNB 0.190901f
C45 Y.n14 VNB 0.078899f
C46 Y.t14 VNB 0.017533f
C47 Y.t7 VNB 0.017533f
C48 Y.n15 VNB 0.074045f
C49 Y.t21 VNB 0.028432f
C50 Y.t19 VNB 0.028432f
C51 Y.n16 VNB 0.061772f
C52 Y.n17 VNB 0.2118f
C53 Y.n18 VNB 0.078908f
C54 Y.t1 VNB 0.017533f
C55 Y.t6 VNB 0.017533f
C56 Y.n19 VNB 0.074551f
C57 Y.t16 VNB 0.028432f
C58 Y.t31 VNB 0.028432f
C59 Y.n20 VNB 0.061808f
C60 Y.n21 VNB 0.2316f
C61 Y.n22 VNB 0.080921f
C62 Y.t0 VNB 0.017533f
C63 Y.t15 VNB 0.017533f
C64 Y.n23 VNB 0.073941f
C65 Y.t25 VNB 0.028432f
C66 Y.t24 VNB 0.028432f
C67 Y.n24 VNB 0.06188f
C68 Y.n25 VNB 0.226892f
C69 Y.n26 VNB 0.075404f
C70 Y.t20 VNB 0.028432f
C71 Y.t30 VNB 0.028432f
C72 Y.n27 VNB 0.061918f
C73 Y.t10 VNB 0.017533f
C74 Y.t5 VNB 0.017533f
C75 Y.n28 VNB 0.075754f
C76 Y.n29 VNB 0.232942f
C77 Y.n30 VNB 0.049674f
C78 VPWR.n0 VNB 0.040808f
C79 VPWR.t4 VNB 0.060735f
C80 VPWR.n1 VNB 0.040808f
C81 VPWR.t10 VNB 0.019433f
C82 VPWR.t6 VNB 0.014574f
C83 VPWR.n2 VNB 0.041719f
C84 VPWR.t5 VNB 0.019433f
C85 VPWR.t11 VNB 0.014574f
C86 VPWR.n3 VNB 0.041545f
C87 VPWR.n4 VNB 0.066913f
C88 VPWR.n5 VNB 0.040808f
C89 VPWR.t13 VNB 0.019433f
C90 VPWR.t14 VNB 0.014574f
C91 VPWR.n6 VNB 0.041545f
C92 VPWR.t8 VNB 0.014574f
C93 VPWR.t7 VNB 0.014574f
C94 VPWR.n7 VNB 0.036609f
C95 VPWR.n8 VNB 0.063369f
C96 VPWR.n9 VNB 0.040808f
C97 VPWR.t1 VNB 0.016518f
C98 VPWR.t9 VNB 0.014574f
C99 VPWR.n10 VNB 0.038784f
C100 VPWR.t15 VNB 0.019433f
C101 VPWR.t0 VNB 0.019433f
C102 VPWR.n11 VNB 0.046714f
C103 VPWR.n12 VNB 0.085896f
C104 VPWR.t3 VNB 0.063115f
C105 VPWR.n13 VNB 0.117088f
C106 VPWR.t2 VNB 0.019433f
C107 VPWR.t12 VNB 0.019433f
C108 VPWR.n14 VNB 0.046714f
C109 VPWR.n15 VNB 0.087431f
C110 VPWR.n16 VNB 0.009881f
C111 VPWR.n17 VNB 0.135007f
C112 VPWR.n18 VNB 0.040808f
C113 VPWR.n19 VNB 0.040808f
C114 VPWR.n20 VNB 0.009881f
C115 VPWR.n21 VNB 0.075195f
C116 VPWR.n22 VNB 0.009734f
C117 VPWR.n23 VNB 0.040808f
C118 VPWR.n24 VNB 0.040808f
C119 VPWR.n25 VNB 0.040808f
C120 VPWR.n26 VNB 0.009881f
C121 VPWR.n27 VNB 0.066913f
C122 VPWR.n28 VNB 0.010323f
C123 VPWR.n29 VNB 0.040808f
C124 VPWR.n30 VNB 0.040808f
C125 VPWR.n31 VNB 0.040808f
C126 VPWR.n32 VNB 0.010323f
C127 VPWR.n33 VNB 0.076386f
C128 VPWR.n34 VNB 0.010176f
C129 VPWR.n35 VNB 0.06762f
C130 VPWR.n36 VNB 0.030606f
C131 A.n0 VNB 0.072399f
C132 A.t10 VNB 0.025933f
C133 A.t15 VNB 0.018017f
C134 A.t9 VNB 0.025933f
C135 A.t7 VNB 0.018017f
C136 A.t0 VNB 0.025933f
C137 A.t30 VNB 0.018017f
C138 A.t29 VNB 0.025933f
C139 A.t5 VNB 0.018017f
C140 A.t21 VNB 0.025933f
C141 A.t28 VNB 0.018017f
C142 A.n1 VNB 0.047273f
C143 A.n2 VNB 0.075212f
C144 A.t26 VNB 0.018017f
C145 A.t16 VNB 0.025933f
C146 A.t13 VNB 0.018017f
C147 A.t14 VNB 0.025933f
C148 A.t4 VNB 0.018017f
C149 A.t6 VNB 0.025933f
C150 A.t27 VNB 0.018017f
C151 A.t8 VNB 0.025933f
C152 A.t19 VNB 0.018017f
C153 A.n3 VNB 0.020083f
C154 A.t31 VNB 0.018017f
C155 A.t3 VNB 0.025933f
C156 A.t23 VNB 0.018017f
C157 A.t2 VNB 0.026728f
C158 A.n4 VNB 0.047024f
C159 A.n5 VNB 0.028282f
C160 A.n6 VNB 0.020264f
C161 A.t22 VNB 0.025933f
C162 A.t12 VNB 0.018017f
C163 A.t24 VNB 0.025933f
C164 A.n7 VNB 0.028282f
C165 A.n8 VNB 0.026446f
C166 A.n9 VNB 0.025372f
C167 A.n10 VNB 0.020992f
C168 A.n11 VNB 0.13885f
C169 A.n12 VNB 0.020153f
C170 A.n13 VNB 0.025554f
C171 A.n14 VNB 0.027537f
C172 A.n15 VNB 0.028282f
C173 A.n16 VNB 0.01881f
C174 A.n17 VNB 0.018227f
C175 A.n18 VNB 0.023191f
C176 A.n19 VNB 0.026446f
C177 A.n20 VNB 0.028282f
C178 A.n21 VNB 0.018446f
C179 A.t18 VNB 0.025933f
C180 A.t17 VNB 0.018017f
C181 A.n22 VNB 0.026446f
C182 A.n23 VNB 0.021372f
C183 A.n24 VNB 0.016946f
C184 A.n25 VNB 0.070133f
C185 A.n26 VNB 0.070458f
C186 A.n27 VNB 0.020192f
C187 A.n28 VNB 0.047637f
C188 A.n29 VNB 0.026446f
C189 A.n30 VNB 0.021918f
C190 A.n31 VNB 0.019546f
C191 A.n32 VNB 0.019719f
C192 A.n33 VNB 0.028282f
C193 A.n34 VNB 0.026446f
C194 A.n35 VNB 0.022282f
C195 A.t25 VNB 0.018017f
C196 A.t20 VNB 0.025933f
C197 A.t11 VNB 0.018017f
C198 A.t1 VNB 0.026728f
C199 A.n36 VNB 0.047024f
C200 A.n37 VNB 0.028282f
C201 A.n38 VNB 0.020083f
C202 A.n39 VNB 0.018927f
C203 A.n40 VNB 0.053993f
.ends


* NGSPICE file created from sky130_fd_sc_hs__sdfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrbp_2 VNB VPB VPWR RESET_B VGND D CLK SCE SCD Q Q_N
X0 VGND.t9 SCE.t0 a_27_79.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=1.39 as=0.1197 ps=1.41 w=0.42 l=0.15
X1 a_2000_74.t0 a_852_74.t2 a_1790_74.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.2165 ps=1.54 w=0.42 l=0.15
X2 a_1790_74.t1 a_852_74.t3 a_1370_289.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.20145 pd=1.64 as=0.15 ps=1.3 w=1 l=0.15
X3 VPWR.t4 a_1790_74.t3 Q_N.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_547_79.t1 SCE.t1 a_388_79.t4 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.13545 ps=1.065 w=0.42 l=0.15
X5 VGND.t8 CLK.t0 a_852_74.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 Q_N.t1 a_1790_74.t4 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1771 ps=1.505 w=1.12 l=0.15
X7 VPWR.t5 a_1790_74.t5 a_2006_373.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1771 pd=1.505 as=0.063 ps=0.72 w=0.42 l=0.15
X8 a_388_79.t1 D.t0 a_310_79.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.13545 pd=1.065 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 a_2006_373.t1 a_1790_74.t6 a_2158_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_310_79.t0 a_27_79.t2 a_223_79.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X11 a_1790_74.t2 a_1025_74.t2 a_1370_289.t2 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.2165 pd=1.54 as=0.0896 ps=0.92 w=0.64 l=0.15
X12 VPWR.t8 SCE.t2 a_27_79.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2576 pd=1.445 as=0.1888 ps=1.87 w=0.64 l=0.15
X13 a_1325_457# a_852_74.t4 a_1223_118# VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X14 VPWR.t7 CLK.t1 a_852_74.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X15 VGND.t10 a_2006_373.t2 a_2000_74.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_1025_74.t0 a_852_74.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_1401_118.t0 a_1370_289.t3 a_1323_118.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X18 VPWR.t10 SCD.t0 a_538_464.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 VGND.t2 RESET_B.t0 a_223_79.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0819 ps=0.81 w=0.42 l=0.15
X20 a_223_79.t2 SCD.t1 a_547_79.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X21 a_2158_74.t0 RESET_B.t1 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 a_1370_289.t1 a_1223_118# VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.350775 ps=1.805 w=0.64 l=0.15
X23 VGND.t0 a_2604_392.t2 Q.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_388_79.t2 D.t1 a_307_464.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1872 pd=1.225 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_2604_392.t1 a_1790_74.t7 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1165 ps=1.065 w=0.64 l=0.15
X26 a_307_464.t1 SCE.t3 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.2576 ps=1.445 w=0.64 l=0.15
X27 a_1025_74.t1 a_852_74.t6 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VGND.t7 a_1790_74.t8 Q_N.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 a_538_464.t0 a_27_79.t3 a_388_79.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1872 ps=1.225 w=0.64 l=0.15
X30 a_1223_118# RESET_B.t2 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.127675 ps=1.14 w=0.42 l=0.15
X31 Q.t2 a_2604_392.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2183 ps=2.07 w=0.74 l=0.15
X32 VPWR.t11 a_2604_392.t4 Q.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X33 a_388_79.t3 RESET_B.t3 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1344 ps=1.06 w=0.64 l=0.15
X34 a_2604_392.t0 a_1790_74.t9 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.1934 ps=1.475 w=1 l=0.15
X35 Q.t0 a_2604_392.t5 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 SCE SCE.t1 458.072
R1 SCE.n0 SCE.t0 404.212
R2 SCE.n5 SCE.t3 163.321
R3 SCE.n0 SCE.t2 152.367
R4 SCE.n6 SCE.n5 152
R5 SCE.n4 SCE.n3 152
R6 SCE.n2 SCE.n1 152
R7 SCE.n5 SCE.n4 49.6611
R8 SCE.n4 SCE.n1 49.6611
R9 SCE.n1 SCE.n0 29.2126
R10 SCE.n3 SCE.n2 13.1884
R11 SCE.n6 SCE 10.4732
R12 SCE SCE.n6 8.14595
R13 SCE.n3 SCE 2.71565
R14 SCE.n2 SCE 2.71565
R15 a_27_79.t0 a_27_79.n1 640.676
R16 a_27_79.n1 a_27_79.t3 480.94
R17 a_27_79.n0 a_27_79.t2 359.063
R18 a_27_79.n0 a_27_79.t1 258.024
R19 a_27_79.n1 a_27_79.n0 60.5666
R20 VGND.n38 VGND.t5 318.723
R21 VGND.n3 VGND.t2 248.468
R22 VGND.n63 VGND.t9 248.468
R23 VGND.n30 VGND.n29 207.498
R24 VGND.n17 VGND.t1 178.623
R25 VGND.n16 VGND.t0 175.919
R26 VGND.n50 VGND.n5 132.637
R27 VGND.n22 VGND.n15 123.335
R28 VGND.n29 VGND.t3 40.0005
R29 VGND.n29 VGND.t10 40.0005
R30 VGND.n18 VGND.n14 36.1417
R31 VGND.n28 VGND.n12 36.1417
R32 VGND.n32 VGND.n31 36.1417
R33 VGND.n32 VGND.n10 36.1417
R34 VGND.n36 VGND.n10 36.1417
R35 VGND.n37 VGND.n36 36.1417
R36 VGND.n43 VGND.n8 36.1417
R37 VGND.n44 VGND.n43 36.1417
R38 VGND.n45 VGND.n44 36.1417
R39 VGND.n45 VGND.n6 36.1417
R40 VGND.n49 VGND.n6 36.1417
R41 VGND.n52 VGND.n51 36.1417
R42 VGND.n56 VGND.n55 36.1417
R43 VGND.n57 VGND.n56 36.1417
R44 VGND.n57 VGND.n1 36.1417
R45 VGND.n61 VGND.n1 36.1417
R46 VGND.n62 VGND.n61 36.1417
R47 VGND.n17 VGND.n16 35.833
R48 VGND.n15 VGND.t6 34.688
R49 VGND.n39 VGND.n37 32.9284
R50 VGND.n23 VGND.n22 29.7417
R51 VGND.n24 VGND.n12 27.4829
R52 VGND.n24 VGND.n23 25.977
R53 VGND.n63 VGND.n62 24.4711
R54 VGND.n22 VGND.n14 22.9652
R55 VGND.n5 VGND.t4 22.7032
R56 VGND.n5 VGND.t8 22.7032
R57 VGND.n15 VGND.t7 22.6611
R58 VGND.n51 VGND.n50 20.7064
R59 VGND.n50 VGND.n49 15.4358
R60 VGND.n30 VGND.n28 10.1652
R61 VGND.n62 VGND.n0 9.3005
R62 VGND.n61 VGND.n60 9.3005
R63 VGND.n59 VGND.n1 9.3005
R64 VGND.n58 VGND.n57 9.3005
R65 VGND.n56 VGND.n2 9.3005
R66 VGND.n55 VGND.n54 9.3005
R67 VGND.n53 VGND.n52 9.3005
R68 VGND.n51 VGND.n4 9.3005
R69 VGND.n49 VGND.n48 9.3005
R70 VGND.n47 VGND.n6 9.3005
R71 VGND.n46 VGND.n45 9.3005
R72 VGND.n44 VGND.n7 9.3005
R73 VGND.n43 VGND.n42 9.3005
R74 VGND.n41 VGND.n8 9.3005
R75 VGND.n40 VGND.n39 9.3005
R76 VGND.n37 VGND.n9 9.3005
R77 VGND.n36 VGND.n35 9.3005
R78 VGND.n34 VGND.n10 9.3005
R79 VGND.n33 VGND.n32 9.3005
R80 VGND.n31 VGND.n11 9.3005
R81 VGND.n28 VGND.n27 9.3005
R82 VGND.n26 VGND.n12 9.3005
R83 VGND.n25 VGND.n24 9.3005
R84 VGND.n23 VGND.n13 9.3005
R85 VGND.n22 VGND.n21 9.3005
R86 VGND.n20 VGND.n14 9.3005
R87 VGND.n19 VGND.n18 9.3005
R88 VGND.n52 VGND.n3 8.28285
R89 VGND.n38 VGND.n8 7.60597
R90 VGND.n64 VGND.n63 7.19894
R91 VGND.n18 VGND.n17 5.64756
R92 VGND.n39 VGND.n38 5.30151
R93 VGND.n55 VGND.n3 3.01226
R94 VGND.n19 VGND.n16 2.11746
R95 VGND.n31 VGND.n30 1.12991
R96 VGND VGND.n64 0.156997
R97 VGND.n64 VGND.n0 0.150766
R98 VGND.n20 VGND.n19 0.122949
R99 VGND.n21 VGND.n20 0.122949
R100 VGND.n21 VGND.n13 0.122949
R101 VGND.n25 VGND.n13 0.122949
R102 VGND.n26 VGND.n25 0.122949
R103 VGND.n27 VGND.n26 0.122949
R104 VGND.n27 VGND.n11 0.122949
R105 VGND.n33 VGND.n11 0.122949
R106 VGND.n34 VGND.n33 0.122949
R107 VGND.n35 VGND.n34 0.122949
R108 VGND.n35 VGND.n9 0.122949
R109 VGND.n40 VGND.n9 0.122949
R110 VGND.n41 VGND.n40 0.122949
R111 VGND.n42 VGND.n41 0.122949
R112 VGND.n42 VGND.n7 0.122949
R113 VGND.n46 VGND.n7 0.122949
R114 VGND.n47 VGND.n46 0.122949
R115 VGND.n48 VGND.n47 0.122949
R116 VGND.n48 VGND.n4 0.122949
R117 VGND.n53 VGND.n4 0.122949
R118 VGND.n54 VGND.n53 0.122949
R119 VGND.n54 VGND.n2 0.122949
R120 VGND.n58 VGND.n2 0.122949
R121 VGND.n59 VGND.n58 0.122949
R122 VGND.n60 VGND.n59 0.122949
R123 VGND.n60 VGND.n0 0.122949
R124 VNB.t12 VNB 28906
R125 VNB.n0 VNB 22645.7
R126 VNB VNB.n1 19482.2
R127 VNB.t4 VNB.t7 4342.26
R128 VNB.t10 VNB.t12 3443.48
R129 VNB.n1 VNB.t4 2402.1
R130 VNB.t13 VNB.t5 2379
R131 VNB.t11 VNB.t2 2263.52
R132 VNB.t0 VNB.t15 2263.52
R133 VNB.t14 VNB.t9 1836.22
R134 VNB.t18 VNB.n0 1454.44
R135 VNB.t5 VNB.t3 1247.24
R136 VNB.n1 VNB.t8 1161.11
R137 VNB.t15 VNB 1143.31
R138 VNB.n0 VNB.t17 1088.04
R139 VNB.t12 VNB.t11 1068.74
R140 VNB.t8 VNB.t18 1051.11
R141 VNB.t16 VNB.t6 1028.26
R142 VNB.t2 VNB.t1 993.177
R143 VNB.t7 VNB.t13 993.177
R144 VNB.t3 VNB.t14 900.788
R145 VNB.t9 VNB.t0 900.788
R146 VNB.t6 VNB.t10 860.87
R147 VNB.t17 VNB.t16 860.87
R148 a_852_74.n0 a_852_74.t3 989.172
R149 a_852_74.t1 a_852_74.n5 893.75
R150 a_852_74.n2 a_852_74.n0 810.563
R151 a_852_74.t3 a_852_74.t2 786.197
R152 a_852_74.n2 a_852_74.n1 277.418
R153 a_852_74.n4 a_852_74.t5 256.264
R154 a_852_74.n3 a_852_74.t6 200.542
R155 a_852_74.n5 a_852_74.t0 194.213
R156 a_852_74.n0 a_852_74.t4 190.659
R157 a_852_74.n5 a_852_74.n4 161.31
R158 a_852_74.n3 a_852_74.n2 59.4472
R159 a_852_74.n4 a_852_74.n3 13.146
R160 a_1790_74.n10 a_1790_74.n9 689.26
R161 a_1790_74.n7 a_1790_74.t5 321.87
R162 a_1790_74.n2 a_1790_74.t9 265.101
R163 a_1790_74.n4 a_1790_74.t3 252.248
R164 a_1790_74.n6 a_1790_74.t4 250.909
R165 a_1790_74.n9 a_1790_74.n0 222.112
R166 a_1790_74.n9 a_1790_74.n8 216.966
R167 a_1790_74.n8 a_1790_74.t6 199.227
R168 a_1790_74.n0 a_1790_74.t2 189.153
R169 a_1790_74.n2 a_1790_74.t7 188.126
R170 a_1790_74.n3 a_1790_74.t8 165.488
R171 a_1790_74.n5 a_1790_74.n1 163.054
R172 a_1790_74.n10 a_1790_74.t1 77.6242
R173 a_1790_74.n8 a_1790_74.n7 67.0667
R174 a_1790_74.n7 a_1790_74.n6 64.0274
R175 a_1790_74.n3 a_1790_74.n2 62.8066
R176 a_1790_74.n0 a_1790_74.t0 55.7148
R177 a_1790_74.n5 a_1790_74.n4 51.3042
R178 a_1790_74.n6 a_1790_74.n5 13.1302
R179 a_1790_74.n4 a_1790_74.n3 10.955
R180 a_1790_74.n11 a_1790_74.n10 4.9255
R181 a_2000_74.t0 a_2000_74.t1 60.0005
R182 a_1370_289.t0 a_1370_289.n3 294.079
R183 a_1370_289.n3 a_1370_289.n1 289.897
R184 a_1370_289.n1 a_1370_289.n0 227
R185 a_1370_289.n1 a_1370_289.t3 226.196
R186 a_1370_289.n3 a_1370_289.n2 185
R187 a_1370_289.n2 a_1370_289.t2 26.2505
R188 a_1370_289.n2 a_1370_289.t1 26.2505
R189 VPB.n0 VPB 6404.84
R190 VPB VPB.n1 3933.25
R191 VPB.t3 VPB.t6 1236.23
R192 VPB.t2 VPB.t1 743.145
R193 VPB.t11 VPB.t10 531.183
R194 VPB.t5 VPB.t16 505.646
R195 VPB.t4 VPB.t2 497.985
R196 VPB.t12 VPB.t13 487.769
R197 VPB.n1 VPB.t3 483.637
R198 VPB.t0 VPB.t9 375.404
R199 VPB.t10 VPB.t14 291.13
R200 VPB.t6 VPB.t7 264.026
R201 VPB.t13 VPB 257.93
R202 VPB.t16 VPB.t15 229.839
R203 VPB.t1 VPB.t11 229.839
R204 VPB.n1 VPB.t4 227.286
R205 VPB.t7 VPB.t8 222.078
R206 VPB.t14 VPB.t0 214.517
R207 VPB.t9 VPB.t12 214.517
R208 VPB.n0 VPB.t5 206.856
R209 VPB.t8 VPB.n0 49.3511
R210 Q_N Q_N.n0 219.493
R211 Q_N.n1 Q_N 197.607
R212 Q_N.n2 Q_N.n1 185
R213 Q_N.n0 Q_N.t2 26.3844
R214 Q_N.n0 Q_N.t1 26.3844
R215 Q_N.n1 Q_N.t0 22.7032
R216 Q_N.n3 Q_N 9.85128
R217 Q_N Q_N.n3 2.2074
R218 Q_N.n3 Q_N.n2 1.93989
R219 Q_N.n2 Q_N 0.970197
R220 VPWR.n40 VPWR.t1 821.179
R221 VPWR.n54 VPWR.n4 606.333
R222 VPWR.n48 VPWR.n7 605.753
R223 VPWR.n61 VPWR.n60 585
R224 VPWR.n63 VPWR.n62 585
R225 VPWR.n19 VPWR.t11 262.053
R226 VPWR.n18 VPWR.t12 250.081
R227 VPWR.n15 VPWR.n14 235.77
R228 VPWR.n22 VPWR.n17 226.459
R229 VPWR.n62 VPWR.n61 140.055
R230 VPWR.n14 VPWR.t5 113.329
R231 VPWR.n4 VPWR.t6 76.9536
R232 VPWR.n62 VPWR.t8 61.563
R233 VPWR.n4 VPWR.t10 52.3286
R234 VPWR.n61 VPWR.t9 46.1724
R235 VPWR.n17 VPWR.t2 40.3855
R236 VPWR.n55 VPWR.n2 36.1417
R237 VPWR.n59 VPWR.n2 36.1417
R238 VPWR.n49 VPWR.n5 36.1417
R239 VPWR.n53 VPWR.n5 36.1417
R240 VPWR.n42 VPWR.n41 36.1417
R241 VPWR.n42 VPWR.n8 36.1417
R242 VPWR.n46 VPWR.n8 36.1417
R243 VPWR.n47 VPWR.n46 36.1417
R244 VPWR.n39 VPWR.n10 36.1417
R245 VPWR.n33 VPWR.n12 36.1417
R246 VPWR.n34 VPWR.n33 36.1417
R247 VPWR.n55 VPWR.n54 35.7652
R248 VPWR.n35 VPWR.n34 33.1299
R249 VPWR.n29 VPWR.n12 32.9329
R250 VPWR.n28 VPWR.n27 32.6412
R251 VPWR.n23 VPWR.n15 29.3652
R252 VPWR.n14 VPWR.t3 28.1447
R253 VPWR.n22 VPWR.n21 27.8593
R254 VPWR.n17 VPWR.t4 27.6909
R255 VPWR.n7 VPWR.t0 26.3844
R256 VPWR.n7 VPWR.t7 26.3844
R257 VPWR.n21 VPWR.n18 25.977
R258 VPWR.n60 VPWR.n59 24.1661
R259 VPWR.n27 VPWR.n15 24.0946
R260 VPWR.n23 VPWR.n22 22.5887
R261 VPWR.n35 VPWR.n10 20.3299
R262 VPWR.n54 VPWR.n53 11.6711
R263 VPWR.n49 VPWR.n48 10.9181
R264 VPWR.n21 VPWR.n20 9.3005
R265 VPWR.n22 VPWR.n16 9.3005
R266 VPWR.n24 VPWR.n23 9.3005
R267 VPWR.n25 VPWR.n15 9.3005
R268 VPWR.n27 VPWR.n26 9.3005
R269 VPWR.n28 VPWR.n13 9.3005
R270 VPWR.n30 VPWR.n29 9.3005
R271 VPWR.n31 VPWR.n12 9.3005
R272 VPWR.n33 VPWR.n32 9.3005
R273 VPWR.n34 VPWR.n11 9.3005
R274 VPWR.n36 VPWR.n35 9.3005
R275 VPWR.n37 VPWR.n10 9.3005
R276 VPWR.n39 VPWR.n38 9.3005
R277 VPWR.n41 VPWR.n9 9.3005
R278 VPWR.n43 VPWR.n42 9.3005
R279 VPWR.n44 VPWR.n8 9.3005
R280 VPWR.n46 VPWR.n45 9.3005
R281 VPWR.n47 VPWR.n6 9.3005
R282 VPWR.n50 VPWR.n49 9.3005
R283 VPWR.n51 VPWR.n5 9.3005
R284 VPWR.n53 VPWR.n52 9.3005
R285 VPWR.n54 VPWR.n3 9.3005
R286 VPWR.n56 VPWR.n55 9.3005
R287 VPWR.n57 VPWR.n2 9.3005
R288 VPWR.n59 VPWR.n58 9.3005
R289 VPWR.n1 VPWR.n0 9.3005
R290 VPWR.n40 VPWR.n39 9.03579
R291 VPWR.n64 VPWR.n63 8.63089
R292 VPWR.n41 VPWR.n40 8.28285
R293 VPWR.n29 VPWR.n28 8.13825
R294 VPWR.n63 VPWR.n1 7.84868
R295 VPWR.n19 VPWR.n18 6.52251
R296 VPWR.n60 VPWR.n1 0.654515
R297 VPWR.n20 VPWR.n19 0.638643
R298 VPWR.n48 VPWR.n47 0.376971
R299 VPWR VPWR.n64 0.161089
R300 VPWR.n64 VPWR.n0 0.146727
R301 VPWR.n20 VPWR.n16 0.122949
R302 VPWR.n24 VPWR.n16 0.122949
R303 VPWR.n25 VPWR.n24 0.122949
R304 VPWR.n26 VPWR.n25 0.122949
R305 VPWR.n26 VPWR.n13 0.122949
R306 VPWR.n30 VPWR.n13 0.122949
R307 VPWR.n31 VPWR.n30 0.122949
R308 VPWR.n32 VPWR.n31 0.122949
R309 VPWR.n32 VPWR.n11 0.122949
R310 VPWR.n36 VPWR.n11 0.122949
R311 VPWR.n37 VPWR.n36 0.122949
R312 VPWR.n38 VPWR.n37 0.122949
R313 VPWR.n38 VPWR.n9 0.122949
R314 VPWR.n43 VPWR.n9 0.122949
R315 VPWR.n44 VPWR.n43 0.122949
R316 VPWR.n45 VPWR.n44 0.122949
R317 VPWR.n45 VPWR.n6 0.122949
R318 VPWR.n50 VPWR.n6 0.122949
R319 VPWR.n51 VPWR.n50 0.122949
R320 VPWR.n52 VPWR.n51 0.122949
R321 VPWR.n52 VPWR.n3 0.122949
R322 VPWR.n56 VPWR.n3 0.122949
R323 VPWR.n57 VPWR.n56 0.122949
R324 VPWR.n58 VPWR.n57 0.122949
R325 VPWR.n58 VPWR.n0 0.122949
R326 a_388_79.n2 a_388_79.n1 679.736
R327 a_388_79.n1 a_388_79.t3 641.742
R328 a_388_79.n1 a_388_79.n0 355.478
R329 a_388_79.n0 a_388_79.t1 141.429
R330 a_388_79.t0 a_388_79.n2 90.8052
R331 a_388_79.n2 a_388_79.t2 89.2661
R332 a_388_79.n0 a_388_79.t4 42.8576
R333 a_547_79.t0 a_547_79.t1 68.5719
R334 CLK.n0 CLK.t1 265.271
R335 CLK CLK.n0 239.121
R336 CLK.n0 CLK.t0 154.24
R337 a_2006_373.n2 a_2006_373.t0 716.1
R338 a_2006_373.n1 a_2006_373.t2 427.642
R339 a_2006_373.t1 a_2006_373.n2 416.661
R340 a_2006_373.n2 a_2006_373.n1 152
R341 a_2006_373.n1 a_2006_373.n0 129.07
R342 RESET_B.n4 RESET_B.n3 428.981
R343 RESET_B.n1 RESET_B.t1 399.284
R344 RESET_B.n2 RESET_B.t0 392.611
R345 RESET_B.n5 RESET_B.n2 220.061
R346 RESET_B RESET_B.n1 166.97
R347 RESET_B.n5 RESET_B.n4 164.726
R348 RESET_B.n4 RESET_B.t2 157.161
R349 RESET_B.n2 RESET_B.t3 152.367
R350 RESET_B.n1 RESET_B.n0 150.492
R351 RESET_B RESET_B.n5 2.42441
R352 D.n0 D.t1 416.127
R353 D D.n0 163.117
R354 D.n0 D.t0 126.927
R355 a_310_79.t0 a_310_79.t1 68.5719
R356 a_2158_74.t0 a_2158_74.t1 60.0005
R357 a_223_79.t0 a_223_79.n0 565.989
R358 a_223_79.n0 a_223_79.t1 71.4291
R359 a_223_79.n0 a_223_79.t2 40.0005
R360 a_1025_74.t0 a_1025_74.n6 884.437
R361 a_1025_74.n1 a_1025_74.t2 442.808
R362 a_1025_74.n2 a_1025_74.n1 355.101
R363 a_1025_74.n5 a_1025_74.n4 344.12
R364 a_1025_74.n1 a_1025_74.n0 322.827
R365 a_1025_74.n5 a_1025_74.n3 217.436
R366 a_1025_74.n6 a_1025_74.n5 170.812
R367 a_1025_74.n2 a_1025_74.t1 135.637
R368 a_1025_74.n6 a_1025_74.n2 48.1191
R369 SCD.n1 SCD.t1 292.413
R370 SCD.n2 SCD.t0 187.178
R371 SCD.n1 SCD.n0 152
R372 SCD.n3 SCD.n2 152
R373 SCD.n2 SCD.n1 49.6611
R374 SCD.n3 SCD.n0 13.1884
R375 SCD.n0 SCD 0.970197
R376 SCD SCD.n3 0.194439
R377 a_538_464.t0 a_538_464.t1 83.1099
R378 a_2604_392.t0 a_2604_392.n3 257.303
R379 a_2604_392.n0 a_2604_392.t4 240.197
R380 a_2604_392.n2 a_2604_392.t5 240.197
R381 a_2604_392.n0 a_2604_392.t2 182.138
R382 a_2604_392.n1 a_2604_392.t3 179.947
R383 a_2604_392.n3 a_2604_392.t1 156.875
R384 a_2604_392.n3 a_2604_392.n2 120.803
R385 a_2604_392.n1 a_2604_392.n0 60.6157
R386 a_2604_392.n2 a_2604_392.n1 5.11262
R387 Q Q.n0 207.26
R388 Q Q.n1 144.24
R389 Q.n0 Q.t1 26.3844
R390 Q.n0 Q.t0 26.3844
R391 Q.n1 Q.t3 22.7032
R392 Q.n1 Q.t2 22.7032
R393 a_307_464.t0 a_307_464.t1 83.1099
C0 VPWR RESET_B 0.38299f
C1 RESET_B VGND 0.203226f
C2 SCE D 0.140736f
C3 VPWR a_1325_457# 0.001699f
C4 VPWR a_1955_471# 0.001255f
C5 SCD D 0.003937f
C6 VPB D 0.063345f
C7 a_1223_118# VPB 0.077959f
C8 VPWR D 0.011551f
C9 a_1223_118# VPWR 0.190565f
C10 VGND D 0.009388f
C11 a_1223_118# VGND 0.021619f
C12 VPB Q 0.006395f
C13 CLK VPB 0.049068f
C14 VPWR Q 0.223149f
C15 CLK VPWR 0.010941f
C16 Q VGND 0.153647f
C17 CLK VGND 0.025257f
C18 RESET_B a_1325_457# 7.31e-19
C19 SCE SCD 0.081865f
C20 a_1955_471# RESET_B 3.65e-19
C21 VPB SCE 0.206854f
C22 VPB SCD 0.073261f
C23 VPWR SCE 0.038669f
C24 RESET_B D 2.45e-19
C25 a_1223_118# RESET_B 0.227113f
C26 VPB Q_N 0.008338f
C27 VPWR SCD 0.01469f
C28 SCE VGND 0.026396f
C29 VPWR Q_N 0.219861f
C30 SCD VGND 0.005762f
C31 VPB VPWR 0.453879f
C32 a_1223_118# a_1325_457# 0.006525f
C33 Q_N VGND 0.116492f
C34 Q RESET_B 1.4e-19
C35 CLK RESET_B 0.076141f
C36 VPB VGND 0.028736f
C37 VPWR VGND 0.151727f
C38 RESET_B SCE 7.23e-19
C39 RESET_B SCD 0.090598f
C40 RESET_B Q_N 0.001027f
C41 VPB RESET_B 0.35955f
C42 Q VNB 0.030236f
C43 Q_N VNB 0.006081f
C44 VGND VNB 1.75338f
C45 VPWR VNB 1.35264f
C46 CLK VNB 0.166764f
C47 RESET_B VNB 0.422465f
C48 SCD VNB 0.119334f
C49 D VNB 0.141631f
C50 SCE VNB 0.333563f
C51 VPB VNB 3.44888f
C52 a_1223_118# VNB 0.133084f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfxbp_2 VNB VPB VPWR VGND SCE CLK D SCD Q Q_N
X0 a_1243_48.t2 a_1021_97.t4 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.2709 pd=1.485 as=0.18955 ps=1.535 w=0.84 l=0.15
X1 VGND.t4 SCD.t0 a_450_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 a_450_74.t1 SCE.t0 a_301_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.12495 ps=1.015 w=0.42 l=0.15
X3 Q.t1 a_1711_48# VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X4 VGND.t9 a_1711_48# a_2322_368.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.1824 ps=1.85 w=0.64 l=0.15
X5 VGND.t0 a_1243_48.t3 a_1173_97.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14435 pd=1.16 as=0.082125 ps=0.885 w=0.42 l=0.15
X6 a_630_74.t0 CLK.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1212 ps=1.1 w=0.74 l=0.15
X7 a_1711_48# a_1511_74.t1 VGND.t12 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1933 ps=1.47 w=0.74 l=0.15
X8 a_828_74.t0 a_630_74.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_1511_74.t0 a_630_74.t3 a_1243_48.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2709 ps=1.485 w=0.84 l=0.15
X10 a_423_453.t1 a_36_74.t2 a_301_74.t4 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1072 pd=0.975 as=0.1136 ps=0.995 w=0.64 l=0.15
X11 VPWR.t9 a_1711_48# Q.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X12 Q_N.t1 a_2322_368.t2 VGND.t11 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.12945 ps=1.1 w=0.74 l=0.15
X13 Q.t2 a_1711_48# VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X14 a_301_74.t2 D.t0 a_238_453.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1136 pd=0.995 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_1021_97.t0 a_630_74.t4 a_301_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1281 pd=1.03 as=0.1155 ps=1.39 w=0.42 l=0.15
X16 VPWR.t7 a_1711_48# a_2322_368.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2046 pd=1.495 as=0.285 ps=2.57 w=1 l=0.15
X17 VGND.t10 a_1711_48# a_1663_74# VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1933 pd=1.47 as=0.0504 ps=0.66 w=0.42 l=0.15
X18 VPWR.t3 SCD.t1 a_423_453.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.259825 pd=1.74 as=0.1072 ps=0.975 w=0.64 l=0.15
X19 a_630_74.t1 CLK.t1 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.5656 pd=3.25 as=0.259825 ps=1.74 w=1.12 l=0.15
X20 a_301_74.t3 D.t1 a_223_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.12495 pd=1.015 as=0.0504 ps=0.66 w=0.42 l=0.15
X21 VGND.t5 SCE.t1 a_36_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X22 VPWR.t6 a_1243_48.t4 a_1217_499.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.18955 pd=1.535 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_1243_48.t1 a_1021_97.t5 VGND.t13 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.14435 ps=1.16 w=0.55 l=0.15
X24 a_1217_499.t1 a_630_74.t5 a_1021_97.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08085 ps=0.805 w=0.42 l=0.15
X25 VPWR a_1711_48# a_1691_508# VPB sky130_fd_pr__pfet_01v8 ad=0.20075 pd=1.59 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND.t7 a_1711_48# Q.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 a_238_453.t0 SCE.t2 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.096 ps=0.94 w=0.64 l=0.15
X28 VPWR.t0 SCE.t3 a_36_74.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.2432 ps=2.04 w=0.64 l=0.15
X29 a_1021_97.t2 a_828_74.t2 a_301_74.t5 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.08085 pd=0.805 as=0.1239 ps=1.43 w=0.42 l=0.15
X30 a_1173_97.t1 a_828_74.t3 a_1021_97.t3 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.082125 pd=0.885 as=0.1281 ps=1.03 w=0.42 l=0.15
X31 a_828_74.t1 a_630_74.t6 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X32 VPWR.t1 a_2322_368.t3 Q_N.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X33 VGND.t3 a_2322_368.t4 Q_N.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1962 pd=2.05 as=0.10915 ps=1.035 w=0.74 l=0.15
X34 a_223_74.t1 a_36_74.t3 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X35 Q_N.t2 a_2322_368.t5 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2046 ps=1.495 w=1.12 l=0.15
R0 a_1021_97.n2 a_1021_97.n0 648.144
R1 a_1021_97.n1 a_1021_97.t5 331.091
R2 a_1021_97.n3 a_1021_97.n2 251.841
R3 a_1021_97.n2 a_1021_97.n1 243.543
R4 a_1021_97.n1 a_1021_97.t4 205.236
R5 a_1021_97.t0 a_1021_97.n3 134.286
R6 a_1021_97.n0 a_1021_97.t1 110.227
R7 a_1021_97.n0 a_1021_97.t2 70.3576
R8 a_1021_97.n3 a_1021_97.t3 40.0005
R9 VPWR.n5 VPWR.t10 875.822
R10 VPWR.n34 VPWR.n33 662.674
R11 VPWR.n47 VPWR.n4 598.867
R12 VPWR.n16 VPWR.t1 349.514
R13 VPWR.n54 VPWR.n1 317.964
R14 VPWR.n21 VPWR.t8 259.171
R15 VPWR.n19 VPWR.t9 250.279
R16 VPWR.n15 VPWR.n14 232.787
R17 VPWR.n33 VPWR.t6 131.333
R18 VPWR.n4 VPWR.t3 86.188
R19 VPWR.n4 VPWR.t5 57.9816
R20 VPWR.n1 VPWR.t4 46.1724
R21 VPWR.n1 VPWR.t0 46.1724
R22 VPWR.n33 VPWR.t11 45.4118
R23 VPWR.n14 VPWR.t7 44.3255
R24 VPWR.n48 VPWR.n2 36.1417
R25 VPWR.n52 VPWR.n2 36.1417
R26 VPWR.n53 VPWR.n52 36.1417
R27 VPWR.n46 VPWR.n45 36.1417
R28 VPWR.n35 VPWR.n7 36.1417
R29 VPWR.n39 VPWR.n7 36.1417
R30 VPWR.n40 VPWR.n39 36.1417
R31 VPWR.n41 VPWR.n40 36.1417
R32 VPWR.n27 VPWR.n9 36.1417
R33 VPWR.n31 VPWR.n9 36.1417
R34 VPWR.n32 VPWR.n31 36.1417
R35 VPWR.n45 VPWR.n5 35.7652
R36 VPWR.n27 VPWR.n26 34.9704
R37 VPWR.n25 VPWR.n11 32.0423
R38 VPWR.n21 VPWR.n20 30.8711
R39 VPWR.n19 VPWR.n18 29.3652
R40 VPWR.n14 VPWR.t2 27.098
R41 VPWR.n18 VPWR.n15 25.977
R42 VPWR.n21 VPWR.n11 22.5887
R43 VPWR.n20 VPWR.n19 18.0711
R44 VPWR.n35 VPWR.n34 11.7447
R45 VPWR.n41 VPWR.n5 11.6711
R46 VPWR.n54 VPWR.n53 10.9181
R47 VPWR.n18 VPWR.n17 9.3005
R48 VPWR.n19 VPWR.n13 9.3005
R49 VPWR.n20 VPWR.n12 9.3005
R50 VPWR.n22 VPWR.n21 9.3005
R51 VPWR.n23 VPWR.n11 9.3005
R52 VPWR.n25 VPWR.n24 9.3005
R53 VPWR.n26 VPWR.n10 9.3005
R54 VPWR.n28 VPWR.n27 9.3005
R55 VPWR.n29 VPWR.n9 9.3005
R56 VPWR.n31 VPWR.n30 9.3005
R57 VPWR.n32 VPWR.n8 9.3005
R58 VPWR.n36 VPWR.n35 9.3005
R59 VPWR.n37 VPWR.n7 9.3005
R60 VPWR.n39 VPWR.n38 9.3005
R61 VPWR.n40 VPWR.n6 9.3005
R62 VPWR.n42 VPWR.n41 9.3005
R63 VPWR.n43 VPWR.n5 9.3005
R64 VPWR.n45 VPWR.n44 9.3005
R65 VPWR.n46 VPWR.n3 9.3005
R66 VPWR.n49 VPWR.n48 9.3005
R67 VPWR.n50 VPWR.n2 9.3005
R68 VPWR.n52 VPWR.n51 9.3005
R69 VPWR.n53 VPWR.n0 9.3005
R70 VPWR.n34 VPWR.n32 8.73298
R71 VPWR.n55 VPWR.n54 8.08026
R72 VPWR.n26 VPWR.n25 8.03187
R73 VPWR.n16 VPWR.n15 6.85135
R74 VPWR.n48 VPWR.n47 2.25932
R75 VPWR.n47 VPWR.n46 2.25932
R76 VPWR.n17 VPWR.n16 0.609796
R77 VPWR VPWR.n55 0.163644
R78 VPWR.n55 VPWR.n0 0.144205
R79 VPWR.n17 VPWR.n13 0.122949
R80 VPWR.n13 VPWR.n12 0.122949
R81 VPWR.n22 VPWR.n12 0.122949
R82 VPWR.n23 VPWR.n22 0.122949
R83 VPWR.n24 VPWR.n23 0.122949
R84 VPWR.n24 VPWR.n10 0.122949
R85 VPWR.n28 VPWR.n10 0.122949
R86 VPWR.n29 VPWR.n28 0.122949
R87 VPWR.n30 VPWR.n29 0.122949
R88 VPWR.n30 VPWR.n8 0.122949
R89 VPWR.n36 VPWR.n8 0.122949
R90 VPWR.n37 VPWR.n36 0.122949
R91 VPWR.n38 VPWR.n37 0.122949
R92 VPWR.n38 VPWR.n6 0.122949
R93 VPWR.n42 VPWR.n6 0.122949
R94 VPWR.n43 VPWR.n42 0.122949
R95 VPWR.n44 VPWR.n43 0.122949
R96 VPWR.n44 VPWR.n3 0.122949
R97 VPWR.n49 VPWR.n3 0.122949
R98 VPWR.n50 VPWR.n49 0.122949
R99 VPWR.n51 VPWR.n50 0.122949
R100 VPWR.n51 VPWR.n0 0.122949
R101 a_1243_48.n2 a_1243_48.n1 645.87
R102 a_1243_48.n0 a_1243_48.t4 385.163
R103 a_1243_48.n1 a_1243_48.t1 241.523
R104 a_1243_48.n1 a_1243_48.n0 188.881
R105 a_1243_48.n0 a_1243_48.t3 180.85
R106 a_1243_48.t0 a_1243_48.n2 112.572
R107 a_1243_48.n2 a_1243_48.t2 38.6969
R108 VPB.t1 VPB.t12 1371.37
R109 VPB.t9 VPB.t15 628.226
R110 VPB.t15 VPB.t14 515.861
R111 VPB.t13 VPB.t11 505.646
R112 VPB.t16 VPB.t1 406.048
R113 VPB.t7 VPB.t9 362.635
R114 VPB VPB.t3 339.651
R115 VPB.t0 VPB.t16 316.668
R116 VPB.t14 VPB.t2 273.253
R117 VPB.t11 VPB.t5 268.146
R118 VPB.t6 VPB.t10 257.93
R119 VPB.t10 VPB.t7 247.715
R120 VPB.t5 VPB.t4 229.839
R121 VPB.t12 VPB.t13 229.839
R122 VPB.t3 VPB.t8 229.839
R123 VPB.t2 VPB.t0 214.517
R124 VPB.t8 VPB.t6 214.517
R125 SCD.n0 SCD.t0 408.094
R126 SCD.n0 SCD.t1 173.788
R127 SCD SCD.n0 152.512
R128 a_450_74.t0 a_450_74.t1 68.5719
R129 VGND.n3 VGND.t2 269.132
R130 VGND.n15 VGND.t3 238.782
R131 VGND.n52 VGND.n49 208.041
R132 VGND.n61 VGND.n60 205.946
R133 VGND.n37 VGND.n36 204.976
R134 VGND.n29 VGND.n28 185
R135 VGND.n27 VGND.n26 185
R136 VGND.n52 VGND.n51 185
R137 VGND.n18 VGND.t7 171.77
R138 VGND.n20 VGND.t8 154.727
R139 VGND.n28 VGND.n27 128.571
R140 VGND.n36 VGND.t13 122.174
R141 VGND.n14 VGND.n13 117.183
R142 VGND.n50 VGND.t4 61.4291
R143 VGND.n60 VGND.t5 60.0005
R144 VGND.t1 VGND.n49 52.5005
R145 VGND.n28 VGND.t10 40.0005
R146 VGND.n36 VGND.t0 40.0005
R147 VGND.n51 VGND.t1 40.0005
R148 VGND.n60 VGND.t6 40.0005
R149 VGND.n13 VGND.t9 38.4442
R150 VGND.n31 VGND.n30 36.1417
R151 VGND.n31 VGND.n7 36.1417
R152 VGND.n35 VGND.n7 36.1417
R153 VGND.n38 VGND.n5 36.1417
R154 VGND.n42 VGND.n5 36.1417
R155 VGND.n43 VGND.n42 36.1417
R156 VGND.n44 VGND.n43 36.1417
R157 VGND.n48 VGND.n47 36.1417
R158 VGND.n54 VGND.n1 36.1417
R159 VGND.n58 VGND.n1 36.1417
R160 VGND.n59 VGND.n58 36.1417
R161 VGND.n25 VGND.n10 34.3629
R162 VGND.n18 VGND.n12 28.6123
R163 VGND.n14 VGND.n12 27.1064
R164 VGND.n53 VGND.n52 26.3685
R165 VGND.n20 VGND.n19 26.3534
R166 VGND.n38 VGND.n37 25.6005
R167 VGND.n19 VGND.n18 24.8476
R168 VGND.n27 VGND.t12 24.5565
R169 VGND.n13 VGND.t11 23.7368
R170 VGND.n30 VGND.n29 23.7229
R171 VGND.n37 VGND.n35 21.8358
R172 VGND.n20 VGND.n10 21.0829
R173 VGND.n61 VGND.n59 15.8123
R174 VGND.n53 VGND.n48 13.177
R175 VGND.n59 VGND.n0 9.3005
R176 VGND.n58 VGND.n57 9.3005
R177 VGND.n56 VGND.n1 9.3005
R178 VGND.n55 VGND.n54 9.3005
R179 VGND.n16 VGND.n12 9.3005
R180 VGND.n18 VGND.n17 9.3005
R181 VGND.n19 VGND.n11 9.3005
R182 VGND.n21 VGND.n20 9.3005
R183 VGND.n22 VGND.n10 9.3005
R184 VGND.n25 VGND.n24 9.3005
R185 VGND.n23 VGND.n9 9.3005
R186 VGND.n30 VGND.n8 9.3005
R187 VGND.n32 VGND.n31 9.3005
R188 VGND.n33 VGND.n7 9.3005
R189 VGND.n35 VGND.n34 9.3005
R190 VGND.n37 VGND.n6 9.3005
R191 VGND.n39 VGND.n38 9.3005
R192 VGND.n40 VGND.n5 9.3005
R193 VGND.n42 VGND.n41 9.3005
R194 VGND.n43 VGND.n4 9.3005
R195 VGND.n45 VGND.n44 9.3005
R196 VGND.n47 VGND.n46 9.3005
R197 VGND.n48 VGND.n2 9.3005
R198 VGND.n62 VGND.n61 7.56047
R199 VGND.n26 VGND.n9 6.6405
R200 VGND.n47 VGND.n3 6.4005
R201 VGND.n15 VGND.n14 6.36273
R202 VGND.n44 VGND.n3 4.89462
R203 VGND.n54 VGND.n53 4.14168
R204 VGND.n50 VGND.n49 1.8755
R205 VGND.n51 VGND.n50 1.42907
R206 VGND.n26 VGND.n25 1.0405
R207 VGND.n16 VGND.n15 0.715227
R208 VGND.n29 VGND.n9 0.5605
R209 VGND VGND.n62 0.161757
R210 VGND.n62 VGND.n0 0.146068
R211 VGND.n17 VGND.n16 0.122949
R212 VGND.n17 VGND.n11 0.122949
R213 VGND.n21 VGND.n11 0.122949
R214 VGND.n22 VGND.n21 0.122949
R215 VGND.n24 VGND.n22 0.122949
R216 VGND.n24 VGND.n23 0.122949
R217 VGND.n23 VGND.n8 0.122949
R218 VGND.n32 VGND.n8 0.122949
R219 VGND.n33 VGND.n32 0.122949
R220 VGND.n34 VGND.n33 0.122949
R221 VGND.n34 VGND.n6 0.122949
R222 VGND.n39 VGND.n6 0.122949
R223 VGND.n40 VGND.n39 0.122949
R224 VGND.n41 VGND.n40 0.122949
R225 VGND.n41 VGND.n4 0.122949
R226 VGND.n45 VGND.n4 0.122949
R227 VGND.n46 VGND.n45 0.122949
R228 VGND.n46 VGND.n2 0.122949
R229 VGND.n55 VGND.n2 0.122949
R230 VGND.n56 VGND.n55 0.122949
R231 VGND.n57 VGND.n56 0.122949
R232 VGND.n57 VGND.n0 0.122949
R233 VNB.t17 VNB.t11 3649.34
R234 VNB.t16 VNB.t13 2448.29
R235 VNB.t10 VNB.t12 2286.61
R236 VNB.t1 VNB.t2 2286.61
R237 VNB.t2 VNB.t3 2228.87
R238 VNB.t11 VNB.t16 2032.55
R239 VNB.t0 VNB.t17 1755.38
R240 VNB.t3 VNB.t15 1755.38
R241 VNB.t6 VNB.t7 1720.73
R242 VNB VNB.t8 1247.24
R243 VNB.t12 VNB.t14 1177.95
R244 VNB.t5 VNB.t1 1177.95
R245 VNB.t15 VNB.t0 1154.86
R246 VNB.t8 VNB.t9 1154.86
R247 VNB.t14 VNB.t4 1027.82
R248 VNB.t13 VNB.t10 993.177
R249 VNB.t7 VNB.t5 900.788
R250 VNB.t9 VNB.t6 900.788
R251 SCE.n1 SCE.n0 401.409
R252 SCE SCE.t0 303.134
R253 SCE.n0 SCE.t2 271.527
R254 SCE SCE.n1 190.732
R255 SCE.n0 SCE.t3 126.927
R256 SCE.n1 SCE.t1 117.028
R257 a_301_74.n1 a_301_74.t5 710.076
R258 a_301_74.n2 a_301_74.n0 380.796
R259 a_301_74.n3 a_301_74.n2 373.426
R260 a_301_74.n1 a_301_74.t1 343.017
R261 a_301_74.n2 a_301_74.n1 100.894
R262 a_301_74.n0 a_301_74.t0 85.7148
R263 a_301_74.n0 a_301_74.t3 84.2862
R264 a_301_74.t2 a_301_74.n3 63.1021
R265 a_301_74.n3 a_301_74.t4 46.1724
R266 Q.n1 Q.n0 270.079
R267 Q.n2 Q.n1 185
R268 Q.n3 Q.n2 185
R269 Q.n0 Q.t3 26.3844
R270 Q.n0 Q.t2 26.3844
R271 Q.n2 Q.t0 22.7032
R272 Q.n2 Q.t1 22.7032
R273 Q.n3 Q 12.6066
R274 Q.n1 Q 4.84898
R275 Q Q.n3 1.74595
R276 a_2322_368.t1 a_2322_368.n3 250.899
R277 a_2322_368.n1 a_2322_368.t5 235.571
R278 a_2322_368.n0 a_2322_368.t3 234.841
R279 a_2322_368.n0 a_2322_368.t4 179.947
R280 a_2322_368.n1 a_2322_368.t2 179.947
R281 a_2322_368.n3 a_2322_368.n2 176.436
R282 a_2322_368.n3 a_2322_368.t0 148.341
R283 a_2322_368.n2 a_2322_368.n0 54.7732
R284 a_2322_368.n2 a_2322_368.n1 10.2247
R285 a_1173_97.n0 a_1173_97.t1 75.059
R286 a_1173_97.n1 a_1173_97.n0 28.8005
R287 a_1173_97.n0 a_1173_97.t0 23.6618
R288 CLK.n0 CLK.t1 244.482
R289 CLK.n0 CLK.t0 228.498
R290 CLK CLK.n0 154.53
R291 a_630_74.t1 a_630_74.n6 745.49
R292 a_630_74.n2 a_630_74.n1 510.902
R293 a_630_74.n1 a_630_74.n0 389.291
R294 a_630_74.n3 a_630_74.n2 304.39
R295 a_630_74.n3 a_630_74.t4 295.627
R296 a_630_74.n5 a_630_74.t2 220.113
R297 a_630_74.n1 a_630_74.t3 211.35
R298 a_630_74.n6 a_630_74.t0 207.262
R299 a_630_74.n4 a_630_74.t6 204.048
R300 a_630_74.n4 a_630_74.n3 181.554
R301 a_630_74.n2 a_630_74.t5 162.542
R302 a_630_74.n6 a_630_74.n5 152
R303 a_630_74.n5 a_630_74.n4 129.994
R304 a_1511_74.t0 a_1511_74.n1 645.755
R305 a_1511_74.n1 a_1511_74.n0 297.195
R306 a_1511_74.n1 a_1511_74.t1 176.964
R307 a_828_74.t1 a_828_74.n5 866.846
R308 a_828_74.n2 a_828_74.n0 583.995
R309 a_828_74.n5 a_828_74.t2 327.192
R310 a_828_74.n3 a_828_74.t3 302.873
R311 a_828_74.n2 a_828_74.n1 296.921
R312 a_828_74.n4 a_828_74.t0 210.457
R313 a_828_74.n3 a_828_74.n2 200.876
R314 a_828_74.n5 a_828_74.n4 118.966
R315 a_828_74.n4 a_828_74.n3 89.224
R316 a_36_74.n0 a_36_74.t3 480.344
R317 a_36_74.n0 a_36_74.t2 438.099
R318 a_36_74.t1 a_36_74.n1 390.195
R319 a_36_74.n1 a_36_74.t0 291.579
R320 a_36_74.n1 a_36_74.n0 8.92171
R321 a_423_453.t0 a_423_453.t1 103.118
R322 Q_N Q_N.n0 217.762
R323 Q_N Q_N.n1 212.52
R324 Q_N.n0 Q_N.t3 26.3844
R325 Q_N.n0 Q_N.t2 26.3844
R326 Q_N.n1 Q_N.t0 24.3248
R327 Q_N.n1 Q_N.t1 23.514
R328 D.n0 D.t1 310.087
R329 D.n0 D.t0 255.46
R330 D D.n0 166.546
R331 a_238_453.t0 a_238_453.t1 83.1099
R332 a_223_74.t0 a_223_74.t1 68.5719
R333 a_1217_499.t0 a_1217_499.t1 126.644
C0 VPB VGND 0.032084f
C1 a_1711_48# a_1663_74# 2.21e-19
C2 SCD VPWR 0.013796f
C3 a_1663_74# VPWR 4.86e-19
C4 VPB Q_N 0.010955f
C5 VPB Q 0.006793f
C6 Q_N VGND 0.083046f
C7 D SCE 0.111272f
C8 VPB SCE 0.140262f
C9 Q VGND 0.165454f
C10 VGND SCE 0.081344f
C11 CLK VPB 0.052227f
C12 VGND a_1691_508# 5.47e-19
C13 VPB a_1711_48# 0.283707f
C14 D VPWR 0.013977f
C15 VPB VPWR 0.416989f
C16 SCD D 0.009302f
C17 CLK VGND 0.015377f
C18 SCD VPB 0.081405f
C19 a_1711_48# VGND 0.262491f
C20 VGND VPWR 0.225355f
C21 SCD VGND 0.019752f
C22 VGND a_1663_74# 0.004859f
C23 a_1711_48# Q_N 0.001237f
C24 Q_N VPWR 0.216676f
C25 a_1711_48# Q 0.10904f
C26 Q VPWR 0.20907f
C27 SCD Q 1.32e-23
C28 VPWR SCE 0.038075f
C29 a_1711_48# a_1691_508# 5.81e-19
C30 SCD SCE 0.038047f
C31 a_1691_508# VPWR 0.006778f
C32 D VPB 0.06524f
C33 CLK VPWR 0.015868f
C34 SCD CLK 0.036429f
C35 a_1711_48# VPWR 0.33396f
C36 SCD a_1711_48# 5.75e-22
C37 D VGND 0.01241f
C38 Q_N VNB 0.065926f
C39 Q VNB 0.013643f
C40 VGND VNB 1.58222f
C41 CLK VNB 0.137511f
C42 SCD VNB 0.130752f
C43 D VNB 0.128908f
C44 SCE VNB 0.365063f
C45 VPWR VNB 1.23084f
C46 VPB VNB 3.08462f
C47 a_1711_48# VNB 0.613926f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfxbp_1 VNB VPB VPWR VGND Q_N Q CLK D SCE SCD
X0 a_1157_100.t0 a_828_74.t2 a_1021_100.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0966 pd=0.88 as=0.1113 ps=0.95 w=0.42 l=0.15
X1 a_296_74.t3 D.t0 a_218_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1134 pd=0.96 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 VGND.t5 SCD.t0 a_434_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1135 pd=1.09 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 VGND.t7 SCE.t0 a_31_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4 a_1243_398.t3 a_1021_100.t4 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.078375 pd=0.835 as=0.1996 ps=1.375 w=0.55 l=0.15
X5 VPWR.t8 SCE.t1 a_31_74.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.1888 ps=1.87 w=0.64 l=0.15
X6 a_1180_496.t0 a_612_74.t2 a_1021_100.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.063 ps=0.72 w=0.42 l=0.15
X7 a_1529_74.t0 a_612_74.t3 a_1243_398.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.3234 ps=1.61 w=0.84 l=0.15
X8 a_828_74.t1 a_612_74.t4 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.2805 ps=2.25 w=0.74 l=0.15
X9 a_1021_100.t2 a_828_74.t3 a_296_74.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X10 VPWR.t6 a_1243_398.t4 a_1180_496.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.18825 pd=1.52 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_1529_74.t1 a_828_74.t4 a_1243_398.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.14435 pd=1.16 as=0.078375 ps=0.835 w=0.55 l=0.15
X12 Q_N.t0 a_2216_94.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1424 ps=1.135 w=0.74 l=0.15
X13 a_1681_74.t1 a_612_74.t5 a_1529_74.t2 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.14435 ps=1.16 w=0.42 l=0.15
X14 a_828_74.t0 a_612_74.t6 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.5264 ps=3.18 w=1.12 l=0.15
X15 a_407_464.t0 a_31_74.t2 a_296_74.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1248 pd=1.03 as=0.096 ps=0.94 w=0.64 l=0.15
X16 VGND.t1 a_1723_48# a_1681_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.148725 pd=1.17 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_434_74.t0 SCE.t2 a_296_74.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1134 ps=0.96 w=0.42 l=0.15
X18 a_296_74.t4 D.t1 a_233_464.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 a_612_74.t1 CLK.t0 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2428 ps=1.68 w=1.12 l=0.15
X20 VPWR.t9 SCD.t1 a_407_464.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2428 pd=1.68 as=0.1248 ps=1.03 w=0.64 l=0.15
X21 a_1243_398.t2 a_1021_100.t5 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3234 pd=1.61 as=0.18825 ps=1.52 w=0.84 l=0.15
X22 a_218_74.t1 a_31_74.t3 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X23 Q.t1 a_1723_48# VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X24 a_1021_100.t0 a_612_74.t7 a_296_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1155 ps=1.39 w=0.42 l=0.15
X25 VPWR a_1723_48# a_1691_508# VPB sky130_fd_pr__pfet_01v8 ad=0.20075 pd=1.59 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND.t0 a_1723_48# a_2216_94.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1424 pd=1.135 as=0.1824 ps=1.85 w=0.64 l=0.15
X27 a_612_74.t0 CLK.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1135 ps=1.09 w=0.74 l=0.15
X28 Q.t0 a_1723_48# VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X29 VPWR.t0 a_1723_48# a_2216_94.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.231 ps=2.23 w=0.84 l=0.15
X30 a_233_464.t0 SCE.t3 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X31 Q_N.t1 a_2216_94.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1862 ps=1.475 w=1.12 l=0.15
R0 a_828_74.t0 a_828_74.n4 866.918
R1 a_828_74.n1 a_828_74.n0 527.206
R2 a_828_74.n1 a_828_74.t4 325.3
R3 a_828_74.n4 a_828_74.t3 324.985
R4 a_828_74.n2 a_828_74.t2 293.572
R5 a_828_74.n3 a_828_74.t1 210.457
R6 a_828_74.n2 a_828_74.n1 201.036
R7 a_828_74.n4 a_828_74.n3 107.596
R8 a_828_74.n3 a_828_74.n2 64.3373
R9 a_1021_100.n2 a_1021_100.n0 650.516
R10 a_1021_100.n1 a_1021_100.t4 322.168
R11 a_1021_100.n2 a_1021_100.n1 247.256
R12 a_1021_100.n3 a_1021_100.n2 242.601
R13 a_1021_100.n1 a_1021_100.t5 205.149
R14 a_1021_100.t0 a_1021_100.n3 111.43
R15 a_1021_100.n0 a_1021_100.t1 70.3576
R16 a_1021_100.n0 a_1021_100.t2 70.3576
R17 a_1021_100.n3 a_1021_100.t3 40.0005
R18 VNB.t2 VNB.t0 4065.09
R19 VNB.t9 VNB.t10 3291.34
R20 VNB.t4 VNB.t13 2494.49
R21 VNB.t0 VNB.t1 2286.61
R22 VNB.t13 VNB.t5 2228.87
R23 VNB.t8 VNB.t14 1755.38
R24 VNB.t6 VNB.t12 1593.7
R25 VNB.t5 VNB.t9 1570.6
R26 VNB.t1 VNB.t3 1258.79
R27 VNB VNB.t11 1189.5
R28 VNB.t7 VNB.t4 1154.86
R29 VNB.t11 VNB.t15 1154.86
R30 VNB.t10 VNB.t8 1004.72
R31 VNB.t12 VNB.t7 900.788
R32 VNB.t15 VNB.t6 900.788
R33 VNB.t14 VNB.t2 831.496
R34 a_1529_74.t0 a_1529_74.n4 459.221
R35 a_1529_74.n2 a_1529_74.n1 259.534
R36 a_1529_74.n4 a_1529_74.n3 245.089
R37 a_1529_74.n2 a_1529_74.n0 188.482
R38 a_1529_74.n3 a_1529_74.t1 122.174
R39 a_1529_74.n4 a_1529_74.n2 91.658
R40 a_1529_74.n3 a_1529_74.t2 40.0005
R41 VGND.n24 VGND.t6 309.115
R42 VGND.n34 VGND.t8 279.212
R43 VGND.n37 VGND.n36 214.696
R44 VGND.n44 VGND.n43 207.498
R45 VGND.n10 VGND.t2 180.233
R46 VGND.n16 VGND.t1 150.585
R47 VGND.n12 VGND.n11 115.859
R48 VGND.n43 VGND.t7 60.0005
R49 VGND.n36 VGND.t5 51.4291
R50 VGND.n43 VGND.t9 40.0005
R51 VGND.n11 VGND.t0 37.025
R52 VGND.n18 VGND.n7 36.1417
R53 VGND.n22 VGND.n7 36.1417
R54 VGND.n23 VGND.n22 36.1417
R55 VGND.n28 VGND.n5 36.1417
R56 VGND.n29 VGND.n28 36.1417
R57 VGND.n30 VGND.n29 36.1417
R58 VGND.n30 VGND.n3 36.1417
R59 VGND.n41 VGND.n1 36.1417
R60 VGND.n42 VGND.n41 36.1417
R61 VGND.n35 VGND.n34 35.7652
R62 VGND.n37 VGND.n1 34.2593
R63 VGND.n36 VGND.t4 33.1279
R64 VGND.n15 VGND.n9 33.0921
R65 VGND.n24 VGND.n5 32.377
R66 VGND.n10 VGND.n9 29.7417
R67 VGND.n11 VGND.t3 29.6851
R68 VGND.n18 VGND.n17 27.6027
R69 VGND.n24 VGND.n23 21.0829
R70 VGND.n37 VGND.n35 19.2005
R71 VGND.n44 VGND.n42 17.6946
R72 VGND.n12 VGND.n10 13.9831
R73 VGND.n34 VGND.n3 10.9181
R74 VGND.n42 VGND.n0 9.3005
R75 VGND.n41 VGND.n40 9.3005
R76 VGND.n39 VGND.n1 9.3005
R77 VGND.n38 VGND.n37 9.3005
R78 VGND.n35 VGND.n2 9.3005
R79 VGND.n34 VGND.n33 9.3005
R80 VGND.n32 VGND.n3 9.3005
R81 VGND.n31 VGND.n30 9.3005
R82 VGND.n29 VGND.n4 9.3005
R83 VGND.n28 VGND.n27 9.3005
R84 VGND.n26 VGND.n5 9.3005
R85 VGND.n25 VGND.n24 9.3005
R86 VGND.n23 VGND.n6 9.3005
R87 VGND.n22 VGND.n21 9.3005
R88 VGND.n20 VGND.n7 9.3005
R89 VGND.n19 VGND.n18 9.3005
R90 VGND.n17 VGND.n8 9.3005
R91 VGND.n15 VGND.n14 9.3005
R92 VGND.n13 VGND.n9 9.3005
R93 VGND.n45 VGND.n44 7.49287
R94 VGND.n16 VGND.n15 4.55231
R95 VGND.n17 VGND.n16 2.2644
R96 VGND.n13 VGND.n12 0.215899
R97 VGND VGND.n45 0.160867
R98 VGND.n45 VGND.n0 0.146947
R99 VGND.n14 VGND.n13 0.122949
R100 VGND.n14 VGND.n8 0.122949
R101 VGND.n19 VGND.n8 0.122949
R102 VGND.n20 VGND.n19 0.122949
R103 VGND.n21 VGND.n20 0.122949
R104 VGND.n21 VGND.n6 0.122949
R105 VGND.n25 VGND.n6 0.122949
R106 VGND.n26 VGND.n25 0.122949
R107 VGND.n27 VGND.n26 0.122949
R108 VGND.n27 VGND.n4 0.122949
R109 VGND.n31 VGND.n4 0.122949
R110 VGND.n32 VGND.n31 0.122949
R111 VGND.n33 VGND.n32 0.122949
R112 VGND.n33 VGND.n2 0.122949
R113 VGND.n38 VGND.n2 0.122949
R114 VGND.n39 VGND.n38 0.122949
R115 VGND.n40 VGND.n39 0.122949
R116 VGND.n40 VGND.n0 0.122949
R117 D.n0 D.t0 305.267
R118 D.n0 D.t1 274.204
R119 D D.n0 165.577
R120 a_218_74.t0 a_218_74.t1 68.5719
R121 a_296_74.n1 a_296_74.t1 709.298
R122 a_296_74.n2 a_296_74.n0 383.204
R123 a_296_74.n3 a_296_74.n2 377.178
R124 a_296_74.n1 a_296_74.t0 349.536
R125 a_296_74.n2 a_296_74.n1 97.8829
R126 a_296_74.n0 a_296_74.t2 77.1434
R127 a_296_74.n0 a_296_74.t3 77.1434
R128 a_296_74.n3 a_296_74.t5 46.1724
R129 a_296_74.t4 a_296_74.n3 46.1724
R130 SCD.n0 SCD.t0 355.074
R131 SCD.n0 SCD.t1 232.7
R132 SCD.n1 SCD.n0 152
R133 SCD.n1 SCD 7.23528
R134 SCD SCD.n1 6.49325
R135 a_434_74.t0 a_434_74.t1 68.5719
R136 SCE.n1 SCE.n0 418.026
R137 SCE SCE.t2 293.315
R138 SCE.n0 SCE.t3 287.594
R139 SCE SCE.n1 191.596
R140 SCE.n1 SCE.t0 144.601
R141 SCE.n0 SCE.t1 126.927
R142 a_31_74.n0 a_31_74.t3 494.366
R143 a_31_74.n0 a_31_74.t2 428.24
R144 a_31_74.t1 a_31_74.n1 375.724
R145 a_31_74.n1 a_31_74.t0 292.875
R146 a_31_74.n1 a_31_74.n0 8.53383
R147 a_1243_398.n4 a_1243_398.n3 645.87
R148 a_1243_398.n2 a_1243_398.t4 429.248
R149 a_1243_398.n3 a_1243_398.n0 201.234
R150 a_1243_398.n3 a_1243_398.n2 185.553
R151 a_1243_398.t0 a_1243_398.n4 136.024
R152 a_1243_398.n2 a_1243_398.n1 126.927
R153 a_1243_398.n4 a_1243_398.t2 44.56
R154 a_1243_398.n0 a_1243_398.t3 31.6369
R155 a_1243_398.n0 a_1243_398.t1 30.546
R156 VPWR.n4 VPWR.t3 772
R157 VPWR.n25 VPWR.n24 660.26
R158 VPWR.n39 VPWR.n38 585
R159 VPWR.n13 VPWR.n11 327.841
R160 VPWR.n46 VPWR.n1 315.832
R161 VPWR.n12 VPWR.t1 250.081
R162 VPWR.n24 VPWR.t6 131.333
R163 VPWR.n38 VPWR.t9 86.188
R164 VPWR.n38 VPWR.t5 68.3788
R165 VPWR.n1 VPWR.t8 61.563
R166 VPWR.n1 VPWR.t7 46.1724
R167 VPWR.n24 VPWR.t4 45.3438
R168 VPWR.n11 VPWR.t2 42.7085
R169 VPWR.n44 VPWR.n2 36.1417
R170 VPWR.n45 VPWR.n44 36.1417
R171 VPWR.n30 VPWR.n6 36.1417
R172 VPWR.n31 VPWR.n30 36.1417
R173 VPWR.n32 VPWR.n31 36.1417
R174 VPWR.n18 VPWR.n8 36.1417
R175 VPWR.n22 VPWR.n8 36.1417
R176 VPWR.n23 VPWR.n22 36.1417
R177 VPWR.n11 VPWR.t0 35.1791
R178 VPWR.n18 VPWR.n17 34.9704
R179 VPWR.n26 VPWR.n6 34.5747
R180 VPWR.n37 VPWR.n36 34.4434
R181 VPWR.n16 VPWR.n10 32.0423
R182 VPWR.n40 VPWR.n2 31.613
R183 VPWR.n12 VPWR.n10 21.0829
R184 VPWR.n25 VPWR.n23 17.3588
R185 VPWR.n36 VPWR.n4 17.3181
R186 VPWR.n32 VPWR.n4 16.9417
R187 VPWR.n46 VPWR.n45 12.8005
R188 VPWR.n14 VPWR.n10 9.3005
R189 VPWR.n16 VPWR.n15 9.3005
R190 VPWR.n17 VPWR.n9 9.3005
R191 VPWR.n19 VPWR.n18 9.3005
R192 VPWR.n20 VPWR.n8 9.3005
R193 VPWR.n22 VPWR.n21 9.3005
R194 VPWR.n23 VPWR.n7 9.3005
R195 VPWR.n27 VPWR.n26 9.3005
R196 VPWR.n28 VPWR.n6 9.3005
R197 VPWR.n30 VPWR.n29 9.3005
R198 VPWR.n31 VPWR.n5 9.3005
R199 VPWR.n33 VPWR.n32 9.3005
R200 VPWR.n34 VPWR.n4 9.3005
R201 VPWR.n36 VPWR.n35 9.3005
R202 VPWR.n37 VPWR.n3 9.3005
R203 VPWR.n41 VPWR.n40 9.3005
R204 VPWR.n42 VPWR.n2 9.3005
R205 VPWR.n44 VPWR.n43 9.3005
R206 VPWR.n45 VPWR.n0 9.3005
R207 VPWR.n17 VPWR.n16 8.03187
R208 VPWR.n47 VPWR.n46 7.65871
R209 VPWR.n13 VPWR.n12 7.20521
R210 VPWR.n39 VPWR.n37 4.95232
R211 VPWR.n40 VPWR.n39 4.01802
R212 VPWR.n26 VPWR.n25 3.11401
R213 VPWR.n14 VPWR.n13 0.227696
R214 VPWR VPWR.n47 0.16305
R215 VPWR.n47 VPWR.n0 0.144791
R216 VPWR.n15 VPWR.n14 0.122949
R217 VPWR.n15 VPWR.n9 0.122949
R218 VPWR.n19 VPWR.n9 0.122949
R219 VPWR.n20 VPWR.n19 0.122949
R220 VPWR.n21 VPWR.n20 0.122949
R221 VPWR.n21 VPWR.n7 0.122949
R222 VPWR.n27 VPWR.n7 0.122949
R223 VPWR.n28 VPWR.n27 0.122949
R224 VPWR.n29 VPWR.n28 0.122949
R225 VPWR.n29 VPWR.n5 0.122949
R226 VPWR.n33 VPWR.n5 0.122949
R227 VPWR.n34 VPWR.n33 0.122949
R228 VPWR.n35 VPWR.n34 0.122949
R229 VPWR.n35 VPWR.n3 0.122949
R230 VPWR.n41 VPWR.n3 0.122949
R231 VPWR.n42 VPWR.n41 0.122949
R232 VPWR.n43 VPWR.n42 0.122949
R233 VPWR.n43 VPWR.n0 0.122949
R234 VPB.t5 VPB.t1 1361.16
R235 VPB.t9 VPB.t3 605.242
R236 VPB.t3 VPB.t7 500.538
R237 VPB.t1 VPB.t0 495.43
R238 VPB.t8 VPB.t5 469.892
R239 VPB.t13 VPB.t9 362.635
R240 VPB.t10 VPB.t8 316.668
R241 VPB VPB.t12 301.344
R242 VPB.t6 VPB.t13 275.807
R243 VPB.t0 VPB.t2 257.93
R244 VPB.t12 VPB.t11 255.376
R245 VPB.t4 VPB.t10 245.161
R246 VPB.t7 VPB.t4 229.839
R247 VPB.t14 VPB.t6 229.839
R248 VPB.t11 VPB.t14 214.517
R249 a_612_74.t1 a_612_74.n5 892.607
R250 a_612_74.n1 a_612_74.n0 506.675
R251 a_612_74.n0 a_612_74.t5 427.543
R252 a_612_74.n2 a_612_74.t7 285.988
R253 a_612_74.n2 a_612_74.n1 259.842
R254 a_612_74.n5 a_612_74.t0 220.471
R255 a_612_74.n4 a_612_74.t4 217.803
R256 a_612_74.n3 a_612_74.t6 204.048
R257 a_612_74.n0 a_612_74.t3 202.75
R258 a_612_74.n3 a_612_74.n2 201.418
R259 a_612_74.n1 a_612_74.t2 170.575
R260 a_612_74.n5 a_612_74.n4 152
R261 a_612_74.n4 a_612_74.n3 100.441
R262 a_1180_496.t0 a_1180_496.t1 154.786
R263 a_2216_94.t1 a_2216_94.n1 429.149
R264 a_2216_94.n0 a_2216_94.t3 285.36
R265 a_2216_94.n1 a_2216_94.t0 234.232
R266 a_2216_94.n1 a_2216_94.n0 178.183
R267 a_2216_94.n0 a_2216_94.t2 177.981
R268 Q_N.n1 Q_N 589.85
R269 Q_N.n1 Q_N.n0 585
R270 Q_N.n2 Q_N.n1 585
R271 Q_N.t0 Q_N.n3 279.738
R272 Q_N.n4 Q_N.t0 246.054
R273 Q_N.n1 Q_N.t1 26.3844
R274 Q_N Q_N.n4 15.5214
R275 Q_N.n2 Q_N 12.9944
R276 Q_N.n3 Q_N 12.2358
R277 Q_N.n0 Q_N 11.249
R278 Q_N.n0 Q_N 3.10353
R279 Q_N.n4 Q_N 1.69462
R280 Q_N.n3 Q_N 1.69462
R281 Q_N Q_N.n2 1.35808
R282 a_1681_74.t0 a_1681_74.t1 60.0005
R283 a_407_464.t0 a_407_464.t1 120.047
R284 a_233_464.t0 a_233_464.t1 83.1099
R285 CLK.n0 CLK.t0 261.62
R286 CLK.n0 CLK.t1 210.766
R287 CLK CLK.n0 184.73
R288 Q.n0 Q.t1 297.19
R289 Q.t0 Q.n0 279.738
R290 Q.n1 Q.t0 279.738
R291 Q.n1 Q 10.0246
R292 Q.n0 Q 3.85592
R293 Q Q.n1 1.38845
C0 VGND VPB 0.029445f
C1 a_1691_508# a_1723_48# 5.77e-19
C2 Q_N a_1723_48# 0.004292f
C3 VGND SCD 0.017164f
C4 a_1691_508# VPWR 0.006778f
C5 Q_N VPWR 0.119481f
C6 SCE VPB 0.142109f
C7 VPB CLK 0.047896f
C8 SCE SCD 0.038515f
C9 Q VPB 0.012569f
C10 SCE VGND 0.074943f
C11 CLK SCD 0.037503f
C12 VGND CLK 0.018756f
C13 VPB a_1723_48# 0.273407f
C14 Q VGND 0.115683f
C15 VPB VPWR 0.3711f
C16 D VPB 0.068224f
C17 VGND a_1723_48# 0.21937f
C18 VPWR SCD 0.016082f
C19 VGND VPWR 0.198162f
C20 D SCD 0.018094f
C21 Q_N VPB 0.014266f
C22 D VGND 0.012536f
C23 VGND a_1691_508# 5.47e-19
C24 Q_N VGND 0.094807f
C25 SCE VPWR 0.043747f
C26 D SCE 0.119402f
C27 Q a_1723_48# 0.08935f
C28 VPWR CLK 0.016322f
C29 Q VPWR 0.12618f
C30 VPWR a_1723_48# 0.321669f
C31 VPB SCD 0.08747f
C32 D VPWR 0.014593f
C33 Q_N VNB 0.111215f
C34 Q VNB 0.016794f
C35 VGND VNB 1.44354f
C36 CLK VNB 0.1502f
C37 SCD VNB 0.136516f
C38 D VNB 0.129052f
C39 SCE VNB 0.354942f
C40 VPWR VNB 1.11603f
C41 VPB VNB 2.87035f
C42 a_1723_48# VNB 0.485832f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfstp_4 VNB VPB VPWR SET_B VGND CLK SCE D SCD Q
X0 VPWR.t9 SCE.t0 a_27_74.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1824 ps=1.85 w=0.64 l=0.15
X1 a_803_74.t0 a_616_74.t2 VPWR.t11 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.3256 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_222_74.t0 a_27_74.t2 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 a_1677_74.t0 a_1017_81.t4 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.172 ps=1.26 w=0.64 l=0.15
X4 a_1445_74.t0 a_1017_81.t5 a_1201_55.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5 VPWR.t15 CLK.t0 a_616_74.t1 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 a_803_74.t1 a_616_74.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 a_417_74.t1 SCE.t1 a_288_464.t4 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.09135 ps=0.855 w=0.42 l=0.15
X8 a_1823_524.t1 a_616_74.t4 a_1620_373.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.195 as=0.126 ps=1.14 w=0.84 l=0.15
X9 VGND.t10 a_2580_74.t3 Q.t5 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.25955 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_1620_373.t0 a_616_74.t5 a_1823_524.t0 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2328 ps=2.27 w=0.84 l=0.15
X11 a_1677_74.t1 a_803_74.t2 a_1823_524.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X12 Q.t4 a_2580_74.t4 VGND.t11 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.16095 pd=1.175 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 VGND.t9 SCE.t2 a_27_74.t0 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.1197 ps=1.41 w=0.42 l=0.15
X14 a_1017_81.t0 a_616_74.t6 a_288_464.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1765 ps=1.73 w=0.42 l=0.15
X15 VGND.t8 CLK.t1 a_616_74.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X16 VPWR.t8 a_2580_74.t5 Q.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_2149_74.t0 a_616_74.t7 a_1823_524.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.10695 ps=1 w=0.42 l=0.15
X18 VPWR.t4 a_1823_524.t6 a_2580_74.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.126 ps=1.14 w=0.84 l=0.15
X19 a_2580_74.t0 a_1823_524.t7 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1302 ps=1.195 w=0.84 l=0.15
X20 a_2103_508.t1 a_803_74.t3 a_1823_524.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1302 ps=1.195 w=0.42 l=0.15
X21 a_288_464.t3 D.t0 a_222_74.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.09135 pd=0.855 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 VGND.t5 a_2580_74.t6 Q.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.16095 ps=1.175 w=0.74 l=0.15
X23 a_1823_524.t5 SET_B.t0 VPWR.t12 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X24 a_288_464.t5 D.t1 a_204_464.t0 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1536 pd=1.12 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 VPWR.t14 a_2191_180.t1 a_2103_508.t0 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.09975 ps=0.895 w=0.42 l=0.15
X26 VGND.t6 a_1823_524.t8 a_2580_74.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X27 a_204_464.t1 SCE.t3 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.096 ps=0.94 w=0.64 l=0.15
X28 VGND.t1 SCD.t0 a_417_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X29 VPWR.t13 SET_B.t1 a_1201_55.t2 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.16695 pd=1.37 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_1201_55.t0 a_1017_81.t6 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.156925 ps=1.24 w=0.42 l=0.15
X31 VPWR.t6 a_2580_74.t7 Q.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X32 VPWR.t3 SCD.t1 a_414_464.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2954 pd=2.4 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 VPWR.t16 a_1201_55.t3 a_1140_495.t1 VPB.t23 sky130_fd_pr__pfet_01v8 ad=0.156925 pd=1.24 as=0.091175 ps=0.965 w=0.42 l=0.15
X34 a_1153_81# a_803_74.t4 a_1017_81.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1113 ps=0.95 w=0.42 l=0.15
X35 Q.t0 a_2580_74.t8 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1862 ps=1.475 w=1.12 l=0.15
X36 a_414_464.t0 a_27_74.t3 a_288_464.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1536 ps=1.12 w=0.64 l=0.15
X37 VGND.t4 SET_B.t2 a_2227_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1092 pd=0.94 as=0.0819 ps=0.81 w=0.42 l=0.15
X38 a_2227_74.t0 a_2191_180.t2 a_2149_74.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X39 VPWR.t1 a_1017_81.t7 a_1620_373.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.23175 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X40 a_1017_81.t3 a_803_74.t5 a_288_464.t2 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.097475 pd=0.995 as=0.1239 ps=1.43 w=0.42 l=0.15
X41 a_1140_495.t0 a_616_74.t8 a_1017_81.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.091175 pd=0.965 as=0.097475 ps=0.995 w=0.42 l=0.15
X42 a_1620_373.t2 a_1017_81.t8 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.16695 ps=1.37 w=0.84 l=0.15
X43 a_2191_180.t0 a_1823_524.t9 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1092 ps=0.94 w=0.42 l=0.15
R0 SCE SCE.t1 463.238
R1 SCE.n1 SCE.t2 314.507
R2 SCE.n0 SCE.t3 153.63
R3 SCE.n0 SCE.t0 152.775
R4 SCE SCE.n1 75.406
R5 SCE.n1 SCE.n0 25.7745
R6 a_27_74.n1 a_27_74.t3 453.644
R7 a_27_74.t1 a_27_74.n1 360.479
R8 a_27_74.n0 a_27_74.t2 342.521
R9 a_27_74.n0 a_27_74.t0 236.008
R10 a_27_74.n1 a_27_74.n0 82.4325
R11 VPWR.n60 VPWR.t3 787.665
R12 VPWR.n9 VPWR.n8 673.53
R13 VPWR.n39 VPWR.t1 658.662
R14 VPWR.n27 VPWR.t5 653.393
R15 VPWR.n45 VPWR.n11 640.718
R16 VPWR.n32 VPWR.n16 611.369
R17 VPWR.n66 VPWR.n1 606.333
R18 VPWR.n58 VPWR.n5 606.333
R19 VPWR.n21 VPWR.t6 342.784
R20 VPWR.n25 VPWR.n20 317.716
R21 VPWR.n22 VPWR.t8 255.333
R22 VPWR.n11 VPWR.t13 178.238
R23 VPWR.n8 VPWR.t0 164.167
R24 VPWR.n8 VPWR.t16 110.227
R25 VPWR.n16 VPWR.t12 70.3576
R26 VPWR.n16 VPWR.t14 70.3576
R27 VPWR.n1 VPWR.t10 46.1724
R28 VPWR.n1 VPWR.t9 46.1724
R29 VPWR.n20 VPWR.t7 43.8979
R30 VPWR.n11 VPWR.t2 38.6969
R31 VPWR.n64 VPWR.n2 36.1417
R32 VPWR.n65 VPWR.n64 36.1417
R33 VPWR.n52 VPWR.n51 36.1417
R34 VPWR.n53 VPWR.n52 36.1417
R35 VPWR.n53 VPWR.n6 36.1417
R36 VPWR.n57 VPWR.n6 36.1417
R37 VPWR.n44 VPWR.n12 36.1417
R38 VPWR.n47 VPWR.n46 36.1417
R39 VPWR.n33 VPWR.n14 36.1417
R40 VPWR.n37 VPWR.n14 36.1417
R41 VPWR.n38 VPWR.n37 36.1417
R42 VPWR.n40 VPWR.n38 36.1417
R43 VPWR.n27 VPWR.n17 36.1417
R44 VPWR.n31 VPWR.n17 36.1417
R45 VPWR.n20 VPWR.t4 35.1791
R46 VPWR.n59 VPWR.n58 33.8829
R47 VPWR.n47 VPWR.n9 32.7534
R48 VPWR.n60 VPWR.n2 30.1181
R49 VPWR.n32 VPWR.n31 28.9887
R50 VPWR.n46 VPWR.n45 27.1064
R51 VPWR.n5 VPWR.t11 26.3844
R52 VPWR.n5 VPWR.t15 26.3844
R53 VPWR.n26 VPWR.n25 25.6005
R54 VPWR.n24 VPWR.n21 25.224
R55 VPWR.n33 VPWR.n32 24.4711
R56 VPWR.n66 VPWR.n65 23.7181
R57 VPWR.n25 VPWR.n24 21.8358
R58 VPWR.n51 VPWR.n9 20.7064
R59 VPWR.n60 VPWR.n59 17.3181
R60 VPWR.n27 VPWR.n26 17.3181
R61 VPWR.n58 VPWR.n57 13.5534
R62 VPWR.n39 VPWR.n12 10.1652
R63 VPWR.n24 VPWR.n23 9.3005
R64 VPWR.n25 VPWR.n19 9.3005
R65 VPWR.n26 VPWR.n18 9.3005
R66 VPWR.n28 VPWR.n27 9.3005
R67 VPWR.n29 VPWR.n17 9.3005
R68 VPWR.n31 VPWR.n30 9.3005
R69 VPWR.n32 VPWR.n15 9.3005
R70 VPWR.n34 VPWR.n33 9.3005
R71 VPWR.n35 VPWR.n14 9.3005
R72 VPWR.n37 VPWR.n36 9.3005
R73 VPWR.n38 VPWR.n13 9.3005
R74 VPWR.n41 VPWR.n40 9.3005
R75 VPWR.n42 VPWR.n12 9.3005
R76 VPWR.n44 VPWR.n43 9.3005
R77 VPWR.n46 VPWR.n10 9.3005
R78 VPWR.n48 VPWR.n47 9.3005
R79 VPWR.n49 VPWR.n9 9.3005
R80 VPWR.n51 VPWR.n50 9.3005
R81 VPWR.n52 VPWR.n7 9.3005
R82 VPWR.n54 VPWR.n53 9.3005
R83 VPWR.n55 VPWR.n6 9.3005
R84 VPWR.n57 VPWR.n56 9.3005
R85 VPWR.n58 VPWR.n4 9.3005
R86 VPWR.n59 VPWR.n3 9.3005
R87 VPWR.n61 VPWR.n60 9.3005
R88 VPWR.n62 VPWR.n2 9.3005
R89 VPWR.n64 VPWR.n63 9.3005
R90 VPWR.n65 VPWR.n0 9.3005
R91 VPWR.n45 VPWR.n44 9.03579
R92 VPWR.n67 VPWR.n66 7.23624
R93 VPWR.n22 VPWR.n21 6.50549
R94 VPWR.n40 VPWR.n39 1.12991
R95 VPWR.n23 VPWR.n22 0.686474
R96 VPWR VPWR.n67 0.157488
R97 VPWR.n67 VPWR.n0 0.150282
R98 VPWR.n23 VPWR.n19 0.122949
R99 VPWR.n19 VPWR.n18 0.122949
R100 VPWR.n28 VPWR.n18 0.122949
R101 VPWR.n29 VPWR.n28 0.122949
R102 VPWR.n30 VPWR.n29 0.122949
R103 VPWR.n30 VPWR.n15 0.122949
R104 VPWR.n34 VPWR.n15 0.122949
R105 VPWR.n35 VPWR.n34 0.122949
R106 VPWR.n36 VPWR.n35 0.122949
R107 VPWR.n36 VPWR.n13 0.122949
R108 VPWR.n41 VPWR.n13 0.122949
R109 VPWR.n42 VPWR.n41 0.122949
R110 VPWR.n43 VPWR.n42 0.122949
R111 VPWR.n43 VPWR.n10 0.122949
R112 VPWR.n48 VPWR.n10 0.122949
R113 VPWR.n49 VPWR.n48 0.122949
R114 VPWR.n50 VPWR.n49 0.122949
R115 VPWR.n50 VPWR.n7 0.122949
R116 VPWR.n54 VPWR.n7 0.122949
R117 VPWR.n55 VPWR.n54 0.122949
R118 VPWR.n56 VPWR.n55 0.122949
R119 VPWR.n56 VPWR.n4 0.122949
R120 VPWR.n4 VPWR.n3 0.122949
R121 VPWR.n61 VPWR.n3 0.122949
R122 VPWR.n62 VPWR.n61 0.122949
R123 VPWR.n63 VPWR.n62 0.122949
R124 VPWR.n63 VPWR.n0 0.122949
R125 VPB.t19 VPB.t7 773.79
R126 VPB.t18 VPB.t17 577.152
R127 VPB.t3 VPB.t22 559.274
R128 VPB.t1 VPB.t16 515.861
R129 VPB.t8 VPB.t11 459.678
R130 VPB.t23 VPB.t0 375.404
R131 VPB.t20 VPB.t2 347.312
R132 VPB.t14 VPB.t5 321.774
R133 VPB.t10 VPB.t21 319.221
R134 VPB.t17 VPB.t4 273.253
R135 VPB.t6 VPB.t9 257.93
R136 VPB.t15 VPB.t10 257.93
R137 VPB.t4 VPB.t23 257.93
R138 VPB VPB.t13 252.823
R139 VPB.t0 VPB.t20 245.161
R140 VPB.t9 VPB.t8 229.839
R141 VPB.t7 VPB.t6 229.839
R142 VPB.t21 VPB.t19 229.839
R143 VPB.t16 VPB.t15 229.839
R144 VPB.t2 VPB.t1 229.839
R145 VPB.t22 VPB.t18 229.839
R146 VPB.t13 VPB.t12 229.839
R147 VPB.t5 VPB.t3 214.517
R148 VPB.t12 VPB.t14 214.517
R149 a_616_74.n1 a_616_74.n0 1222.35
R150 a_616_74.t1 a_616_74.n5 862.136
R151 a_616_74.t4 a_616_74.t7 788.874
R152 a_616_74.n2 a_616_74.n1 771.447
R153 a_616_74.n2 a_616_74.t6 367.928
R154 a_616_74.n0 a_616_74.t4 299.447
R155 a_616_74.n3 a_616_74.t2 226.809
R156 a_616_74.n5 a_616_74.t0 212.448
R157 a_616_74.n5 a_616_74.n4 199.399
R158 a_616_74.n3 a_616_74.t3 198.935
R159 a_616_74.n0 a_616_74.t5 159.06
R160 a_616_74.n1 a_616_74.t8 91.5805
R161 a_616_74.n4 a_616_74.n2 58.4247
R162 a_616_74.n4 a_616_74.n3 13.146
R163 a_803_74.n6 a_803_74.n5 726.782
R164 a_803_74.n0 a_803_74.t1 471.89
R165 a_803_74.n4 a_803_74.t3 440.779
R166 a_803_74.n4 a_803_74.n3 383.361
R167 a_803_74.n5 a_803_74.n4 343.8
R168 a_803_74.n1 a_803_74.t4 321.041
R169 a_803_74.n3 a_803_74.n2 265.101
R170 a_803_74.n0 a_803_74.t5 220.113
R171 a_803_74.n5 a_803_74.n1 214.839
R172 a_803_74.n6 a_803_74.t0 167.374
R173 a_803_74.n3 a_803_74.t2 126.927
R174 a_803_74.n1 a_803_74.n0 115.972
R175 VGND.n55 VGND.t1 246.139
R176 VGND.n18 VGND.t5 232.721
R177 VGND.n62 VGND.n61 206.139
R178 VGND.n13 VGND.n12 198.185
R179 VGND.n17 VGND.t10 156.154
R180 VGND.n16 VGND.n15 116.644
R181 VGND.n53 VGND.n4 116.288
R182 VGND.n8 VGND.t2 98.9807
R183 VGND.n12 VGND.t7 84.2862
R184 VGND.n12 VGND.t4 64.2862
R185 VGND.n61 VGND.t9 60.0005
R186 VGND.n61 VGND.t3 51.4291
R187 VGND.n24 VGND.n23 36.1417
R188 VGND.n25 VGND.n24 36.1417
R189 VGND.n30 VGND.n29 36.1417
R190 VGND.n31 VGND.n30 36.1417
R191 VGND.n31 VGND.n10 36.1417
R192 VGND.n35 VGND.n10 36.1417
R193 VGND.n42 VGND.n41 36.1417
R194 VGND.n47 VGND.n6 36.1417
R195 VGND.n48 VGND.n47 36.1417
R196 VGND.n49 VGND.n48 36.1417
R197 VGND.n49 VGND.n3 36.1417
R198 VGND.n59 VGND.n1 36.1417
R199 VGND.n60 VGND.n59 36.1417
R200 VGND.n15 VGND.t6 34.0546
R201 VGND.n4 VGND.t8 34.0546
R202 VGND.n19 VGND.n16 33.8829
R203 VGND.n54 VGND.n53 33.1299
R204 VGND.n43 VGND.n42 31.624
R205 VGND.n37 VGND.n36 29.3652
R206 VGND.n29 VGND.n13 27.8593
R207 VGND.n55 VGND.n54 25.6005
R208 VGND.n15 VGND.t11 22.7032
R209 VGND.n4 VGND.t0 22.7032
R210 VGND.n55 VGND.n1 21.8358
R211 VGND.n62 VGND.n60 19.2005
R212 VGND.n36 VGND.n35 18.0711
R213 VGND.n19 VGND.n18 17.6946
R214 VGND.n43 VGND.n6 15.8123
R215 VGND.n53 VGND.n3 14.3064
R216 VGND.n23 VGND.n16 13.5534
R217 VGND.n41 VGND.n8 11.2946
R218 VGND.n37 VGND.n8 10.5417
R219 VGND.n60 VGND.n0 9.3005
R220 VGND.n59 VGND.n58 9.3005
R221 VGND.n57 VGND.n1 9.3005
R222 VGND.n56 VGND.n55 9.3005
R223 VGND.n54 VGND.n2 9.3005
R224 VGND.n53 VGND.n52 9.3005
R225 VGND.n51 VGND.n3 9.3005
R226 VGND.n50 VGND.n49 9.3005
R227 VGND.n48 VGND.n5 9.3005
R228 VGND.n47 VGND.n46 9.3005
R229 VGND.n45 VGND.n6 9.3005
R230 VGND.n44 VGND.n43 9.3005
R231 VGND.n42 VGND.n7 9.3005
R232 VGND.n41 VGND.n40 9.3005
R233 VGND.n39 VGND.n8 9.3005
R234 VGND.n38 VGND.n37 9.3005
R235 VGND.n36 VGND.n9 9.3005
R236 VGND.n35 VGND.n34 9.3005
R237 VGND.n33 VGND.n10 9.3005
R238 VGND.n32 VGND.n31 9.3005
R239 VGND.n30 VGND.n11 9.3005
R240 VGND.n29 VGND.n28 9.3005
R241 VGND.n27 VGND.n13 9.3005
R242 VGND.n26 VGND.n25 9.3005
R243 VGND.n24 VGND.n14 9.3005
R244 VGND.n23 VGND.n22 9.3005
R245 VGND.n20 VGND.n19 9.3005
R246 VGND.n21 VGND.n16 9.3005
R247 VGND.n63 VGND.n62 7.43488
R248 VGND.n18 VGND.n17 6.96039
R249 VGND.n25 VGND.n13 6.77697
R250 VGND.n20 VGND.n17 0.594857
R251 VGND VGND.n63 0.160103
R252 VGND.n63 VGND.n0 0.1477
R253 VGND.n21 VGND.n20 0.122949
R254 VGND.n22 VGND.n21 0.122949
R255 VGND.n22 VGND.n14 0.122949
R256 VGND.n26 VGND.n14 0.122949
R257 VGND.n27 VGND.n26 0.122949
R258 VGND.n28 VGND.n27 0.122949
R259 VGND.n28 VGND.n11 0.122949
R260 VGND.n32 VGND.n11 0.122949
R261 VGND.n33 VGND.n32 0.122949
R262 VGND.n34 VGND.n33 0.122949
R263 VGND.n34 VGND.n9 0.122949
R264 VGND.n38 VGND.n9 0.122949
R265 VGND.n39 VGND.n38 0.122949
R266 VGND.n40 VGND.n39 0.122949
R267 VGND.n40 VGND.n7 0.122949
R268 VGND.n44 VGND.n7 0.122949
R269 VGND.n45 VGND.n44 0.122949
R270 VGND.n46 VGND.n45 0.122949
R271 VGND.n46 VGND.n5 0.122949
R272 VGND.n50 VGND.n5 0.122949
R273 VGND.n51 VGND.n50 0.122949
R274 VGND.n52 VGND.n51 0.122949
R275 VGND.n52 VGND.n2 0.122949
R276 VGND.n56 VGND.n2 0.122949
R277 VGND.n57 VGND.n56 0.122949
R278 VGND.n58 VGND.n57 0.122949
R279 VGND.n58 VGND.n0 0.122949
R280 a_222_74.t0 a_222_74.t1 68.5719
R281 VNB.t8 VNB.t5 3372.18
R282 VNB.t4 VNB.t9 3279.79
R283 VNB.t5 VNB.t4 2679.26
R284 VNB.t2 VNB.t1 2471.39
R285 VNB.t3 VNB.t14 2402.1
R286 VNB.t13 VNB.t12 2286.61
R287 VNB.t9 VNB.t0 2171.13
R288 VNB.t10 VNB.t18 2148.03
R289 VNB.t1 VNB.t8 1570.6
R290 VNB.t7 VNB.t13 1547.51
R291 VNB.t19 VNB.t10 1351.18
R292 VNB.t15 VNB.t17 1351.18
R293 VNB.t11 VNB.t7 1247.24
R294 VNB.t16 VNB.t6 1247.24
R295 VNB.t12 VNB.t19 1154.86
R296 VNB.t14 VNB.t2 1154.86
R297 VNB VNB.t16 1143.31
R298 VNB.t0 VNB.t11 900.788
R299 VNB.t17 VNB.t3 900.788
R300 VNB.t6 VNB.t15 900.788
R301 a_1017_81.n9 a_1017_81.n8 660.039
R302 a_1017_81.n3 a_1017_81.t7 274.204
R303 a_1017_81.n4 a_1017_81.t8 261.06
R304 a_1017_81.n6 a_1017_81.n4 235.103
R305 a_1017_81.n5 a_1017_81.t5 232.968
R306 a_1017_81.n0 a_1017_81.t6 230.825
R307 a_1017_81.n10 a_1017_81.n9 216.806
R308 a_1017_81.n2 a_1017_81.n1 183.161
R309 a_1017_81.n7 a_1017_81.n0 155.685
R310 a_1017_81.n6 a_1017_81.n5 152
R311 a_1017_81.n8 a_1017_81.t1 148.975
R312 a_1017_81.n2 a_1017_81.t4 137.881
R313 a_1017_81.t0 a_1017_81.n10 111.43
R314 a_1017_81.n9 a_1017_81.n7 86.5887
R315 a_1017_81.n8 a_1017_81.t3 72.295
R316 a_1017_81.n5 a_1017_81.n0 49.6611
R317 a_1017_81.n10 a_1017_81.t2 40.0005
R318 a_1017_81.n4 a_1017_81.n3 19.7187
R319 a_1017_81.n3 a_1017_81.n2 18.2581
R320 a_1017_81.n7 a_1017_81.n6 9.50353
R321 a_1677_74.t0 a_1677_74.t1 495.474
R322 a_1201_55.n1 a_1201_55.n0 827.918
R323 a_1201_55.t1 a_1201_55.n3 429.923
R324 a_1201_55.n3 a_1201_55.n1 213.688
R325 a_1201_55.n1 a_1201_55.t3 142.458
R326 a_1201_55.n3 a_1201_55.n2 126.927
R327 a_1201_55.n0 a_1201_55.t0 84.4291
R328 a_1201_55.n0 a_1201_55.t2 70.3576
R329 CLK.n0 CLK.t0 285.719
R330 CLK.n0 CLK.t1 178.34
R331 CLK CLK.n0 158.054
R332 a_288_464.n1 a_288_464.t2 660.409
R333 a_288_464.n3 a_288_464.n2 616.745
R334 a_288_464.n2 a_288_464.n0 340.32
R335 a_288_464.n1 a_288_464.t0 338.577
R336 a_288_464.n2 a_288_464.n1 164.894
R337 a_288_464.t1 a_288_464.n3 73.8755
R338 a_288_464.n3 a_288_464.t5 73.8755
R339 a_288_464.n0 a_288_464.t4 62.8576
R340 a_288_464.n0 a_288_464.t3 61.4291
R341 a_417_74.t0 a_417_74.t1 68.5719
R342 a_1620_373.n1 a_1620_373.n0 683.327
R343 a_1620_373.n0 a_1620_373.t1 35.1791
R344 a_1620_373.n0 a_1620_373.t0 35.1791
R345 a_1620_373.n1 a_1620_373.t3 35.1791
R346 a_1620_373.t2 a_1620_373.n1 35.1791
R347 a_1823_524.n8 a_1823_524.t0 681.774
R348 a_1823_524.n6 a_1823_524.t5 669.128
R349 a_1823_524.n9 a_1823_524.n8 585
R350 a_1823_524.n1 a_1823_524.t8 369.534
R351 a_1823_524.n5 a_1823_524.t9 271.664
R352 a_1823_524.n1 a_1823_524.t6 228.821
R353 a_1823_524.n4 a_1823_524.n3 211.673
R354 a_1823_524.n0 a_1823_524.t4 191.082
R355 a_1823_524.n0 a_1823_524.t2 159.369
R356 a_1823_524.n2 a_1823_524.t7 159.06
R357 a_1823_524.n4 a_1823_524.n2 132.421
R358 a_1823_524.n7 a_1823_524.n0 122.99
R359 a_1823_524.n6 a_1823_524.n5 118.188
R360 a_1823_524.n2 a_1823_524.n1 72.9743
R361 a_1823_524.n9 a_1823_524.t3 72.7029
R362 a_1823_524.t1 a_1823_524.n9 63.3219
R363 a_1823_524.n8 a_1823_524.n7 62.141
R364 a_1823_524.n7 a_1823_524.n6 41.7887
R365 a_1823_524.n5 a_1823_524.n4 22.592
R366 a_2580_74.n14 a_2580_74.n13 348.807
R367 a_2580_74.n3 a_2580_74.t5 302.322
R368 a_2580_74.n4 a_2580_74.n2 234.841
R369 a_2580_74.n7 a_2580_74.t7 234.841
R370 a_2580_74.n10 a_2580_74.t8 234.841
R371 a_2580_74.n11 a_2580_74.t4 199.519
R372 a_2580_74.n3 a_2580_74.t3 186.374
R373 a_2580_74.n8 a_2580_74.t6 186.374
R374 a_2580_74.n5 a_2580_74.n1 186.374
R375 a_2580_74.n6 a_2580_74.n0 165.189
R376 a_2580_74.n13 a_2580_74.t2 164.47
R377 a_2580_74.n12 a_2580_74.n11 152
R378 a_2580_74.n9 a_2580_74.n0 152
R379 a_2580_74.n4 a_2580_74.n3 109.546
R380 a_2580_74.n6 a_2580_74.n5 46.0096
R381 a_2580_74.t1 a_2580_74.n14 35.1791
R382 a_2580_74.n14 a_2580_74.t0 35.1791
R383 a_2580_74.n10 a_2580_74.n9 29.9429
R384 a_2580_74.n13 a_2580_74.n12 23.0793
R385 a_2580_74.n9 a_2580_74.n8 22.6399
R386 a_2580_74.n11 a_2580_74.n10 19.7187
R387 a_2580_74.n7 a_2580_74.n6 13.8763
R388 a_2580_74.n12 a_2580_74.n0 13.1884
R389 a_2580_74.n8 a_2580_74.n7 13.146
R390 a_2580_74.n5 a_2580_74.n4 5.84292
R391 Q.n1 Q.n0 237.351
R392 Q.n1 Q.t2 232.788
R393 Q.n3 Q.n2 150.994
R394 Q.n3 Q.t5 148.827
R395 Q Q.n3 43.3472
R396 Q Q.n1 37.6476
R397 Q.n2 Q.t4 36.487
R398 Q.n2 Q.t3 34.0546
R399 Q.n0 Q.t1 26.3844
R400 Q.n0 Q.t0 26.3844
R401 a_2191_180.t0 a_2191_180.n0 474.623
R402 a_2191_180.n0 a_2191_180.t1 446.387
R403 a_2191_180.n0 a_2191_180.t2 126.927
R404 a_2149_74.t0 a_2149_74.t1 68.5719
R405 a_2103_508.t0 a_2103_508.t1 222.798
R406 D.n0 D.t0 422.553
R407 D.n0 D.t1 176.466
R408 D D.n0 163.442
R409 SET_B.n0 SET_B.t2 325.837
R410 SET_B.n2 SET_B.n1 298.497
R411 SET_B.n2 SET_B.t1 225.661
R412 SET_B.n0 SET_B.t0 219.55
R413 SET_B SET_B.n2 168.113
R414 SET_B SET_B.n0 78.4174
R415 a_204_464.t0 a_204_464.t1 83.1099
R416 SCD.n2 SCD.t0 181.959
R417 SCD.n4 SCD.t1 177.942
R418 SCD.n3 SCD.n0 152
R419 SCD.n2 SCD.n1 152
R420 SCD.n5 SCD.n4 152
R421 SCD.n4 SCD.n3 30.6323
R422 SCD.n3 SCD.n2 30.6323
R423 SCD.n5 SCD.n0 15.5434
R424 SCD.n1 SCD 14.4005
R425 SCD.n1 SCD 2.51479
R426 SCD SCD.n0 1.14336
R427 SCD SCD.n5 0.229071
R428 a_414_464.t0 a_414_464.t1 83.1099
R429 a_1140_495.n0 a_1140_495.t1 140.409
R430 a_1140_495.n1 a_1140_495.n0 70.6231
R431 a_1140_495.n0 a_1140_495.t0 13.117
R432 a_2227_74.t0 a_2227_74.t1 111.43
C0 VPWR a_1153_81# 4.97e-19
C1 VGND VPB 0.025875f
C2 D SCD 0.004868f
C3 SCE SCD 0.061333f
C4 VPWR VPB 0.408291f
C5 VGND CLK 0.037189f
C6 VGND Q 0.357339f
C7 VGND SCD 0.038212f
C8 D SET_B 2.79e-20
C9 SCE SET_B 9.05e-20
C10 CLK VPWR 0.015542f
C11 VPWR Q 0.395904f
C12 VPWR SCD 0.017174f
C13 CLK VPB 0.033627f
C14 VGND SET_B 0.172881f
C15 Q VPB 0.014713f
C16 SCD VPB 0.104014f
C17 SCE D 0.182182f
C18 VPWR SET_B 0.15371f
C19 VGND D 0.013074f
C20 CLK SCD 0.027907f
C21 VGND SCE 0.035793f
C22 SET_B VPB 0.201214f
C23 VPWR D 0.012797f
C24 VPWR SCE 0.033689f
C25 D VPB 0.071904f
C26 VGND a_1153_81# 0.004492f
C27 CLK SET_B 8.73e-20
C28 Q SET_B 1.78e-19
C29 SCE VPB 0.13131f
C30 SCD SET_B 1.12e-19
C31 VGND VPWR 0.179005f
C32 Q VNB 0.057038f
C33 VGND VNB 1.85776f
C34 SET_B VNB 0.293546f
C35 CLK VNB 0.114114f
C36 VPWR VNB 1.42372f
C37 SCD VNB 0.168388f
C38 D VNB 0.117336f
C39 SCE VNB 0.328257f
C40 VPB VNB 3.6203f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfstp_2 VNB VPB VPWR SET_B VGND CLK SCE D SCD Q
X0 VPWR.t10 SCD.t0 a_416_464.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.2749 pd=2.35 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_2186_367.t0 a_1804_424.t5 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.14385 ps=1.105 w=0.42 l=0.15
X2 a_416_464.t0 a_27_74.t2 a_290_464.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1536 ps=1.12 w=0.64 l=0.15
X3 a_403_74.t0 SCE.t0 a_290_464.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VGND.t0 CLK.t0 a_608_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_795_74.t1 a_608_74.t2 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3076 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_991_81.t1 a_608_74.t3 a_290_464.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1281 pd=1.03 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 VPWR.t7 a_1804_424.t6 a_2611_98.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR.t1 CLK.t1 a_608_74.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X9 VPWR.t4 SET_B.t0 a_1185_55.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.325 as=0.07245 ps=0.765 w=0.42 l=0.15
X10 VGND.t8 SCE.t1 a_27_74.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.09975 pd=0.895 as=0.1197 ps=1.41 w=0.42 l=0.15
X11 a_1117_483.t0 a_608_74.t4 a_991_81.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0857 pd=0.89 as=0.092225 ps=0.935 w=0.42 l=0.15
X12 VPWR.t15 a_1185_55.t3 a_1117_483.t1 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.11235 pd=0.955 as=0.0857 ps=0.89 w=0.42 l=0.15
X13 a_2141_508.t1 a_795_74.t2 a_1804_424.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.17955 ps=1.43 w=0.42 l=0.15
X14 VPWR.t11 SCE.t2 a_27_74.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1888 ps=1.87 w=0.64 l=0.15
X15 a_290_464.t3 D.t0 a_239_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X16 Q.t1 a_2611_98.t2 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1345 ps=1.115 w=0.74 l=0.15
X17 VGND.t9 SCD.t1 a_403_74.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0672 ps=0.74 w=0.42 l=0.15
X18 a_991_81.t2 a_795_74.t3 a_290_464.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.092225 pd=0.935 as=0.1239 ps=1.43 w=0.42 l=0.15
X19 a_1804_424.t0 a_608_74.t5 a_1584_379.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.17955 pd=1.43 as=0.126 ps=1.14 w=0.84 l=0.15
X20 a_1429_74.t0 a_991_81.t3 a_1185_55.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X21 VPWR.t8 a_1804_424.t7 a_2186_367.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.15
X22 a_2219_74.t0 a_2186_367.t2 a_2141_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 VPWR.t6 a_991_81.t4 a_1584_379.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=2.24 as=0.126 ps=1.14 w=0.84 l=0.15
X24 a_2141_74.t1 a_608_74.t6 a_1804_424.t4 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X25 VGND.t7 a_2611_98.t3 Q.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=2.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 a_1641_74.t0 a_991_81.t5 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1367 ps=1.16 w=0.64 l=0.15
X27 a_1584_379.t1 a_991_81.t6 VPWR.t13 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1638 ps=1.325 w=0.84 l=0.15
X28 a_1185_55.t0 a_991_81.t7 VPWR.t14 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.07245 pd=0.765 as=0.11235 ps=0.955 w=0.42 l=0.15
X29 VGND.t3 a_1804_424.t8 a_2611_98.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1345 pd=1.115 as=0.1824 ps=1.85 w=0.64 l=0.15
X30 a_795_74.t0 a_608_74.t7 VGND.t10 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1295 ps=1.09 w=0.74 l=0.15
X31 a_290_464.t4 D.t1 a_206_464.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1536 pd=1.12 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 a_239_74.t0 a_27_74.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.09975 ps=0.895 w=0.42 l=0.15
X33 a_1804_424.t2 a_795_74.t4 a_1641_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.101 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X34 VGND.t5 SET_B.t1 a_2219_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.14385 pd=1.105 as=0.0882 ps=0.84 w=0.42 l=0.15
X35 a_1804_424.t3 SET_B.t2 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X36 VPWR.t2 a_2611_98.t4 Q.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X37 a_206_464.t0 SCE.t3 VPWR.t12 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.096 ps=0.94 w=0.64 l=0.15
X38 VPWR.t0 a_2186_367.t3 a_2141_508.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X39 Q.t2 a_2611_98.t5 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1934 ps=1.475 w=1.12 l=0.15
R0 SCD.n2 SCD.t1 196.013
R1 SCD.n0 SCD.t0 168.433
R2 SCD SCD.n0 153.992
R3 SCD.n4 SCD.n3 152
R4 SCD.n2 SCD.n1 152
R5 SCD.n3 SCD.n0 33.1076
R6 SCD.n3 SCD.n2 33.1076
R7 SCD SCD.n4 17.3516
R8 SCD.n1 SCD 15.6449
R9 SCD.n1 SCD 5.40494
R10 SCD.n4 SCD 3.69828
R11 a_416_464.t0 a_416_464.t1 83.1099
R12 VPWR.n38 VPWR.t6 809.846
R13 VPWR.n57 VPWR.t10 801.591
R14 VPWR.n25 VPWR.t8 675.333
R15 VPWR.n9 VPWR.n8 622.889
R16 VPWR.n17 VPWR.n16 611.625
R17 VPWR.n63 VPWR.n1 606.333
R18 VPWR.n55 VPWR.n5 606.333
R19 VPWR.n12 VPWR.n11 349.587
R20 VPWR.n22 VPWR.t2 349.481
R21 VPWR.n21 VPWR.n20 227.151
R22 VPWR.n8 VPWR.t14 178.238
R23 VPWR.n11 VPWR.t4 157.131
R24 VPWR.n8 VPWR.t15 72.7029
R25 VPWR.n16 VPWR.t9 70.3576
R26 VPWR.n16 VPWR.t0 70.3576
R27 VPWR.n1 VPWR.t12 46.1724
R28 VPWR.n1 VPWR.t11 46.1724
R29 VPWR.n20 VPWR.t7 39.4005
R30 VPWR.n61 VPWR.n2 36.1417
R31 VPWR.n62 VPWR.n61 36.1417
R32 VPWR.n49 VPWR.n48 36.1417
R33 VPWR.n50 VPWR.n49 36.1417
R34 VPWR.n50 VPWR.n6 36.1417
R35 VPWR.n54 VPWR.n6 36.1417
R36 VPWR.n40 VPWR.n39 36.1417
R37 VPWR.n44 VPWR.n43 36.1417
R38 VPWR.n45 VPWR.n44 36.1417
R39 VPWR.n32 VPWR.n31 36.1417
R40 VPWR.n33 VPWR.n32 36.1417
R41 VPWR.n33 VPWR.n14 36.1417
R42 VPWR.n37 VPWR.n14 36.1417
R43 VPWR.n27 VPWR.n26 36.1417
R44 VPWR.n11 VPWR.t13 35.1791
R45 VPWR.n27 VPWR.n17 32.377
R46 VPWR.n56 VPWR.n55 32.0005
R47 VPWR.n57 VPWR.n2 30.1181
R48 VPWR.n20 VPWR.t3 28.5357
R49 VPWR.n25 VPWR.n24 27.1064
R50 VPWR.n5 VPWR.t5 26.3844
R51 VPWR.n5 VPWR.t1 26.3844
R52 VPWR.n24 VPWR.n21 25.6005
R53 VPWR.n63 VPWR.n62 22.9652
R54 VPWR.n40 VPWR.n12 22.5887
R55 VPWR.n31 VPWR.n17 21.0829
R56 VPWR.n26 VPWR.n25 20.3299
R57 VPWR.n57 VPWR.n56 17.3181
R58 VPWR.n55 VPWR.n54 15.4358
R59 VPWR.n38 VPWR.n37 14.6829
R60 VPWR.n43 VPWR.n12 13.5534
R61 VPWR.n45 VPWR.n9 10.1652
R62 VPWR.n24 VPWR.n23 9.3005
R63 VPWR.n25 VPWR.n19 9.3005
R64 VPWR.n26 VPWR.n18 9.3005
R65 VPWR.n28 VPWR.n27 9.3005
R66 VPWR.n29 VPWR.n17 9.3005
R67 VPWR.n31 VPWR.n30 9.3005
R68 VPWR.n32 VPWR.n15 9.3005
R69 VPWR.n34 VPWR.n33 9.3005
R70 VPWR.n35 VPWR.n14 9.3005
R71 VPWR.n37 VPWR.n36 9.3005
R72 VPWR.n39 VPWR.n13 9.3005
R73 VPWR.n41 VPWR.n40 9.3005
R74 VPWR.n43 VPWR.n42 9.3005
R75 VPWR.n44 VPWR.n10 9.3005
R76 VPWR.n46 VPWR.n45 9.3005
R77 VPWR.n48 VPWR.n47 9.3005
R78 VPWR.n49 VPWR.n7 9.3005
R79 VPWR.n51 VPWR.n50 9.3005
R80 VPWR.n52 VPWR.n6 9.3005
R81 VPWR.n54 VPWR.n53 9.3005
R82 VPWR.n55 VPWR.n4 9.3005
R83 VPWR.n56 VPWR.n3 9.3005
R84 VPWR.n58 VPWR.n57 9.3005
R85 VPWR.n59 VPWR.n2 9.3005
R86 VPWR.n61 VPWR.n60 9.3005
R87 VPWR.n62 VPWR.n0 9.3005
R88 VPWR.n64 VPWR.n63 7.27223
R89 VPWR.n48 VPWR.n9 7.15344
R90 VPWR.n22 VPWR.n21 6.71896
R91 VPWR.n39 VPWR.n38 2.63579
R92 VPWR.n23 VPWR.n22 0.636081
R93 VPWR VPWR.n64 0.157962
R94 VPWR.n64 VPWR.n0 0.149814
R95 VPWR.n23 VPWR.n19 0.122949
R96 VPWR.n19 VPWR.n18 0.122949
R97 VPWR.n28 VPWR.n18 0.122949
R98 VPWR.n29 VPWR.n28 0.122949
R99 VPWR.n30 VPWR.n29 0.122949
R100 VPWR.n30 VPWR.n15 0.122949
R101 VPWR.n34 VPWR.n15 0.122949
R102 VPWR.n35 VPWR.n34 0.122949
R103 VPWR.n36 VPWR.n35 0.122949
R104 VPWR.n36 VPWR.n13 0.122949
R105 VPWR.n41 VPWR.n13 0.122949
R106 VPWR.n42 VPWR.n41 0.122949
R107 VPWR.n42 VPWR.n10 0.122949
R108 VPWR.n46 VPWR.n10 0.122949
R109 VPWR.n47 VPWR.n46 0.122949
R110 VPWR.n47 VPWR.n7 0.122949
R111 VPWR.n51 VPWR.n7 0.122949
R112 VPWR.n52 VPWR.n51 0.122949
R113 VPWR.n53 VPWR.n52 0.122949
R114 VPWR.n53 VPWR.n4 0.122949
R115 VPWR.n4 VPWR.n3 0.122949
R116 VPWR.n58 VPWR.n3 0.122949
R117 VPWR.n59 VPWR.n58 0.122949
R118 VPWR.n60 VPWR.n59 0.122949
R119 VPWR.n60 VPWR.n0 0.122949
R120 VPB.t11 VPB.t5 814.652
R121 VPB.t16 VPB.t1 541.399
R122 VPB.t10 VPB.t7 531.183
R123 VPB.t13 VPB.t12 500.538
R124 VPB.t14 VPB.t13 500.538
R125 VPB.t5 VPB.t6 377.957
R126 VPB.t21 VPB.t20 349.866
R127 VPB.t9 VPB.t19 324.329
R128 VPB.t15 VPB.t8 321.774
R129 VPB.t7 VPB.t4 273.253
R130 VPB.t4 VPB.t21 265.591
R131 VPB.t12 VPB.t3 257.93
R132 VPB VPB.t17 257.93
R133 VPB.t20 VPB.t9 252.823
R134 VPB.t3 VPB.t2 229.839
R135 VPB.t0 VPB.t14 229.839
R136 VPB.t19 VPB.t11 229.839
R137 VPB.t1 VPB.t10 229.839
R138 VPB.t17 VPB.t18 229.839
R139 VPB.t8 VPB.t16 214.517
R140 VPB.t18 VPB.t15 214.517
R141 VPB.t6 VPB.t0 199.195
R142 a_1804_424.n8 a_1804_424.t3 666.024
R143 a_1804_424.n10 a_1804_424.n9 635.183
R144 a_1804_424.n9 a_1804_424.n0 304.604
R145 a_1804_424.n2 a_1804_424.t6 283.426
R146 a_1804_424.n6 a_1804_424.t7 198.388
R147 a_1804_424.n3 a_1804_424.t5 197.941
R148 a_1804_424.n3 a_1804_424.n1 165.189
R149 a_1804_424.n7 a_1804_424.n6 152
R150 a_1804_424.n5 a_1804_424.n1 152
R151 a_1804_424.n4 a_1804_424.n2 136.316
R152 a_1804_424.n10 a_1804_424.t1 133.679
R153 a_1804_424.n2 a_1804_424.t8 126.927
R154 a_1804_424.t0 a_1804_424.n10 112.572
R155 a_1804_424.n0 a_1804_424.t2 47.7237
R156 a_1804_424.n6 a_1804_424.n5 43.7018
R157 a_1804_424.n0 a_1804_424.t4 40.0005
R158 a_1804_424.n5 a_1804_424.n4 34.7045
R159 a_1804_424.n8 a_1804_424.n7 27.9916
R160 a_1804_424.n9 a_1804_424.n8 18.25
R161 a_1804_424.n7 a_1804_424.n1 13.1884
R162 a_1804_424.n4 a_1804_424.n3 8.99783
R163 VGND.n8 VGND.t2 270.193
R164 VGND.n54 VGND.t9 246.139
R165 VGND.n61 VGND.n60 199.488
R166 VGND.n21 VGND.n20 185
R167 VGND.n23 VGND.n22 185
R168 VGND.n16 VGND.t7 178.162
R169 VGND.n15 VGND.n14 125.314
R170 VGND.n52 VGND.n4 116.288
R171 VGND.n22 VGND.n21 102.858
R172 VGND.n60 VGND.t8 77.1434
R173 VGND.n60 VGND.t1 58.5719
R174 VGND.n22 VGND.t4 52.8576
R175 VGND.n14 VGND.t3 43.1255
R176 VGND.n21 VGND.t5 40.0005
R177 VGND.n19 VGND.n18 36.1417
R178 VGND.n29 VGND.n28 36.1417
R179 VGND.n30 VGND.n29 36.1417
R180 VGND.n30 VGND.n10 36.1417
R181 VGND.n34 VGND.n10 36.1417
R182 VGND.n41 VGND.n40 36.1417
R183 VGND.n42 VGND.n41 36.1417
R184 VGND.n46 VGND.n6 36.1417
R185 VGND.n47 VGND.n46 36.1417
R186 VGND.n48 VGND.n47 36.1417
R187 VGND.n48 VGND.n3 36.1417
R188 VGND.n58 VGND.n1 36.1417
R189 VGND.n59 VGND.n58 36.1417
R190 VGND.n4 VGND.t0 34.0546
R191 VGND.n24 VGND.n19 31.047
R192 VGND.n53 VGND.n52 30.1181
R193 VGND.n36 VGND.n8 29.3652
R194 VGND.n28 VGND.n12 29.3487
R195 VGND.n18 VGND.n15 26.7299
R196 VGND.n35 VGND.n34 25.6005
R197 VGND.n54 VGND.n53 24.8476
R198 VGND.n4 VGND.t10 22.7032
R199 VGND.n54 VGND.n1 22.5887
R200 VGND.n14 VGND.t6 21.8669
R201 VGND.n36 VGND.n35 21.8358
R202 VGND.n42 VGND.n6 20.7868
R203 VGND.n52 VGND.n3 17.3181
R204 VGND.n61 VGND.n59 9.78874
R205 VGND.n59 VGND.n0 9.3005
R206 VGND.n58 VGND.n57 9.3005
R207 VGND.n56 VGND.n1 9.3005
R208 VGND.n55 VGND.n54 9.3005
R209 VGND.n53 VGND.n2 9.3005
R210 VGND.n52 VGND.n51 9.3005
R211 VGND.n50 VGND.n3 9.3005
R212 VGND.n49 VGND.n48 9.3005
R213 VGND.n47 VGND.n5 9.3005
R214 VGND.n46 VGND.n45 9.3005
R215 VGND.n44 VGND.n6 9.3005
R216 VGND.n43 VGND.n42 9.3005
R217 VGND.n41 VGND.n7 9.3005
R218 VGND.n40 VGND.n39 9.3005
R219 VGND.n38 VGND.n8 9.3005
R220 VGND.n37 VGND.n36 9.3005
R221 VGND.n35 VGND.n9 9.3005
R222 VGND.n34 VGND.n33 9.3005
R223 VGND.n32 VGND.n10 9.3005
R224 VGND.n31 VGND.n30 9.3005
R225 VGND.n29 VGND.n11 9.3005
R226 VGND.n28 VGND.n27 9.3005
R227 VGND.n26 VGND.n12 9.3005
R228 VGND.n25 VGND.n24 9.3005
R229 VGND.n19 VGND.n13 9.3005
R230 VGND.n18 VGND.n17 9.3005
R231 VGND.n62 VGND.n61 7.43488
R232 VGND.n16 VGND.n15 6.87704
R233 VGND.n23 VGND.n20 6.72751
R234 VGND.n40 VGND.n8 5.27109
R235 VGND.n24 VGND.n23 1.40196
R236 VGND.n20 VGND.n12 0.841376
R237 VGND.n17 VGND.n16 0.561413
R238 VGND VGND.n62 0.160103
R239 VGND.n62 VGND.n0 0.1477
R240 VGND.n17 VGND.n13 0.122949
R241 VGND.n25 VGND.n13 0.122949
R242 VGND.n26 VGND.n25 0.122949
R243 VGND.n27 VGND.n26 0.122949
R244 VGND.n27 VGND.n11 0.122949
R245 VGND.n31 VGND.n11 0.122949
R246 VGND.n32 VGND.n31 0.122949
R247 VGND.n33 VGND.n32 0.122949
R248 VGND.n33 VGND.n9 0.122949
R249 VGND.n37 VGND.n9 0.122949
R250 VGND.n38 VGND.n37 0.122949
R251 VGND.n39 VGND.n38 0.122949
R252 VGND.n39 VGND.n7 0.122949
R253 VGND.n43 VGND.n7 0.122949
R254 VGND.n44 VGND.n43 0.122949
R255 VGND.n45 VGND.n44 0.122949
R256 VGND.n45 VGND.n5 0.122949
R257 VGND.n49 VGND.n5 0.122949
R258 VGND.n50 VGND.n49 0.122949
R259 VGND.n51 VGND.n50 0.122949
R260 VGND.n51 VGND.n2 0.122949
R261 VGND.n55 VGND.n2 0.122949
R262 VGND.n56 VGND.n55 0.122949
R263 VGND.n57 VGND.n56 0.122949
R264 VGND.n57 VGND.n0 0.122949
R265 a_2186_367.n1 a_2186_367.t1 809.619
R266 a_2186_367.n0 a_2186_367.t3 478.788
R267 a_2186_367.n1 a_2186_367.n0 251.606
R268 a_2186_367.t0 a_2186_367.n1 237.381
R269 a_2186_367.n0 a_2186_367.t2 126.927
R270 VNB.t4 VNB.t3 5058.27
R271 VNB.t5 VNB.t6 4619.42
R272 VNB.t3 VNB.t5 2448.29
R273 VNB.t9 VNB.t8 2286.61
R274 VNB.t15 VNB.t0 2286.61
R275 VNB.t17 VNB.t4 2263.52
R276 VNB.t10 VNB.t9 1928.61
R277 VNB.t14 VNB.t1 1443.57
R278 VNB.t2 VNB.t10 1316.54
R279 VNB.t8 VNB.t11 1212.6
R280 VNB.t6 VNB.t16 1154.86
R281 VNB.t0 VNB.t17 1154.86
R282 VNB VNB.t14 1143.31
R283 VNB.t13 VNB.t15 1085.56
R284 VNB.t11 VNB.t12 993.177
R285 VNB.t7 VNB.t13 993.177
R286 VNB.t16 VNB.t2 900.788
R287 VNB.t1 VNB.t7 900.788
R288 SET_B.n0 SET_B.t1 306.122
R289 SET_B.n2 SET_B.t0 294.173
R290 SET_B.n0 SET_B.t2 289.786
R291 SET_B.n2 SET_B.n1 226.424
R292 SET_B SET_B.n0 171.468
R293 SET_B SET_B.n2 168.484
R294 a_27_74.n1 a_27_74.t2 454.45
R295 a_27_74.t1 a_27_74.n1 357.098
R296 a_27_74.n0 a_27_74.t3 309.182
R297 a_27_74.n0 a_27_74.t0 237.412
R298 a_27_74.n1 a_27_74.n0 89.2852
R299 a_290_464.n1 a_290_464.t0 661.952
R300 a_290_464.n3 a_290_464.n2 616.232
R301 a_290_464.n2 a_290_464.n0 338.132
R302 a_290_464.n1 a_290_464.t1 337.925
R303 a_290_464.n2 a_290_464.n1 178.071
R304 a_290_464.t2 a_290_464.n3 73.8755
R305 a_290_464.n3 a_290_464.t4 73.8755
R306 a_290_464.n0 a_290_464.t5 40.0005
R307 a_290_464.n0 a_290_464.t3 40.0005
R308 SCE SCE.t0 475.632
R309 SCE.n1 SCE.t1 324.161
R310 SCE.n0 SCE.t3 194.407
R311 SCE.n0 SCE.t2 164.314
R312 SCE SCE.n1 72.034
R313 SCE.n1 SCE.n0 30.4479
R314 a_403_74.t0 a_403_74.t1 91.4291
R315 CLK.n0 CLK.t1 285.719
R316 CLK.n0 CLK.t0 178.34
R317 CLK CLK.n0 157.399
R318 a_608_74.n2 a_608_74.n1 1227.83
R319 a_608_74.n0 a_608_74.t6 931.063
R320 a_608_74.t1 a_608_74.n6 871.861
R321 a_608_74.n3 a_608_74.n2 750.313
R322 a_608_74.n3 a_608_74.t3 334.188
R323 a_608_74.n1 a_608_74.t5 299.447
R324 a_608_74.n4 a_608_74.t2 226.809
R325 a_608_74.n6 a_608_74.t0 213.397
R326 a_608_74.n4 a_608_74.t7 201.125
R327 a_608_74.n6 a_608_74.n5 200.679
R328 a_608_74.n1 a_608_74.n0 159.06
R329 a_608_74.n2 a_608_74.t4 155.847
R330 a_608_74.n5 a_608_74.n3 54.7732
R331 a_608_74.n5 a_608_74.n4 16.7975
R332 a_795_74.n7 a_795_74.n6 742.817
R333 a_795_74.n0 a_795_74.t0 477.616
R334 a_795_74.n5 a_795_74.n4 457.267
R335 a_795_74.n5 a_795_74.t2 417.332
R336 a_795_74.n6 a_795_74.n5 348.021
R337 a_795_74.n2 a_795_74.n1 303.904
R338 a_795_74.n4 a_795_74.t4 265.101
R339 a_795_74.n0 a_795_74.t3 220.113
R340 a_795_74.n6 a_795_74.n2 196.159
R341 a_795_74.n7 a_795_74.t1 190.561
R342 a_795_74.n4 a_795_74.n3 126.927
R343 a_795_74.n2 a_795_74.n0 120.793
R344 a_991_81.n9 a_991_81.n0 660.024
R345 a_991_81.t1 a_991_81.n9 362.55
R346 a_991_81.n7 a_991_81.t7 295.091
R347 a_991_81.n3 a_991_81.t4 254.121
R348 a_991_81.n5 a_991_81.n4 248.879
R349 a_991_81.n4 a_991_81.t6 240.976
R350 a_991_81.n2 a_991_81.n1 183.161
R351 a_991_81.n6 a_991_81.t3 170.892
R352 a_991_81.n8 a_991_81.n7 152
R353 a_991_81.n6 a_991_81.n5 152
R354 a_991_81.n2 a_991_81.t5 137.881
R355 a_991_81.n0 a_991_81.t0 131.252
R356 a_991_81.n9 a_991_81.n8 74.4162
R357 a_991_81.n0 a_991_81.t2 71.409
R358 a_991_81.n7 a_991_81.n6 49.6611
R359 a_991_81.n3 a_991_81.n2 33.5944
R360 a_991_81.n4 a_991_81.n3 19.7187
R361 a_991_81.n8 a_991_81.n5 13.1884
R362 a_2611_98.t1 a_2611_98.n2 255.618
R363 a_2611_98.n1 a_2611_98.t4 234.841
R364 a_2611_98.n0 a_2611_98.t5 234.841
R365 a_2611_98.n0 a_2611_98.t2 179.947
R366 a_2611_98.n2 a_2611_98.n0 178.207
R367 a_2611_98.n1 a_2611_98.t3 173.788
R368 a_2611_98.n2 a_2611_98.t0 151.95
R369 a_2611_98.n0 a_2611_98.n1 65.7278
R370 a_1185_55.n1 a_1185_55.n0 843.183
R371 a_1185_55.t1 a_1185_55.n3 430.459
R372 a_1185_55.n1 a_1185_55.t3 185.303
R373 a_1185_55.n3 a_1185_55.n1 171.913
R374 a_1185_55.n3 a_1185_55.n2 127.275
R375 a_1185_55.n0 a_1185_55.t2 91.4648
R376 a_1185_55.n0 a_1185_55.t0 70.3576
R377 a_1117_483.n0 a_1117_483.t1 127.963
R378 a_1117_483.n0 a_1117_483.t0 40.447
R379 a_1117_483.n1 a_1117_483.n0 37.1703
R380 a_2141_508.t0 a_2141_508.t1 112.572
R381 D.n0 D.t0 422.553
R382 D.n0 D.t1 176.466
R383 D D.n0 163.831
R384 a_239_74.t0 a_239_74.t1 68.5719
R385 Q Q.n0 210.031
R386 Q Q.n1 138.899
R387 Q.n0 Q.t3 26.3844
R388 Q.n0 Q.t2 26.3844
R389 Q.n1 Q.t0 22.7032
R390 Q.n1 Q.t1 22.7032
R391 a_1584_379.t0 a_1584_379.n0 729.187
R392 a_1584_379.n0 a_1584_379.t2 35.1791
R393 a_1584_379.n0 a_1584_379.t1 35.1791
R394 a_2141_74.t0 a_2141_74.t1 68.5719
R395 a_2219_74.t0 a_2219_74.t1 120.001
R396 a_1641_74.t0 a_1641_74.t1 446.587
R397 a_206_464.t0 a_206_464.t1 83.1099
C0 D SCE 0.181297f
C1 VPB SCD 0.100454f
C2 VPB VPWR 0.389279f
C3 D VPB 0.076159f
C4 VPB SCE 0.132438f
C5 VGND a_1143_81# 0.003473f
C6 VPWR a_1143_81# 4.35e-19
C7 Q VGND 0.192228f
C8 Q SET_B 1.99e-19
C9 VGND SET_B 0.205212f
C10 VGND CLK 0.040642f
C11 VPWR Q 0.224193f
C12 SCD VGND 0.035485f
C13 VPWR VGND 0.162721f
C14 D VGND 0.012595f
C15 SCE VGND 0.034432f
C16 CLK SET_B 1.26e-19
C17 VPB Q 0.011338f
C18 VPB VGND 0.026673f
C19 SCD SET_B 1.1e-19
C20 VPWR SET_B 0.127488f
C21 D SET_B 3.3e-20
C22 SCE SET_B 6.83e-20
C23 SCD CLK 0.028788f
C24 VPWR CLK 0.016255f
C25 VPB SET_B 0.180791f
C26 VPWR SCD 0.016929f
C27 D SCD 0.005333f
C28 VPB CLK 0.033702f
C29 D VPWR 0.012867f
C30 SCD SCE 0.054643f
C31 VPWR SCE 0.03256f
C32 Q VNB 0.052629f
C33 VGND VNB 1.74286f
C34 SET_B VNB 0.312746f
C35 CLK VNB 0.114926f
C36 VPWR VNB 1.34344f
C37 SCD VNB 0.16237f
C38 D VNB 0.115232f
C39 SCE VNB 0.323656f
C40 VPB VNB 3.40603f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfstp_1 VNB VPB VPWR SET_B VGND Q SCD CLK SCE D
X0 a_1958_48.t1 a_1764_74.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0882 ps=0.84 w=0.42 l=0.15
X1 Q.t1 a_2395_94.t2 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X2 a_402_74.t1 SCE.t0 a_289_464.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_1764_74.t1 SET_B.t0 VPWR.t8 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4 VPWR.t4 SCE.t1 a_27_464.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1856 ps=1.86 w=0.64 l=0.15
X5 a_800_74.t0 a_599_74.t2 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3076 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_800_74.t1 a_599_74.t3 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X7 VPWR.t6 CLK.t0 a_599_74.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8 VPWR.t12 a_1958_48.t2 a_1721_374.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 VPWR.t1 a_1764_74.t6 a_1958_48.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X10 a_1686_74.t0 a_998_81.t4 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.23495 ps=1.4 w=0.64 l=0.15
X11 VGND.t6 SET_B.t1 a_1988_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.1596 ps=1.18 w=0.42 l=0.15
X12 VGND.t2 a_1764_74.t7 a_2395_94.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.448 ps=2.68 w=0.64 l=0.15
X13 a_1988_74.t1 a_1958_48.t3 a_1910_74.t1 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1596 pd=1.18 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 a_289_464.t2 D.t0 a_238_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X15 a_1610_341.t0 a_998_81.t5 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.18815 ps=1.53 w=1 l=0.15
X16 a_1910_74.t0 a_599_74.t4 a_1764_74.t4 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.17735 ps=1.22 w=0.42 l=0.15
X17 VGND.t10 SCE.t2 a_27_464.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.1197 ps=1.41 w=0.42 l=0.15
X18 a_1128_457.t0 a_599_74.t5 a_998_81.t1 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.0735 ps=0.77 w=0.42 l=0.15
X19 VGND.t5 SCD.t0 a_402_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X20 a_1764_74.t0 a_800_74.t2 a_1686_74.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.17735 pd=1.22 as=0.0768 ps=0.88 w=0.64 l=0.15
X21 a_289_464.t1 D.t1 a_205_464.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1536 pd=1.12 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1610_341.t1 a_599_74.t6 a_1764_74.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.28 pd=2.56 as=0.16295 ps=1.41 w=1 l=0.15
X23 VGND.t3 SET_B.t2 a_1426_118.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.23495 pd=1.4 as=0.0504 ps=0.66 w=0.42 l=0.15
X24 a_998_81.t2 a_800_74.t3 a_289_464.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X25 a_205_464.t1 SCE.t3 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.096 ps=0.94 w=0.64 l=0.15
X26 VGND.t4 a_1198_55.t3 a_1150_81.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 VPWR.t5 SCD.t1 a_415_464.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2954 pd=2.4 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_1150_81.t0 a_800_74.t4 a_998_81.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1281 ps=1.03 w=0.42 l=0.15
X29 VGND.t11 CLK.t1 a_599_74.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X30 a_998_81.t0 a_599_74.t7 a_289_464.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1281 pd=1.03 as=0.1197 ps=1.41 w=0.42 l=0.15
X31 a_1426_118.t0 a_998_81.t6 a_1198_55.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X32 a_1198_55.t0 a_998_81.t7 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1649 ps=1.295 w=0.42 l=0.15
X33 VPWR.t9 SET_B.t3 a_1198_55.t2 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.18815 pd=1.53 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1764_74.t3 a_800_74.t5 a_1721_374.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.16295 pd=1.41 as=0.2584 ps=3.07 w=0.42 l=0.15
X35 VPWR.t0 a_1764_74.t8 a_2395_94.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2394 ps=2.25 w=0.84 l=0.15
X36 Q.t0 a_2395_94.t3 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1862 ps=1.475 w=1.12 l=0.15
X37 a_415_464.t0 a_27_464.t2 a_289_464.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1536 ps=1.12 w=0.64 l=0.15
X38 a_238_74.t0 a_27_464.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
R0 a_1764_74.n3 a_1764_74.t1 670.753
R1 a_1764_74.n6 a_1764_74.n5 599.429
R2 a_1764_74.n0 a_1764_74.t7 321.334
R3 a_1764_74.n2 a_1764_74.t5 303.356
R4 a_1764_74.n1 a_1764_74.n0 248.477
R5 a_1764_74.n1 a_1764_74.t6 215.561
R6 a_1764_74.n0 a_1764_74.t8 213.688
R7 a_1764_74.n5 a_1764_74.n3 155.482
R8 a_1764_74.n5 a_1764_74.n4 151.436
R9 a_1764_74.n6 a_1764_74.t3 119.608
R10 a_1764_74.n2 a_1764_74.n1 89.7775
R11 a_1764_74.n3 a_1764_74.n2 88.9365
R12 a_1764_74.n4 a_1764_74.t4 69.2416
R13 a_1764_74.n4 a_1764_74.t0 46.8755
R14 a_1764_74.t2 a_1764_74.n6 35.9765
R15 VGND.n30 VGND.t4 247.304
R16 VGND.n43 VGND.t5 246.333
R17 VGND.n16 VGND.n15 207.498
R18 VGND.n50 VGND.n49 206.721
R19 VGND.n14 VGND.n13 121.847
R20 VGND.n41 VGND.n4 115.659
R21 VGND.n15 VGND.t1 80.0005
R22 VGND.n9 VGND.n8 60.6604
R23 VGND.n49 VGND.t10 60.0005
R24 VGND.n49 VGND.t0 51.4291
R25 VGND.n13 VGND.t2 41.2505
R26 VGND.n15 VGND.t6 40.0005
R27 VGND.n18 VGND.n17 36.1417
R28 VGND.n18 VGND.n11 36.1417
R29 VGND.n22 VGND.n11 36.1417
R30 VGND.n23 VGND.n22 36.1417
R31 VGND.n24 VGND.n23 36.1417
R32 VGND.n29 VGND.n28 36.1417
R33 VGND.n31 VGND.n29 36.1417
R34 VGND.n35 VGND.n6 36.1417
R35 VGND.n36 VGND.n35 36.1417
R36 VGND.n37 VGND.n36 36.1417
R37 VGND.n37 VGND.n3 36.1417
R38 VGND.n47 VGND.n1 36.1417
R39 VGND.n48 VGND.n47 36.1417
R40 VGND.n4 VGND.t7 34.0546
R41 VGND.n4 VGND.t11 34.0546
R42 VGND.n43 VGND.n42 31.2476
R43 VGND.n13 VGND.t9 30.2643
R44 VGND.n8 VGND.t3 29.7074
R45 VGND.n42 VGND.n41 26.7299
R46 VGND.n41 VGND.n3 20.7064
R47 VGND.n16 VGND.n14 17.0486
R48 VGND.n43 VGND.n1 16.1887
R49 VGND.n50 VGND.n48 13.177
R50 VGND.n8 VGND.t8 9.50606
R51 VGND.n48 VGND.n0 9.3005
R52 VGND.n47 VGND.n46 9.3005
R53 VGND.n45 VGND.n1 9.3005
R54 VGND.n44 VGND.n43 9.3005
R55 VGND.n42 VGND.n2 9.3005
R56 VGND.n41 VGND.n40 9.3005
R57 VGND.n17 VGND.n12 9.3005
R58 VGND.n19 VGND.n18 9.3005
R59 VGND.n20 VGND.n11 9.3005
R60 VGND.n22 VGND.n21 9.3005
R61 VGND.n23 VGND.n10 9.3005
R62 VGND.n25 VGND.n24 9.3005
R63 VGND.n26 VGND.n9 9.3005
R64 VGND.n28 VGND.n27 9.3005
R65 VGND.n29 VGND.n7 9.3005
R66 VGND.n32 VGND.n31 9.3005
R67 VGND.n33 VGND.n6 9.3005
R68 VGND.n35 VGND.n34 9.3005
R69 VGND.n36 VGND.n5 9.3005
R70 VGND.n38 VGND.n37 9.3005
R71 VGND.n39 VGND.n3 9.3005
R72 VGND.n30 VGND.n6 8.65932
R73 VGND.n51 VGND.n50 7.64704
R74 VGND.n24 VGND.n9 7.15344
R75 VGND.n31 VGND.n30 2.63579
R76 VGND.n17 VGND.n16 1.88285
R77 VGND.n28 VGND.n9 1.12991
R78 VGND.n14 VGND.n12 0.163003
R79 VGND VGND.n51 0.162897
R80 VGND.n51 VGND.n0 0.144943
R81 VGND.n19 VGND.n12 0.122949
R82 VGND.n20 VGND.n19 0.122949
R83 VGND.n21 VGND.n20 0.122949
R84 VGND.n21 VGND.n10 0.122949
R85 VGND.n25 VGND.n10 0.122949
R86 VGND.n26 VGND.n25 0.122949
R87 VGND.n27 VGND.n26 0.122949
R88 VGND.n27 VGND.n7 0.122949
R89 VGND.n32 VGND.n7 0.122949
R90 VGND.n33 VGND.n32 0.122949
R91 VGND.n34 VGND.n33 0.122949
R92 VGND.n34 VGND.n5 0.122949
R93 VGND.n38 VGND.n5 0.122949
R94 VGND.n39 VGND.n38 0.122949
R95 VGND.n40 VGND.n39 0.122949
R96 VGND.n40 VGND.n2 0.122949
R97 VGND.n44 VGND.n2 0.122949
R98 VGND.n45 VGND.n44 0.122949
R99 VGND.n46 VGND.n45 0.122949
R100 VGND.n46 VGND.n0 0.122949
R101 a_1958_48.n1 a_1958_48.t0 758.232
R102 a_1958_48.n0 a_1958_48.t2 465.521
R103 a_1958_48.t1 a_1958_48.n1 242.579
R104 a_1958_48.n1 a_1958_48.n0 129.361
R105 a_1958_48.n0 a_1958_48.t3 118.513
R106 VNB.n1 VNB 19667.2
R107 VNB.t2 VNB.t1 3245.14
R108 VNB VNB.n1 2656.6
R109 VNB.t18 VNB.t6 2379
R110 VNB.t16 VNB.t4 2286.61
R111 VNB.t11 VNB.t8 2286.61
R112 VNB.t17 VNB.t7 2101.84
R113 VNB.t14 VNB.t11 1755.38
R114 VNB.t9 VNB.t19 1686.09
R115 VNB.t1 VNB.t13 1339.63
R116 VNB.t15 VNB 1328.08
R117 VNB.t7 VNB.t2 1316.54
R118 VNB.t8 VNB.t18 1316.54
R119 VNB.t0 VNB.t15 1247.24
R120 VNB.t12 VNB.t5 993.177
R121 VNB.t19 VNB.t17 900.788
R122 VNB.t3 VNB.t16 900.788
R123 VNB.t4 VNB.t14 900.788
R124 VNB.t6 VNB.t12 900.788
R125 VNB.t5 VNB.t0 900.788
R126 VNB.n1 VNB.t9 531.235
R127 VNB.n0 VNB.t10 137.894
R128 VNB.n0 VNB.t3 15.3466
R129 VNB.n1 VNB.n0 6.97627
R130 a_2395_94.t0 a_2395_94.n1 432.712
R131 a_2395_94.n0 a_2395_94.t3 279.293
R132 a_2395_94.n1 a_2395_94.n0 175.856
R133 a_2395_94.n0 a_2395_94.t2 171.913
R134 a_2395_94.n1 a_2395_94.t1 158.899
R135 Q.n3 Q 591.4
R136 Q.n3 Q.n0 585
R137 Q.n4 Q.n3 585
R138 Q.t1 Q.n1 279.738
R139 Q.n2 Q.t1 246.054
R140 Q.n3 Q.t0 26.3844
R141 Q Q.n4 17.1525
R142 Q Q.n0 14.8485
R143 Q Q.n2 13.0477
R144 Q.n1 Q 9.56372
R145 Q Q.n0 4.0965
R146 Q.n4 Q 1.7925
R147 Q.n2 Q 1.32464
R148 Q.n1 Q 1.32464
R149 SCE.n3 SCE.t0 472.548
R150 SCE.n0 SCE.t3 283.844
R151 SCE.n2 SCE.t2 249.034
R152 SCE.n0 SCE.t1 216.876
R153 SCE SCE.n1 158.4
R154 SCE.n3 SCE.n2 154.499
R155 SCE.n2 SCE.n1 49.6611
R156 SCE.n1 SCE.n0 13.146
R157 SCE SCE.n3 1.71757
R158 a_289_464.n1 a_289_464.t4 663.539
R159 a_289_464.n3 a_289_464.n2 616.489
R160 a_289_464.n1 a_289_464.t5 348.86
R161 a_289_464.n2 a_289_464.n0 338.144
R162 a_289_464.n2 a_289_464.n1 169.774
R163 a_289_464.t0 a_289_464.n3 73.8755
R164 a_289_464.n3 a_289_464.t1 73.8755
R165 a_289_464.n0 a_289_464.t3 40.0005
R166 a_289_464.n0 a_289_464.t2 40.0005
R167 a_402_74.t0 a_402_74.t1 68.5719
R168 SET_B.n0 SET_B.t1 302.38
R169 SET_B.n0 SET_B.t0 248.524
R170 SET_B.n1 SET_B.t2 242.929
R171 SET_B.n1 SET_B.t3 213.206
R172 SET_B SET_B.n1 170.553
R173 SET_B SET_B.n0 77.7595
R174 VPWR.n8 VPWR.t11 872.244
R175 VPWR.n50 VPWR.t5 787.665
R176 VPWR.n19 VPWR.t1 684.029
R177 VPWR.n11 VPWR.n10 626.729
R178 VPWR.n25 VPWR.n15 620.765
R179 VPWR.n56 VPWR.n1 606.333
R180 VPWR.n48 VPWR.n5 606.333
R181 VPWR.n18 VPWR.n17 327.507
R182 VPWR.n10 VPWR.t9 178.238
R183 VPWR.n15 VPWR.t8 70.3576
R184 VPWR.n15 VPWR.t12 70.3576
R185 VPWR.n17 VPWR.t0 46.9053
R186 VPWR.n1 VPWR.t3 46.1724
R187 VPWR.n1 VPWR.t4 46.1724
R188 VPWR.n54 VPWR.n2 36.1417
R189 VPWR.n55 VPWR.n54 36.1417
R190 VPWR.n42 VPWR.n41 36.1417
R191 VPWR.n43 VPWR.n42 36.1417
R192 VPWR.n43 VPWR.n6 36.1417
R193 VPWR.n47 VPWR.n6 36.1417
R194 VPWR.n37 VPWR.n36 36.1417
R195 VPWR.n38 VPWR.n37 36.1417
R196 VPWR.n20 VPWR.n16 36.1417
R197 VPWR.n24 VPWR.n16 36.1417
R198 VPWR.n27 VPWR.n26 36.1417
R199 VPWR.n27 VPWR.n13 36.1417
R200 VPWR.n31 VPWR.n13 36.1417
R201 VPWR.n32 VPWR.n31 36.1417
R202 VPWR.n33 VPWR.n32 36.1417
R203 VPWR.n49 VPWR.n48 34.2593
R204 VPWR.n10 VPWR.t7 33.6312
R205 VPWR.n17 VPWR.t10 30.9824
R206 VPWR.n50 VPWR.n2 30.4946
R207 VPWR.n26 VPWR.n25 29.7417
R208 VPWR.n5 VPWR.t2 26.3844
R209 VPWR.n5 VPWR.t6 26.3844
R210 VPWR.n56 VPWR.n55 23.3417
R211 VPWR.n20 VPWR.n19 23.3417
R212 VPWR.n50 VPWR.n49 16.9417
R213 VPWR.n41 VPWR.n8 16.9417
R214 VPWR.n36 VPWR.n11 16.9417
R215 VPWR.n48 VPWR.n47 13.177
R216 VPWR.n21 VPWR.n20 9.3005
R217 VPWR.n22 VPWR.n16 9.3005
R218 VPWR.n24 VPWR.n23 9.3005
R219 VPWR.n26 VPWR.n14 9.3005
R220 VPWR.n28 VPWR.n27 9.3005
R221 VPWR.n29 VPWR.n13 9.3005
R222 VPWR.n31 VPWR.n30 9.3005
R223 VPWR.n32 VPWR.n12 9.3005
R224 VPWR.n34 VPWR.n33 9.3005
R225 VPWR.n36 VPWR.n35 9.3005
R226 VPWR.n37 VPWR.n9 9.3005
R227 VPWR.n39 VPWR.n38 9.3005
R228 VPWR.n41 VPWR.n40 9.3005
R229 VPWR.n42 VPWR.n7 9.3005
R230 VPWR.n44 VPWR.n43 9.3005
R231 VPWR.n45 VPWR.n6 9.3005
R232 VPWR.n47 VPWR.n46 9.3005
R233 VPWR.n48 VPWR.n4 9.3005
R234 VPWR.n49 VPWR.n3 9.3005
R235 VPWR.n51 VPWR.n50 9.3005
R236 VPWR.n52 VPWR.n2 9.3005
R237 VPWR.n54 VPWR.n53 9.3005
R238 VPWR.n55 VPWR.n0 9.3005
R239 VPWR.n57 VPWR.n56 7.25439
R240 VPWR.n19 VPWR.n18 7.08122
R241 VPWR.n25 VPWR.n24 6.4005
R242 VPWR.n21 VPWR.n18 0.490447
R243 VPWR.n38 VPWR.n8 0.376971
R244 VPWR.n33 VPWR.n11 0.376971
R245 VPWR VPWR.n57 0.157727
R246 VPWR.n57 VPWR.n0 0.150046
R247 VPWR.n22 VPWR.n21 0.122949
R248 VPWR.n23 VPWR.n22 0.122949
R249 VPWR.n23 VPWR.n14 0.122949
R250 VPWR.n28 VPWR.n14 0.122949
R251 VPWR.n29 VPWR.n28 0.122949
R252 VPWR.n30 VPWR.n29 0.122949
R253 VPWR.n30 VPWR.n12 0.122949
R254 VPWR.n34 VPWR.n12 0.122949
R255 VPWR.n35 VPWR.n34 0.122949
R256 VPWR.n35 VPWR.n9 0.122949
R257 VPWR.n39 VPWR.n9 0.122949
R258 VPWR.n40 VPWR.n39 0.122949
R259 VPWR.n40 VPWR.n7 0.122949
R260 VPWR.n44 VPWR.n7 0.122949
R261 VPWR.n45 VPWR.n44 0.122949
R262 VPWR.n46 VPWR.n45 0.122949
R263 VPWR.n46 VPWR.n4 0.122949
R264 VPWR.n4 VPWR.n3 0.122949
R265 VPWR.n51 VPWR.n3 0.122949
R266 VPWR.n52 VPWR.n51 0.122949
R267 VPWR.n53 VPWR.n52 0.122949
R268 VPWR.n53 VPWR.n0 0.122949
R269 VPB.t18 VPB.t16 638.442
R270 VPB.t4 VPB.t8 561.828
R271 VPB.t7 VPB.t9 559.274
R272 VPB.t2 VPB.t1 505.646
R273 VPB.t13 VPB.t2 505.646
R274 VPB.t11 VPB.t17 503.091
R275 VPB.t10 VPB.t15 495.43
R276 VPB.t12 VPB.t10 347.312
R277 VPB.t3 VPB.t0 321.774
R278 VPB.t15 VPB.t11 286.022
R279 VPB.t1 VPB.t14 257.93
R280 VPB.t8 VPB.t18 255.376
R281 VPB VPB.t6 255.376
R282 VPB.t16 VPB.t12 245.161
R283 VPB.t17 VPB.t13 229.839
R284 VPB.t9 VPB.t4 229.839
R285 VPB.t6 VPB.t5 229.839
R286 VPB.t0 VPB.t7 214.517
R287 VPB.t5 VPB.t3 214.517
R288 a_27_464.n1 a_27_464.t2 454.039
R289 a_27_464.t0 a_27_464.n1 358.76
R290 a_27_464.n0 a_27_464.t3 325.663
R291 a_27_464.n0 a_27_464.t1 237.946
R292 a_27_464.n1 a_27_464.n0 96.9605
R293 a_599_74.n0 a_599_74.t6 1447.87
R294 a_599_74.t0 a_599_74.n4 862.136
R295 a_599_74.n1 a_599_74.n0 729.025
R296 a_599_74.t6 a_599_74.t4 546.638
R297 a_599_74.n1 a_599_74.t7 335.793
R298 a_599_74.n2 a_599_74.t2 226.809
R299 a_599_74.n2 a_599_74.t3 203.141
R300 a_599_74.n4 a_599_74.n3 199.143
R301 a_599_74.n4 a_599_74.t1 197.165
R302 a_599_74.n0 a_599_74.t5 190.659
R303 a_599_74.n3 a_599_74.n1 59.155
R304 a_599_74.n3 a_599_74.n2 12.4157
R305 a_800_74.n4 a_800_74.n3 740.482
R306 a_800_74.n3 a_800_74.n2 495.719
R307 a_800_74.n0 a_800_74.t1 379.26
R308 a_800_74.n1 a_800_74.t4 330.098
R309 a_800_74.n2 a_800_74.t5 205.752
R310 a_800_74.n4 a_800_74.t0 190.561
R311 a_800_74.n3 a_800_74.n1 188.518
R312 a_800_74.n0 a_800_74.t3 160.042
R313 a_800_74.n2 a_800_74.t2 159.963
R314 a_800_74.n1 a_800_74.n0 130.34
R315 CLK.n0 CLK.t0 285.719
R316 CLK.n0 CLK.t1 178.34
R317 CLK CLK.n0 157.601
R318 a_1721_374.t0 a_1721_374.t1 2149.81
R319 a_998_81.n4 a_998_81.n0 664.322
R320 a_998_81.n1 a_998_81.t6 274.74
R321 a_998_81.n2 a_998_81.t5 251.27
R322 a_998_81.n5 a_998_81.n4 223.144
R323 a_998_81.n1 a_998_81.t7 216.097
R324 a_998_81.n2 a_998_81.t4 170.507
R325 a_998_81.n3 a_998_81.n1 158.738
R326 a_998_81.n3 a_998_81.n2 152.12
R327 a_998_81.t0 a_998_81.n5 134.286
R328 a_998_81.n0 a_998_81.t2 93.81
R329 a_998_81.n4 a_998_81.n3 70.9709
R330 a_998_81.n0 a_998_81.t1 70.3576
R331 a_998_81.n5 a_998_81.t3 40.0005
R332 a_1686_74.t0 a_1686_74.t1 45.0005
R333 a_1988_74.t0 a_1988_74.t1 217.143
R334 a_1910_74.t0 a_1910_74.t1 68.5719
R335 D.n0 D.t0 422.553
R336 D.n0 D.t1 176.466
R337 D D.n0 163.637
R338 a_238_74.t0 a_238_74.t1 68.5719
R339 a_1610_341.t0 a_1610_341.t1 793.298
R340 SCD.n2 SCD.t0 175.952
R341 SCD.n0 SCD.t1 169.179
R342 SCD SCD.n0 153.792
R343 SCD.n4 SCD.n3 152
R344 SCD.n2 SCD.n1 152
R345 SCD.n3 SCD.n0 33.7902
R346 SCD.n3 SCD.n2 33.7902
R347 SCD SCD.n4 15.6165
R348 SCD.n1 SCD 14.0805
R349 SCD.n1 SCD 4.8645
R350 SCD.n4 SCD 3.3285
R351 a_205_464.t0 a_205_464.t1 83.1099
R352 a_1426_118.t0 a_1426_118.t1 68.5719
R353 a_1198_55.n2 a_1198_55.n1 821.24
R354 a_1198_55.t1 a_1198_55.n3 404.541
R355 a_1198_55.n3 a_1198_55.n2 216.81
R356 a_1198_55.n3 a_1198_55.t3 157.745
R357 a_1198_55.n2 a_1198_55.n0 136.744
R358 a_1198_55.n1 a_1198_55.t0 84.4291
R359 a_1198_55.n1 a_1198_55.t2 70.3576
R360 a_1150_81.t0 a_1150_81.t1 68.5719
R361 a_415_464.t0 a_415_464.t1 83.1099
C0 VGND CLK 0.044973f
C1 Q VGND 0.107057f
C2 SCD VGND 0.037448f
C3 SET_B VGND 0.138784f
C4 SCD CLK 0.028626f
C5 SCE VGND 0.035791f
C6 VGND VPWR 0.158341f
C7 SET_B CLK 8.75e-20
C8 VPWR CLK 0.01542f
C9 Q SET_B 1.36e-19
C10 SCD SET_B 1.12e-19
C11 D VGND 0.012897f
C12 SCE SCD 0.057112f
C13 Q VPWR 0.108466f
C14 SCD VPWR 0.017175f
C15 SCE SET_B 8.56e-20
C16 VPB VGND 0.027662f
C17 SET_B VPWR 0.125005f
C18 VPB CLK 0.03383f
C19 SCE VPWR 0.032723f
C20 D SCD 0.004923f
C21 D SET_B 2.43e-20
C22 VPB Q 0.013767f
C23 VPB SCD 0.104047f
C24 SCE D 0.182694f
C25 D VPWR 0.012836f
C26 VPB SET_B 0.195007f
C27 VPB SCE 0.13725f
C28 VPB VPWR 0.363031f
C29 VPB D 0.074965f
C30 Q VNB 0.116881f
C31 VGND VNB 1.63993f
C32 SET_B VNB 0.253536f
C33 CLK VNB 0.115926f
C34 VPWR VNB 1.23671f
C35 SCD VNB 0.174554f
C36 D VNB 0.114174f
C37 SCE VNB 0.330168f
C38 VPB VNB 3.20893f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfsbp_2 VNB VPB SET_B VPWR VGND SCD Q_N Q CLK D SCE
X0 a_1789_424.t2 a_1069_81.t4 VPWR.t15 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X1 VPWR.t12 a_2067_74.t6 a_2513_258.t0 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.1841 pd=1.505 as=0.1239 ps=1.43 w=0.42 l=0.15
X2 a_2513_258.t1 a_2067_74.t7 VGND.t14 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0756 ps=0.78 w=0.42 l=0.15
X3 VPWR.t11 SCE.t0 a_27_74.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.1888 ps=1.87 w=0.64 l=0.15
X4 VGND.t6 SCD.t0 a_495_74.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5 VPWR.t14 a_1069_81.t5 a_1789_424.t1 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2898 ps=2.37 w=0.84 l=0.15
X6 a_2067_74.t2 a_871_74.t2 a_2277_455.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.126 ps=1.44 w=0.42 l=0.15
X7 a_2067_74.t3 SET_B.t0 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X8 a_1252_376# a_1069_81.t6 VPWR.t13 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.084 pd=0.82 as=0.19635 ps=1.355 w=0.42 l=0.15
X9 VPWR.t5 a_2513_258.t2 a_2277_455.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X10 a_1069_81.t0 a_871_74.t3 a_304_464.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X11 Q_N.t1 a_2067_74.t8 VGND.t13 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.2479 ps=2.15 w=0.74 l=0.15
X12 a_304_464.t0 D.t0 a_229_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1659 pd=1.21 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 VGND.t1 a_1252_376# a_1274_81.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.58 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 VGND.t4 SCE.t1 a_27_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.08925 pd=0.845 as=0.1197 ps=1.41 w=0.42 l=0.15
X15 a_304_464.t1 D.t1 a_220_464.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 VPWR.t8 SCD.t1 a_418_464.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.91 as=0.0864 ps=0.91 w=0.64 l=0.15
X17 a_871_74.t1 a_619_368.t2 VGND.t9 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 VGND.t7 SET_B.t1 a_2579_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X19 a_220_464.t0 SCE.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X20 VPWR.t7 a_3177_368.t2 Q.t2 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_418_464.t1 a_27_74.t2 a_304_464.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1344 ps=1.06 w=0.64 l=0.15
X22 VPWR.t0 CLK.t0 a_619_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.3304 ps=2.83 w=1.12 l=0.15
X23 Q_N.t2 a_2067_74.t9 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1841 ps=1.505 w=1.12 l=0.15
X24 VGND.t0 SET_B.t2 a_1567_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.189 pd=1.74 as=0.0504 ps=0.66 w=0.42 l=0.15
X25 Q.t1 a_3177_368.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.14705 ps=1.155 w=0.74 l=0.15
X26 VPWR.t1 SET_B.t3 a_1252_376# VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2457 pd=2.01 as=0.084 ps=0.82 w=0.42 l=0.15
X27 VGND.t11 a_2067_74.t10 a_3177_368.t0 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.14705 pd=1.155 as=0.1824 ps=1.85 w=0.64 l=0.15
X28 a_495_74.t1 SCE.t3 a_304_464.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1659 ps=1.21 w=0.42 l=0.15
X29 VGND.t5 CLK.t1 a_619_368.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X30 a_1794_74# a_1069_81.t7 VGND.t8 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.096 ps=0.94 w=0.64 l=0.15
X31 a_1789_424.t3 a_619_368.t3 a_2067_74.t5 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X32 VGND.t10 a_3177_368.t4 Q.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 a_2067_74.t1 a_619_368.t4 a_1789_424.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X34 VPWR.t2 a_1252_376# a_1201_463.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.19635 pd=1.355 as=0.0567 ps=0.69 w=0.42 l=0.15
X35 a_229_74.t1 a_27_74.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.08925 ps=0.845 w=0.42 l=0.15
X36 a_1794_74# a_871_74.t4 a_2067_74.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.112 ps=0.99 w=0.64 l=0.15
X37 a_1201_463.t1 a_619_368.t5 a_1069_81.t2 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0735 ps=0.77 w=0.42 l=0.15
X38 a_1274_81.t1 a_871_74.t5 a_1069_81.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.18375 ps=1.295 w=0.42 l=0.15
X39 a_2579_74.t1 a_2513_258.t3 a_2501_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X40 a_871_74.t0 a_619_368.t6 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3696 pd=2.9 as=0.3808 ps=1.8 w=1.12 l=0.15
X41 a_1069_81.t3 a_619_368.t7 a_304_464.t5 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.18375 pd=1.295 as=0.1197 ps=1.41 w=0.42 l=0.15
X42 VPWR.t3 a_2067_74.t11 a_3177_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2177 pd=1.52 as=0.295 ps=2.59 w=1 l=0.15
X43 a_2501_74.t0 a_619_368.t8 a_2067_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.3759 ps=2.63 w=0.42 l=0.15
X44 VGND.t12 a_2067_74.t12 Q_N.t0 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.2442 pd=2.14 as=0.111 ps=1.04 w=0.74 l=0.15
R0 a_1069_81.n8 a_1069_81.n7 711.981
R1 a_1069_81.n6 a_1069_81.n3 373.524
R2 a_1069_81.n0 a_1069_81.t4 355.877
R3 a_1069_81.n1 a_1069_81.t5 355.877
R4 a_1069_81.n5 a_1069_81.t6 303.283
R5 a_1069_81.n5 a_1069_81.n4 230.923
R6 a_1069_81.n0 a_1069_81.t7 195.21
R7 a_1069_81.n9 a_1069_81.n8 185
R8 a_1069_81.n9 a_1069_81.t3 182.857
R9 a_1069_81.n6 a_1069_81.n5 152
R10 a_1069_81.n3 a_1069_81.n2 147.011
R11 a_1069_81.n8 a_1069_81.n6 132.911
R12 a_1069_81.n7 a_1069_81.t0 93.81
R13 a_1069_81.n1 a_1069_81.n0 86.7605
R14 a_1069_81.n7 a_1069_81.t2 70.3576
R15 a_1069_81.t1 a_1069_81.n9 67.1434
R16 a_1069_81.n3 a_1069_81.n1 40.1672
R17 VPWR.n50 VPWR.t1 820.861
R18 VPWR.n70 VPWR.t8 713.279
R19 VPWR.n17 VPWR.n16 622.271
R20 VPWR.n12 VPWR.n11 615.976
R21 VPWR.n55 VPWR.n8 601.473
R22 VPWR.n62 VPWR.n4 585
R23 VPWR.n64 VPWR.n63 585
R24 VPWR.n76 VPWR.n1 315.736
R25 VPWR.n8 VPWR.t13 311.918
R26 VPWR.n23 VPWR.t3 282.038
R27 VPWR.n24 VPWR.t7 266.248
R28 VPWR.n20 VPWR.n19 243.916
R29 VPWR.n8 VPWR.t2 126.644
R30 VPWR.n19 VPWR.t12 110.227
R31 VPWR.n16 VPWR.t10 70.3576
R32 VPWR.n16 VPWR.t5 70.3576
R33 VPWR.n63 VPWR.n62 64.2014
R34 VPWR.n1 VPWR.t11 61.563
R35 VPWR.n1 VPWR.t4 46.1724
R36 VPWR.n74 VPWR.n2 36.1417
R37 VPWR.n75 VPWR.n74 36.1417
R38 VPWR.n56 VPWR.n6 36.1417
R39 VPWR.n60 VPWR.n6 36.1417
R40 VPWR.n61 VPWR.n60 36.1417
R41 VPWR.n54 VPWR.n9 36.1417
R42 VPWR.n49 VPWR.n48 36.1417
R43 VPWR.n29 VPWR.n28 36.1417
R44 VPWR.n33 VPWR.n32 36.1417
R45 VPWR.n34 VPWR.n33 36.1417
R46 VPWR.n38 VPWR.n37 36.1417
R47 VPWR.n39 VPWR.n38 36.1417
R48 VPWR.n39 VPWR.n14 36.1417
R49 VPWR.n43 VPWR.n14 36.1417
R50 VPWR.n44 VPWR.n43 36.1417
R51 VPWR.n45 VPWR.n44 36.1417
R52 VPWR.n11 VPWR.t15 35.1791
R53 VPWR.n11 VPWR.t14 35.1791
R54 VPWR.n55 VPWR.n54 34.2593
R55 VPWR.n27 VPWR.n26 33.5064
R56 VPWR.n69 VPWR.n68 31.7495
R57 VPWR.n50 VPWR.n9 31.2476
R58 VPWR.n56 VPWR.n55 30.8711
R59 VPWR.n32 VPWR.n20 30.8711
R60 VPWR.n63 VPWR.t9 29.0228
R61 VPWR.n65 VPWR.n61 27.943
R62 VPWR.n62 VPWR.t0 26.3844
R63 VPWR.n19 VPWR.t6 25.9146
R64 VPWR.n70 VPWR.n2 25.224
R65 VPWR.n26 VPWR.n23 25.224
R66 VPWR.n37 VPWR.n17 22.9652
R67 VPWR.n70 VPWR.n69 20.7064
R68 VPWR.n76 VPWR.n75 17.6946
R69 VPWR.n50 VPWR.n49 16.1887
R70 VPWR.n28 VPWR.n27 13.9299
R71 VPWR.n34 VPWR.n17 13.177
R72 VPWR.n45 VPWR.n12 12.424
R73 VPWR.n26 VPWR.n25 9.3005
R74 VPWR.n27 VPWR.n22 9.3005
R75 VPWR.n28 VPWR.n21 9.3005
R76 VPWR.n30 VPWR.n29 9.3005
R77 VPWR.n32 VPWR.n31 9.3005
R78 VPWR.n33 VPWR.n18 9.3005
R79 VPWR.n35 VPWR.n34 9.3005
R80 VPWR.n37 VPWR.n36 9.3005
R81 VPWR.n38 VPWR.n15 9.3005
R82 VPWR.n40 VPWR.n39 9.3005
R83 VPWR.n41 VPWR.n14 9.3005
R84 VPWR.n43 VPWR.n42 9.3005
R85 VPWR.n44 VPWR.n13 9.3005
R86 VPWR.n46 VPWR.n45 9.3005
R87 VPWR.n48 VPWR.n47 9.3005
R88 VPWR.n49 VPWR.n10 9.3005
R89 VPWR.n51 VPWR.n50 9.3005
R90 VPWR.n52 VPWR.n9 9.3005
R91 VPWR.n54 VPWR.n53 9.3005
R92 VPWR.n57 VPWR.n56 9.3005
R93 VPWR.n58 VPWR.n6 9.3005
R94 VPWR.n60 VPWR.n59 9.3005
R95 VPWR.n61 VPWR.n5 9.3005
R96 VPWR.n66 VPWR.n65 9.3005
R97 VPWR.n68 VPWR.n67 9.3005
R98 VPWR.n69 VPWR.n3 9.3005
R99 VPWR.n71 VPWR.n70 9.3005
R100 VPWR.n72 VPWR.n2 9.3005
R101 VPWR.n74 VPWR.n73 9.3005
R102 VPWR.n75 VPWR.n0 9.3005
R103 VPWR.n77 VPWR.n76 7.49287
R104 VPWR.n24 VPWR.n23 6.95806
R105 VPWR.n64 VPWR.n4 6.10769
R106 VPWR.n29 VPWR.n20 5.27109
R107 VPWR.n48 VPWR.n12 4.89462
R108 VPWR.n55 VPWR.n7 4.62059
R109 VPWR.n68 VPWR.n4 1.50638
R110 VPWR.n25 VPWR.n24 0.546775
R111 VPWR.n65 VPWR.n64 0.418801
R112 VPWR.n53 VPWR.n7 0.184273
R113 VPWR.n57 VPWR.n7 0.184273
R114 VPWR VPWR.n77 0.160867
R115 VPWR.n77 VPWR.n0 0.146947
R116 VPWR.n25 VPWR.n22 0.122949
R117 VPWR.n22 VPWR.n21 0.122949
R118 VPWR.n30 VPWR.n21 0.122949
R119 VPWR.n31 VPWR.n30 0.122949
R120 VPWR.n31 VPWR.n18 0.122949
R121 VPWR.n35 VPWR.n18 0.122949
R122 VPWR.n36 VPWR.n35 0.122949
R123 VPWR.n36 VPWR.n15 0.122949
R124 VPWR.n40 VPWR.n15 0.122949
R125 VPWR.n41 VPWR.n40 0.122949
R126 VPWR.n42 VPWR.n41 0.122949
R127 VPWR.n42 VPWR.n13 0.122949
R128 VPWR.n46 VPWR.n13 0.122949
R129 VPWR.n47 VPWR.n46 0.122949
R130 VPWR.n47 VPWR.n10 0.122949
R131 VPWR.n51 VPWR.n10 0.122949
R132 VPWR.n52 VPWR.n51 0.122949
R133 VPWR.n53 VPWR.n52 0.122949
R134 VPWR.n58 VPWR.n57 0.122949
R135 VPWR.n59 VPWR.n58 0.122949
R136 VPWR.n59 VPWR.n5 0.122949
R137 VPWR.n66 VPWR.n5 0.122949
R138 VPWR.n67 VPWR.n66 0.122949
R139 VPWR.n67 VPWR.n3 0.122949
R140 VPWR.n71 VPWR.n3 0.122949
R141 VPWR.n72 VPWR.n71 0.122949
R142 VPWR.n73 VPWR.n72 0.122949
R143 VPWR.n73 VPWR.n0 0.122949
R144 a_1789_424.n0 a_1789_424.t1 437.637
R145 a_1789_424.n0 a_1789_424.t3 409.474
R146 a_1789_424.n1 a_1789_424.n0 285.627
R147 a_1789_424.n1 a_1789_424.t0 35.1791
R148 a_1789_424.t2 a_1789_424.n1 35.1791
R149 VPB.t11 VPB.t4 745.699
R150 VPB.t2 VPB.t20 704.84
R151 VPB.t14 VPB.t9 579.705
R152 VPB.t3 VPB.t19 554.168
R153 VPB.t22 VPB.t8 533.737
R154 VPB.t8 VPB.t10 531.183
R155 VPB.t13 VPB.t0 526.076
R156 VPB.t15 VPB.t18 515.861
R157 VPB.t4 VPB.t12 510.753
R158 VPB.t0 VPB.t14 423.925
R159 VPB.t1 VPB.t5 291.13
R160 VPB.t19 VPB.t2 280.914
R161 VPB.t18 VPB.t11 273.253
R162 VPB VPB.t16 268.146
R163 VPB.t9 VPB.t17 255.376
R164 VPB.t16 VPB.t6 255.376
R165 VPB.t10 VPB.t15 229.839
R166 VPB.t7 VPB.t22 229.839
R167 VPB.t21 VPB.t7 229.839
R168 VPB.t20 VPB.t21 229.839
R169 VPB.t17 VPB.t3 214.517
R170 VPB.t5 VPB.t13 214.517
R171 VPB.t6 VPB.t1 214.517
R172 a_2067_74.n10 a_2067_74.n9 699.023
R173 a_2067_74.n6 a_2067_74.t3 675.721
R174 a_2067_74.n9 a_2067_74.t2 655.357
R175 a_2067_74.n2 a_2067_74.n1 308.481
R176 a_2067_74.n3 a_2067_74.t9 308.481
R177 a_2067_74.n7 a_2067_74.t4 303.139
R178 a_2067_74.n0 a_2067_74.t11 289.2
R179 a_2067_74.n2 a_2067_74.n0 266.707
R180 a_2067_74.n5 a_2067_74.t6 245.364
R181 a_2067_74.n4 a_2067_74.t7 242.315
R182 a_2067_74.n4 a_2067_74.n3 234.573
R183 a_2067_74.n2 a_2067_74.t12 200.03
R184 a_2067_74.n3 a_2067_74.t8 200.03
R185 a_2067_74.n0 a_2067_74.t10 183.964
R186 a_2067_74.n7 a_2067_74.t0 157.032
R187 a_2067_74.n8 a_2067_74.n7 119.999
R188 a_2067_74.n3 a_2067_74.n2 86.7605
R189 a_2067_74.n8 a_2067_74.n6 73.0358
R190 a_2067_74.n5 a_2067_74.n4 54.3774
R191 a_2067_74.n6 a_2067_74.n5 44.3142
R192 a_2067_74.n10 a_2067_74.t5 35.1791
R193 a_2067_74.t1 a_2067_74.n10 35.1791
R194 a_2067_74.n9 a_2067_74.n8 4.4568
R195 a_2513_258.n1 a_2513_258.t0 772.977
R196 a_2513_258.n0 a_2513_258.t2 273.271
R197 a_2513_258.n0 a_2513_258.t3 272.825
R198 a_2513_258.t1 a_2513_258.n1 243.036
R199 a_2513_258.n1 a_2513_258.n0 150.231
R200 VGND.n64 VGND.t6 246.916
R201 VGND.n52 VGND.t1 245.442
R202 VGND.n47 VGND.t0 244.976
R203 VGND.n26 VGND.t13 240.054
R204 VGND.n10 VGND.t8 234.136
R205 VGND.n29 VGND.n28 207.109
R206 VGND.n72 VGND.n71 201.278
R207 VGND.n18 VGND.t10 178.81
R208 VGND.n22 VGND.t12 165.3
R209 VGND.n20 VGND.n19 124.466
R210 VGND.n4 VGND.n3 115.272
R211 VGND.n71 VGND.t4 70.0005
R212 VGND.n28 VGND.t14 62.8576
R213 VGND.n71 VGND.t2 51.4291
R214 VGND.n19 VGND.t11 51.3826
R215 VGND.n28 VGND.t7 40.0005
R216 VGND.n30 VGND.n27 36.1417
R217 VGND.n34 VGND.n14 36.1417
R218 VGND.n35 VGND.n34 36.1417
R219 VGND.n36 VGND.n35 36.1417
R220 VGND.n36 VGND.n12 36.1417
R221 VGND.n40 VGND.n12 36.1417
R222 VGND.n41 VGND.n40 36.1417
R223 VGND.n42 VGND.n41 36.1417
R224 VGND.n46 VGND.n45 36.1417
R225 VGND.n51 VGND.n8 36.1417
R226 VGND.n53 VGND.n6 36.1417
R227 VGND.n57 VGND.n6 36.1417
R228 VGND.n58 VGND.n57 36.1417
R229 VGND.n59 VGND.n58 36.1417
R230 VGND.n65 VGND.n1 36.1417
R231 VGND.n69 VGND.n1 36.1417
R232 VGND.n70 VGND.n69 36.1417
R233 VGND.n3 VGND.t9 34.0546
R234 VGND.n26 VGND.n16 33.1299
R235 VGND.n64 VGND.n63 32.377
R236 VGND.n22 VGND.n21 32.0005
R237 VGND.n59 VGND.n4 30.1181
R238 VGND.n21 VGND.n20 28.2358
R239 VGND.n47 VGND.n46 26.3534
R240 VGND.n53 VGND.n52 25.224
R241 VGND.n3 VGND.t5 22.7032
R242 VGND.n52 VGND.n51 21.8358
R243 VGND.n22 VGND.n16 21.4593
R244 VGND.n19 VGND.t3 21.1849
R245 VGND.n47 VGND.n8 21.0829
R246 VGND.n63 VGND.n4 17.3181
R247 VGND.n65 VGND.n64 15.0593
R248 VGND.n27 VGND.n26 14.3064
R249 VGND.n72 VGND.n70 13.5534
R250 VGND.n70 VGND.n0 9.3005
R251 VGND.n69 VGND.n68 9.3005
R252 VGND.n67 VGND.n1 9.3005
R253 VGND.n66 VGND.n65 9.3005
R254 VGND.n64 VGND.n2 9.3005
R255 VGND.n63 VGND.n62 9.3005
R256 VGND.n61 VGND.n4 9.3005
R257 VGND.n60 VGND.n59 9.3005
R258 VGND.n58 VGND.n5 9.3005
R259 VGND.n57 VGND.n56 9.3005
R260 VGND.n55 VGND.n6 9.3005
R261 VGND.n54 VGND.n53 9.3005
R262 VGND.n52 VGND.n7 9.3005
R263 VGND.n51 VGND.n50 9.3005
R264 VGND.n49 VGND.n8 9.3005
R265 VGND.n48 VGND.n47 9.3005
R266 VGND.n46 VGND.n9 9.3005
R267 VGND.n45 VGND.n44 9.3005
R268 VGND.n43 VGND.n42 9.3005
R269 VGND.n41 VGND.n11 9.3005
R270 VGND.n40 VGND.n39 9.3005
R271 VGND.n38 VGND.n12 9.3005
R272 VGND.n37 VGND.n36 9.3005
R273 VGND.n35 VGND.n13 9.3005
R274 VGND.n34 VGND.n33 9.3005
R275 VGND.n32 VGND.n14 9.3005
R276 VGND.n31 VGND.n30 9.3005
R277 VGND.n27 VGND.n15 9.3005
R278 VGND.n26 VGND.n25 9.3005
R279 VGND.n24 VGND.n16 9.3005
R280 VGND.n21 VGND.n17 9.3005
R281 VGND.n23 VGND.n22 9.3005
R282 VGND.n73 VGND.n72 7.43488
R283 VGND.n20 VGND.n18 6.79022
R284 VGND.n30 VGND.n29 6.77697
R285 VGND.n45 VGND.n10 6.77697
R286 VGND.n29 VGND.n14 4.51815
R287 VGND.n42 VGND.n10 4.51815
R288 VGND.n18 VGND.n17 0.5771
R289 VGND VGND.n73 0.160103
R290 VGND.n73 VGND.n0 0.1477
R291 VGND.n23 VGND.n17 0.122949
R292 VGND.n24 VGND.n23 0.122949
R293 VGND.n25 VGND.n24 0.122949
R294 VGND.n25 VGND.n15 0.122949
R295 VGND.n31 VGND.n15 0.122949
R296 VGND.n32 VGND.n31 0.122949
R297 VGND.n33 VGND.n32 0.122949
R298 VGND.n33 VGND.n13 0.122949
R299 VGND.n37 VGND.n13 0.122949
R300 VGND.n38 VGND.n37 0.122949
R301 VGND.n39 VGND.n38 0.122949
R302 VGND.n39 VGND.n11 0.122949
R303 VGND.n43 VGND.n11 0.122949
R304 VGND.n44 VGND.n43 0.122949
R305 VGND.n44 VGND.n9 0.122949
R306 VGND.n48 VGND.n9 0.122949
R307 VGND.n49 VGND.n48 0.122949
R308 VGND.n50 VGND.n49 0.122949
R309 VGND.n50 VGND.n7 0.122949
R310 VGND.n54 VGND.n7 0.122949
R311 VGND.n55 VGND.n54 0.122949
R312 VGND.n56 VGND.n55 0.122949
R313 VGND.n56 VGND.n5 0.122949
R314 VGND.n60 VGND.n5 0.122949
R315 VGND.n61 VGND.n60 0.122949
R316 VGND.n62 VGND.n61 0.122949
R317 VGND.n62 VGND.n2 0.122949
R318 VGND.n66 VGND.n2 0.122949
R319 VGND.n67 VGND.n66 0.122949
R320 VGND.n68 VGND.n67 0.122949
R321 VGND.n68 VGND.n0 0.122949
R322 VNB.t1 VNB.t14 3880.31
R323 VNB.t12 VNB.t4 3857.22
R324 VNB.t2 VNB.t1 3383.73
R325 VNB.t21 VNB.t20 2448.29
R326 VNB.t18 VNB.t19 2402.1
R327 VNB.t15 VNB.t13 2367.45
R328 VNB.t16 VNB.t15 2286.61
R329 VNB.t9 VNB.t7 2286.61
R330 VNB.t0 VNB.t10 2171.13
R331 VNB.t14 VNB.t12 2148.03
R332 VNB.t6 VNB.t3 1328.08
R333 VNB.t19 VNB.t5 1304.99
R334 VNB.t11 VNB.t21 1177.95
R335 VNB.t7 VNB.t16 1154.86
R336 VNB VNB.t6 1143.31
R337 VNB.t20 VNB.t18 1039.37
R338 VNB.t5 VNB.t17 993.177
R339 VNB.t8 VNB.t11 900.788
R340 VNB.t4 VNB.t8 900.788
R341 VNB.t13 VNB.t2 900.788
R342 VNB.t10 VNB.t9 900.788
R343 VNB.t3 VNB.t0 900.788
R344 SCE.n0 SCE.t2 334.454
R345 SCE.n1 SCE.t1 327.014
R346 SCE.n0 SCE.t0 318.389
R347 SCE.n2 SCE.t3 201.508
R348 SCE.n2 SCE.n1 157.887
R349 SCE.n1 SCE.n0 22.152
R350 SCE SCE.n2 3.41394
R351 a_27_74.n1 a_27_74.t2 436.18
R352 a_27_74.t1 a_27_74.n1 367.668
R353 a_27_74.n0 a_27_74.t3 299.678
R354 a_27_74.n0 a_27_74.t0 242.244
R355 a_27_74.n1 a_27_74.n0 64.448
R356 SCD.n0 SCD.t1 406.094
R357 SCD.n0 SCD.t0 154.923
R358 SCD SCD.n0 70.0255
R359 a_495_74.t0 a_495_74.t1 68.5719
R360 a_871_74.t0 a_871_74.n7 944.889
R361 a_871_74.n7 a_871_74.n4 448
R362 a_871_74.n0 a_871_74.t2 393.979
R363 a_871_74.n5 a_871_74.t1 326.125
R364 a_871_74.n3 a_871_74.n2 221.376
R365 a_871_74.n5 a_871_74.t3 213.02
R366 a_871_74.n6 a_871_74.n5 195.871
R367 a_871_74.n1 a_871_74.t4 163.881
R368 a_871_74.n4 a_871_74.n3 152
R369 a_871_74.n6 a_871_74.t5 151.421
R370 a_871_74.n7 a_871_74.n6 119.383
R371 a_871_74.n4 a_871_74.n0 83.6776
R372 a_871_74.n1 a_871_74.n0 30.9964
R373 a_871_74.n3 a_871_74.n1 24.6743
R374 a_2277_455.t0 a_2277_455.t1 1402.16
R375 SET_B.n1 SET_B.t2 335.793
R376 SET_B.n0 SET_B.t1 277.072
R377 SET_B.n0 SET_B.t0 269.545
R378 SET_B.n1 SET_B.t3 212.081
R379 SET_B SET_B.n1 171.298
R380 SET_B SET_B.n0 77.7214
R381 a_304_464.n1 a_304_464.t3 663.357
R382 a_304_464.n3 a_304_464.n2 341.76
R383 a_304_464.n1 a_304_464.t5 330.421
R384 a_304_464.n2 a_304_464.n0 326.587
R385 a_304_464.n0 a_304_464.t0 177.143
R386 a_304_464.n2 a_304_464.n1 176.941
R387 a_304_464.n3 a_304_464.t4 64.6411
R388 a_304_464.t1 a_304_464.n3 64.6411
R389 a_304_464.n0 a_304_464.t2 48.5719
R390 Q_N Q_N.t2 268.099
R391 Q_N.n2 Q_N.n1 185
R392 Q_N.n1 Q_N.n0 185
R393 Q_N.n1 Q_N.t1 25.9464
R394 Q_N.n1 Q_N.t0 22.7032
R395 Q_N.n0 Q_N 10.8057
R396 Q_N Q_N.n2 8.14595
R397 Q_N.n2 Q_N 4.15634
R398 Q_N.n0 Q_N 1.4966
R399 D.n0 D.t1 435.675
R400 D D.n0 159.024
R401 D.n0 D.t0 126.927
R402 a_229_74.t0 a_229_74.t1 68.5719
R403 a_1274_81.t0 a_1274_81.t1 68.5719
R404 a_220_464.t0 a_220_464.t1 83.1099
R405 a_418_464.t0 a_418_464.t1 83.1099
R406 a_619_368.n2 a_619_368.n1 1870.25
R407 a_619_368.n1 a_619_368.n0 1420.29
R408 a_619_368.t0 a_619_368.n6 846.808
R409 a_619_368.n3 a_619_368.n2 766.38
R410 a_619_368.n3 a_619_368.t7 322.94
R411 a_619_368.n0 a_619_368.t4 303.661
R412 a_619_368.n6 a_619_368.n5 232.696
R413 a_619_368.n4 a_619_368.t6 226.809
R414 a_619_368.n4 a_619_368.t2 198.204
R415 a_619_368.n6 a_619_368.t1 185.407
R416 a_619_368.n2 a_619_368.t5 182.625
R417 a_619_368.n0 a_619_368.t3 159.06
R418 a_619_368.n1 a_619_368.t8 137.881
R419 a_619_368.n5 a_619_368.n3 43.0884
R420 a_619_368.n5 a_619_368.n4 37.9763
R421 a_2579_74.t0 a_2579_74.t1 68.5719
R422 a_3177_368.t1 a_3177_368.n4 251.756
R423 a_3177_368.n1 a_3177_368.t2 240.994
R424 a_3177_368.n3 a_3177_368.n0 240.197
R425 a_3177_368.n4 a_3177_368.n3 183.81
R426 a_3177_368.n1 a_3177_368.t4 182.109
R427 a_3177_368.n2 a_3177_368.t3 179.947
R428 a_3177_368.n4 a_3177_368.t0 150.452
R429 a_3177_368.n2 a_3177_368.n1 60.6419
R430 a_3177_368.n3 a_3177_368.n2 4.38232
R431 Q.n0 Q.t2 293.426
R432 Q.n1 Q.n0 185
R433 Q.n2 Q.n1 185
R434 Q.n1 Q.t0 22.7032
R435 Q.n1 Q.t1 22.7032
R436 Q.n2 Q 12.2358
R437 Q.n0 Q 4.70638
R438 Q Q.n2 1.69462
R439 CLK.n0 CLK.t0 307.628
R440 CLK CLK.n0 163.97
R441 CLK.n0 CLK.t1 154.24
R442 a_1201_463.t0 a_1201_463.t1 126.644
R443 a_2501_74.t0 a_2501_74.t1 68.5719
C0 Q_N SET_B 3.93e-19
C1 CLK SET_B 3.74e-21
C2 VPB Q_N 0.006153f
C3 VPB CLK 0.049509f
C4 D SET_B 3.04e-20
C5 VPB SET_B 0.183086f
C6 VPB D 0.05662f
C7 a_1252_376# SET_B 0.02559f
C8 a_1252_376# VPB 0.129013f
C9 VGND Q_N 0.149388f
C10 CLK VGND 0.055231f
C11 VGND SET_B 0.187003f
C12 Q_N VPWR 0.21216f
C13 Q SET_B 5.97e-20
C14 SCD SET_B 5.87e-20
C15 VPWR SET_B 0.177582f
C16 SCD CLK 0.042278f
C17 CLK VPWR 0.018279f
C18 VPB Q 0.007028f
C19 VPB VGND 0.034506f
C20 D VGND 0.055069f
C21 VPB SCD 0.109093f
C22 VPB VPWR 0.474051f
C23 SCE SET_B 6.98e-20
C24 D SCD 0.003254f
C25 D VPWR 0.014267f
C26 SET_B a_1794_74# 0.018987f
C27 VPB SCE 0.148993f
C28 SCE D 0.18402f
C29 a_1252_376# VGND 0.130168f
C30 a_1252_376# SCD 4.12e-21
C31 a_1252_376# VPWR 0.025123f
C32 a_1252_376# a_1794_74# 0.004016f
C33 VGND Q 0.166542f
C34 SCD VGND 0.053237f
C35 VGND VPWR 0.226266f
C36 Q VPWR 0.227139f
C37 SCD VPWR 0.018026f
C38 SCE VGND 0.038265f
C39 SCE SCD 0.069333f
C40 SCE VPWR 0.041828f
C41 VGND a_1794_74# 0.317642f
C42 Q VNB 0.030869f
C43 Q_N VNB 0.015446f
C44 VGND VNB 2.09541f
C45 SET_B VNB 0.278691f
C46 VPWR VNB 1.60417f
C47 CLK VNB 0.143091f
C48 SCD VNB 0.170939f
C49 D VNB 0.144947f
C50 SCE VNB 0.36562f
C51 VPB VNB 4.04885f
C52 a_1794_74# VNB 0.031235f
C53 a_1252_376# VNB 0.185835f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfsbp_1 VNB VPB VPWR VGND SET_B Q Q_N SCD CLK SCE D
X0 VPWR.t3 SCD.t0 a_416_464.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.93 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 VGND.t9 CLK.t0 a_594_74.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 a_416_464.t1 a_27_74.t2 a_290_464.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1536 ps=1.12 w=0.64 l=0.15
X3 a_781_74.t0 a_594_74.t2 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t11 CLK.t1 a_594_74.t0 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
X5 VGND.t8 SET_B.t0 a_1954_74.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1323 pd=1.05 as=0.0819 ps=0.81 w=0.42 l=0.15
X6 a_995_74.t2 a_781_74.t2 a_290_464.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.10585 pd=0.95 as=0.1197 ps=1.41 w=0.42 l=0.15
X7 a_290_464.t4 D.t0 a_228_74.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X8 VGND.t10 SCE.t0 a_27_74.t0 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 a_1684_74.t1 a_995_74.t3 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.25575 ps=1.465 w=0.64 l=0.15
X10 a_995_74.t1 a_594_74.t3 a_290_464.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0945 pd=0.87 as=0.18665 ps=1.8 w=0.42 l=0.15
X11 VPWR.t10 SET_B.t1 a_1163_48# VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.15875 pd=1.39 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VPWR.t13 SCE.t1 a_27_74.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1888 ps=1.87 w=0.64 l=0.15
X13 a_1133_478.t1 a_594_74.t4 a_995_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0837 pd=0.865 as=0.10585 ps=0.95 w=0.42 l=0.15
X14 VPWR.t6 a_1163_48# a_1133_478.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.11235 pd=0.955 as=0.0837 ps=0.865 w=0.42 l=0.15
X15 VGND.t3 SCD.t1 a_392_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X16 a_1762_74# SET_B.t2 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.063 ps=0.72 w=0.42 l=0.15
X17 VPWR.t14 a_1924_48.t2 a_1712_374# VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X18 Q_N.t0 a_1762_74# VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.1673 ps=1.475 w=1.12 l=0.15
X19 a_1163_48# a_995_74.t4 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0924 pd=0.86 as=0.11235 ps=0.955 w=0.42 l=0.15
X20 a_1876_74.t0 a_594_74.t5 a_1762_74# VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.11955 ps=1.06 w=0.42 l=0.15
X21 VGND.t7 SET_B.t3 a_1411_74# VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.25575 pd=1.465 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 a_1924_48.t1 a_1762_74# VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1323 ps=1.05 w=0.42 l=0.15
X23 VGND.t1 a_1762_74# a_2556_94.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.21455 pd=1.355 as=0.1824 ps=1.85 w=0.64 l=0.15
X24 a_1600_347# a_995_74.t5 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.15875 ps=1.39 w=1 l=0.15
X25 VPWR.t2 a_1762_74# a_2556_94.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2436 ps=2.26 w=0.84 l=0.15
X26 a_1762_74# a_781_74.t3 a_1684_74.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.11955 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
X27 Q.t0 a_2556_94.t2 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.1862 ps=1.475 w=1.12 l=0.15
X28 Q_N.t1 a_1762_74# VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X29 a_228_74.t1 a_27_74.t3 VGND.t11 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0882 ps=0.84 w=0.42 l=0.15
X30 a_781_74.t1 a_594_74.t6 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X31 VGND.t4 a_1163_48# a_1115_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.17255 pd=1.68 as=0.0504 ps=0.66 w=0.42 l=0.15
X32 VPWR.t0 a_1762_74# a_1924_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1673 pd=1.475 as=0.1218 ps=1.42 w=0.42 l=0.15
X33 a_290_464.t0 D.t1 a_206_464.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1536 pd=1.12 as=0.0864 ps=0.91 w=0.64 l=0.15
X34 Q.t1 a_2556_94.t3 VGND.t12 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.21455 ps=1.355 w=0.74 l=0.15
X35 a_206_464.t1 SCE.t2 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.096 ps=0.94 w=0.64 l=0.15
X36 a_392_74.t1 SCE.t3 a_290_464.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 a_1954_74.t0 a_1924_48.t3 a_1876_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 SCD.n2 SCD.t1 201.87
R1 SCD.n0 SCD.t0 171.781
R2 SCD SCD.n0 154.133
R3 SCD.n4 SCD.n3 152
R4 SCD.n2 SCD.n1 152
R5 SCD.n3 SCD.n0 35.2435
R6 SCD.n3 SCD.n2 35.2435
R7 SCD SCD.n4 18.591
R8 SCD.n1 SCD 16.7624
R9 SCD.n1 SCD 5.79098
R10 SCD.n4 SCD 3.9624
R11 a_416_464.t0 a_416_464.t1 83.1099
R12 VPWR.n52 VPWR.t3 721.532
R13 VPWR.n12 VPWR.n11 639.212
R14 VPWR.n9 VPWR.n8 622.889
R15 VPWR.n27 VPWR.n16 622.271
R16 VPWR.n21 VPWR.n20 607.497
R17 VPWR.n50 VPWR.n5 606.333
R18 VPWR.n58 VPWR.n1 605.365
R19 VPWR.n19 VPWR.n18 327.846
R20 VPWR.n8 VPWR.t4 178.238
R21 VPWR.n11 VPWR.t10 112.572
R22 VPWR.n8 VPWR.t6 72.7029
R23 VPWR.n20 VPWR.t1 72.2026
R24 VPWR.n16 VPWR.t9 70.3576
R25 VPWR.n16 VPWR.t14 70.3576
R26 VPWR.n20 VPWR.t0 70.3576
R27 VPWR.n1 VPWR.t12 46.1724
R28 VPWR.n1 VPWR.t13 46.1724
R29 VPWR.n18 VPWR.t7 42.7085
R30 VPWR.n56 VPWR.n2 36.1417
R31 VPWR.n57 VPWR.n56 36.1417
R32 VPWR.n44 VPWR.n43 36.1417
R33 VPWR.n45 VPWR.n44 36.1417
R34 VPWR.n45 VPWR.n6 36.1417
R35 VPWR.n49 VPWR.n6 36.1417
R36 VPWR.n22 VPWR.n17 36.1417
R37 VPWR.n26 VPWR.n17 36.1417
R38 VPWR.n29 VPWR.n28 36.1417
R39 VPWR.n29 VPWR.n14 36.1417
R40 VPWR.n33 VPWR.n14 36.1417
R41 VPWR.n34 VPWR.n33 36.1417
R42 VPWR.n35 VPWR.n34 36.1417
R43 VPWR.n39 VPWR.n38 36.1417
R44 VPWR.n40 VPWR.n39 36.1417
R45 VPWR.n18 VPWR.t2 35.1791
R46 VPWR.n51 VPWR.n50 34.2593
R47 VPWR.n11 VPWR.t5 33.6312
R48 VPWR.n52 VPWR.n2 29.7417
R49 VPWR.n5 VPWR.t8 26.3844
R50 VPWR.n5 VPWR.t11 26.3844
R51 VPWR.n28 VPWR.n27 25.977
R52 VPWR.n58 VPWR.n57 22.9652
R53 VPWR.n52 VPWR.n51 22.5887
R54 VPWR.n38 VPWR.n12 19.577
R55 VPWR.n35 VPWR.n12 16.5652
R56 VPWR.n22 VPWR.n21 14.3064
R57 VPWR.n43 VPWR.n9 13.177
R58 VPWR.n50 VPWR.n49 13.177
R59 VPWR.n27 VPWR.n26 10.1652
R60 VPWR.n23 VPWR.n22 9.3005
R61 VPWR.n24 VPWR.n17 9.3005
R62 VPWR.n26 VPWR.n25 9.3005
R63 VPWR.n28 VPWR.n15 9.3005
R64 VPWR.n30 VPWR.n29 9.3005
R65 VPWR.n31 VPWR.n14 9.3005
R66 VPWR.n33 VPWR.n32 9.3005
R67 VPWR.n34 VPWR.n13 9.3005
R68 VPWR.n36 VPWR.n35 9.3005
R69 VPWR.n38 VPWR.n37 9.3005
R70 VPWR.n39 VPWR.n10 9.3005
R71 VPWR.n41 VPWR.n40 9.3005
R72 VPWR.n43 VPWR.n42 9.3005
R73 VPWR.n44 VPWR.n7 9.3005
R74 VPWR.n46 VPWR.n45 9.3005
R75 VPWR.n47 VPWR.n6 9.3005
R76 VPWR.n49 VPWR.n48 9.3005
R77 VPWR.n50 VPWR.n4 9.3005
R78 VPWR.n51 VPWR.n3 9.3005
R79 VPWR.n53 VPWR.n52 9.3005
R80 VPWR.n54 VPWR.n2 9.3005
R81 VPWR.n56 VPWR.n55 9.3005
R82 VPWR.n57 VPWR.n0 9.3005
R83 VPWR.n21 VPWR.n19 7.48727
R84 VPWR.n59 VPWR.n58 7.27223
R85 VPWR.n40 VPWR.n9 4.14168
R86 VPWR.n23 VPWR.n19 0.214419
R87 VPWR VPWR.n59 0.157962
R88 VPWR.n59 VPWR.n0 0.149814
R89 VPWR.n24 VPWR.n23 0.122949
R90 VPWR.n25 VPWR.n24 0.122949
R91 VPWR.n25 VPWR.n15 0.122949
R92 VPWR.n30 VPWR.n15 0.122949
R93 VPWR.n31 VPWR.n30 0.122949
R94 VPWR.n32 VPWR.n31 0.122949
R95 VPWR.n32 VPWR.n13 0.122949
R96 VPWR.n36 VPWR.n13 0.122949
R97 VPWR.n37 VPWR.n36 0.122949
R98 VPWR.n37 VPWR.n10 0.122949
R99 VPWR.n41 VPWR.n10 0.122949
R100 VPWR.n42 VPWR.n41 0.122949
R101 VPWR.n42 VPWR.n7 0.122949
R102 VPWR.n46 VPWR.n7 0.122949
R103 VPWR.n47 VPWR.n46 0.122949
R104 VPWR.n48 VPWR.n47 0.122949
R105 VPWR.n48 VPWR.n4 0.122949
R106 VPWR.n4 VPWR.n3 0.122949
R107 VPWR.n53 VPWR.n3 0.122949
R108 VPWR.n54 VPWR.n53 0.122949
R109 VPWR.n55 VPWR.n54 0.122949
R110 VPWR.n55 VPWR.n0 0.122949
R111 VPB.t7 VPB.t18 1284.54
R112 VPB.t5 VPB.t14 556.721
R113 VPB.t11 VPB.t9 520.968
R114 VPB.t2 VPB.t1 510.753
R115 VPB.t12 VPB.t0 510.753
R116 VPB.t8 VPB.t6 349.866
R117 VPB.t4 VPB.t15 321.774
R118 VPB.t9 VPB.t3 309.005
R119 VPB.t6 VPB.t13 301.344
R120 VPB.t13 VPB.t7 275.807
R121 VPB.t3 VPB.t8 265.591
R122 VPB.t1 VPB.t10 257.93
R123 VPB.t0 VPB.t2 257.93
R124 VPB VPB.t17 257.93
R125 VPB.t18 VPB.t12 229.839
R126 VPB.t14 VPB.t11 229.839
R127 VPB.t17 VPB.t16 229.839
R128 VPB.t15 VPB.t5 214.517
R129 VPB.t16 VPB.t4 214.517
R130 CLK.n0 CLK.t1 283.195
R131 CLK.n0 CLK.t0 178.34
R132 CLK CLK.n0 157.091
R133 a_594_74.n1 a_594_74.n0 1418.95
R134 a_594_74.t0 a_594_74.n5 866.914
R135 a_594_74.n2 a_594_74.n1 819.4
R136 a_594_74.n0 a_594_74.t5 551.087
R137 a_594_74.n2 a_594_74.t3 294.021
R138 a_594_74.n3 a_594_74.t2 261.62
R139 a_594_74.n5 a_594_74.n4 210.946
R140 a_594_74.n5 a_594_74.t1 198.566
R141 a_594_74.n3 a_594_74.t6 181.196
R142 a_594_74.n1 a_594_74.t4 162.542
R143 a_594_74.n4 a_594_74.n2 62.0763
R144 a_594_74.n4 a_594_74.n3 12.4157
R145 VGND.n37 VGND.t4 268.269
R146 VGND.n50 VGND.t3 246.333
R147 VGND.n57 VGND.n56 206.916
R148 VGND.n21 VGND.n20 185
R149 VGND.n19 VGND.n18 185
R150 VGND.n30 VGND.n8 185
R151 VGND.n31 VGND.n30 185
R152 VGND.n14 VGND.t0 154.727
R153 VGND.n15 VGND.n13 122.15
R154 VGND.n48 VGND.n4 115.272
R155 VGND.n20 VGND.n19 100.001
R156 VGND.n13 VGND.t1 75.938
R157 VGND.n56 VGND.t11 60.0005
R158 VGND.n56 VGND.t10 60.0005
R159 VGND.n19 VGND.t2 40.0005
R160 VGND.n20 VGND.t8 40.0005
R161 VGND.n23 VGND.n10 36.1417
R162 VGND.n27 VGND.n10 36.1417
R163 VGND.n28 VGND.n27 36.1417
R164 VGND.n36 VGND.n35 36.1417
R165 VGND.n38 VGND.n36 36.1417
R166 VGND.n42 VGND.n6 36.1417
R167 VGND.n43 VGND.n42 36.1417
R168 VGND.n44 VGND.n43 36.1417
R169 VGND.n44 VGND.n3 36.1417
R170 VGND.n54 VGND.n1 36.1417
R171 VGND.n55 VGND.n54 36.1417
R172 VGND.n50 VGND.n49 35.0123
R173 VGND.n23 VGND.n22 34.092
R174 VGND.n4 VGND.t5 34.0546
R175 VGND.n18 VGND.n12 30.5783
R176 VGND.n13 VGND.t12 30.2643
R177 VGND.n48 VGND.n3 27.8593
R178 VGND.n14 VGND.n12 25.977
R179 VGND.n4 VGND.t9 22.7032
R180 VGND.n29 VGND.t7 21.4291
R181 VGND.n49 VGND.n48 19.577
R182 VGND.n57 VGND.n55 19.2005
R183 VGND.n29 VGND.t6 17.6005
R184 VGND.n50 VGND.n1 12.424
R185 VGND.n31 VGND.n28 10.482
R186 VGND.n55 VGND.n0 9.3005
R187 VGND.n54 VGND.n53 9.3005
R188 VGND.n52 VGND.n1 9.3005
R189 VGND.n51 VGND.n50 9.3005
R190 VGND.n49 VGND.n2 9.3005
R191 VGND.n48 VGND.n47 9.3005
R192 VGND.n46 VGND.n3 9.3005
R193 VGND.n45 VGND.n44 9.3005
R194 VGND.n43 VGND.n5 9.3005
R195 VGND.n42 VGND.n41 9.3005
R196 VGND.n40 VGND.n6 9.3005
R197 VGND.n39 VGND.n38 9.3005
R198 VGND.n36 VGND.n7 9.3005
R199 VGND.n35 VGND.n34 9.3005
R200 VGND.n33 VGND.n32 9.3005
R201 VGND.n28 VGND.n9 9.3005
R202 VGND.n27 VGND.n26 9.3005
R203 VGND.n25 VGND.n10 9.3005
R204 VGND.n24 VGND.n23 9.3005
R205 VGND.n22 VGND.n11 9.3005
R206 VGND.n18 VGND.n17 9.3005
R207 VGND.n16 VGND.n12 9.3005
R208 VGND.n38 VGND.n37 8.28285
R209 VGND.n58 VGND.n57 7.43488
R210 VGND.n15 VGND.n14 7.00747
R211 VGND.n21 VGND.n18 5.85671
R212 VGND.n35 VGND.n8 5.84498
R213 VGND.n32 VGND.n8 5.22977
R214 VGND.n32 VGND.n31 3.27855
R215 VGND.n22 VGND.n21 2.17566
R216 VGND.n30 VGND.n29 1.6005
R217 VGND.n37 VGND.n6 1.50638
R218 VGND.n16 VGND.n15 0.173805
R219 VGND VGND.n58 0.160103
R220 VGND.n58 VGND.n0 0.1477
R221 VGND.n17 VGND.n16 0.122949
R222 VGND.n17 VGND.n11 0.122949
R223 VGND.n24 VGND.n11 0.122949
R224 VGND.n25 VGND.n24 0.122949
R225 VGND.n26 VGND.n25 0.122949
R226 VGND.n26 VGND.n9 0.122949
R227 VGND.n33 VGND.n9 0.122949
R228 VGND.n34 VGND.n33 0.122949
R229 VGND.n34 VGND.n7 0.122949
R230 VGND.n39 VGND.n7 0.122949
R231 VGND.n40 VGND.n39 0.122949
R232 VGND.n41 VGND.n40 0.122949
R233 VGND.n41 VGND.n5 0.122949
R234 VGND.n45 VGND.n5 0.122949
R235 VGND.n46 VGND.n45 0.122949
R236 VGND.n47 VGND.n46 0.122949
R237 VGND.n47 VGND.n2 0.122949
R238 VGND.n51 VGND.n2 0.122949
R239 VGND.n52 VGND.n51 0.122949
R240 VGND.n53 VGND.n52 0.122949
R241 VGND.n53 VGND.n0 0.122949
R242 VNB.n0 VNB 19563.3
R243 VNB.t12 VNB.t6 3418.37
R244 VNB.t9 VNB.t7 2471.39
R245 VNB.t0 VNB.t1 2459.84
R246 VNB.t2 VNB.t0 2448.29
R247 VNB.t15 VNB.t3 2436.75
R248 VNB VNB.t12 2396.24
R249 VNB.t6 VNB.t9 2286.61
R250 VNB.t13 VNB.t2 1801.57
R251 VNB.t1 VNB.t18 1766.93
R252 VNB.t10 VNB.t8 1316.54
R253 VNB.t17 VNB.t16 1316.54
R254 VNB.t5 VNB.t13 1247.24
R255 VNB.t7 VNB.t15 1154.86
R256 VNB.t16 VNB 1143.31
R257 VNB.t4 VNB.t14 993.177
R258 VNB.t8 VNB.t5 900.788
R259 VNB.t3 VNB.t4 900.788
R260 VNB.t14 VNB.t17 900.788
R261 VNB.n0 VNB.t10 612.073
R262 VNB.n0 VNB.t11 144.601
R263 VNB.t12 VNB.n0 64.1137
R264 a_27_74.n1 a_27_74.t2 452.914
R265 a_27_74.t1 a_27_74.n1 359.966
R266 a_27_74.n0 a_27_74.t3 321.952
R267 a_27_74.n0 a_27_74.t0 239.352
R268 a_27_74.n1 a_27_74.n0 65.2495
R269 a_290_464.n1 a_290_464.t3 670.163
R270 a_290_464.n3 a_290_464.n2 632.163
R271 a_290_464.n1 a_290_464.t2 352.433
R272 a_290_464.n2 a_290_464.n0 329.108
R273 a_290_464.n2 a_290_464.n1 160.995
R274 a_290_464.n3 a_290_464.t5 73.8755
R275 a_290_464.t0 a_290_464.n3 73.8755
R276 a_290_464.n0 a_290_464.t1 40.0005
R277 a_290_464.n0 a_290_464.t4 40.0005
R278 a_781_74.t0 a_781_74.n5 1000.91
R279 a_781_74.n5 a_781_74.n4 514.165
R280 a_781_74.n2 a_781_74.n0 356.68
R281 a_781_74.n1 a_781_74.t1 343.483
R282 a_781_74.n4 a_781_74.t3 236.18
R283 a_781_74.n5 a_781_74.n2 185.895
R284 a_781_74.n1 a_781_74.t2 176.542
R285 a_781_74.n4 a_781_74.n3 132.477
R286 a_781_74.n2 a_781_74.n1 126.666
R287 SET_B.n0 SET_B.t0 332.377
R288 SET_B.n1 SET_B.t1 293.752
R289 SET_B.n0 SET_B.t2 272.611
R290 SET_B.n1 SET_B.t3 237.787
R291 SET_B SET_B.n1 173.186
R292 SET_B SET_B.n0 121.01
R293 a_1954_74.t0 a_1954_74.t1 111.43
R294 a_995_74.n5 a_995_74.n4 660.335
R295 a_995_74.t1 a_995_74.n5 317.348
R296 a_995_74.n2 a_995_74.t4 308.481
R297 a_995_74.n0 a_995_74.t5 251.956
R298 a_995_74.n3 a_995_74.n0 238.327
R299 a_995_74.n2 a_995_74.n1 220.113
R300 a_995_74.n0 a_995_74.t3 188.565
R301 a_995_74.n3 a_995_74.n2 152
R302 a_995_74.n4 a_995_74.t0 112.469
R303 a_995_74.n4 a_995_74.t2 110.124
R304 a_995_74.n5 a_995_74.n3 102.4
R305 D.n0 D.t0 412.913
R306 D.n0 D.t1 184.5
R307 D D.n0 163.831
R308 a_228_74.t0 a_228_74.t1 68.5719
R309 SCE.n2 SCE.t3 478.036
R310 SCE.n1 SCE.t2 313.033
R311 SCE.n0 SCE.t0 303.514
R312 SCE.n0 SCE.t1 232.7
R313 SCE.n2 SCE.n1 152
R314 SCE.n1 SCE.n0 24.1005
R315 SCE SCE.n2 1.1205
R316 a_1684_74.t0 a_1684_74.t1 45.0005
R317 a_1133_478.n0 a_1133_478.t1 102.627
R318 a_1133_478.n0 a_1133_478.t0 43.5989
R319 a_1133_478.n1 a_1133_478.n0 29.7363
R320 a_392_74.t0 a_392_74.t1 68.5719
R321 a_1924_48.n1 a_1924_48.t0 847.628
R322 a_1924_48.n0 a_1924_48.t2 605.348
R323 a_1924_48.n1 a_1924_48.n0 242.353
R324 a_1924_48.t1 a_1924_48.n1 240.709
R325 a_1924_48.n0 a_1924_48.t3 120.793
R326 Q_N.n0 Q_N.t0 297.089
R327 Q_N.t1 Q_N.n0 279.738
R328 Q_N.n1 Q_N.t1 279.738
R329 Q_N.n1 Q_N 8.40454
R330 Q_N.n0 Q_N 3.23282
R331 Q_N Q_N.n1 1.16414
R332 a_1876_74.t0 a_1876_74.t1 68.5719
R333 a_2556_94.t0 a_2556_94.n1 424.053
R334 a_2556_94.n0 a_2556_94.t2 276.485
R335 a_2556_94.n1 a_2556_94.t1 224.958
R336 a_2556_94.n1 a_2556_94.n0 171.006
R337 a_2556_94.n0 a_2556_94.t3 169.106
R338 Q.n3 Q 589.777
R339 Q.n3 Q.n0 585
R340 Q.n4 Q.n3 585
R341 Q.n2 Q.t1 279.738
R342 Q.t1 Q.n1 279.738
R343 Q.n3 Q.t0 26.3844
R344 Q Q.n4 12.8005
R345 Q.n1 Q 12.4184
R346 Q Q.n0 11.0811
R347 Q Q.n2 9.36169
R348 Q.n2 Q 4.77662
R349 Q Q.n0 3.05722
R350 Q.n1 Q 1.7199
R351 Q.n4 Q 1.33781
R352 a_206_464.t0 a_206_464.t1 83.1099
C0 SET_B a_1762_74# 0.285842f
C1 SET_B a_1712_374# 0.004653f
C2 VPB a_1762_74# 0.333316f
C3 VPB a_1712_374# 0.028224f
C4 a_1411_74# a_1762_74# 9.89e-20
C5 a_1762_74# a_1600_347# 0.084982f
C6 a_1712_374# a_1600_347# 0.112427f
C7 a_1762_74# a_1712_374# 0.032959f
C8 VGND Q 0.097701f
C9 VPWR Q 0.12168f
C10 VGND VPWR 0.18472f
C11 SCE VGND 0.035819f
C12 VGND SCD 0.034944f
C13 SCE VPWR 0.032579f
C14 VPWR SCD 0.017977f
C15 SCE SCD 0.055567f
C16 VGND a_1163_48# 0.136898f
C17 VPWR a_1163_48# 0.021227f
C18 VGND Q_N 0.125308f
C19 SET_B Q 7.39e-20
C20 SET_B VGND 0.117791f
C21 VPWR Q_N 0.077997f
C22 VPB Q 0.014268f
C23 VGND CLK 0.053575f
C24 SET_B VPWR 0.097759f
C25 SCE SET_B 1.01e-19
C26 SET_B SCD 1.13e-19
C27 VGND D 0.012851f
C28 VPB VGND 0.030722f
C29 CLK VPWR 0.015181f
C30 VPWR D 0.012857f
C31 CLK SCD 0.029934f
C32 VPB VPWR 0.371039f
C33 SCE D 0.181025f
C34 VPB SCE 0.132696f
C35 D SCD 0.004653f
C36 VPB SCD 0.10153f
C37 VGND a_1411_74# 0.005462f
C38 VGND a_1600_347# 3.88e-19
C39 a_1411_74# VPWR 4.86e-19
C40 a_1762_74# Q 0.003061f
C41 VPWR a_1600_347# 0.075186f
C42 SET_B a_1163_48# 0.017637f
C43 VGND a_1762_74# 0.140608f
C44 VGND a_1712_374# 5.31e-19
C45 VPB a_1163_48# 0.09468f
C46 VPWR a_1762_74# 0.16323f
C47 VPWR a_1712_374# 0.255861f
C48 a_1411_74# a_1163_48# 0.002876f
C49 a_1163_48# a_1600_347# 6.65e-19
C50 a_1762_74# a_1163_48# 0.00206f
C51 a_1712_374# a_1163_48# 6.62e-20
C52 SET_B Q_N 9.7e-20
C53 VPB Q_N 0.006643f
C54 SET_B CLK 9.24e-20
C55 SET_B D 2.25e-20
C56 VPB SET_B 0.214054f
C57 VPB CLK 0.036741f
C58 VPB D 0.073675f
C59 SET_B a_1600_347# 0.016963f
C60 a_1762_74# Q_N 0.052957f
C61 VPB a_1600_347# 0.021572f
C62 Q VNB 0.11043f
C63 Q_N VNB 0.028908f
C64 VGND VNB 1.6853f
C65 SET_B VNB 0.337867f
C66 VPWR VNB 1.28937f
C67 CLK VNB 0.118748f
C68 SCD VNB 0.177184f
C69 D VNB 0.115547f
C70 SCE VNB 0.320356f
C71 VPB VNB 3.31231f
C72 a_1600_347# VNB 0.001881f
C73 a_1163_48# VNB 0.197882f
C74 a_1762_74# VNB 0.521671f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrtp_4 VNB VPB VPWR RESET_B VGND D SCE SCD CLK Q
X0 Q.t2 a_2339_74.t3 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3293 ps=1.63 w=0.74 l=0.15
X1 VPWR.t7 a_2003_48.t3 a_1982_508.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.11235 pd=0.955 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR.t11 a_1745_74.t3 a_2003_48.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.17955 pd=1.535 as=0.08085 ps=0.805 w=0.42 l=0.15
X3 a_2003_48.t2 RESET_B.t0 VPWR.t15 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.08085 pd=0.805 as=0.11235 ps=0.955 w=0.42 l=0.15
X4 a_225_81.t0 SCD.t0 a_572_81.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X5 a_1397_138.t0 a_1367_112.t4 a_1319_138# VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X6 a_1233_138# a_1034_74.t2 a_415_81.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X7 a_312_81.t0 a_27_74.t2 a_225_81.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.07665 pd=0.785 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 VGND.t3 SCE.t0 a_27_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 a_1745_74.t0 a_1034_74.t3 a_1367_112.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2165 pd=1.54 as=0.1165 ps=1.065 w=0.64 l=0.15
X10 VGND.t6 a_2339_74.t4 Q.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.3293 pd=1.63 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VGND.t0 CLK.t0 a_855_368.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 a_1233_138# a_855_368.t2 a_415_81.t5 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X13 a_1982_508.t1 a_1034_74.t4 a_1745_74.t2 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.214125 ps=1.785 w=0.42 l=0.15
X14 VPWR.t3 SCE.t1 a_27_74.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3104 pd=1.61 as=0.1888 ps=1.87 w=0.64 l=0.15
X15 a_1745_74.t1 a_855_368.t3 a_1367_112.t3 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.214125 pd=1.785 as=0.15 ps=1.3 w=1 l=0.15
X16 VGND.t9 a_1745_74.t4 a_2339_74.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X17 VPWR.t13 CLK.t1 a_855_368.t1 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X18 a_1233_138# RESET_B.t1 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.139325 ps=1.145 w=0.42 l=0.15
X19 a_1367_112.t1 a_1233_138# VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X20 VGND.t4 RESET_B.t2 a_225_81.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_514_464.t1 a_27_74.t3 a_415_81.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1248 pd=1.03 as=0.096 ps=0.94 w=0.64 l=0.15
X22 a_1034_74.t1 a_855_368.t4 VPWR.t16 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_415_81.t3 D.t0 a_340_464.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 VPWR.t6 SCD.t1 a_514_464.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.1248 ps=1.03 w=0.64 l=0.15
X25 VPWR.t0 a_1367_112.t5 a_1342_463.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.139325 pd=1.145 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 VPWR.t10 a_2339_74.t5 Q.t5 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X27 VPWR.t9 a_2339_74.t6 Q.t4 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 VGND.t2 a_2003_48.t4 a_1955_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X29 a_2141_74.t1 RESET_B.t3 VGND.t10 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X30 Q.t3 a_2339_74.t7 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.203 ps=1.505 w=1.12 l=0.15
X31 VGND.t5 a_2339_74.t8 Q.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 a_572_81.t1 SCE.t2 a_415_81.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.13335 ps=1.055 w=0.42 l=0.15
X33 VPWR.t12 a_1745_74.t5 a_2339_74.t2 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.126 ps=1.14 w=0.84 l=0.15
X34 a_340_464.t0 SCE.t3 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.3104 ps=1.61 w=0.64 l=0.15
X35 a_2339_74.t0 a_1745_74.t6 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.17955 ps=1.535 w=0.84 l=0.15
X36 a_2003_48.t0 a_1745_74.t7 a_2141_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1512 pd=1.56 as=0.0441 ps=0.63 w=0.42 l=0.15
X37 a_415_81.t6 D.t1 a_312_81.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.13335 pd=1.055 as=0.07665 ps=0.785 w=0.42 l=0.15
X38 a_1367_112.t0 a_1233_138# VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.2838 ps=1.655 w=0.74 l=0.15
X39 a_1342_463.t1 a_855_368.t5 a_1233_138# VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X40 a_1034_74.t0 a_855_368.t6 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X41 a_415_81.t4 RESET_B.t4 VPWR.t14 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1344 ps=1.06 w=0.64 l=0.15
R0 a_2339_74.n14 a_2339_74.n13 312.673
R1 a_2339_74.n10 a_2339_74.n9 279.56
R2 a_2339_74.n2 a_2339_74.t5 249.148
R3 a_2339_74.n4 a_2339_74.n1 248.231
R4 a_2339_74.n6 a_2339_74.t6 248.231
R5 a_2339_74.n8 a_2339_74.t7 248.231
R6 a_2339_74.n13 a_2339_74.t1 187.306
R7 a_2339_74.n5 a_2339_74.n0 165.189
R8 a_2339_74.n2 a_2339_74.t8 157.745
R9 a_2339_74.n10 a_2339_74.t4 155.847
R10 a_2339_74.n3 a_2339_74.t3 155.847
R11 a_2339_74.n12 a_2339_74.n11 152
R12 a_2339_74.n7 a_2339_74.n0 152
R13 a_2339_74.n3 a_2339_74.n2 53.3701
R14 a_2339_74.n8 a_2339_74.n7 41.1312
R15 a_2339_74.n14 a_2339_74.t2 35.1791
R16 a_2339_74.t0 a_2339_74.n14 35.1791
R17 a_2339_74.n5 a_2339_74.n4 30.8485
R18 a_2339_74.n13 a_2339_74.n12 28.7035
R19 a_2339_74.n6 a_2339_74.n5 26.9925
R20 a_2339_74.n7 a_2339_74.n6 16.7098
R21 a_2339_74.n12 a_2339_74.n0 13.1884
R22 a_2339_74.n11 a_2339_74.n10 11.5685
R23 a_2339_74.n4 a_2339_74.n3 3.8565
R24 a_2339_74.n11 a_2339_74.n8 2.57117
R25 VGND.n38 VGND.t1 285.514
R26 VGND.n3 VGND.t4 268.467
R27 VGND.n64 VGND.t3 246.528
R28 VGND.n51 VGND.n50 213.161
R29 VGND.n31 VGND.n30 199.982
R30 VGND.n16 VGND.n13 185
R31 VGND.n18 VGND.n17 185
R32 VGND.n15 VGND.t5 169.025
R33 VGND.n24 VGND.t9 167.998
R34 VGND.n17 VGND.n16 98.9194
R35 VGND.n30 VGND.t10 55.7148
R36 VGND.n30 VGND.t2 55.7148
R37 VGND.n25 VGND.n11 36.1417
R38 VGND.n29 VGND.n11 36.1417
R39 VGND.n32 VGND.n9 36.1417
R40 VGND.n36 VGND.n9 36.1417
R41 VGND.n37 VGND.n36 36.1417
R42 VGND.n39 VGND.n37 36.1417
R43 VGND.n44 VGND.n43 36.1417
R44 VGND.n45 VGND.n44 36.1417
R45 VGND.n45 VGND.n5 36.1417
R46 VGND.n49 VGND.n5 36.1417
R47 VGND.n53 VGND.n52 36.1417
R48 VGND.n57 VGND.n56 36.1417
R49 VGND.n58 VGND.n57 36.1417
R50 VGND.n58 VGND.n1 36.1417
R51 VGND.n62 VGND.n1 36.1417
R52 VGND.n63 VGND.n62 36.1417
R53 VGND.n43 VGND.n7 35.6473
R54 VGND.n24 VGND.n23 26.7299
R55 VGND.n18 VGND.n15 26.5843
R56 VGND.n25 VGND.n24 25.977
R57 VGND.n23 VGND.n13 25.1572
R58 VGND.n64 VGND.n63 24.4711
R59 VGND.n17 VGND.t7 22.7032
R60 VGND.n16 VGND.t6 22.7032
R61 VGND.n50 VGND.t8 22.7032
R62 VGND.n50 VGND.t0 22.7032
R63 VGND.n32 VGND.n31 22.5887
R64 VGND.n31 VGND.n29 16.5652
R65 VGND.n39 VGND.n38 16.3142
R66 VGND.n52 VGND.n51 11.6711
R67 VGND.n56 VGND.n3 9.41227
R68 VGND.n63 VGND.n0 9.3005
R69 VGND.n62 VGND.n61 9.3005
R70 VGND.n60 VGND.n1 9.3005
R71 VGND.n59 VGND.n58 9.3005
R72 VGND.n57 VGND.n2 9.3005
R73 VGND.n56 VGND.n55 9.3005
R74 VGND.n54 VGND.n53 9.3005
R75 VGND.n52 VGND.n4 9.3005
R76 VGND.n49 VGND.n48 9.3005
R77 VGND.n47 VGND.n5 9.3005
R78 VGND.n46 VGND.n45 9.3005
R79 VGND.n44 VGND.n6 9.3005
R80 VGND.n43 VGND.n42 9.3005
R81 VGND.n41 VGND.n7 9.3005
R82 VGND.n40 VGND.n39 9.3005
R83 VGND.n37 VGND.n8 9.3005
R84 VGND.n36 VGND.n35 9.3005
R85 VGND.n34 VGND.n9 9.3005
R86 VGND.n33 VGND.n32 9.3005
R87 VGND.n31 VGND.n10 9.3005
R88 VGND.n29 VGND.n28 9.3005
R89 VGND.n27 VGND.n11 9.3005
R90 VGND.n26 VGND.n25 9.3005
R91 VGND.n24 VGND.n12 9.3005
R92 VGND.n19 VGND.n14 9.3005
R93 VGND.n21 VGND.n20 9.3005
R94 VGND.n23 VGND.n22 9.3005
R95 VGND.n20 VGND.n19 7.27151
R96 VGND.n65 VGND.n64 7.19894
R97 VGND.n51 VGND.n49 5.64756
R98 VGND.n38 VGND.n7 4.00858
R99 VGND.n15 VGND.n14 2.34593
R100 VGND.n53 VGND.n3 1.88285
R101 VGND.n20 VGND.n13 1.06085
R102 VGND.n19 VGND.n18 0.909376
R103 VGND VGND.n65 0.156997
R104 VGND.n65 VGND.n0 0.150766
R105 VGND.n21 VGND.n14 0.122949
R106 VGND.n22 VGND.n21 0.122949
R107 VGND.n22 VGND.n12 0.122949
R108 VGND.n26 VGND.n12 0.122949
R109 VGND.n27 VGND.n26 0.122949
R110 VGND.n28 VGND.n27 0.122949
R111 VGND.n28 VGND.n10 0.122949
R112 VGND.n33 VGND.n10 0.122949
R113 VGND.n34 VGND.n33 0.122949
R114 VGND.n35 VGND.n34 0.122949
R115 VGND.n35 VGND.n8 0.122949
R116 VGND.n40 VGND.n8 0.122949
R117 VGND.n41 VGND.n40 0.122949
R118 VGND.n42 VGND.n41 0.122949
R119 VGND.n42 VGND.n6 0.122949
R120 VGND.n46 VGND.n6 0.122949
R121 VGND.n47 VGND.n46 0.122949
R122 VGND.n48 VGND.n47 0.122949
R123 VGND.n48 VGND.n4 0.122949
R124 VGND.n54 VGND.n4 0.122949
R125 VGND.n55 VGND.n54 0.122949
R126 VGND.n55 VGND.n2 0.122949
R127 VGND.n59 VGND.n2 0.122949
R128 VGND.n60 VGND.n59 0.122949
R129 VGND.n61 VGND.n60 0.122949
R130 VGND.n61 VGND.n0 0.122949
R131 Q.n1 Q.n0 265.611
R132 Q.n3 Q.t1 242.561
R133 Q.n1 Q.t5 237.27
R134 Q.n3 Q.n2 99.7039
R135 Q.n0 Q.t4 26.3844
R136 Q.n0 Q.t3 26.3844
R137 Q.n2 Q.t0 22.7032
R138 Q.n2 Q.t2 22.7032
R139 Q Q.n1 22.4539
R140 Q Q.n3 20.4086
R141 VNB.n0 VNB 22277.2
R142 VNB VNB.n1 19861.1
R143 VNB.n1 VNB.t14 2806.3
R144 VNB.t3 VNB.t15 2459.84
R145 VNB.t1 VNB.t8 2448.29
R146 VNB.t6 VNB.n0 2432.22
R147 VNB.t11 VNB.t12 2402.1
R148 VNB.t17 VNB.t13 2298.16
R149 VNB.t5 VNB.t7 2286.61
R150 VNB.t15 VNB.t11 1986.35
R151 VNB.t14 VNB.t17 1893.96
R152 VNB.t0 VNB.t18 1813.12
R153 VNB.t4 VNB.t16 1247.24
R154 VNB.t18 VNB.t5 1189.5
R155 VNB.t2 VNB.t6 1161.11
R156 VNB.t7 VNB 1143.31
R157 VNB.n0 VNB.t4 1027.82
R158 VNB.t12 VNB.t10 993.177
R159 VNB.t13 VNB.t1 993.177
R160 VNB.t8 VNB.t9 993.177
R161 VNB.t9 VNB.t0 900.788
R162 VNB.t16 VNB.t3 831.496
R163 VNB.n1 VNB.t2 59.3797
R164 a_2003_48.n2 a_2003_48.n0 666.581
R165 a_2003_48.n1 a_2003_48.t3 359.358
R166 a_2003_48.t0 a_2003_48.n2 314.733
R167 a_2003_48.n1 a_2003_48.t4 231.361
R168 a_2003_48.n2 a_2003_48.n1 226.166
R169 a_2003_48.n0 a_2003_48.t1 110.227
R170 a_2003_48.n0 a_2003_48.t2 70.3576
R171 a_1982_508.t0 a_1982_508.t1 126.644
R172 VPWR.n43 VPWR.n11 660.663
R173 VPWR.n30 VPWR.n29 607.497
R174 VPWR.n57 VPWR.n4 605.946
R175 VPWR.n51 VPWR.n7 604.976
R176 VPWR.n27 VPWR.n17 355.945
R177 VPWR.n20 VPWR.t10 353.757
R178 VPWR.n21 VPWR.t9 352.005
R179 VPWR.n66 VPWR.n65 292.5
R180 VPWR.n64 VPWR.n63 292.5
R181 VPWR.n37 VPWR.t1 287.534
R182 VPWR.n17 VPWR.t11 262.885
R183 VPWR.n19 VPWR.n18 242.994
R184 VPWR.n65 VPWR.n64 190.845
R185 VPWR.n29 VPWR.t7 140.714
R186 VPWR.n11 VPWR.t5 114.918
R187 VPWR.n11 VPWR.t0 114.918
R188 VPWR.n29 VPWR.t15 110.227
R189 VPWR.n4 VPWR.t14 83.1099
R190 VPWR.n65 VPWR.t3 61.563
R191 VPWR.n18 VPWR.t12 55.1136
R192 VPWR.n17 VPWR.t2 51.8752
R193 VPWR.n64 VPWR.t4 46.1724
R194 VPWR.n4 VPWR.t6 46.1724
R195 VPWR.n58 VPWR.n2 36.1417
R196 VPWR.n62 VPWR.n2 36.1417
R197 VPWR.n52 VPWR.n5 36.1417
R198 VPWR.n56 VPWR.n5 36.1417
R199 VPWR.n45 VPWR.n44 36.1417
R200 VPWR.n45 VPWR.n8 36.1417
R201 VPWR.n49 VPWR.n8 36.1417
R202 VPWR.n50 VPWR.n49 36.1417
R203 VPWR.n35 VPWR.n14 36.1417
R204 VPWR.n36 VPWR.n35 36.1417
R205 VPWR.n38 VPWR.n36 36.1417
R206 VPWR.n42 VPWR.n12 36.1417
R207 VPWR.n31 VPWR.n28 36.1417
R208 VPWR.n58 VPWR.n57 34.2593
R209 VPWR.n38 VPWR.n37 32.377
R210 VPWR.n22 VPWR.n21 31.2476
R211 VPWR.n43 VPWR.n42 30.1181
R212 VPWR.n26 VPWR.n19 29.7417
R213 VPWR.n18 VPWR.t8 29.6087
R214 VPWR.n28 VPWR.n27 27.8593
R215 VPWR.n7 VPWR.t16 26.3844
R216 VPWR.n7 VPWR.t13 26.3844
R217 VPWR.n27 VPWR.n26 25.6005
R218 VPWR.n22 VPWR.n19 23.7181
R219 VPWR.n44 VPWR.n43 15.8123
R220 VPWR.n57 VPWR.n56 13.177
R221 VPWR.n52 VPWR.n51 10.9181
R222 VPWR.n30 VPWR.n14 10.9181
R223 VPWR.n63 VPWR.n62 10.6332
R224 VPWR.n23 VPWR.n22 9.3005
R225 VPWR.n24 VPWR.n19 9.3005
R226 VPWR.n26 VPWR.n25 9.3005
R227 VPWR.n27 VPWR.n16 9.3005
R228 VPWR.n28 VPWR.n15 9.3005
R229 VPWR.n32 VPWR.n31 9.3005
R230 VPWR.n33 VPWR.n14 9.3005
R231 VPWR.n35 VPWR.n34 9.3005
R232 VPWR.n36 VPWR.n13 9.3005
R233 VPWR.n39 VPWR.n38 9.3005
R234 VPWR.n40 VPWR.n12 9.3005
R235 VPWR.n42 VPWR.n41 9.3005
R236 VPWR.n43 VPWR.n10 9.3005
R237 VPWR.n44 VPWR.n9 9.3005
R238 VPWR.n46 VPWR.n45 9.3005
R239 VPWR.n47 VPWR.n8 9.3005
R240 VPWR.n49 VPWR.n48 9.3005
R241 VPWR.n50 VPWR.n6 9.3005
R242 VPWR.n53 VPWR.n52 9.3005
R243 VPWR.n54 VPWR.n5 9.3005
R244 VPWR.n56 VPWR.n55 9.3005
R245 VPWR.n57 VPWR.n3 9.3005
R246 VPWR.n59 VPWR.n58 9.3005
R247 VPWR.n60 VPWR.n2 9.3005
R248 VPWR.n62 VPWR.n61 9.3005
R249 VPWR.n1 VPWR.n0 9.3005
R250 VPWR.n67 VPWR.n66 8.20125
R251 VPWR.n21 VPWR.n20 6.54868
R252 VPWR.n66 VPWR.n1 5.0248
R253 VPWR.n37 VPWR.n12 3.76521
R254 VPWR.n63 VPWR.n1 2.39302
R255 VPWR.n23 VPWR.n20 0.651178
R256 VPWR.n51 VPWR.n50 0.376971
R257 VPWR.n31 VPWR.n30 0.376971
R258 VPWR VPWR.n67 0.160743
R259 VPWR.n67 VPWR.n0 0.147068
R260 VPWR.n24 VPWR.n23 0.122949
R261 VPWR.n25 VPWR.n24 0.122949
R262 VPWR.n25 VPWR.n16 0.122949
R263 VPWR.n16 VPWR.n15 0.122949
R264 VPWR.n32 VPWR.n15 0.122949
R265 VPWR.n33 VPWR.n32 0.122949
R266 VPWR.n34 VPWR.n33 0.122949
R267 VPWR.n34 VPWR.n13 0.122949
R268 VPWR.n39 VPWR.n13 0.122949
R269 VPWR.n40 VPWR.n39 0.122949
R270 VPWR.n41 VPWR.n40 0.122949
R271 VPWR.n41 VPWR.n10 0.122949
R272 VPWR.n10 VPWR.n9 0.122949
R273 VPWR.n46 VPWR.n9 0.122949
R274 VPWR.n47 VPWR.n46 0.122949
R275 VPWR.n48 VPWR.n47 0.122949
R276 VPWR.n48 VPWR.n6 0.122949
R277 VPWR.n53 VPWR.n6 0.122949
R278 VPWR.n54 VPWR.n53 0.122949
R279 VPWR.n55 VPWR.n54 0.122949
R280 VPWR.n55 VPWR.n3 0.122949
R281 VPWR.n59 VPWR.n3 0.122949
R282 VPWR.n60 VPWR.n59 0.122949
R283 VPWR.n61 VPWR.n60 0.122949
R284 VPWR.n61 VPWR.n0 0.122949
R285 VPB.t5 VPB.t6 572.043
R286 VPB.t22 VPB.t7 531.183
R287 VPB.t20 VPB.t18 531.183
R288 VPB.t8 VPB.t1 515.861
R289 VPB.t13 VPB.t14 459.678
R290 VPB.t17 VPB.t19 362.635
R291 VPB.t11 VPB.t21 349.866
R292 VPB.t0 VPB.t8 326.882
R293 VPB.t9 VPB.t20 291.13
R294 VPB.t15 VPB.t3 288.575
R295 VPB.t2 VPB.t9 275.807
R296 VPB.t16 VPB.t12 273.253
R297 VPB.t21 VPB.t15 273.253
R298 VPB VPB.t5 257.93
R299 VPB.t7 VPB.t4 255.376
R300 VPB.t1 VPB.t17 229.839
R301 VPB.t12 VPB.t13 229.839
R302 VPB.t3 VPB.t16 229.839
R303 VPB.t18 VPB.t22 229.839
R304 VPB.t10 VPB.t2 229.839
R305 VPB.t19 VPB.t11 214.517
R306 VPB.t6 VPB.t10 214.517
R307 VPB.t4 VPB.t0 199.195
R308 a_1745_74.n5 a_1745_74.n4 752.188
R309 a_1745_74.n2 a_1745_74.t3 407.022
R310 a_1745_74.n4 a_1745_74.t0 388.582
R311 a_1745_74.n0 a_1745_74.t5 298.841
R312 a_1745_74.t1 a_1745_74.n5 275.111
R313 a_1745_74.n4 a_1745_74.n3 252.142
R314 a_1745_74.n2 a_1745_74.n1 175.405
R315 a_1745_74.n0 a_1745_74.t6 163.881
R316 a_1745_74.n1 a_1745_74.t4 142.994
R317 a_1745_74.n5 a_1745_74.t2 115.278
R318 a_1745_74.n3 a_1745_74.t7 112.799
R319 a_1745_74.n1 a_1745_74.n0 89.9738
R320 a_1745_74.n3 a_1745_74.n2 42.1062
R321 RESET_B.n0 RESET_B.t3 415.197
R322 RESET_B.n1 RESET_B.t2 390.421
R323 RESET_B.n3 RESET_B.n2 380.274
R324 RESET_B.n4 RESET_B.n1 220.061
R325 RESET_B.n0 RESET_B.t0 192.673
R326 RESET_B.n4 RESET_B.n3 163.627
R327 RESET_B RESET_B.n0 163.286
R328 RESET_B.n1 RESET_B.t4 149.689
R329 RESET_B.n3 RESET_B.t1 129.633
R330 RESET_B RESET_B.n4 2.42441
R331 SCD.n1 SCD.t0 289.2
R332 SCD.n2 SCD.t1 187.178
R333 SCD.n1 SCD.n0 152
R334 SCD.n3 SCD.n2 152
R335 SCD.n2 SCD.n1 49.6611
R336 SCD.n3 SCD.n0 13.1884
R337 SCD.n0 SCD 0.970197
R338 SCD SCD.n3 0.194439
R339 a_572_81.t0 a_572_81.t1 68.5719
R340 a_225_81.n0 a_225_81.t1 561.649
R341 a_225_81.n0 a_225_81.t2 40.0005
R342 a_225_81.t0 a_225_81.n0 40.0005
R343 a_1367_112.n2 a_1367_112.n0 264.161
R344 a_1367_112.n3 a_1367_112.n2 257.245
R345 a_1367_112.n0 a_1367_112.t4 245.048
R346 a_1367_112.n0 a_1367_112.t5 185.869
R347 a_1367_112.n2 a_1367_112.n1 185
R348 a_1367_112.n1 a_1367_112.t0 31.0986
R349 a_1367_112.n3 a_1367_112.t3 29.5505
R350 a_1367_112.t1 a_1367_112.n3 29.5505
R351 a_1367_112.n1 a_1367_112.t2 26.2505
R352 a_1034_74.t1 a_1034_74.n4 823.63
R353 a_1034_74.n0 a_1034_74.t3 442.808
R354 a_1034_74.n0 a_1034_74.t4 374.731
R355 a_1034_74.n3 a_1034_74.n2 326.445
R356 a_1034_74.n1 a_1034_74.n0 322.88
R357 a_1034_74.n3 a_1034_74.t2 202.708
R358 a_1034_74.n4 a_1034_74.n3 172.559
R359 a_1034_74.n1 a_1034_74.t0 131.226
R360 a_1034_74.n4 a_1034_74.n1 47.8405
R361 a_415_81.n1 a_415_81.t0 657.298
R362 a_415_81.n1 a_415_81.t5 386.289
R363 a_415_81.n3 a_415_81.n0 374.014
R364 a_415_81.n0 a_415_81.n2 361.589
R365 a_415_81.n0 a_415_81.t4 353.688
R366 a_415_81.n0 a_415_81.n1 133.619
R367 a_415_81.n2 a_415_81.t6 121.43
R368 a_415_81.n2 a_415_81.t1 60.0005
R369 a_415_81.t2 a_415_81.n3 46.1724
R370 a_415_81.n3 a_415_81.t3 46.1724
R371 a_27_74.n1 a_27_74.t3 477.228
R372 a_27_74.n0 a_27_74.t2 418.296
R373 a_27_74.t0 a_27_74.n1 368.841
R374 a_27_74.n0 a_27_74.t1 243.177
R375 a_27_74.n1 a_27_74.n0 60.5666
R376 a_312_81.t0 a_312_81.t1 104.287
R377 SCE SCE.t2 420.082
R378 SCE.n4 SCE.t0 298.695
R379 SCE.n2 SCE.t3 262.276
R380 SCE.n4 SCE.t1 236.716
R381 SCE.n2 SCE.n1 152
R382 SCE.n3 SCE.n0 152
R383 SCE.n6 SCE.n5 152
R384 SCE.n3 SCE.n2 49.6611
R385 SCE.n5 SCE.n3 49.6611
R386 SCE.n5 SCE.n4 38.7066
R387 SCE.n6 SCE.n0 12.615
R388 SCE.n1 SCE 12.4295
R389 SCE.n1 SCE 5.38021
R390 SCE SCE.n6 5.0092
R391 SCE SCE.n0 0.186007
R392 CLK.n0 CLK.t1 250.909
R393 CLK.n0 CLK.t0 170.016
R394 CLK.n1 CLK.n0 118.308
R395 CLK.n1 CLK 13.6005
R396 CLK CLK.n1 3.29747
R397 a_855_368.n1 a_855_368.t3 1018.09
R398 a_855_368.t1 a_855_368.n5 889.902
R399 a_855_368.n2 a_855_368.n1 854.747
R400 a_855_368.t3 a_855_368.n0 668.374
R401 a_855_368.n4 a_855_368.t4 279.024
R402 a_855_368.n2 a_855_368.t2 247.428
R403 a_855_368.n5 a_855_368.t0 191.552
R404 a_855_368.n1 a_855_368.t5 182.625
R405 a_855_368.n3 a_855_368.t6 157.161
R406 a_855_368.n5 a_855_368.n4 152
R407 a_855_368.n3 a_855_368.n2 107.647
R408 a_855_368.n4 a_855_368.n3 20.449
R409 a_514_464.t0 a_514_464.t1 120.047
R410 D.n0 D.t0 411.139
R411 D D.n0 161.565
R412 D.n0 D.t1 124.617
R413 a_340_464.t0 a_340_464.t1 83.1099
R414 a_1342_463.t0 a_1342_463.t1 112.572
R415 a_2141_74.t0 a_2141_74.t1 60.0005
C0 VPWR RESET_B 0.367027f
C1 VPWR Q 0.425582f
C2 RESET_B Q 4.24e-19
C3 D RESET_B 1.06e-19
C4 VPWR D 0.013211f
C5 RESET_B VPB 0.37366f
C6 VPB Q 0.01534f
C7 VPWR VPB 0.437056f
C8 D VPB 0.054783f
C9 RESET_B a_1233_138# 0.241243f
C10 VPWR a_1233_138# 0.182081f
C11 a_1233_138# VPB 0.089295f
C12 VGND Q 0.390302f
C13 VPWR VGND 0.13085f
C14 VPWR SCD 0.014715f
C15 CLK RESET_B 0.071236f
C16 RESET_B VGND 0.19764f
C17 SCD RESET_B 0.100666f
C18 CLK VPWR 0.010458f
C19 D VGND 0.010334f
C20 SCE RESET_B 1.16e-19
C21 VPWR SCE 0.045732f
C22 D SCD 0.005546f
C23 SCE D 0.157424f
C24 VPB VGND 0.024108f
C25 SCD VPB 0.074674f
C26 CLK VPB 0.051401f
C27 SCE VPB 0.204602f
C28 RESET_B a_1319_138# 6.47e-19
C29 a_1233_138# VGND 0.018185f
C30 SCE a_1233_138# 2.96e-21
C31 a_1233_138# a_1319_138# 0.005862f
C32 SCD VGND 0.005743f
C33 CLK VGND 0.028423f
C34 SCE VGND 0.026623f
C35 SCE SCD 0.07669f
C36 CLK SCE 1.39e-19
C37 a_1319_138# VGND 8.94e-19
C38 Q VNB 0.05796f
C39 VGND VNB 1.72563f
C40 VPWR VNB 1.34198f
C41 CLK VNB 0.162749f
C42 RESET_B VNB 0.412995f
C43 SCD VNB 0.11682f
C44 D VNB 0.153917f
C45 SCE VNB 0.387895f
C46 VPB VNB 3.42518f
C47 a_1233_138# VNB 0.144755f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrtp_2 VNB VPB RESET_B VPWR VGND D SCE SCD CLK Q
X0 a_1242_457.t3 a_855_368.t2 a_390_81.t5 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1 a_547_81.t1 SCE.t0 a_390_81.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.13335 ps=1.055 w=0.42 l=0.15
X2 VGND.t8 RESET_B.t0 a_1432_138.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.367875 pd=1.845 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 a_2492_392.t0 a_1824_74# VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.1914 ps=1.435 w=1 l=0.15
X4 a_2078_74.t1 a_855_368.t3 a_1824_74# VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.2752 ps=1.86 w=0.42 l=0.15
X5 a_312_81.t0 a_27_74.t2 a_225_81.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X6 VGND.t3 SCE.t1 a_27_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X7 a_1034_368.t1 a_855_368.t4 VGND.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 VPWR.t10 SCE.t2 a_27_74.t0 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.3104 pd=1.61 as=0.1888 ps=1.87 w=0.64 l=0.15
X9 a_2242_74.t0 RESET_B.t1 VGND.t7 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VPWR.t5 CLK.t0 a_855_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X11 a_514_464.t0 a_27_74.t3 a_390_81.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1248 pd=1.03 as=0.096 ps=0.94 w=0.64 l=0.15
X12 a_1034_368.t0 a_855_368.t5 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t6 RESET_B.t2 a_225_81.t0 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.08295 ps=0.815 w=0.42 l=0.15
X14 a_390_81.t2 D.t0 a_340_464.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 VPWR.t9 SCD.t0 a_514_464.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.1248 ps=1.03 w=0.64 l=0.15
X16 VPWR.t0 a_1383_349# a_1332_457.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.138825 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_2082_446.t1 a_1824_74# a_2242_74.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 VPWR.t1 a_2082_446.t3 a_2037_508.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.12 as=0.0504 ps=0.66 w=0.42 l=0.15
X19 a_225_81.t2 SCD.t1 a_547_81.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.08295 pd=0.815 as=0.0504 ps=0.66 w=0.42 l=0.15
X20 a_1432_138.t0 a_1383_349# a_1354_138.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X21 VGND.t4 a_2082_446.t4 a_2078_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 Q.t2 a_2492_392.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X23 VPWR.t6 a_1824_74# a_2082_446.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1914 pd=1.435 as=0.063 ps=0.72 w=0.42 l=0.15
X24 VGND.t2 CLK.t1 a_855_368.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X25 a_1354_138.t1 a_1034_368.t2 a_1242_457.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X26 a_390_81.t1 D.t1 a_312_81.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.13335 pd=1.055 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 a_2082_446.t0 RESET_B.t3 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.147 ps=1.12 w=0.42 l=0.15
X28 a_1824_74# a_1034_368.t3 a_1383_349# VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2752 pd=1.86 as=0.13135 ps=1.095 w=0.74 l=0.15
X29 a_340_464.t1 SCE.t3 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.3104 ps=1.61 w=0.64 l=0.15
X30 a_1242_457.t4 RESET_B.t4 VPWR.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.138825 ps=1.16 w=0.42 l=0.15
X31 a_1332_457.t1 a_855_368.t6 a_1242_457.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X32 VGND.t1 a_2492_392.t2 Q.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 Q.t0 a_2492_392.t3 VPWR.t12 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X34 a_1242_457.t0 a_1034_368.t4 a_390_81.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X35 a_390_81.t6 RESET_B.t5 VPWR.t4 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1344 ps=1.06 w=0.64 l=0.15
X36 a_2037_508.t1 a_1034_368.t5 a_1824_74# VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.223625 ps=1.83 w=0.42 l=0.15
R0 a_855_368.n1 a_855_368.n0 1052.1
R1 a_855_368.t1 a_855_368.n5 886.754
R2 a_855_368.n2 a_855_368.n1 822.614
R3 a_855_368.n0 a_855_368.t3 794.497
R4 a_855_368.n2 a_855_368.t2 297.233
R5 a_855_368.n4 a_855_368.t5 265.637
R6 a_855_368.n5 a_855_368.t0 194.052
R7 a_855_368.n1 a_855_368.t6 190.659
R8 a_855_368.n3 a_855_368.t4 173.228
R9 a_855_368.n5 a_855_368.n4 152
R10 a_855_368.n3 a_855_368.n2 99.6138
R11 a_855_368.n4 a_855_368.n3 20.449
R12 a_390_81.n1 a_390_81.t3 656.381
R13 a_390_81.n3 a_390_81.n0 374.014
R14 a_390_81.n1 a_390_81.t5 363.592
R15 a_390_81.n0 a_390_81.n2 360.33
R16 a_390_81.n0 a_390_81.t6 353.688
R17 a_390_81.n2 a_390_81.t1 140
R18 a_390_81.n0 a_390_81.n1 133.619
R19 a_390_81.n3 a_390_81.t4 46.1724
R20 a_390_81.t2 a_390_81.n3 46.1724
R21 a_390_81.n2 a_390_81.t0 41.4291
R22 a_1242_457.n3 a_1242_457.t4 669.607
R23 a_1242_457.n5 a_1242_457.n4 617.091
R24 a_1242_457.n6 a_1242_457.n5 296.56
R25 a_1242_457.n3 a_1242_457.n2 277.557
R26 a_1242_457.n2 a_1242_457.n1 221.738
R27 a_1242_457.n2 a_1242_457.n0 162.274
R28 a_1242_457.n4 a_1242_457.t2 70.3576
R29 a_1242_457.n4 a_1242_457.t0 70.3576
R30 a_1242_457.n6 a_1242_457.t3 60.0005
R31 a_1242_457.n5 a_1242_457.n3 52.7064
R32 a_1242_457.t1 a_1242_457.n6 40.0005
R33 VNB.n0 VNB 22589
R34 VNB VNB.n1 19848.9
R35 VNB.t12 VNB.t0 4573.23
R36 VNB.t3 VNB.t16 2529.13
R37 VNB.t15 VNB.t13 2321.26
R38 VNB.t11 VNB.t5 2286.61
R39 VNB.n1 VNB.t10 2261.11
R40 VNB.t4 VNB.t6 1813.12
R41 VNB.t10 VNB.n0 1796.67
R42 VNB.n1 VNB.t18 1489.76
R43 VNB.t16 VNB.t7 1258.79
R44 VNB.n0 VNB.t14 1235.7
R45 VNB.t9 VNB.t15 1154.86
R46 VNB.t13 VNB.t3 1154.86
R47 VNB.t5 VNB 1143.31
R48 VNB.t0 VNB.t1 993.177
R49 VNB.t8 VNB.t17 993.177
R50 VNB.t14 VNB.t8 900.788
R51 VNB.t18 VNB.t2 900.788
R52 VNB.t2 VNB.t9 900.788
R53 VNB.t7 VNB.t4 900.788
R54 VNB.t6 VNB.t11 900.788
R55 VNB.t17 VNB.t12 831.496
R56 VGND.n32 VGND.t8 294.558
R57 VGND.n3 VGND.t6 268.856
R58 VGND.n56 VGND.t3 246.528
R59 VGND.n24 VGND.n13 207.498
R60 VGND.n43 VGND.n6 206.333
R61 VGND.n16 VGND.t1 178.81
R62 VGND.n15 VGND.t0 171.77
R63 VGND.n13 VGND.t7 40.0005
R64 VGND.n13 VGND.t4 40.0005
R65 VGND.n20 VGND.n12 36.1417
R66 VGND.n26 VGND.n25 36.1417
R67 VGND.n26 VGND.n10 36.1417
R68 VGND.n30 VGND.n10 36.1417
R69 VGND.n31 VGND.n30 36.1417
R70 VGND.n37 VGND.n8 36.1417
R71 VGND.n38 VGND.n37 36.1417
R72 VGND.n39 VGND.n38 36.1417
R73 VGND.n39 VGND.n5 36.1417
R74 VGND.n45 VGND.n44 36.1417
R75 VGND.n49 VGND.n48 36.1417
R76 VGND.n50 VGND.n49 36.1417
R77 VGND.n50 VGND.n1 36.1417
R78 VGND.n54 VGND.n1 36.1417
R79 VGND.n55 VGND.n54 36.1417
R80 VGND.n6 VGND.t5 34.0546
R81 VGND.n43 VGND.n5 33.8829
R82 VGND.n25 VGND.n24 32.7534
R83 VGND.n18 VGND.n15 28.2358
R84 VGND.n33 VGND.n31 28.232
R85 VGND.n20 VGND.n19 25.977
R86 VGND.n56 VGND.n55 24.4711
R87 VGND.n6 VGND.t2 22.7032
R88 VGND.n19 VGND.n18 21.4593
R89 VGND.n32 VGND.n8 18.5008
R90 VGND.n24 VGND.n12 14.6829
R91 VGND.n44 VGND.n43 13.5534
R92 VGND.n55 VGND.n0 9.3005
R93 VGND.n54 VGND.n53 9.3005
R94 VGND.n52 VGND.n1 9.3005
R95 VGND.n51 VGND.n50 9.3005
R96 VGND.n49 VGND.n2 9.3005
R97 VGND.n48 VGND.n47 9.3005
R98 VGND.n46 VGND.n45 9.3005
R99 VGND.n44 VGND.n4 9.3005
R100 VGND.n43 VGND.n42 9.3005
R101 VGND.n41 VGND.n5 9.3005
R102 VGND.n40 VGND.n39 9.3005
R103 VGND.n38 VGND.n7 9.3005
R104 VGND.n37 VGND.n36 9.3005
R105 VGND.n35 VGND.n8 9.3005
R106 VGND.n34 VGND.n33 9.3005
R107 VGND.n31 VGND.n9 9.3005
R108 VGND.n30 VGND.n29 9.3005
R109 VGND.n28 VGND.n10 9.3005
R110 VGND.n27 VGND.n26 9.3005
R111 VGND.n25 VGND.n11 9.3005
R112 VGND.n24 VGND.n23 9.3005
R113 VGND.n22 VGND.n12 9.3005
R114 VGND.n21 VGND.n20 9.3005
R115 VGND.n19 VGND.n14 9.3005
R116 VGND.n18 VGND.n17 9.3005
R117 VGND.n48 VGND.n3 8.65932
R118 VGND.n57 VGND.n56 7.19894
R119 VGND.n16 VGND.n15 6.79022
R120 VGND.n45 VGND.n3 2.63579
R121 VGND.n33 VGND.n32 2.06919
R122 VGND.n17 VGND.n16 0.5771
R123 VGND VGND.n57 0.156997
R124 VGND.n57 VGND.n0 0.150766
R125 VGND.n17 VGND.n14 0.122949
R126 VGND.n21 VGND.n14 0.122949
R127 VGND.n22 VGND.n21 0.122949
R128 VGND.n23 VGND.n22 0.122949
R129 VGND.n23 VGND.n11 0.122949
R130 VGND.n27 VGND.n11 0.122949
R131 VGND.n28 VGND.n27 0.122949
R132 VGND.n29 VGND.n28 0.122949
R133 VGND.n29 VGND.n9 0.122949
R134 VGND.n34 VGND.n9 0.122949
R135 VGND.n35 VGND.n34 0.122949
R136 VGND.n36 VGND.n35 0.122949
R137 VGND.n36 VGND.n7 0.122949
R138 VGND.n40 VGND.n7 0.122949
R139 VGND.n41 VGND.n40 0.122949
R140 VGND.n42 VGND.n41 0.122949
R141 VGND.n42 VGND.n4 0.122949
R142 VGND.n46 VGND.n4 0.122949
R143 VGND.n47 VGND.n46 0.122949
R144 VGND.n47 VGND.n2 0.122949
R145 VGND.n51 VGND.n2 0.122949
R146 VGND.n52 VGND.n51 0.122949
R147 VGND.n53 VGND.n52 0.122949
R148 VGND.n53 VGND.n0 0.122949
R149 SCE SCE.t0 437.724
R150 SCE.n4 SCE.t1 298.695
R151 SCE.n2 SCE.t3 262.276
R152 SCE.n4 SCE.t2 236.716
R153 SCE.n2 SCE.n1 152
R154 SCE.n3 SCE.n0 152
R155 SCE.n6 SCE.n5 152
R156 SCE.n3 SCE.n2 49.6611
R157 SCE.n5 SCE.n3 49.6611
R158 SCE.n5 SCE.n4 38.7066
R159 SCE.n6 SCE.n0 12.615
R160 SCE.n1 SCE 12.4295
R161 SCE.n1 SCE 5.38021
R162 SCE SCE.n6 5.0092
R163 SCE SCE.n0 0.186007
R164 a_547_81.t0 a_547_81.t1 68.5719
R165 a_2492_392.t0 a_2492_392.n3 463.115
R166 a_2492_392.n1 a_2492_392.n0 240.197
R167 a_2492_392.n3 a_2492_392.t3 240.197
R168 a_2492_392.n1 a_2492_392.t2 190.006
R169 a_2492_392.n2 a_2492_392.t1 179.947
R170 a_2492_392.n2 a_2492_392.n1 54.0429
R171 a_2492_392.n3 a_2492_392.n2 11.6853
R172 VPB.t13 VPB.t6 1266.67
R173 VPB.t16 VPB.t15 572.043
R174 VPB.t11 VPB.t5 531.183
R175 VPB.t12 VPB.t3 531.183
R176 VPB.t9 VPB.t17 515.861
R177 VPB.t2 VPB.t0 434.14
R178 VPB.t1 VPB.t13 319.221
R179 VPB.t8 VPB.t9 298.791
R180 VPB.t14 VPB.t12 291.13
R181 VPB.t7 VPB.t14 275.807
R182 VPB VPB.t16 257.93
R183 VPB.t0 VPB.t8 229.839
R184 VPB.t5 VPB.t10 229.839
R185 VPB.t3 VPB.t11 229.839
R186 VPB.t4 VPB.t7 229.839
R187 VPB.t10 VPB.t1 214.517
R188 VPB.t15 VPB.t4 214.517
R189 VPB.t6 VPB.t2 199.195
R190 RESET_B.n0 RESET_B.t1 446.985
R191 RESET_B.n1 RESET_B.t2 391.882
R192 RESET_B.n2 RESET_B.t0 294.021
R193 RESET_B.n3 RESET_B.n2 224.825
R194 RESET_B.n3 RESET_B.n1 220.489
R195 RESET_B.n0 RESET_B.t3 177.269
R196 RESET_B RESET_B.n0 162.704
R197 RESET_B.n1 RESET_B.t5 149.689
R198 RESET_B.n2 RESET_B.t4 116.532
R199 RESET_B RESET_B.n3 2.42441
R200 a_1432_138.t0 a_1432_138.t1 68.5719
R201 VPWR.n37 VPWR.n11 684.432
R202 VPWR.n51 VPWR.n4 605.946
R203 VPWR.n45 VPWR.n7 604.976
R204 VPWR.n25 VPWR.n24 585
R205 VPWR.n23 VPWR.n22 585
R206 VPWR.n60 VPWR.n59 292.5
R207 VPWR.n58 VPWR.n57 292.5
R208 VPWR.n18 VPWR.t12 255.73
R209 VPWR.n17 VPWR.n16 223.417
R210 VPWR.n59 VPWR.n58 190.845
R211 VPWR.n24 VPWR.n23 164.167
R212 VPWR.n16 VPWR.t6 117.725
R213 VPWR.n11 VPWR.t3 112.572
R214 VPWR.n11 VPWR.t0 110.227
R215 VPWR.n23 VPWR.t2 93.81
R216 VPWR.n4 VPWR.t4 83.1099
R217 VPWR.n24 VPWR.t1 70.3576
R218 VPWR.n59 VPWR.t10 61.563
R219 VPWR.n58 VPWR.t11 46.1724
R220 VPWR.n4 VPWR.t9 46.1724
R221 VPWR.n16 VPWR.t7 38.5539
R222 VPWR.n52 VPWR.n2 36.1417
R223 VPWR.n56 VPWR.n2 36.1417
R224 VPWR.n46 VPWR.n5 36.1417
R225 VPWR.n50 VPWR.n5 36.1417
R226 VPWR.n39 VPWR.n38 36.1417
R227 VPWR.n39 VPWR.n8 36.1417
R228 VPWR.n43 VPWR.n8 36.1417
R229 VPWR.n44 VPWR.n43 36.1417
R230 VPWR.n30 VPWR.n14 36.1417
R231 VPWR.n31 VPWR.n30 36.1417
R232 VPWR.n32 VPWR.n31 36.1417
R233 VPWR.n21 VPWR.n20 36.1417
R234 VPWR.n52 VPWR.n51 34.2593
R235 VPWR.n37 VPWR.n36 32.7534
R236 VPWR.n7 VPWR.t8 26.3844
R237 VPWR.n7 VPWR.t5 26.3844
R238 VPWR.n36 VPWR.n12 24.8476
R239 VPWR.n32 VPWR.n12 22.5887
R240 VPWR.n25 VPWR.n14 21.1543
R241 VPWR.n38 VPWR.n37 14.3064
R242 VPWR.n20 VPWR.n17 13.9299
R243 VPWR.n51 VPWR.n50 13.177
R244 VPWR.n46 VPWR.n45 10.9181
R245 VPWR.n57 VPWR.n56 10.6332
R246 VPWR.n20 VPWR.n19 9.3005
R247 VPWR.n21 VPWR.n15 9.3005
R248 VPWR.n27 VPWR.n26 9.3005
R249 VPWR.n28 VPWR.n14 9.3005
R250 VPWR.n30 VPWR.n29 9.3005
R251 VPWR.n31 VPWR.n13 9.3005
R252 VPWR.n33 VPWR.n32 9.3005
R253 VPWR.n34 VPWR.n12 9.3005
R254 VPWR.n36 VPWR.n35 9.3005
R255 VPWR.n37 VPWR.n10 9.3005
R256 VPWR.n38 VPWR.n9 9.3005
R257 VPWR.n40 VPWR.n39 9.3005
R258 VPWR.n41 VPWR.n8 9.3005
R259 VPWR.n43 VPWR.n42 9.3005
R260 VPWR.n44 VPWR.n6 9.3005
R261 VPWR.n47 VPWR.n46 9.3005
R262 VPWR.n48 VPWR.n5 9.3005
R263 VPWR.n50 VPWR.n49 9.3005
R264 VPWR.n51 VPWR.n3 9.3005
R265 VPWR.n53 VPWR.n52 9.3005
R266 VPWR.n54 VPWR.n2 9.3005
R267 VPWR.n56 VPWR.n55 9.3005
R268 VPWR.n1 VPWR.n0 9.3005
R269 VPWR.n61 VPWR.n60 8.20125
R270 VPWR.n18 VPWR.n17 7.21174
R271 VPWR.n22 VPWR.n21 6.09548
R272 VPWR.n26 VPWR.n22 5.13919
R273 VPWR.n60 VPWR.n1 5.0248
R274 VPWR.n57 VPWR.n1 2.39302
R275 VPWR.n26 VPWR.n25 1.40196
R276 VPWR.n19 VPWR.n18 0.481592
R277 VPWR.n45 VPWR.n44 0.376971
R278 VPWR VPWR.n61 0.160743
R279 VPWR.n61 VPWR.n0 0.147068
R280 VPWR.n19 VPWR.n15 0.122949
R281 VPWR.n27 VPWR.n15 0.122949
R282 VPWR.n28 VPWR.n27 0.122949
R283 VPWR.n29 VPWR.n28 0.122949
R284 VPWR.n29 VPWR.n13 0.122949
R285 VPWR.n33 VPWR.n13 0.122949
R286 VPWR.n34 VPWR.n33 0.122949
R287 VPWR.n35 VPWR.n34 0.122949
R288 VPWR.n35 VPWR.n10 0.122949
R289 VPWR.n10 VPWR.n9 0.122949
R290 VPWR.n40 VPWR.n9 0.122949
R291 VPWR.n41 VPWR.n40 0.122949
R292 VPWR.n42 VPWR.n41 0.122949
R293 VPWR.n42 VPWR.n6 0.122949
R294 VPWR.n47 VPWR.n6 0.122949
R295 VPWR.n48 VPWR.n47 0.122949
R296 VPWR.n49 VPWR.n48 0.122949
R297 VPWR.n49 VPWR.n3 0.122949
R298 VPWR.n53 VPWR.n3 0.122949
R299 VPWR.n54 VPWR.n53 0.122949
R300 VPWR.n55 VPWR.n54 0.122949
R301 VPWR.n55 VPWR.n0 0.122949
R302 a_2078_74.t0 a_2078_74.t1 68.5719
R303 a_27_74.n1 a_27_74.t3 477.228
R304 a_27_74.n0 a_27_74.t2 418.296
R305 a_27_74.t0 a_27_74.n1 368.841
R306 a_27_74.n0 a_27_74.t1 243.177
R307 a_27_74.n1 a_27_74.n0 60.5666
R308 a_225_81.n0 a_225_81.t1 562.837
R309 a_225_81.n0 a_225_81.t2 72.8576
R310 a_225_81.t0 a_225_81.n0 40.0005
R311 a_312_81.t0 a_312_81.t1 68.5719
R312 a_1034_368.t0 a_1034_368.n3 822.225
R313 a_1034_368.n0 a_1034_368.t3 458.873
R314 a_1034_368.n1 a_1034_368.n0 355.43
R315 a_1034_368.n0 a_1034_368.t5 349.457
R316 a_1034_368.n2 a_1034_368.t2 343.007
R317 a_1034_368.n2 a_1034_368.t4 181.286
R318 a_1034_368.n3 a_1034_368.n2 171.589
R319 a_1034_368.n1 a_1034_368.t1 135.911
R320 a_1034_368.n3 a_1034_368.n1 50.4489
R321 a_2242_74.t0 a_2242_74.t1 60.0005
R322 CLK.n0 CLK.t0 250.909
R323 CLK.n0 CLK.t1 173.667
R324 CLK.n1 CLK.n0 117.234
R325 CLK.n1 CLK 13.6005
R326 CLK CLK.n1 3.29747
R327 a_514_464.t0 a_514_464.t1 120.047
R328 D.n0 D.t0 411.139
R329 D D.n0 161.565
R330 D.n0 D.t1 124.617
R331 a_340_464.t0 a_340_464.t1 83.1099
R332 SCD.n1 SCD.t1 302.053
R333 SCD.n0 SCD.t0 176.466
R334 SCD SCD.n0 153.358
R335 SCD.n2 SCD.n1 152
R336 SCD.n1 SCD.n0 49.6611
R337 SCD SCD.n2 11.8308
R338 SCD.n2 SCD 2.52171
R339 a_1332_457.t0 a_1332_457.t1 126.644
R340 a_2082_446.n2 a_2082_446.n1 649.308
R341 a_2082_446.t1 a_2082_446.n6 401.69
R342 a_2082_446.n5 a_2082_446.t4 273.252
R343 a_2082_446.n6 a_2082_446.n5 157.738
R344 a_2082_446.n3 a_2082_446.n2 152
R345 a_2082_446.n4 a_2082_446.n0 152
R346 a_2082_446.n3 a_2082_446.t3 133.834
R347 a_2082_446.n1 a_2082_446.t2 70.3576
R348 a_2082_446.n1 a_2082_446.t0 70.3576
R349 a_2082_446.n4 a_2082_446.n3 39.9712
R350 a_2082_446.n5 a_2082_446.n4 39.9712
R351 a_2082_446.n2 a_2082_446.n0 15.0074
R352 a_2082_446.n6 a_2082_446.n0 9.26947
R353 a_2037_508.t0 a_2037_508.t1 112.572
R354 a_1354_138.t0 a_1354_138.t1 68.5719
R355 Q Q.t0 268.443
R356 Q.n2 Q.n1 185
R357 Q.n1 Q.n0 185
R358 Q.n1 Q.t1 22.7032
R359 Q.n1 Q.t2 22.7032
R360 Q.n0 Q 12.6066
R361 Q Q.n2 9.50353
R362 Q.n2 Q 4.84898
R363 Q.n0 Q 1.74595
C0 CLK VGND 0.030215f
C1 VGND SCD 0.005176f
C2 SCE VGND 0.026018f
C3 CLK SCE 1.38e-19
C4 SCE SCD 0.078077f
C5 VGND a_1824_74# 0.177959f
C6 VGND a_1383_349# 0.037986f
C7 a_1824_74# a_1383_349# 0.070416f
C8 VPWR Q 0.22103f
C9 Q RESET_B 2.83e-19
C10 Q VPB 0.006542f
C11 VPWR RESET_B 0.374581f
C12 VPWR D 0.013211f
C13 VPWR VPB 0.424249f
C14 VPB RESET_B 0.359763f
C15 D RESET_B 1.06e-19
C16 D VPB 0.054783f
C17 VGND Q 0.164626f
C18 VPWR VGND 0.126168f
C19 VGND RESET_B 0.21106f
C20 VGND VPB 0.026073f
C21 D VGND 0.010379f
C22 CLK VPWR 0.010531f
C23 VPWR SCD 0.014553f
C24 CLK RESET_B 0.069335f
C25 SCD RESET_B 0.08917f
C26 CLK VPB 0.052356f
C27 VPWR SCE 0.045579f
C28 VPB SCD 0.074634f
C29 SCE RESET_B 1.16e-19
C30 D SCD 0.005234f
C31 SCE VPB 0.201965f
C32 SCE D 0.161738f
C33 Q a_1824_74# 8.48e-19
C34 VPWR a_1824_74# 0.150318f
C35 a_1824_74# RESET_B 0.194395f
C36 a_1824_74# VPB 0.172449f
C37 VPWR a_1383_349# 0.075526f
C38 RESET_B a_1383_349# 0.187204f
C39 VPB a_1383_349# 0.087272f
C40 Q VNB 0.030387f
C41 VGND VNB 1.70534f
C42 VPWR VNB 1.30653f
C43 CLK VNB 0.166579f
C44 RESET_B VNB 0.401299f
C45 SCD VNB 0.118151f
C46 D VNB 0.151214f
C47 SCE VNB 0.374606f
C48 VPB VNB 3.31981f
C49 a_1824_74# VNB 0.34925f
C50 a_1383_349# VNB 0.114432f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrtp_1 VNB VPB VPWR RESET_B VGND Q SCE CLK SCD D
X0 a_2399_424.t0 a_1745_74.t4 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.1595 ps=1.68 w=0.55 l=0.15
X1 a_1745_74.t2 a_855_368.t2 a_1367_92.t2 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.221475 pd=1.82 as=0.15 ps=1.3 w=1 l=0.15
X2 a_545_81.t0 SCE.t0 a_300_464.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.13125 ps=1.045 w=0.42 l=0.15
X3 a_1367_92.t1 a_1233_118# VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X4 VPWR.t4 a_1745_74.t5 a_1997_272.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.275 as=0.063 ps=0.72 w=0.42 l=0.15
X5 a_2399_424.t1 a_1745_74.t6 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1638 ps=1.275 w=0.84 l=0.15
X6 a_312_81.t0 a_27_88.t2 a_225_81.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7 a_1993_508.t1 a_1034_368.t2 a_1745_74.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.221475 ps=1.82 w=0.42 l=0.15
X8 a_1745_74.t0 a_1034_368.t3 a_1367_92.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.23435 pd=1.625 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 VGND.t3 CLK.t0 a_855_368.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 VGND.t0 SCE.t1 a_27_88.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X11 a_2135_74.t1 RESET_B.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.06405 ps=0.725 w=0.42 l=0.15
X12 VPWR.t0 SCE.t2 a_27_88.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.1888 ps=1.87 w=0.64 l=0.15
X13 Q.t1 a_2399_424.t2 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X14 VPWR.t2 CLK.t1 a_855_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X15 a_1233_118# RESET_B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.135875 ps=1.14 w=0.42 l=0.15
X16 a_1972_74.t1 a_855_368.t3 a_1745_74.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.23435 ps=1.625 w=0.42 l=0.15
X17 a_1034_368.t1 a_855_368.t4 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_1997_272.t0 a_1745_74.t7 a_2135_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 VPWR.t5 SCD.t0 a_538_464.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VGND.t5 RESET_B.t2 a_225_81.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.09765 ps=0.885 w=0.42 l=0.15
X21 a_300_464.t2 D.t0 a_216_464.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3328 pd=1.68 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 Q.t0 a_2399_424.t3 VGND.t2 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X23 a_225_81.t1 SCD.t1 a_545_81.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.09765 pd=0.885 as=0.0504 ps=0.66 w=0.42 l=0.15
X24 a_216_464.t0 SCE.t3 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X25 a_300_464.t1 D.t1 a_312_81.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.13125 pd=1.045 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 a_1397_118.t0 a_1367_92.t3 a_1319_118# VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 VGND.t6 a_1997_272.t2 a_1972_74.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_1034_368.t0 a_855_368.t5 VGND.t7 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10545 ps=1.025 w=0.74 l=0.15
X29 a_538_464.t0 a_27_88.t3 a_300_464.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.3328 ps=1.68 w=0.64 l=0.15
X30 a_1233_118# a_1034_368.t4 a_300_464.t6 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0763 pd=0.795 as=0.1239 ps=1.43 w=0.42 l=0.15
X31 VPWR.t9 a_1997_272.t3 a_1993_508.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 a_1233_118# a_855_368.t6 a_300_464.t5 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X33 a_300_464.t4 RESET_B.t3 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1344 ps=1.06 w=0.64 l=0.15
R0 a_1745_74.n5 a_1745_74.n4 737.106
R1 a_1745_74.n2 a_1745_74.t4 358.288
R2 a_1745_74.n1 a_1745_74.t6 324.012
R3 a_1745_74.t2 a_1745_74.n5 295.317
R4 a_1745_74.n4 a_1745_74.n3 268.769
R5 a_1745_74.n1 a_1745_74.t5 238.858
R6 a_1745_74.n0 a_1745_74.t0 229.153
R7 a_1745_74.n4 a_1745_74.n0 217.151
R8 a_1745_74.n2 a_1745_74.n1 188.492
R9 a_1745_74.n3 a_1745_74.t7 174.25
R10 a_1745_74.n5 a_1745_74.t1 119.608
R11 a_1745_74.n0 a_1745_74.t3 40.0005
R12 a_1745_74.n3 a_1745_74.n2 13.146
R13 VGND.n3 VGND.t5 261.142
R14 VGND.n50 VGND.t0 250.213
R15 VGND.n12 VGND.t4 235.742
R16 VGND.n37 VGND.n36 213.161
R17 VGND.n18 VGND.n17 207.498
R18 VGND.n13 VGND.t2 177.618
R19 VGND.n17 VGND.t1 47.1434
R20 VGND.n17 VGND.t6 40.0005
R21 VGND.n16 VGND.n11 36.1417
R22 VGND.n19 VGND.n9 36.1417
R23 VGND.n23 VGND.n9 36.1417
R24 VGND.n24 VGND.n23 36.1417
R25 VGND.n25 VGND.n24 36.1417
R26 VGND.n30 VGND.n29 36.1417
R27 VGND.n31 VGND.n30 36.1417
R28 VGND.n31 VGND.n5 36.1417
R29 VGND.n35 VGND.n5 36.1417
R30 VGND.n39 VGND.n38 36.1417
R31 VGND.n43 VGND.n42 36.1417
R32 VGND.n44 VGND.n43 36.1417
R33 VGND.n44 VGND.n1 36.1417
R34 VGND.n48 VGND.n1 36.1417
R35 VGND.n49 VGND.n48 36.1417
R36 VGND.n29 VGND.n7 35.6473
R37 VGND.n19 VGND.n18 26.7299
R38 VGND.n50 VGND.n49 24.4711
R39 VGND.n36 VGND.t7 23.514
R40 VGND.n36 VGND.t3 22.7032
R41 VGND.n12 VGND.n11 21.8358
R42 VGND.n18 VGND.n16 20.7064
R43 VGND.n42 VGND.n3 20.3299
R44 VGND.n25 VGND.n7 20.3223
R45 VGND.n39 VGND.n3 15.8123
R46 VGND.n38 VGND.n37 11.6711
R47 VGND.n49 VGND.n0 9.3005
R48 VGND.n48 VGND.n47 9.3005
R49 VGND.n46 VGND.n1 9.3005
R50 VGND.n45 VGND.n44 9.3005
R51 VGND.n43 VGND.n2 9.3005
R52 VGND.n42 VGND.n41 9.3005
R53 VGND.n40 VGND.n39 9.3005
R54 VGND.n38 VGND.n4 9.3005
R55 VGND.n35 VGND.n34 9.3005
R56 VGND.n33 VGND.n5 9.3005
R57 VGND.n32 VGND.n31 9.3005
R58 VGND.n30 VGND.n6 9.3005
R59 VGND.n29 VGND.n28 9.3005
R60 VGND.n27 VGND.n7 9.3005
R61 VGND.n26 VGND.n25 9.3005
R62 VGND.n24 VGND.n8 9.3005
R63 VGND.n23 VGND.n22 9.3005
R64 VGND.n21 VGND.n9 9.3005
R65 VGND.n20 VGND.n19 9.3005
R66 VGND.n18 VGND.n10 9.3005
R67 VGND.n16 VGND.n15 9.3005
R68 VGND.n14 VGND.n11 9.3005
R69 VGND.n51 VGND.n50 7.19894
R70 VGND.n13 VGND.n12 6.82733
R71 VGND.n37 VGND.n35 5.64756
R72 VGND.n14 VGND.n13 0.530796
R73 VGND VGND.n51 0.156997
R74 VGND.n51 VGND.n0 0.150766
R75 VGND.n15 VGND.n14 0.122949
R76 VGND.n15 VGND.n10 0.122949
R77 VGND.n20 VGND.n10 0.122949
R78 VGND.n21 VGND.n20 0.122949
R79 VGND.n22 VGND.n21 0.122949
R80 VGND.n22 VGND.n8 0.122949
R81 VGND.n26 VGND.n8 0.122949
R82 VGND.n27 VGND.n26 0.122949
R83 VGND.n28 VGND.n27 0.122949
R84 VGND.n28 VGND.n6 0.122949
R85 VGND.n32 VGND.n6 0.122949
R86 VGND.n33 VGND.n32 0.122949
R87 VGND.n34 VGND.n33 0.122949
R88 VGND.n34 VGND.n4 0.122949
R89 VGND.n40 VGND.n4 0.122949
R90 VGND.n41 VGND.n40 0.122949
R91 VGND.n41 VGND.n2 0.122949
R92 VGND.n45 VGND.n2 0.122949
R93 VGND.n46 VGND.n45 0.122949
R94 VGND.n47 VGND.n46 0.122949
R95 VGND.n47 VGND.n0 0.122949
R96 a_2399_424.t1 a_2399_424.n1 423.303
R97 a_2399_424.n1 a_2399_424.t0 249.082
R98 a_2399_424.n0 a_2399_424.t2 240.197
R99 a_2399_424.n0 a_2399_424.t3 182.138
R100 a_2399_424.n1 a_2399_424.n0 125.391
R101 VNB.n0 VNB 22323.4
R102 VNB VNB.n1 19910
R103 VNB.n1 VNB.t13 2852.49
R104 VNB.t2 VNB.n0 2481.11
R105 VNB.t5 VNB.t10 2332.81
R106 VNB.t7 VNB.t8 2298.16
R107 VNB.t8 VNB.t11 2286.61
R108 VNB.t16 VNB.t15 2286.61
R109 VNB.t4 VNB.t1 2286.61
R110 VNB.t13 VNB.t16 1893.96
R111 VNB.t0 VNB.t9 1790.03
R112 VNB.t10 VNB.t6 1420.47
R113 VNB.n1 VNB.t2 1234.44
R114 VNB.t1 VNB 1143.31
R115 VNB.t12 VNB.t3 1050.92
R116 VNB.t15 VNB.t5 1004.72
R117 VNB.t6 VNB.t0 900.788
R118 VNB.t9 VNB.t4 900.788
R119 VNB.t3 VNB.t7 831.496
R120 VNB.t14 VNB.t12 831.496
R121 VNB.n0 VNB.t14 277.166
R122 a_855_368.n1 a_855_368.t2 1022.91
R123 a_855_368.t0 a_855_368.n5 886.183
R124 a_855_368.n2 a_855_368.n1 859.567
R125 a_855_368.t2 a_855_368.t3 644.514
R126 a_855_368.n2 a_855_368.t6 276.348
R127 a_855_368.n4 a_855_368.t4 264.298
R128 a_855_368.n5 a_855_368.t1 196.117
R129 a_855_368.n1 a_855_368.n0 185.303
R130 a_855_368.n3 a_855_368.t5 153.948
R131 a_855_368.n5 a_855_368.n4 152
R132 a_855_368.n3 a_855_368.n2 107.647
R133 a_855_368.n4 a_855_368.n3 29.9429
R134 a_1367_92.n3 a_1367_92.n2 275.752
R135 a_1367_92.n2 a_1367_92.n1 256.976
R136 a_1367_92.n1 a_1367_92.t3 232.344
R137 a_1367_92.n1 a_1367_92.n0 220.828
R138 a_1367_92.n2 a_1367_92.t0 211.25
R139 a_1367_92.n3 a_1367_92.t2 29.5505
R140 a_1367_92.t1 a_1367_92.n3 29.5505
R141 VPB.t15 VPB.t1 791.668
R142 VPB.t6 VPB.t8 607.797
R143 VPB.t13 VPB.t15 531.183
R144 VPB.t11 VPB.t2 531.183
R145 VPB.t12 VPB.t4 523.521
R146 VPB.t3 VPB.t7 515.861
R147 VPB.t1 VPB.t10 515.861
R148 VPB.t14 VPB.t9 380.512
R149 VPB.t4 VPB.t3 298.791
R150 VPB.t5 VPB.t11 291.13
R151 VPB VPB.t0 257.93
R152 VPB.t0 VPB.t16 255.376
R153 VPB.t10 VPB.t14 229.839
R154 VPB.t2 VPB.t13 229.839
R155 VPB.t9 VPB.t12 214.517
R156 VPB.t8 VPB.t5 214.517
R157 VPB.t16 VPB.t6 214.517
R158 VPWR.n32 VPWR.t1 783.648
R159 VPWR.n19 VPWR.t9 701.471
R160 VPWR.n46 VPWR.n4 605.946
R161 VPWR.n40 VPWR.n7 604.976
R162 VPWR.n17 VPWR.n16 317.613
R163 VPWR.n53 VPWR.n1 315.832
R164 VPWR.n26 VPWR.t7 287.534
R165 VPWR.n15 VPWR.t6 255.805
R166 VPWR.n16 VPWR.t4 115.874
R167 VPWR.n4 VPWR.t8 83.1099
R168 VPWR.n1 VPWR.t0 61.563
R169 VPWR.n16 VPWR.t3 47.0087
R170 VPWR.n1 VPWR.t11 46.1724
R171 VPWR.n4 VPWR.t5 46.1724
R172 VPWR.n47 VPWR.n2 36.1417
R173 VPWR.n51 VPWR.n2 36.1417
R174 VPWR.n52 VPWR.n51 36.1417
R175 VPWR.n41 VPWR.n5 36.1417
R176 VPWR.n45 VPWR.n5 36.1417
R177 VPWR.n34 VPWR.n33 36.1417
R178 VPWR.n34 VPWR.n8 36.1417
R179 VPWR.n38 VPWR.n8 36.1417
R180 VPWR.n39 VPWR.n38 36.1417
R181 VPWR.n24 VPWR.n13 36.1417
R182 VPWR.n25 VPWR.n24 36.1417
R183 VPWR.n27 VPWR.n25 36.1417
R184 VPWR.n31 VPWR.n11 36.1417
R185 VPWR.n20 VPWR.n18 36.1417
R186 VPWR.n47 VPWR.n46 34.2593
R187 VPWR.n27 VPWR.n26 30.8711
R188 VPWR.n32 VPWR.n31 28.6123
R189 VPWR.n7 VPWR.t10 26.3844
R190 VPWR.n7 VPWR.t2 26.3844
R191 VPWR.n53 VPWR.n52 19.2005
R192 VPWR.n33 VPWR.n32 18.4476
R193 VPWR.n18 VPWR.n17 15.0593
R194 VPWR.n46 VPWR.n45 13.177
R195 VPWR.n19 VPWR.n13 12.424
R196 VPWR.n41 VPWR.n40 10.9181
R197 VPWR.n18 VPWR.n14 9.3005
R198 VPWR.n21 VPWR.n20 9.3005
R199 VPWR.n22 VPWR.n13 9.3005
R200 VPWR.n24 VPWR.n23 9.3005
R201 VPWR.n25 VPWR.n12 9.3005
R202 VPWR.n28 VPWR.n27 9.3005
R203 VPWR.n29 VPWR.n11 9.3005
R204 VPWR.n31 VPWR.n30 9.3005
R205 VPWR.n32 VPWR.n10 9.3005
R206 VPWR.n33 VPWR.n9 9.3005
R207 VPWR.n35 VPWR.n34 9.3005
R208 VPWR.n36 VPWR.n8 9.3005
R209 VPWR.n38 VPWR.n37 9.3005
R210 VPWR.n39 VPWR.n6 9.3005
R211 VPWR.n42 VPWR.n41 9.3005
R212 VPWR.n43 VPWR.n5 9.3005
R213 VPWR.n45 VPWR.n44 9.3005
R214 VPWR.n46 VPWR.n3 9.3005
R215 VPWR.n48 VPWR.n47 9.3005
R216 VPWR.n49 VPWR.n2 9.3005
R217 VPWR.n51 VPWR.n50 9.3005
R218 VPWR.n52 VPWR.n0 9.3005
R219 VPWR.n54 VPWR.n53 7.43488
R220 VPWR.n17 VPWR.n15 7.17443
R221 VPWR.n26 VPWR.n11 5.27109
R222 VPWR.n20 VPWR.n19 4.89462
R223 VPWR.n15 VPWR.n14 0.48133
R224 VPWR.n40 VPWR.n39 0.376971
R225 VPWR VPWR.n54 0.160103
R226 VPWR.n54 VPWR.n0 0.1477
R227 VPWR.n21 VPWR.n14 0.122949
R228 VPWR.n22 VPWR.n21 0.122949
R229 VPWR.n23 VPWR.n22 0.122949
R230 VPWR.n23 VPWR.n12 0.122949
R231 VPWR.n28 VPWR.n12 0.122949
R232 VPWR.n29 VPWR.n28 0.122949
R233 VPWR.n30 VPWR.n29 0.122949
R234 VPWR.n30 VPWR.n10 0.122949
R235 VPWR.n10 VPWR.n9 0.122949
R236 VPWR.n35 VPWR.n9 0.122949
R237 VPWR.n36 VPWR.n35 0.122949
R238 VPWR.n37 VPWR.n36 0.122949
R239 VPWR.n37 VPWR.n6 0.122949
R240 VPWR.n42 VPWR.n6 0.122949
R241 VPWR.n43 VPWR.n42 0.122949
R242 VPWR.n44 VPWR.n43 0.122949
R243 VPWR.n44 VPWR.n3 0.122949
R244 VPWR.n48 VPWR.n3 0.122949
R245 VPWR.n49 VPWR.n48 0.122949
R246 VPWR.n50 VPWR.n49 0.122949
R247 VPWR.n50 VPWR.n0 0.122949
R248 SCE SCE.t0 441.238
R249 SCE.n2 SCE.t1 276.171
R250 SCE.n1 SCE.t3 243.288
R251 SCE.n2 SCE.t2 238.672
R252 SCE SCE.n3 152.558
R253 SCE.n1 SCE.n0 152
R254 SCE.n3 SCE.n1 49.6611
R255 SCE.n3 SCE.n2 16.8278
R256 SCE SCE.n0 12.0585
R257 SCE.n0 SCE 5.75122
R258 a_300_464.n1 a_300_464.t6 656.381
R259 a_300_464.n1 a_300_464.t5 395.135
R260 a_300_464.n3 a_300_464.n0 360.995
R261 a_300_464.n2 a_300_464.t4 354.103
R262 a_300_464.n4 a_300_464.n3 142.03
R263 a_300_464.n0 a_300_464.t1 138.571
R264 a_300_464.n2 a_300_464.n1 137.984
R265 a_300_464.t2 a_300_464.n4 130.774
R266 a_300_464.n4 a_300_464.t3 126.668
R267 a_300_464.n0 a_300_464.t0 40.0005
R268 a_300_464.n3 a_300_464.n2 11.2791
R269 a_545_81.t0 a_545_81.t1 68.5719
R270 a_1997_272.n1 a_1997_272.t1 731.564
R271 a_1997_272.t0 a_1997_272.n1 329.579
R272 a_1997_272.n0 a_1997_272.t3 313.808
R273 a_1997_272.n0 a_1997_272.t2 274.74
R274 a_1997_272.n1 a_1997_272.n0 232.251
R275 a_27_88.n1 a_27_88.t3 377.115
R276 a_27_88.t1 a_27_88.n1 368.841
R277 a_27_88.n0 a_27_88.t2 361.158
R278 a_27_88.n0 a_27_88.t0 250.857
R279 a_27_88.n1 a_27_88.n0 64.6471
R280 a_225_81.t0 a_225_81.n0 549.854
R281 a_225_81.n0 a_225_81.t2 67.1434
R282 a_225_81.n0 a_225_81.t1 65.7148
R283 a_312_81.t0 a_312_81.t1 68.5719
R284 RESET_B.n1 RESET_B.t0 401.277
R285 RESET_B.n4 RESET_B.n3 399.038
R286 RESET_B.n2 RESET_B.t2 390.421
R287 RESET_B.n5 RESET_B.n2 212.758
R288 RESET_B.n5 RESET_B.n4 210.367
R289 RESET_B.n1 RESET_B.n0 199.671
R290 RESET_B RESET_B.n1 163.286
R291 RESET_B.n2 RESET_B.t3 156.131
R292 RESET_B.n4 RESET_B.t1 114.341
R293 RESET_B RESET_B.n5 2.42441
R294 a_1034_368.t1 a_1034_368.n4 866.264
R295 a_1034_368.n2 a_1034_368.t3 442.808
R296 a_1034_368.n2 a_1034_368.t2 384.587
R297 a_1034_368.n1 a_1034_368.n0 350.985
R298 a_1034_368.n3 a_1034_368.n2 344.704
R299 a_1034_368.n1 a_1034_368.t4 205.387
R300 a_1034_368.n4 a_1034_368.n1 169.262
R301 a_1034_368.n3 a_1034_368.t0 136.871
R302 a_1034_368.n4 a_1034_368.n3 54.1615
R303 a_1993_508.t0 a_1993_508.t1 126.644
R304 CLK.n0 CLK.t1 250.909
R305 CLK.n0 CLK.t0 170.016
R306 CLK.n1 CLK.n0 117.77
R307 CLK.n1 CLK 13.6005
R308 CLK CLK.n1 3.29747
R309 a_2135_74.t0 a_2135_74.t1 60.0005
R310 Q.n1 Q 591.274
R311 Q.n1 Q.n0 585
R312 Q.n2 Q.n1 585
R313 Q.t0 Q.n3 279.738
R314 Q.n4 Q.t0 279.738
R315 Q.n1 Q.t1 26.3844
R316 Q.n2 Q 16.8162
R317 Q.n0 Q 14.5574
R318 Q.n4 Q 12.6066
R319 Q.n3 Q 10.4162
R320 Q.n3 Q 4.84898
R321 Q.n0 Q 4.01619
R322 Q Q.n2 1.75736
R323 Q Q.n4 1.74595
R324 a_1972_74.t0 a_1972_74.t1 60.0005
R325 SCD.n1 SCD.t1 289.2
R326 SCD.n2 SCD.t0 187.178
R327 SCD.n1 SCD.n0 152
R328 SCD.n3 SCD.n2 152
R329 SCD.n2 SCD.n1 49.6611
R330 SCD.n3 SCD.n0 13.1884
R331 SCD.n0 SCD 0.970197
R332 SCD SCD.n3 0.194439
R333 a_538_464.t0 a_538_464.t1 83.1099
R334 D.n0 D.t0 494.587
R335 D D.n0 161.565
R336 D.n0 D.t1 126.927
R337 a_216_464.t0 a_216_464.t1 83.1099
C0 a_1233_118# VGND 0.019108f
C1 RESET_B Q 2.89e-19
C2 VPB VGND 0.02548f
C3 SCE VPWR 0.041126f
C4 D VPWR 0.014528f
C5 SCD SCE 0.081634f
C6 D SCD 0.003639f
C7 RESET_B VPWR 0.358405f
C8 VPB Q 0.013733f
C9 SCD RESET_B 0.07716f
C10 a_1343_461# VPWR 6.3e-19
C11 RESET_B CLK 0.076051f
C12 a_1233_118# VPWR 0.173685f
C13 VPB VPWR 0.394626f
C14 D SCE 0.133293f
C15 SCD VPB 0.075307f
C16 VPB CLK 0.051196f
C17 SCE RESET_B 9.07e-20
C18 a_1319_118# RESET_B 7.06e-19
C19 D RESET_B 6.74e-20
C20 VGND Q 0.100718f
C21 a_1233_118# a_1319_118# 0.005793f
C22 a_1343_461# RESET_B 4.36e-19
C23 a_1233_118# RESET_B 0.247657f
C24 VPB SCE 0.150182f
C25 D VPB 0.092838f
C26 VPWR VGND 0.104847f
C27 a_1233_118# a_1343_461# 0.006779f
C28 SCD VGND 0.005873f
C29 VPB RESET_B 0.361036f
C30 CLK VGND 0.025909f
C31 VPWR Q 0.121768f
C32 VPB a_1233_118# 0.092298f
C33 SCE VGND 0.02701f
C34 a_1319_118# VGND 0.001081f
C35 D VGND 0.012397f
C36 SCD VPWR 0.014663f
C37 RESET_B VGND 0.200476f
C38 CLK VPWR 0.01046f
C39 Q VNB 0.11184f
C40 VGND VNB 1.56223f
C41 VPWR VNB 1.20007f
C42 CLK VNB 0.161482f
C43 RESET_B VNB 0.428338f
C44 SCD VNB 0.122695f
C45 D VNB 0.16909f
C46 SCE VNB 0.34783f
C47 VPB VNB 3.10378f
C48 a_1233_118# VNB 0.152935f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrtn_1 VNB VPB VPWR RESET_B VGND Q CLK_N SCD SCE D
X0 VGND RESET_B a_1489_131# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.164 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 a_2087_410.t1 a_1827_144# a_2265_74.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.21 pd=1.84 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 VPWR.t0 a_2087_410.t3 a_2042_508.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.13125 pd=1.045 as=0.0546 ps=0.68 w=0.42 l=0.15
X3 a_1489_131# a_1429_308.t2 a_1411_131.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4 a_1272_131.t0 RESET_B.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X5 VGND.t3 SCE.t0 a_27_88.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.1197 ps=1.41 w=0.42 l=0.15
X6 VPWR.t9 a_1429_308.t3 a_1384_508.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_324_81.t1 a_27_88.t2 a_239_81.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1155 ps=1.39 w=0.42 l=0.15
X8 a_239_81.t2 SCD.t0 a_538_81.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0609 pd=0.71 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 VPWR.t8 SCE.t1 a_27_88.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1888 ps=1.87 w=0.64 l=0.15
X10 a_2073_74.t1 a_1074_88.t2 a_1827_144# VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0525 pd=0.67 as=0.312825 ps=2.13 w=0.42 l=0.15
X11 Q.t1 a_2492_424.t1 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.2282 ps=1.55 w=1.12 l=0.15
X12 VPWR.t12 a_1827_144# a_2492_424.t0 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.2282 pd=1.55 as=0.2478 ps=2.27 w=0.84 l=0.15
X13 Q.t0 a_2492_424.t2 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X14 a_1384_508.t0 a_1074_88.t3 a_1272_131.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X15 a_284_464.t3 D.t0 a_324_81.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1176 pd=0.98 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_1272_131.t3 a_854_74.t2 a_284_464.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X17 a_1429_308.t0 a_1272_131.t4 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3925 pd=1.785 as=0.285 ps=2.57 w=1 l=0.15
X18 a_1429_308.t1 a_1272_131.t5 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1792 pd=1.2 as=0.164 ps=1.41 w=0.64 l=0.15
X19 a_1074_88.t1 a_854_74.t3 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X20 a_2265_74.t0 RESET_B.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0861 ps=0.83 w=0.42 l=0.15
X21 VPWR.t11 a_1827_144# a_2087_410.t2 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.1449 pd=1.53 as=0.063 ps=0.72 w=0.42 l=0.15
X22 a_284_464.t0 RESET_B.t2 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.184475 ps=1.345 w=0.64 l=0.15
X23 a_1074_88.t0 a_854_74.t4 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.3899 ps=2.88 w=0.74 l=0.15
X24 a_854_74.t1 CLK_N.t0 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.4144 ps=2.98 w=1.12 l=0.15
X25 a_2087_410.t0 RESET_B.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.13125 ps=1.045 w=0.42 l=0.15
X26 a_1272_131.t2 a_1074_88.t4 a_284_464.t6 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.11445 pd=0.965 as=0.1197 ps=1.41 w=0.42 l=0.15
X27 VGND.t5 a_2087_410.t4 a_2073_74.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0861 pd=0.83 as=0.0525 ps=0.67 w=0.42 l=0.15
X28 a_284_464.t2 D.t1 a_206_464.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.2512 pd=1.425 as=0.0768 ps=0.88 w=0.64 l=0.15
X29 a_2042_508.t1 a_854_74.t5 a_1827_144# VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0546 pd=0.68 as=0.1564 ps=1.365 w=0.42 l=0.15
X30 VPWR.t5 SCD.t1 a_471_464.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.184475 pd=1.345 as=0.0768 ps=0.88 w=0.64 l=0.15
X31 a_538_81.t0 SCE.t2 a_284_464.t4 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1176 ps=0.98 w=0.42 l=0.15
X32 a_854_74.t0 CLK_N.t1 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.223675 ps=1.575 w=0.74 l=0.15
X33 a_471_464.t0 a_27_88.t3 a_284_464.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.2512 ps=1.425 w=0.64 l=0.15
X34 a_206_464.t1 SCE.t3 VPWR.t13 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.096 ps=0.94 w=0.64 l=0.15
X35 VGND.t0 RESET_B.t4 a_239_81.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.223675 pd=1.575 as=0.0609 ps=0.71 w=0.42 l=0.15
R0 RESET_B.n0 RESET_B.t3 393.873
R1 RESET_B.n2 RESET_B.t0 296.966
R2 RESET_B.n4 RESET_B.t4 279.123
R3 RESET_B.n4 RESET_B.t2 240.803
R4 RESET_B.n0 RESET_B.t1 226.541
R5 RESET_B.n2 RESET_B.n1 218.507
R6 RESET_B.n3 RESET_B.n0 177.48
R7 RESET_B.n3 RESET_B.n2 164.016
R8 RESET_B.n5 RESET_B.n4 78.7626
R9 RESET_B.n5 RESET_B.n3 3.75632
R10 RESET_B RESET_B.n5 0.0466957
R11 VGND.n33 VGND.t6 359.281
R12 VGND.n22 VGND.t2 345.849
R13 VGND.n46 VGND.t3 270.212
R14 VGND.n4 VGND.n3 210.333
R15 VGND.n14 VGND.n13 199.026
R16 VGND.n12 VGND.t7 153.27
R17 VGND.n3 VGND.t0 80.7697
R18 VGND.n3 VGND.t4 66.4246
R19 VGND.n13 VGND.t1 60.0005
R20 VGND.n13 VGND.t5 57.1434
R21 VGND.n16 VGND.n15 36.1417
R22 VGND.n16 VGND.n10 36.1417
R23 VGND.n20 VGND.n10 36.1417
R24 VGND.n21 VGND.n20 36.1417
R25 VGND.n26 VGND.n8 36.1417
R26 VGND.n27 VGND.n26 36.1417
R27 VGND.n28 VGND.n27 36.1417
R28 VGND.n28 VGND.n6 36.1417
R29 VGND.n35 VGND.n34 36.1417
R30 VGND.n40 VGND.n39 36.1417
R31 VGND.n40 VGND.n1 36.1417
R32 VGND.n44 VGND.n1 36.1417
R33 VGND.n45 VGND.n44 36.1417
R34 VGND.n39 VGND.n38 34.9784
R35 VGND.n22 VGND.n8 33.8829
R36 VGND.n15 VGND.n14 30.8711
R37 VGND.n32 VGND.n6 30.3254
R38 VGND.n34 VGND.n33 23.6251
R39 VGND.n46 VGND.n45 19.2005
R40 VGND.n22 VGND.n21 13.5534
R41 VGND.n45 VGND.n0 9.3005
R42 VGND.n44 VGND.n43 9.3005
R43 VGND.n42 VGND.n1 9.3005
R44 VGND.n41 VGND.n40 9.3005
R45 VGND.n39 VGND.n2 9.3005
R46 VGND.n38 VGND.n37 9.3005
R47 VGND.n36 VGND.n35 9.3005
R48 VGND.n34 VGND.n5 9.3005
R49 VGND.n32 VGND.n31 9.3005
R50 VGND.n30 VGND.n6 9.3005
R51 VGND.n29 VGND.n28 9.3005
R52 VGND.n27 VGND.n7 9.3005
R53 VGND.n26 VGND.n25 9.3005
R54 VGND.n24 VGND.n8 9.3005
R55 VGND.n23 VGND.n22 9.3005
R56 VGND.n21 VGND.n9 9.3005
R57 VGND.n20 VGND.n19 9.3005
R58 VGND.n18 VGND.n10 9.3005
R59 VGND.n17 VGND.n16 9.3005
R60 VGND.n15 VGND.n11 9.3005
R61 VGND.n35 VGND.n4 8.1771
R62 VGND.n47 VGND.n46 7.43488
R63 VGND.n38 VGND.n4 6.32859
R64 VGND.n14 VGND.n12 5.49636
R65 VGND.n33 VGND.n32 1.58252
R66 VGND.n12 VGND.n11 0.187568
R67 VGND VGND.n47 0.160103
R68 VGND.n47 VGND.n0 0.1477
R69 VGND.n17 VGND.n11 0.122949
R70 VGND.n18 VGND.n17 0.122949
R71 VGND.n19 VGND.n18 0.122949
R72 VGND.n19 VGND.n9 0.122949
R73 VGND.n23 VGND.n9 0.122949
R74 VGND.n24 VGND.n23 0.122949
R75 VGND.n25 VGND.n24 0.122949
R76 VGND.n25 VGND.n7 0.122949
R77 VGND.n29 VGND.n7 0.122949
R78 VGND.n30 VGND.n29 0.122949
R79 VGND.n31 VGND.n30 0.122949
R80 VGND.n31 VGND.n5 0.122949
R81 VGND.n36 VGND.n5 0.122949
R82 VGND.n37 VGND.n36 0.122949
R83 VGND.n37 VGND.n2 0.122949
R84 VGND.n41 VGND.n2 0.122949
R85 VGND.n42 VGND.n41 0.122949
R86 VGND.n43 VGND.n42 0.122949
R87 VGND.n43 VGND.n0 0.122949
R88 VNB.n0 VNB 22461.9
R89 VNB VNB.n1 13026.2
R90 VNB.t14 VNB.t12 4122.83
R91 VNB.t4 VNB.n0 2987.65
R92 VNB.t11 VNB.t8 2540.68
R93 VNB.t5 VNB.t6 2425.2
R94 VNB.t13 VNB.t9 2357.53
R95 VNB.t9 VNB.t4 2129.38
R96 VNB.t8 VNB.t2 1732.28
R97 VNB.t15 VNB.t1 1639.9
R98 VNB.n1 VNB.t11 1616.8
R99 VNB.n0 VNB.t0 1304.99
R100 VNB.t10 VNB.t3 1293.44
R101 VNB.t6 VNB 1143.31
R102 VNB.t2 VNB.t7 1016.27
R103 VNB.t0 VNB.t10 923.885
R104 VNB.t3 VNB.t14 900.788
R105 VNB.t7 VNB.t15 900.788
R106 VNB.t1 VNB.t5 831.496
R107 VNB.n1 VNB.t13 630.124
R108 a_2265_74.t0 a_2265_74.t1 68.5719
R109 a_2087_410.n2 a_2087_410.n1 599.545
R110 a_2087_410.n0 a_2087_410.t4 496.461
R111 a_2087_410.t1 a_2087_410.n2 417.575
R112 a_2087_410.n2 a_2087_410.n0 212.522
R113 a_2087_410.n0 a_2087_410.t3 138.441
R114 a_2087_410.n1 a_2087_410.t2 70.3576
R115 a_2087_410.n1 a_2087_410.t0 70.3576
R116 a_2042_508.t0 a_2042_508.t1 121.953
R117 VPWR.n40 VPWR.t7 878.966
R118 VPWR.n4 VPWR.t10 823.467
R119 VPWR.n14 VPWR.t11 699.173
R120 VPWR.n48 VPWR.n47 649.534
R121 VPWR.n33 VPWR.n9 612.393
R122 VPWR.n55 VPWR.n1 605.365
R123 VPWR.n21 VPWR.n20 585
R124 VPWR.n10 VPWR.t4 345.288
R125 VPWR.n16 VPWR.n15 235.579
R126 VPWR.n20 VPWR.t1 159.476
R127 VPWR.n20 VPWR.t0 133.679
R128 VPWR.n47 VPWR.t3 72.3364
R129 VPWR.n47 VPWR.t5 72.3364
R130 VPWR.n9 VPWR.t2 70.3576
R131 VPWR.n9 VPWR.t9 70.3576
R132 VPWR.n15 VPWR.t12 56.8374
R133 VPWR.n1 VPWR.t13 46.1724
R134 VPWR.n1 VPWR.t8 46.1724
R135 VPWR.n49 VPWR.n2 36.1417
R136 VPWR.n53 VPWR.n2 36.1417
R137 VPWR.n54 VPWR.n53 36.1417
R138 VPWR.n35 VPWR.n34 36.1417
R139 VPWR.n35 VPWR.n6 36.1417
R140 VPWR.n39 VPWR.n6 36.1417
R141 VPWR.n26 VPWR.n12 36.1417
R142 VPWR.n27 VPWR.n26 36.1417
R143 VPWR.n28 VPWR.n27 36.1417
R144 VPWR.n19 VPWR.n18 36.1417
R145 VPWR.n15 VPWR.t6 36.1099
R146 VPWR.n46 VPWR.n45 34.9784
R147 VPWR.n41 VPWR.n40 32.7534
R148 VPWR.n32 VPWR.n10 28.2358
R149 VPWR.n33 VPWR.n32 28.2358
R150 VPWR.n34 VPWR.n33 25.224
R151 VPWR.n22 VPWR.n12 24.7221
R152 VPWR.n41 VPWR.n4 24.0946
R153 VPWR.n45 VPWR.n4 23.3417
R154 VPWR.n55 VPWR.n54 22.9652
R155 VPWR.n28 VPWR.n10 19.2005
R156 VPWR.n49 VPWR.n48 17.923
R157 VPWR.n40 VPWR.n39 14.6829
R158 VPWR.n21 VPWR.n19 10.3744
R159 VPWR.n16 VPWR.n14 9.54324
R160 VPWR.n18 VPWR.n17 9.3005
R161 VPWR.n19 VPWR.n13 9.3005
R162 VPWR.n23 VPWR.n22 9.3005
R163 VPWR.n24 VPWR.n12 9.3005
R164 VPWR.n26 VPWR.n25 9.3005
R165 VPWR.n27 VPWR.n11 9.3005
R166 VPWR.n29 VPWR.n28 9.3005
R167 VPWR.n30 VPWR.n10 9.3005
R168 VPWR.n32 VPWR.n31 9.3005
R169 VPWR.n33 VPWR.n8 9.3005
R170 VPWR.n34 VPWR.n7 9.3005
R171 VPWR.n36 VPWR.n35 9.3005
R172 VPWR.n37 VPWR.n6 9.3005
R173 VPWR.n39 VPWR.n38 9.3005
R174 VPWR.n40 VPWR.n5 9.3005
R175 VPWR.n42 VPWR.n41 9.3005
R176 VPWR.n43 VPWR.n4 9.3005
R177 VPWR.n45 VPWR.n44 9.3005
R178 VPWR.n46 VPWR.n3 9.3005
R179 VPWR.n50 VPWR.n49 9.3005
R180 VPWR.n51 VPWR.n2 9.3005
R181 VPWR.n53 VPWR.n52 9.3005
R182 VPWR.n54 VPWR.n0 9.3005
R183 VPWR.n18 VPWR.n14 9.03579
R184 VPWR.n56 VPWR.n55 7.27223
R185 VPWR.n48 VPWR.n46 4.02747
R186 VPWR.n22 VPWR.n21 1.75736
R187 VPWR.n17 VPWR.n16 0.491584
R188 VPWR VPWR.n56 0.157962
R189 VPWR.n56 VPWR.n0 0.149814
R190 VPWR.n17 VPWR.n13 0.122949
R191 VPWR.n23 VPWR.n13 0.122949
R192 VPWR.n24 VPWR.n23 0.122949
R193 VPWR.n25 VPWR.n24 0.122949
R194 VPWR.n25 VPWR.n11 0.122949
R195 VPWR.n29 VPWR.n11 0.122949
R196 VPWR.n30 VPWR.n29 0.122949
R197 VPWR.n31 VPWR.n30 0.122949
R198 VPWR.n31 VPWR.n8 0.122949
R199 VPWR.n8 VPWR.n7 0.122949
R200 VPWR.n36 VPWR.n7 0.122949
R201 VPWR.n37 VPWR.n36 0.122949
R202 VPWR.n38 VPWR.n37 0.122949
R203 VPWR.n38 VPWR.n5 0.122949
R204 VPWR.n42 VPWR.n5 0.122949
R205 VPWR.n43 VPWR.n42 0.122949
R206 VPWR.n44 VPWR.n43 0.122949
R207 VPWR.n44 VPWR.n3 0.122949
R208 VPWR.n50 VPWR.n3 0.122949
R209 VPWR.n51 VPWR.n50 0.122949
R210 VPWR.n52 VPWR.n51 0.122949
R211 VPWR.n52 VPWR.n0 0.122949
R212 VPB.n0 VPB 4967.07
R213 VPB VPB.n1 3273.13
R214 VPB.t4 VPB.n0 567.817
R215 VPB.t13 VPB.t2 554.168
R216 VPB.t3 VPB.t4 545.977
R217 VPB.t16 VPB.t17 541.399
R218 VPB.t9 VPB.t13 515.861
R219 VPB.t6 VPB.t15 477.555
R220 VPB.t0 VPB.t1 395.834
R221 VPB.t2 VPB.t5 316.668
R222 VPB.n1 VPB.t9 311.56
R223 VPB.t17 VPB.t7 296.238
R224 VPB.t10 VPB 257.93
R225 VPB.t11 VPB.t3 245.69
R226 VPB.t8 VPB.t12 245.69
R227 VPB.t1 VPB.t16 229.839
R228 VPB.t18 VPB.t10 229.839
R229 VPB.n1 VPB.t8 218.392
R230 VPB.t12 VPB.t11 212.931
R231 VPB.t14 VPB.t0 209.41
R232 VPB.n0 VPB.t14 209.41
R233 VPB.t5 VPB.t6 199.195
R234 VPB.t15 VPB.t18 199.195
R235 a_1429_308.n0 a_1429_308.t3 275.009
R236 a_1429_308.n1 a_1429_308.n0 263.618
R237 a_1429_308.n0 a_1429_308.t2 241
R238 a_1429_308.t0 a_1429_308.n1 237.786
R239 a_1429_308.n1 a_1429_308.t1 237.5
R240 a_854_74.n1 a_854_74.n0 1097.35
R241 a_854_74.n0 a_854_74.t5 898.957
R242 a_854_74.t1 a_854_74.n5 876.971
R243 a_854_74.n2 a_854_74.t2 477.18
R244 a_854_74.n2 a_854_74.n1 461.113
R245 a_854_74.n5 a_854_74.t0 339.904
R246 a_854_74.n3 a_854_74.t3 242.875
R247 a_854_74.n5 a_854_74.n4 193.627
R248 a_854_74.n3 a_854_74.n2 164.173
R249 a_854_74.n4 a_854_74.t4 154.24
R250 a_854_74.n4 a_854_74.n3 13.146
R251 a_1272_131.n1 a_1272_131.t0 670.485
R252 a_1272_131.n3 a_1272_131.n2 613.771
R253 a_1272_131.t2 a_1272_131.n3 394.675
R254 a_1272_131.n0 a_1272_131.t4 250.617
R255 a_1272_131.n1 a_1272_131.n0 201.381
R256 a_1272_131.n0 a_1272_131.t5 144.017
R257 a_1272_131.n2 a_1272_131.t1 70.3576
R258 a_1272_131.n2 a_1272_131.t3 70.3576
R259 a_1272_131.n3 a_1272_131.n1 67.7652
R260 a_2492_424.t0 a_2492_424.n0 679.817
R261 a_2492_424.n0 a_2492_424.t1 225.47
R262 a_2492_424.n0 a_2492_424.t2 199.811
R263 SCE SCE.t2 303.568
R264 SCE.n1 SCE.t0 277.899
R265 SCE.n0 SCE.t3 191.194
R266 SCE.n0 SCE.t1 180.496
R267 SCE SCE.n1 159.712
R268 SCE.n1 SCE.n0 26.9332
R269 a_27_88.n1 a_27_88.t3 562.431
R270 a_27_88.n0 a_27_88.t2 393.178
R271 a_27_88.t1 a_27_88.n1 359.966
R272 a_27_88.n0 a_27_88.t0 234.216
R273 a_27_88.n1 a_27_88.n0 79.1045
R274 a_1384_508.t0 a_1384_508.t1 112.572
R275 a_239_81.n0 a_239_81.t1 547.617
R276 a_239_81.t0 a_239_81.n0 41.4291
R277 a_239_81.n0 a_239_81.t2 41.4291
R278 a_324_81.t0 a_324_81.t1 60.0005
R279 SCD.n0 SCD.t0 316.514
R280 SCD.n0 SCD.t1 294.021
R281 SCD.n1 SCD.n0 152
R282 SCD SCD.n1 7.65107
R283 SCD.n1 SCD 3.23728
R284 a_538_81.t0 a_538_81.t1 68.5719
R285 a_1074_88.t1 a_1074_88.n4 843.654
R286 a_1074_88.n4 a_1074_88.t3 431.38
R287 a_1074_88.n1 a_1074_88.n0 384.262
R288 a_1074_88.n2 a_1074_88.n1 382.423
R289 a_1074_88.n3 a_1074_88.t0 291.955
R290 a_1074_88.n2 a_1074_88.t4 284.769
R291 a_1074_88.n1 a_1074_88.t2 259.259
R292 a_1074_88.n3 a_1074_88.n2 113.085
R293 a_1074_88.n4 a_1074_88.n3 24.2429
R294 a_2073_74.t0 a_2073_74.t1 71.4291
R295 Q.n3 Q 589.85
R296 Q.n3 Q.n0 585
R297 Q.n4 Q.n3 585
R298 Q.n2 Q.t0 279.738
R299 Q.t0 Q.n1 279.738
R300 Q.n3 Q.t1 27.2639
R301 Q Q.n4 12.9944
R302 Q.n1 Q 12.6066
R303 Q Q.n0 11.249
R304 Q Q.n2 9.50353
R305 Q.n2 Q 4.84898
R306 Q Q.n0 3.10353
R307 Q.n1 Q 1.74595
R308 Q.n4 Q 1.35808
R309 D.n0 D.t0 387.5
R310 D.n0 D.t1 276.348
R311 D D.n0 160.282
R312 a_284_464.n4 a_284_464.t5 825.324
R313 a_284_464.t0 a_284_464.n1 706.985
R314 a_284_464.t0 a_284_464.n5 701.865
R315 a_284_464.n3 a_284_464.t6 405.707
R316 a_284_464.n1 a_284_464.n0 361.486
R317 a_284_464.n3 a_284_464.n2 334.082
R318 a_284_464.n0 a_284_464.t2 113.538
R319 a_284_464.n0 a_284_464.t1 111.441
R320 a_284_464.n4 a_284_464.n3 83.9534
R321 a_284_464.n2 a_284_464.t4 80.0005
R322 a_284_464.n2 a_284_464.t3 80.0005
R323 a_284_464.n5 a_284_464.n4 26.7708
R324 a_284_464.n5 a_284_464.n1 12.8005
R325 CLK_N.n0 CLK_N.t0 278.017
R326 CLK_N.n0 CLK_N.t1 170.638
R327 CLK_N CLK_N.n0 157.601
R328 a_206_464.t0 a_206_464.t1 73.8755
R329 a_471_464.t0 a_471_464.t1 73.8755
C0 SCE SCD 0.045493f
C1 VPB Q 0.013631f
C2 CLK_N VPB 0.04529f
C3 VPB SCD 0.088636f
C4 SCE VPB 0.131676f
C5 VGND Q 0.10291f
C6 CLK_N VGND 0.011554f
C7 RESET_B Q 2.48e-19
C8 SCD VGND 0.006408f
C9 RESET_B CLK_N 0.048448f
C10 RESET_B SCD 0.146756f
C11 VPWR Q 0.134174f
C12 SCE VGND 0.029159f
C13 D SCD 0.004627f
C14 RESET_B SCE 0.004248f
C15 CLK_N VPWR 0.016021f
C16 SCE D 0.193031f
C17 VPWR SCD 0.014749f
C18 VPB VGND 0.01685f
C19 VPWR SCE 0.034415f
C20 RESET_B VPB 0.31907f
C21 a_1489_131# VGND 0.001392f
C22 VPB D 0.113158f
C23 RESET_B a_1489_131# 8.87e-19
C24 VPWR VPB 0.408116f
C25 a_1827_144# Q 0.002004f
C26 VPB a_1827_144# 0.234208f
C27 a_1489_131# a_1827_144# 1.23e-19
C28 RESET_B VGND 0.261576f
C29 D VGND 0.006149f
C30 RESET_B D 2.73e-19
C31 VPWR VGND 0.107905f
C32 RESET_B VPWR 0.277657f
C33 VPWR D 0.014656f
C34 a_1827_144# VGND 0.242893f
C35 RESET_B a_1827_144# 0.327064f
C36 VPWR a_1827_144# 0.098048f
C37 Q VNB 0.110216f
C38 VGND VNB 1.5908f
C39 CLK_N VNB 0.139524f
C40 RESET_B VNB 0.442874f
C41 SCD VNB 0.126665f
C42 D VNB 0.134184f
C43 SCE VNB 0.351846f
C44 VPWR VNB 1.2258f
C45 VPB VNB 3.13805f
C46 a_1827_144# VNB 0.376852f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdlclkp_1 VNB VPB VPWR VGND GCLK CLK GATE SCE
X0 a_566_74.t2 a_318_74.t2 a_114_112.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.155475 pd=1.37 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VPWR.t6 a_709_54.t2 a_1238_94.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.126 ps=1.14 w=0.84 l=0.15
X2 a_1238_94.t0 CLK.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.281825 ps=1.675 w=0.84 l=0.15
X3 GCLK.t0 a_1238_94.t3 VPWR.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.4256 pd=3 as=0.1862 ps=1.475 w=1.12 l=0.15
X4 a_114_112.t3 GATE.t0 a_116_424.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1008 ps=1.08 w=0.84 l=0.15
X5 a_709_54.t0 a_566_74.t4 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1513 ps=1.27 w=0.74 l=0.15
X6 a_318_74.t0 a_288_48.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.4033 ps=3.02 w=0.84 l=0.15
X7 GCLK.t1 a_1238_94.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.2664 ps=2.2 w=0.74 l=0.15
X8 VPWR.t3 CLK.t1 a_288_48.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.281825 pd=1.675 as=0.2478 ps=2.27 w=0.84 l=0.15
X9 a_318_74.t1 a_288_48.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.189025 ps=1.41 w=0.74 l=0.15
X10 VPWR.t5 a_709_54.t3 a_722_492.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1673 pd=1.475 as=0.0504 ps=0.66 w=0.42 l=0.15
X11 a_1166_94.t0 CLK.t2 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1165 ps=1.065 w=0.64 l=0.15
X12 a_116_424.t1 SCE.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1008 pd=1.08 as=0.2478 ps=2.27 w=0.84 l=0.15
X13 a_722_492.t1 a_288_48.t4 a_566_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.155475 ps=1.37 w=0.42 l=0.15
X14 a_1238_94.t1 a_709_54.t4 a_1166_94.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0672 ps=0.85 w=0.64 l=0.15
X15 VGND.t5 CLK.t3 a_288_48.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.2072 ps=2.04 w=0.74 l=0.15
X16 VGND.t2 GATE.t1 a_114_112.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.189025 pd=1.41 as=0.077 ps=0.83 w=0.55 l=0.15
X17 a_566_74.t3 a_288_48.t5 a_114_112.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0923 pd=0.905 as=0.29425 ps=2.17 w=0.55 l=0.15
X18 a_667_80.t0 a_318_74.t3 a_566_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0923 ps=0.905 w=0.42 l=0.15
X19 a_114_112.t2 SCE.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.15675 ps=1.67 w=0.55 l=0.15
X20 a_709_54.t1 a_566_74.t5 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1673 ps=1.475 w=1.12 l=0.15
X21 VGND.t6 a_709_54.t5 a_667_80.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1513 pd=1.27 as=0.0441 ps=0.63 w=0.42 l=0.15
R0 a_318_74.t0 a_318_74.n1 768.644
R1 a_318_74.n1 a_318_74.t1 323.784
R2 a_318_74.n0 a_318_74.t3 287.01
R3 a_318_74.n1 a_318_74.n0 211.012
R4 a_318_74.n0 a_318_74.t2 187.178
R5 a_114_112.t1 a_114_112.n2 470.13
R6 a_114_112.n1 a_114_112.t4 376.086
R7 a_114_112.n2 a_114_112.t3 350.803
R8 a_114_112.n1 a_114_112.n0 185
R9 a_114_112.n2 a_114_112.n1 144.189
R10 a_114_112.n0 a_114_112.t0 30.546
R11 a_114_112.n0 a_114_112.t2 30.546
R12 a_566_74.n3 a_566_74.n2 344.921
R13 a_566_74.n0 a_566_74.t5 255.202
R14 a_566_74.n2 a_566_74.n1 217.298
R15 a_566_74.n2 a_566_74.n0 187.88
R16 a_566_74.n0 a_566_74.t4 169.246
R17 a_566_74.n3 a_566_74.t0 157.856
R18 a_566_74.n1 a_566_74.t1 61.4291
R19 a_566_74.t2 a_566_74.n3 28.7722
R20 a_566_74.n1 a_566_74.t3 22.2729
R21 VPB.t8 VPB.t0 559.274
R22 VPB.t9 VPB.t5 515.861
R23 VPB.t0 VPB.t4 515.861
R24 VPB.t5 VPB.t1 354.974
R25 VPB.t4 VPB.t3 273.253
R26 VPB.t2 VPB.t10 257.93
R27 VPB.t7 VPB.t9 257.93
R28 VPB VPB.t6 257.93
R29 VPB.t1 VPB.t2 229.839
R30 VPB.t3 VPB.t7 199.195
R31 VPB.t6 VPB.t8 199.195
R32 a_709_54.n0 a_709_54.t5 396.096
R33 a_709_54.n2 a_709_54.t2 378.37
R34 a_709_54.n3 a_709_54.n2 326.048
R35 a_709_54.n1 a_709_54.t0 265.964
R36 a_709_54.t1 a_709_54.n3 218.153
R37 a_709_54.n1 a_709_54.n0 179.621
R38 a_709_54.n0 a_709_54.t3 179.463
R39 a_709_54.n2 a_709_54.t4 162.274
R40 a_709_54.n3 a_709_54.n1 10.7353
R41 a_1238_94.n2 a_1238_94.n1 330.048
R42 a_1238_94.n0 a_1238_94.t3 250.565
R43 a_1238_94.n0 a_1238_94.t4 181.554
R44 a_1238_94.n1 a_1238_94.n0 172.171
R45 a_1238_94.n1 a_1238_94.t1 151.831
R46 a_1238_94.n2 a_1238_94.t2 35.1791
R47 a_1238_94.t0 a_1238_94.n2 35.1791
R48 VPWR.n1 VPWR.t0 920.826
R49 VPWR.n9 VPWR.n8 663.26
R50 VPWR.n15 VPWR.n5 610.601
R51 VPWR.n27 VPWR.t4 404.334
R52 VPWR.n10 VPWR.n7 326.707
R53 VPWR.n5 VPWR.t7 72.2026
R54 VPWR.n5 VPWR.t5 70.3576
R55 VPWR.n8 VPWR.t1 64.4945
R56 VPWR.n8 VPWR.t3 63.3219
R57 VPWR.n7 VPWR.t6 46.9053
R58 VPWR.n26 VPWR.n25 36.1417
R59 VPWR.n19 VPWR.n3 36.1417
R60 VPWR.n20 VPWR.n19 36.1417
R61 VPWR.n21 VPWR.n20 36.1417
R62 VPWR.n13 VPWR.n6 36.1417
R63 VPWR.n14 VPWR.n13 36.1417
R64 VPWR.n7 VPWR.t2 30.9824
R65 VPWR.n15 VPWR.n3 28.9887
R66 VPWR.n25 VPWR.n1 23.7181
R67 VPWR.n21 VPWR.n1 23.7181
R68 VPWR.n27 VPWR.n26 20.7064
R69 VPWR.n15 VPWR.n14 18.4476
R70 VPWR.n10 VPWR.n9 12.5175
R71 VPWR.n9 VPWR.n6 9.30841
R72 VPWR.n11 VPWR.n6 9.3005
R73 VPWR.n13 VPWR.n12 9.3005
R74 VPWR.n14 VPWR.n4 9.3005
R75 VPWR.n16 VPWR.n15 9.3005
R76 VPWR.n17 VPWR.n3 9.3005
R77 VPWR.n19 VPWR.n18 9.3005
R78 VPWR.n20 VPWR.n2 9.3005
R79 VPWR.n22 VPWR.n21 9.3005
R80 VPWR.n23 VPWR.n1 9.3005
R81 VPWR.n25 VPWR.n24 9.3005
R82 VPWR.n26 VPWR.n0 9.3005
R83 VPWR.n28 VPWR.n27 9.3005
R84 VPWR.n11 VPWR.n10 0.528998
R85 VPWR.n12 VPWR.n11 0.122949
R86 VPWR.n12 VPWR.n4 0.122949
R87 VPWR.n16 VPWR.n4 0.122949
R88 VPWR.n17 VPWR.n16 0.122949
R89 VPWR.n18 VPWR.n17 0.122949
R90 VPWR.n18 VPWR.n2 0.122949
R91 VPWR.n22 VPWR.n2 0.122949
R92 VPWR.n23 VPWR.n22 0.122949
R93 VPWR.n24 VPWR.n23 0.122949
R94 VPWR.n24 VPWR.n0 0.122949
R95 VPWR.n28 VPWR.n0 0.122949
R96 VPWR VPWR.n28 0.0617245
R97 CLK.n0 CLK.t0 302.432
R98 CLK.n1 CLK.t3 229.024
R99 CLK.n0 CLK.t2 205.654
R100 CLK.n0 CLK.t1 187.413
R101 CLK CLK.n1 153.808
R102 CLK.n1 CLK.n0 13.8763
R103 GCLK.n1 GCLK 589.572
R104 GCLK.n1 GCLK.n0 585
R105 GCLK.n2 GCLK.n1 585
R106 GCLK GCLK.t1 207.599
R107 GCLK.n1 GCLK.t0 41.3353
R108 GCLK GCLK.n2 12.2519
R109 GCLK GCLK.n0 10.6062
R110 GCLK GCLK.n0 2.92621
R111 GCLK.n2 GCLK 1.2805
R112 GATE.n0 GATE.t1 279.56
R113 GATE.n0 GATE.t0 205.922
R114 GATE GATE.n0 156.133
R115 a_116_424.t0 a_116_424.t1 56.2862
R116 VGND.n27 VGND.t3 258.041
R117 VGND.n2 VGND.n1 242.279
R118 VGND.n15 VGND.n6 219.636
R119 VGND.n10 VGND.t1 168.186
R120 VGND.n9 VGND.n8 128.262
R121 VGND.n6 VGND.t7 94.4201
R122 VGND.n1 VGND.t2 55.6369
R123 VGND.n6 VGND.t6 40.0005
R124 VGND.n13 VGND.n7 36.1417
R125 VGND.n14 VGND.n13 36.1417
R126 VGND.n16 VGND.n4 36.1417
R127 VGND.n20 VGND.n4 36.1417
R128 VGND.n21 VGND.n20 36.1417
R129 VGND.n22 VGND.n21 36.1417
R130 VGND.n8 VGND.t4 34.688
R131 VGND.n1 VGND.t0 30.0005
R132 VGND.n26 VGND.n25 29.3032
R133 VGND.n9 VGND.n7 27.8593
R134 VGND.n22 VGND.n2 26.854
R135 VGND.n27 VGND.n26 26.7299
R136 VGND.n8 VGND.t5 22.6611
R137 VGND.n15 VGND.n14 18.4476
R138 VGND.n16 VGND.n15 17.6946
R139 VGND.n28 VGND.n27 9.3005
R140 VGND.n11 VGND.n7 9.3005
R141 VGND.n13 VGND.n12 9.3005
R142 VGND.n14 VGND.n5 9.3005
R143 VGND.n17 VGND.n16 9.3005
R144 VGND.n18 VGND.n4 9.3005
R145 VGND.n20 VGND.n19 9.3005
R146 VGND.n21 VGND.n3 9.3005
R147 VGND.n23 VGND.n22 9.3005
R148 VGND.n25 VGND.n24 9.3005
R149 VGND.n26 VGND.n0 9.3005
R150 VGND.n10 VGND.n9 7.17905
R151 VGND.n25 VGND.n2 0.563137
R152 VGND.n11 VGND.n10 0.219196
R153 VGND.n12 VGND.n11 0.122949
R154 VGND.n12 VGND.n5 0.122949
R155 VGND.n17 VGND.n5 0.122949
R156 VGND.n18 VGND.n17 0.122949
R157 VGND.n19 VGND.n18 0.122949
R158 VGND.n19 VGND.n3 0.122949
R159 VGND.n23 VGND.n3 0.122949
R160 VGND.n24 VGND.n23 0.122949
R161 VGND.n24 VGND.n0 0.122949
R162 VGND.n28 VGND.n0 0.122949
R163 VGND VGND.n28 0.0617245
R164 VNB.n0 VNB 11502.4
R165 VNB VNB.n1 9426.85
R166 VNB.t9 VNB.t0 2864.04
R167 VNB.t8 VNB.t1 2482.94
R168 VNB.t10 VNB.n0 1639.45
R169 VNB.t0 VNB.t3 1362.73
R170 VNB.t2 VNB.t9 1166.4
R171 VNB.t4 VNB 1143.31
R172 VNB.t5 VNB.t6 1097.11
R173 VNB.t3 VNB.t4 993.177
R174 VNB.n1 VNB.t10 940.274
R175 VNB.t6 VNB.t8 831.496
R176 VNB.t7 VNB.t2 831.496
R177 VNB.n0 VNB.t5 692.913
R178 VNB.n1 VNB.t7 669.817
R179 a_288_48.t1 a_288_48.n2 854.054
R180 a_288_48.t2 a_288_48.t4 847.25
R181 a_288_48.n2 a_288_48.n1 474.83
R182 a_288_48.n0 a_288_48.t2 287.594
R183 a_288_48.n0 a_288_48.t3 274.74
R184 a_288_48.n1 a_288_48.t5 243.51
R185 a_288_48.n2 a_288_48.t0 136.482
R186 a_288_48.n1 a_288_48.n0 23.3962
R187 a_722_492.t0 a_722_492.t1 112.572
R188 a_1166_94.t0 a_1166_94.t1 39.3755
R189 SCE.n0 SCE.t0 222.381
R190 SCE.n0 SCE.t1 186.433
R191 SCE SCE.n0 68.9943
R192 a_667_80.t0 a_667_80.t1 60.0005
C0 GCLK VGND 0.10297f
C1 GCLK GATE 6.38e-21
C2 VPWR VGND 0.12394f
C3 SCE VGND 0.040567f
C4 GATE VPWR 0.021606f
C5 SCE GATE 0.108757f
C6 GCLK VPB 0.014765f
C7 VPB VPWR 0.238445f
C8 SCE VPB 0.061925f
C9 GCLK VPWR 0.112376f
C10 CLK VGND 0.05857f
C11 CLK GATE 6.84e-20
C12 SCE VPWR 0.054002f
C13 CLK VPB 0.118531f
C14 CLK VPWR 0.025319f
C15 GATE VGND 0.006389f
C16 VPB VGND 0.018746f
C17 GATE VPB 0.070379f
C18 GCLK VNB 0.111925f
C19 CLK VNB 0.216642f
C20 VGND VNB 0.957552f
C21 VPWR VNB 0.744094f
C22 GATE VNB 0.111932f
C23 SCE VNB 0.176884f
C24 VPB VNB 1.80926f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdlclkp_2 VNB VPB VPWR VGND GCLK CLK GATE SCE
X0 VGND.t5 a_706_317.t2 a_685_81.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1513 pd=1.27 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 a_708_451.t0 a_288_48.t2 a_580_74.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.1386 ps=1.215 w=0.42 l=0.15
X2 a_706_317.t0 a_580_74.t4 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1513 ps=1.27 w=0.74 l=0.15
X3 a_1195_374# CLK VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.2575 pd=1.515 as=0.194175 ps=1.51 w=1 l=0.15
X4 VPWR a_1195_374# GCLK VPB sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VGND.t7 a_1195_374# GCLK.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 GCLK.t0 a_1195_374# VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.237 ps=1.555 w=1.12 l=0.15
X7 a_114_424.t1 SCE.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1008 pd=1.08 as=0.2394 ps=2.25 w=0.84 l=0.15
X8 a_1195_374# a_706_317.t3 a_1198_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.0777 ps=0.95 w=0.74 l=0.15
X9 a_318_74.t1 a_288_48.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.189025 ps=1.41 w=0.74 l=0.15
X10 a_580_74.t2 a_288_48.t4 a_114_112.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.097375 pd=0.925 as=0.33275 ps=2.31 w=0.55 l=0.15
X11 GCLK.t1 a_1195_374# VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2035 ps=2.03 w=0.74 l=0.15
X12 a_706_317.t1 a_580_74.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1785 ps=1.495 w=1.12 l=0.15
X13 VPWR.t4 a_706_317.t4 a_1195_374# VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.555 as=0.2575 ps=1.515 w=1 l=0.15
X14 a_685_81.t0 a_318_74.t2 a_580_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.097375 ps=0.925 w=0.42 l=0.15
X15 a_1198_74.t0 CLK.t0 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.13135 ps=1.095 w=0.74 l=0.15
X16 VPWR.t3 CLK.t1 a_288_48.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.194175 pd=1.51 as=0.2394 ps=2.25 w=0.84 l=0.15
X17 a_114_112.t0 GATE.t0 a_114_424.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2394 pd=2.25 as=0.1008 ps=1.08 w=0.84 l=0.15
X18 VGND.t8 GATE.t1 a_114_112.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.189025 pd=1.41 as=0.077 ps=0.83 w=0.55 l=0.15
X19 a_318_74.t0 a_288_48.t5 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2394 pd=2.25 as=0.3807 ps=2.98 w=0.84 l=0.15
X20 VGND.t3 CLK.t2 a_288_48.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.13135 pd=1.095 as=0.2109 ps=2.05 w=0.74 l=0.15
X21 a_114_112.t3 SCE.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.15675 ps=1.67 w=0.55 l=0.15
X22 a_580_74.t3 a_318_74.t3 a_114_112.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.215 as=0.2394 ps=2.25 w=0.84 l=0.15
X23 VPWR.t5 a_706_317.t5 a_708_451.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1785 pd=1.495 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_706_317.n0 a_706_317.t2 330.858
R1 a_706_317.n3 a_706_317.n2 300.327
R2 a_706_317.n1 a_706_317.t0 272.901
R3 a_706_317.n2 a_706_317.t4 246.429
R4 a_706_317.t1 a_706_317.n3 220.625
R5 a_706_317.n1 a_706_317.n0 201.882
R6 a_706_317.n2 a_706_317.t3 197.427
R7 a_706_317.n0 a_706_317.t5 181.706
R8 a_706_317.n3 a_706_317.n1 11.0875
R9 a_685_81.t0 a_685_81.t1 68.5719
R10 VGND.n9 VGND.t6 288.366
R11 VGND.n34 VGND.t0 258.041
R12 VGND.n2 VGND.n1 242.279
R13 VGND.n22 VGND.n6 220.766
R14 VGND.n10 VGND.t7 180.566
R15 VGND.n15 VGND.n14 116.288
R16 VGND.n6 VGND.t4 95.9851
R17 VGND.n1 VGND.t8 55.6369
R18 VGND.n6 VGND.t5 40.0005
R19 VGND.n13 VGND.n12 36.1417
R20 VGND.n16 VGND.n7 36.1417
R21 VGND.n20 VGND.n7 36.1417
R22 VGND.n21 VGND.n20 36.1417
R23 VGND.n23 VGND.n4 36.1417
R24 VGND.n27 VGND.n4 36.1417
R25 VGND.n28 VGND.n27 36.1417
R26 VGND.n29 VGND.n28 36.1417
R27 VGND.n14 VGND.t3 34.0546
R28 VGND.n1 VGND.t1 30.0005
R29 VGND.n33 VGND.n32 29.3032
R30 VGND.n12 VGND.n9 28.9887
R31 VGND.n29 VGND.n2 26.854
R32 VGND.n23 VGND.n22 26.7299
R33 VGND.n34 VGND.n33 26.7299
R34 VGND.n14 VGND.t2 23.514
R35 VGND.n15 VGND.n13 10.5417
R36 VGND.n22 VGND.n21 9.41227
R37 VGND.n35 VGND.n34 9.3005
R38 VGND.n12 VGND.n11 9.3005
R39 VGND.n13 VGND.n8 9.3005
R40 VGND.n17 VGND.n16 9.3005
R41 VGND.n18 VGND.n7 9.3005
R42 VGND.n20 VGND.n19 9.3005
R43 VGND.n21 VGND.n5 9.3005
R44 VGND.n24 VGND.n23 9.3005
R45 VGND.n25 VGND.n4 9.3005
R46 VGND.n27 VGND.n26 9.3005
R47 VGND.n28 VGND.n3 9.3005
R48 VGND.n30 VGND.n29 9.3005
R49 VGND.n32 VGND.n31 9.3005
R50 VGND.n33 VGND.n0 9.3005
R51 VGND.n10 VGND.n9 6.75343
R52 VGND.n16 VGND.n15 0.753441
R53 VGND.n11 VGND.n10 0.577955
R54 VGND.n32 VGND.n2 0.563137
R55 VGND.n11 VGND.n8 0.122949
R56 VGND.n17 VGND.n8 0.122949
R57 VGND.n18 VGND.n17 0.122949
R58 VGND.n19 VGND.n18 0.122949
R59 VGND.n19 VGND.n5 0.122949
R60 VGND.n24 VGND.n5 0.122949
R61 VGND.n25 VGND.n24 0.122949
R62 VGND.n26 VGND.n25 0.122949
R63 VGND.n26 VGND.n3 0.122949
R64 VGND.n30 VGND.n3 0.122949
R65 VGND.n31 VGND.n30 0.122949
R66 VGND.n31 VGND.n0 0.122949
R67 VGND.n35 VGND.n0 0.122949
R68 VGND VGND.n35 0.0617245
R69 VNB.n0 VNB 13604.2
R70 VNB VNB.n1 9360.67
R71 VNB.t3 VNB.t2 3025.72
R72 VNB.t6 VNB.t5 2413.3
R73 VNB.t7 VNB.t9 2240.42
R74 VNB.n1 VNB.t6 1413.85
R75 VNB.t2 VNB.t11 1362.73
R76 VNB.t1 VNB.t3 1212.6
R77 VNB.t5 VNB.n0 1170.08
R78 VNB.t0 VNB 1143.31
R79 VNB.t9 VNB.t10 993.177
R80 VNB.t11 VNB.t0 993.177
R81 VNB.t8 VNB.t1 900.788
R82 VNB.t4 VNB.t7 831.496
R83 VNB.n1 VNB.t8 230.971
R84 VNB.n0 VNB.t4 29.6501
R85 a_288_48.t5 a_288_48.t2 892.504
R86 a_288_48.t0 a_288_48.n2 845.019
R87 a_288_48.n2 a_288_48.n1 478.959
R88 a_288_48.n0 a_288_48.t5 287.594
R89 a_288_48.n0 a_288_48.t3 261.887
R90 a_288_48.n1 a_288_48.t4 245.117
R91 a_288_48.n2 a_288_48.t1 132.03
R92 a_288_48.n1 a_288_48.n0 57.1362
R93 a_580_74.n3 a_580_74.n2 654.919
R94 a_580_74.n1 a_580_74.t5 259.572
R95 a_580_74.n2 a_580_74.n0 226.638
R96 a_580_74.n2 a_580_74.n1 224.471
R97 a_580_74.n1 a_580_74.t4 177.631
R98 a_580_74.n3 a_580_74.t1 105.537
R99 a_580_74.n0 a_580_74.t0 64.2862
R100 a_580_74.n4 a_580_74.t3 30.9603
R101 a_580_74.n0 a_580_74.t2 23.2811
R102 a_580_74.n5 a_580_74.n4 20.7373
R103 a_580_74.n4 a_580_74.n3 4.69098
R104 a_708_451.t0 a_708_451.t1 112.572
R105 VPB.n0 VPB 3008.33
R106 VPB.t4 VPB.t1 543.952
R107 VPB.t9 VPB.t4 505.646
R108 VPB.n0 VPB.t7 344.759
R109 VPB.t7 VPB.t8 298.791
R110 VPB.t5 VPB.t9 268.146
R111 VPB.t2 VPB 252.823
R112 VPB VPB.n0 229.391
R113 VPB.t1 VPB.t2 199.195
R114 VPB.n0 VPB.t5 191.532
R115 VPB.t0 VPB.t3 83.4151
R116 VPB.t6 VPB.t0 57.9273
R117 VPB.n0 VPB.t6 6.76688
R118 CLK.n1 CLK.n0 250.373
R119 CLK.n2 CLK.t1 195.697
R120 CLK CLK.n3 158.788
R121 CLK.n1 CLK.t0 156.431
R122 CLK.n2 CLK.t2 154.24
R123 CLK.n3 CLK.n1 58.4247
R124 CLK.n3 CLK.n2 13.146
R125 VPWR.n1 VPWR.t2 940.218
R126 VPWR.n6 VPWR.t3 924.703
R127 VPWR.n24 VPWR.t1 407.38
R128 VPWR.n12 VPWR.n5 341.337
R129 VPWR.n8 VPWR.n7 323.219
R130 VPWR.n5 VPWR.t5 106.68
R131 VPWR.n7 VPWR.t4 46.2955
R132 VPWR.n23 VPWR.n22 36.1417
R133 VPWR.n16 VPWR.n3 36.1417
R134 VPWR.n17 VPWR.n16 36.1417
R135 VPWR.n18 VPWR.n17 36.1417
R136 VPWR.n11 VPWR.n10 36.1417
R137 VPWR.n10 VPWR.n6 35.3887
R138 VPWR.n7 VPWR.t6 34.1481
R139 VPWR.n12 VPWR.n3 29.3652
R140 VPWR.n5 VPWR.t0 29.2495
R141 VPWR.n18 VPWR.n1 25.977
R142 VPWR.n12 VPWR.n11 24.0946
R143 VPWR.n22 VPWR.n1 21.4593
R144 VPWR.n24 VPWR.n23 21.4593
R145 VPWR.n10 VPWR.n9 9.3005
R146 VPWR.n11 VPWR.n4 9.3005
R147 VPWR.n13 VPWR.n12 9.3005
R148 VPWR.n14 VPWR.n3 9.3005
R149 VPWR.n16 VPWR.n15 9.3005
R150 VPWR.n17 VPWR.n2 9.3005
R151 VPWR.n19 VPWR.n18 9.3005
R152 VPWR.n20 VPWR.n1 9.3005
R153 VPWR.n22 VPWR.n21 9.3005
R154 VPWR.n23 VPWR.n0 9.3005
R155 VPWR.n25 VPWR.n24 9.3005
R156 VPWR.n8 VPWR.n6 6.16751
R157 VPWR.n9 VPWR.n8 0.286599
R158 VPWR.n9 VPWR.n4 0.122949
R159 VPWR.n13 VPWR.n4 0.122949
R160 VPWR.n14 VPWR.n13 0.122949
R161 VPWR.n15 VPWR.n14 0.122949
R162 VPWR.n15 VPWR.n2 0.122949
R163 VPWR.n19 VPWR.n2 0.122949
R164 VPWR.n20 VPWR.n19 0.122949
R165 VPWR.n21 VPWR.n20 0.122949
R166 VPWR.n21 VPWR.n0 0.122949
R167 VPWR.n25 VPWR.n0 0.122949
R168 VPWR VPWR.n25 0.0617245
R169 GCLK.n2 GCLK 589.508
R170 GCLK.n2 GCLK.n0 585
R171 GCLK.n3 GCLK.n2 585
R172 GCLK GCLK.n1 159.708
R173 GCLK.n2 GCLK.t0 26.3844
R174 GCLK.n1 GCLK.t2 22.7032
R175 GCLK.n1 GCLK.t1 22.7032
R176 GCLK GCLK.n3 12.0794
R177 GCLK GCLK.n0 10.4568
R178 GCLK GCLK.n0 2.88501
R179 GCLK.n3 GCLK 1.26247
R180 SCE.n0 SCE.t0 223.423
R181 SCE.n0 SCE.t1 187.47
R182 SCE SCE.n0 68.7345
R183 a_114_424.t0 a_114_424.t1 56.2862
R184 a_1198_74.t0 a_1198_74.t1 34.0546
R185 a_318_74.t0 a_318_74.n1 775.088
R186 a_318_74.n1 a_318_74.t1 335.356
R187 a_318_74.n0 a_318_74.t2 264.762
R188 a_318_74.n1 a_318_74.n0 200.66
R189 a_318_74.n0 a_318_74.t3 187.178
R190 a_114_112.n2 a_114_112.t1 467.647
R191 a_114_112.n1 a_114_112.t2 391.825
R192 a_114_112.t0 a_114_112.n2 352.685
R193 a_114_112.n1 a_114_112.n0 185
R194 a_114_112.n2 a_114_112.n1 144.784
R195 a_114_112.n0 a_114_112.t4 30.546
R196 a_114_112.n0 a_114_112.t3 30.546
R197 GATE.n0 GATE.t1 279.56
R198 GATE.n0 GATE.t0 205.922
R199 GATE GATE.n0 155.815
C0 VPWR GCLK 0.208654f
C1 VPWR SCE 0.053172f
C2 VGND a_1195_374# 0.163665f
C3 CLK a_1195_374# 0.012129f
C4 a_1195_374# GATE 1.2e-20
C5 VPB a_1195_374# 0.085583f
C6 CLK VGND 0.05319f
C7 VGND GATE 0.006436f
C8 VPB VGND 0.022745f
C9 CLK VPB 0.090857f
C10 VPB GATE 0.070858f
C11 GCLK a_1195_374# 0.160211f
C12 VPWR a_1195_374# 0.195394f
C13 GCLK VGND 0.138763f
C14 VPWR VGND 0.142946f
C15 CLK GCLK 9.74e-20
C16 VPWR CLK 0.02375f
C17 GCLK GATE 8.68e-21
C18 VGND SCE 0.040466f
C19 VPWR GATE 0.021789f
C20 VPB GCLK 0.00607f
C21 VPWR VPB 0.27935f
C22 SCE GATE 0.108966f
C23 VPB SCE 0.061074f
C24 VGND VNB 1.04505f
C25 GCLK VNB 0.029869f
C26 CLK VNB 0.197795f
C27 VPWR VNB 0.831112f
C28 GATE VNB 0.112665f
C29 SCE VNB 0.176901f
C30 VPB VNB 1.93073f
C31 a_1195_374# VNB 0.267998f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfxtp_1 VNB VPB VPWR VGND SCE Q CLK SCD D
X0 VGND.t6 SCD.t0 a_450_74.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 a_450_74.t0 SCE.t0 a_301_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.12495 ps=1.015 w=0.42 l=0.15
X2 VPWR.t0 SCE.t1 a_35_74.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.1888 ps=1.87 w=0.64 l=0.15
X3 a_630_74.t0 CLK.t0 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1212 ps=1.1 w=0.74 l=0.15
X4 VPWR.t6 a_1736_74.t1 a_1688_508.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1806 pd=1.435 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_1018_100.t1 a_630_74.t2 a_301_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 a_1202_508.t0 a_630_74.t3 a_1018_100.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0525 pd=0.67 as=0.0735 ps=0.77 w=0.42 l=0.15
X7 a_828_74.t0 a_630_74.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 a_1688_508.t1 a_828_74.t2 a_1520_74# VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.19635 ps=1.395 w=0.42 l=0.15
X9 a_412_464.t0 a_35_74.t2 a_301_74.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1248 pd=1.03 as=0.096 ps=0.94 w=0.64 l=0.15
X10 a_301_74.t1 D.t0 a_238_464.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 a_630_74.t1 CLK.t1 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2428 ps=1.68 w=1.12 l=0.15
X12 VPWR.t5 a_1239_74# a_1202_508.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.52 as=0.0525 ps=0.67 w=0.42 l=0.15
X13 a_301_74.t3 D.t1 a_223_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12495 pd=1.015 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 VPWR.t8 SCD.t1 a_412_464.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.2428 pd=1.68 as=0.1248 ps=1.03 w=0.64 l=0.15
X15 a_828_74.t1 a_630_74.t5 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.532 ps=3.19 w=1.12 l=0.15
X16 a_1154_100.t1 a_828_74.t3 a_1018_100.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.08925 pd=0.845 as=0.1113 ps=0.95 w=0.42 l=0.15
X17 a_1018_100.t3 a_828_74.t4 a_301_74.t4 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X18 VGND.t8 SCE.t2 a_35_74.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.07455 pd=0.775 as=0.1197 ps=1.41 w=0.42 l=0.15
X19 Q.t0 a_1736_74.t2 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1998 ps=2.02 w=0.74 l=0.15
X20 a_1520_74# a_828_74.t5 a_1239_74# VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.16115 pd=1.24 as=0.078375 ps=0.835 w=0.55 l=0.15
X21 a_1239_74# a_1018_100.t4 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.1848 ps=1.52 w=0.84 l=0.15
X22 Q.t1 a_1736_74.t3 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.3304 ps=2.83 w=1.12 l=0.15
X23 a_1736_74.t0 a_1520_74# VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1806 ps=1.435 w=0.84 l=0.15
X24 a_238_464.t0 SCE.t3 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X25 VGND.t5 a_1736_74.t4 a_1688_100.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1622 pd=1.245 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 VGND.t2 a_1239_74# a_1154_100.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.201375 pd=1.38 as=0.08925 ps=0.845 w=0.42 l=0.15
X27 a_1239_74# a_1018_100.t5 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.078375 pd=0.835 as=0.201375 ps=1.38 w=0.55 l=0.15
X28 a_1688_100.t1 a_630_74.t6 a_1520_74# VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.16115 ps=1.24 w=0.42 l=0.15
X29 a_223_74.t0 a_35_74.t3 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.07455 ps=0.775 w=0.42 l=0.15
R0 SCD.n0 SCD.t0 330.675
R1 SCD.n0 SCD.t1 201.492
R2 SCD SCD.n0 70.5016
R3 a_450_74.t0 a_450_74.t1 68.5719
R4 VGND.n4 VGND.t0 295.89
R5 VGND.n33 VGND.n3 226.256
R6 VGND.n21 VGND.n20 209.721
R7 VGND.n41 VGND.n40 206.916
R8 VGND.n11 VGND.t4 181.332
R9 VGND.n10 VGND.t5 150.793
R10 VGND.n20 VGND.t3 100.365
R11 VGND.n3 VGND.t6 62.2404
R12 VGND.n40 VGND.t1 61.4291
R13 VGND.n20 VGND.t2 50.8836
R14 VGND.n40 VGND.t8 40.0005
R15 VGND.n15 VGND.n14 36.1417
R16 VGND.n15 VGND.n8 36.1417
R17 VGND.n19 VGND.n8 36.1417
R18 VGND.n22 VGND.n6 36.1417
R19 VGND.n26 VGND.n6 36.1417
R20 VGND.n27 VGND.n26 36.1417
R21 VGND.n28 VGND.n27 36.1417
R22 VGND.n32 VGND.n31 36.1417
R23 VGND.n34 VGND.n1 36.1417
R24 VGND.n38 VGND.n1 36.1417
R25 VGND.n39 VGND.n38 36.1417
R26 VGND.n14 VGND.n13 31.5672
R27 VGND.n22 VGND.n21 28.9887
R28 VGND.n21 VGND.n19 24.4711
R29 VGND.n3 VGND.t7 22.7037
R30 VGND.n41 VGND.n39 21.4593
R31 VGND.n33 VGND.n32 19.577
R32 VGND.n34 VGND.n33 16.5652
R33 VGND.n11 VGND.n10 10.6313
R34 VGND.n39 VGND.n0 9.3005
R35 VGND.n38 VGND.n37 9.3005
R36 VGND.n36 VGND.n1 9.3005
R37 VGND.n35 VGND.n34 9.3005
R38 VGND.n32 VGND.n2 9.3005
R39 VGND.n31 VGND.n30 9.3005
R40 VGND.n29 VGND.n28 9.3005
R41 VGND.n27 VGND.n5 9.3005
R42 VGND.n26 VGND.n25 9.3005
R43 VGND.n24 VGND.n6 9.3005
R44 VGND.n23 VGND.n22 9.3005
R45 VGND.n21 VGND.n7 9.3005
R46 VGND.n19 VGND.n18 9.3005
R47 VGND.n17 VGND.n8 9.3005
R48 VGND.n16 VGND.n15 9.3005
R49 VGND.n14 VGND.n9 9.3005
R50 VGND.n13 VGND.n12 9.3005
R51 VGND.n42 VGND.n41 7.34058
R52 VGND.n31 VGND.n4 6.4005
R53 VGND.n28 VGND.n4 4.89462
R54 VGND.n13 VGND.n10 3.21591
R55 VGND.n12 VGND.n11 0.490927
R56 VGND VGND.n42 0.158861
R57 VGND.n42 VGND.n0 0.148926
R58 VGND.n12 VGND.n9 0.122949
R59 VGND.n16 VGND.n9 0.122949
R60 VGND.n17 VGND.n16 0.122949
R61 VGND.n18 VGND.n17 0.122949
R62 VGND.n18 VGND.n7 0.122949
R63 VGND.n23 VGND.n7 0.122949
R64 VGND.n24 VGND.n23 0.122949
R65 VGND.n25 VGND.n24 0.122949
R66 VGND.n25 VGND.n5 0.122949
R67 VGND.n29 VGND.n5 0.122949
R68 VGND.n30 VGND.n29 0.122949
R69 VGND.n30 VGND.n2 0.122949
R70 VGND.n35 VGND.n2 0.122949
R71 VGND.n36 VGND.n35 0.122949
R72 VGND.n37 VGND.n36 0.122949
R73 VGND.n37 VGND.n0 0.122949
R74 VNB.t10 VNB.t9 4157.48
R75 VNB.t12 VNB.t1 2286.61
R76 VNB.t1 VNB.t3 2194.23
R77 VNB.t14 VNB.t2 1940.16
R78 VNB.t6 VNB.t7 1893.96
R79 VNB.t5 VNB.t8 1720.73
R80 VNB.t3 VNB.t0 1570.6
R81 VNB.t0 VNB.t6 1328.08
R82 VNB VNB.t13 1235.7
R83 VNB.t11 VNB.t12 1177.95
R84 VNB.t13 VNB.t4 1166.4
R85 VNB.t7 VNB.t14 1004.72
R86 VNB.t2 VNB.t10 900.788
R87 VNB.t8 VNB.t11 900.788
R88 VNB.t4 VNB.t5 900.788
R89 SCE.n2 SCE.n1 491.933
R90 SCE.n0 SCE.t0 308.351
R91 SCE.n1 SCE.t3 287.594
R92 SCE SCE.n2 172.197
R93 SCE.n2 SCE.t2 144.601
R94 SCE.n1 SCE.t1 126.927
R95 SCE.n0 SCE 12.0894
R96 SCE SCE.n0 2.82647
R97 a_301_74.n1 a_301_74.t4 715.915
R98 a_301_74.n3 a_301_74.n2 379.43
R99 a_301_74.n2 a_301_74.n0 354.822
R100 a_301_74.n1 a_301_74.t2 353.014
R101 a_301_74.n0 a_301_74.t3 88.5719
R102 a_301_74.n0 a_301_74.t0 81.4291
R103 a_301_74.n2 a_301_74.n1 75.7614
R104 a_301_74.n3 a_301_74.t5 46.1724
R105 a_301_74.t1 a_301_74.n3 46.1724
R106 a_35_74.n0 a_35_74.t3 548.847
R107 a_35_74.t1 a_35_74.n1 362.56
R108 a_35_74.n0 a_35_74.t2 352.512
R109 a_35_74.n1 a_35_74.t0 292.719
R110 a_35_74.n1 a_35_74.n0 7.25383
R111 VPWR.n5 VPWR.t4 770.042
R112 VPWR.n22 VPWR.n21 629.155
R113 VPWR.n34 VPWR.n4 598.053
R114 VPWR.n13 VPWR.n12 585
R115 VPWR.n41 VPWR.n1 315.832
R116 VPWR.n11 VPWR.t7 265.065
R117 VPWR.n12 VPWR.t6 126.644
R118 VPWR.n12 VPWR.t3 120.781
R119 VPWR.n21 VPWR.t5 110.227
R120 VPWR.n4 VPWR.t8 98.5005
R121 VPWR.n21 VPWR.t2 78.566
R122 VPWR.n1 VPWR.t0 61.563
R123 VPWR.n4 VPWR.t9 56.0664
R124 VPWR.n1 VPWR.t1 46.1724
R125 VPWR.n35 VPWR.n2 36.1417
R126 VPWR.n39 VPWR.n2 36.1417
R127 VPWR.n40 VPWR.n39 36.1417
R128 VPWR.n23 VPWR.n7 36.1417
R129 VPWR.n27 VPWR.n7 36.1417
R130 VPWR.n28 VPWR.n27 36.1417
R131 VPWR.n29 VPWR.n28 36.1417
R132 VPWR.n15 VPWR.n9 36.1417
R133 VPWR.n19 VPWR.n9 36.1417
R134 VPWR.n20 VPWR.n19 36.1417
R135 VPWR.n15 VPWR.n14 34.092
R136 VPWR.n34 VPWR.n33 32.0005
R137 VPWR.n33 VPWR.n5 19.2005
R138 VPWR.n22 VPWR.n20 15.1
R139 VPWR.n29 VPWR.n5 14.6829
R140 VPWR.n13 VPWR.n11 11.0346
R141 VPWR.n41 VPWR.n40 10.9181
R142 VPWR.n14 VPWR.n10 9.3005
R143 VPWR.n16 VPWR.n15 9.3005
R144 VPWR.n17 VPWR.n9 9.3005
R145 VPWR.n19 VPWR.n18 9.3005
R146 VPWR.n20 VPWR.n8 9.3005
R147 VPWR.n24 VPWR.n23 9.3005
R148 VPWR.n25 VPWR.n7 9.3005
R149 VPWR.n27 VPWR.n26 9.3005
R150 VPWR.n28 VPWR.n6 9.3005
R151 VPWR.n30 VPWR.n29 9.3005
R152 VPWR.n31 VPWR.n5 9.3005
R153 VPWR.n33 VPWR.n32 9.3005
R154 VPWR.n34 VPWR.n3 9.3005
R155 VPWR.n36 VPWR.n35 9.3005
R156 VPWR.n37 VPWR.n2 9.3005
R157 VPWR.n39 VPWR.n38 9.3005
R158 VPWR.n40 VPWR.n0 9.3005
R159 VPWR.n42 VPWR.n41 8.08026
R160 VPWR.n14 VPWR.n13 4.18351
R161 VPWR.n23 VPWR.n22 3.80591
R162 VPWR.n35 VPWR.n34 2.25932
R163 VPWR.n11 VPWR.n10 0.480487
R164 VPWR VPWR.n42 0.163644
R165 VPWR.n42 VPWR.n0 0.144205
R166 VPWR.n16 VPWR.n10 0.122949
R167 VPWR.n17 VPWR.n16 0.122949
R168 VPWR.n18 VPWR.n17 0.122949
R169 VPWR.n18 VPWR.n8 0.122949
R170 VPWR.n24 VPWR.n8 0.122949
R171 VPWR.n25 VPWR.n24 0.122949
R172 VPWR.n26 VPWR.n25 0.122949
R173 VPWR.n26 VPWR.n6 0.122949
R174 VPWR.n30 VPWR.n6 0.122949
R175 VPWR.n31 VPWR.n30 0.122949
R176 VPWR.n32 VPWR.n31 0.122949
R177 VPWR.n32 VPWR.n3 0.122949
R178 VPWR.n36 VPWR.n3 0.122949
R179 VPWR.n37 VPWR.n36 0.122949
R180 VPWR.n38 VPWR.n37 0.122949
R181 VPWR.n38 VPWR.n0 0.122949
R182 VPB.t4 VPB.t3 720.162
R183 VPB.t13 VPB.t7 607.797
R184 VPB.t5 VPB.t11 515.861
R185 VPB.t7 VPB.t14 515.861
R186 VPB.t10 VPB.t5 380.512
R187 VPB.t12 VPB.t13 362.635
R188 VPB.t9 VPB.t4 316.668
R189 VPB VPB.t1 314.113
R190 VPB.t8 VPB.t12 275.807
R191 VPB.t14 VPB.t6 255.376
R192 VPB.t1 VPB.t0 255.376
R193 VPB.t2 VPB.t8 229.839
R194 VPB.t3 VPB.t10 214.517
R195 VPB.t0 VPB.t2 214.517
R196 VPB.t6 VPB.t9 204.302
R197 CLK.n0 CLK.t1 279.902
R198 CLK.n0 CLK.t0 186.543
R199 CLK CLK.n0 157.149
R200 a_630_74.t1 a_630_74.n6 881.284
R201 a_630_74.n2 a_630_74.n1 500.329
R202 a_630_74.n1 a_630_74.t6 400.353
R203 a_630_74.n3 a_630_74.n2 290.077
R204 a_630_74.n4 a_630_74.t5 260.281
R205 a_630_74.n3 a_630_74.t2 247.428
R206 a_630_74.n1 a_630_74.n0 213.954
R207 a_630_74.n5 a_630_74.t4 202.671
R208 a_630_74.n6 a_630_74.t0 191.245
R209 a_630_74.n2 a_630_74.t3 186.642
R210 a_630_74.n4 a_630_74.n3 160.667
R211 a_630_74.n6 a_630_74.n5 152
R212 a_630_74.n5 a_630_74.n4 75.0548
R213 a_1736_74.n0 a_1736_74.t1 451.474
R214 a_1736_74.t0 a_1736_74.n2 438.394
R215 a_1736_74.n1 a_1736_74.t3 234.841
R216 a_1736_74.n2 a_1736_74.n1 219.71
R217 a_1736_74.n2 a_1736_74.n0 212.532
R218 a_1736_74.n1 a_1736_74.t2 182.138
R219 a_1736_74.n0 a_1736_74.t4 147.046
R220 a_1688_508.t0 a_1688_508.t1 126.644
R221 a_1018_100.n2 a_1018_100.n0 660.91
R222 a_1018_100.n1 a_1018_100.t5 322.168
R223 a_1018_100.n2 a_1018_100.n1 244.999
R224 a_1018_100.n3 a_1018_100.n2 242.601
R225 a_1018_100.n1 a_1018_100.t4 205.149
R226 a_1018_100.n3 a_1018_100.t1 111.43
R227 a_1018_100.n0 a_1018_100.t3 93.81
R228 a_1018_100.n0 a_1018_100.t2 70.3576
R229 a_1018_100.t0 a_1018_100.n3 40.0005
R230 a_1202_508.t0 a_1202_508.t1 117.263
R231 a_828_74.t1 a_828_74.n3 860.985
R232 a_828_74.n0 a_828_74.t2 355.274
R233 a_828_74.n3 a_828_74.t4 329.805
R234 a_828_74.n0 a_828_74.t5 306.019
R235 a_828_74.n1 a_828_74.t3 298.12
R236 a_828_74.n2 a_828_74.t0 210.272
R237 a_828_74.n1 a_828_74.n0 196.894
R238 a_828_74.n3 a_828_74.n2 123.129
R239 a_828_74.n2 a_828_74.n1 75.5054
R240 a_412_464.t0 a_412_464.t1 120.047
R241 D.n0 D.t1 305.267
R242 D.n0 D.t0 274.204
R243 D D.n0 166.546
R244 a_238_464.t0 a_238_464.t1 83.1099
R245 a_223_74.t0 a_223_74.t1 68.5719
R246 a_1154_100.t0 a_1154_100.t1 121.43
R247 Q.n3 Q 589.777
R248 Q.n3 Q.n0 585
R249 Q.n4 Q.n3 585
R250 Q.n2 Q.t0 283.183
R251 Q.t0 Q.n1 283.183
R252 Q.n3 Q.t1 26.3844
R253 Q Q.n4 12.8005
R254 Q.n1 Q 11.6542
R255 Q Q.n0 11.0811
R256 Q Q.n2 8.59751
R257 Q.n2 Q 5.5408
R258 Q Q.n0 3.05722
R259 Q.n1 Q 2.48408
R260 Q.n4 Q 1.33781
R261 a_1688_100.t0 a_1688_100.t1 68.5719
C0 SCD VGND 0.008384f
C1 SCE VGND 0.083875f
C2 VPB VGND 0.025525f
C3 SCD SCE 0.038574f
C4 SCD VPB 0.084348f
C5 SCE VPB 0.149196f
C6 a_1239_74# VGND 0.02568f
C7 SCD a_1239_74# 1.3e-20
C8 a_1239_74# VPB 0.085984f
C9 Q VGND 0.101079f
C10 SCD Q 6.91e-22
C11 CLK VGND 0.01405f
C12 D VGND 0.012311f
C13 Q VPB 0.014051f
C14 SCD CLK 0.038587f
C15 VPWR VGND 0.180238f
C16 VPB CLK 0.046701f
C17 D SCD 0.003978f
C18 D SCE 0.11271f
C19 SCD VPWR 0.015011f
C20 VPWR SCE 0.042191f
C21 D VPB 0.067614f
C22 a_1520_74# VGND 0.095046f
C23 VPWR VPB 0.318428f
C24 SCD a_1520_74# 2.05e-20
C25 a_1520_74# VPB 0.101487f
C26 VPWR a_1239_74# 0.026096f
C27 a_1239_74# a_1520_74# 0.002102f
C28 VPWR Q 0.127488f
C29 VPWR CLK 0.017539f
C30 D VPWR 0.014497f
C31 Q a_1520_74# 9.27e-19
C32 VPWR a_1520_74# 0.121942f
C33 Q VNB 0.109281f
C34 VGND VNB 1.29371f
C35 CLK VNB 0.141261f
C36 SCD VNB 0.134264f
C37 D VNB 0.126573f
C38 SCE VNB 0.360563f
C39 VPWR VNB 0.998157f
C40 VPB VNB 2.54894f
C41 a_1520_74# VNB 0.160569f
C42 a_1239_74# VNB 0.159187f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfxtp_2 VNB VPB VPWR VGND SCE CLK D SCD Q
X0 a_634_74.t0 CLK.t0 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.28755 ps=1.85 w=1.12 l=0.15
X1 VPWR.t4 a_1829_398.t2 a_1704_496.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.21335 pd=1.65 as=0.1344 ps=1.06 w=0.42 l=0.15
X2 VPWR.t2 a_1287_320.t4 a_1210_508.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.16695 pd=1.37 as=0.084 ps=0.82 w=0.42 l=0.15
X3 a_634_74.t1 CLK.t1 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1338 ps=1.16 w=0.74 l=0.15
X4 a_1044_100.t1 a_634_74.t2 a_300_453.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.15225 pd=1.145 as=0.1197 ps=1.41 w=0.42 l=0.15
X5 a_1829_398.t0 a_1592_424.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1135 ps=1.09 w=0.74 l=0.15
X6 VGND.t6 a_1287_320.t5 a_1219_100# VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.225725 pd=1.45 as=0.0882 ps=0.84 w=0.42 l=0.15
X7 a_1287_320.t2 a_1044_100.t3 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.18975 pd=1.24 as=0.225725 ps=1.45 w=0.55 l=0.15
X8 a_1592_424.t1 a_846_74.t2 a_1287_320.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.094125 pd=0.91 as=0.18975 ps=1.24 w=0.55 l=0.15
X9 VGND.t5 SCD.t0 a_442_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1338 pd=1.16 as=0.0504 ps=0.66 w=0.42 l=0.15
X10 VPWR.t0 SCE.t0 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.1888 ps=1.87 w=0.64 l=0.15
X11 a_439_453.t1 a_27_74.t2 a_300_453.t5 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1744 ps=1.185 w=0.64 l=0.15
X12 VGND.t1 a_1829_398.t3 a_1787_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1135 pd=1.09 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 a_300_453.t0 D.t0 a_223_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=0.975 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 VGND.t4 SCE.t1 a_27_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1386 ps=1.5 w=0.42 l=0.15
X15 a_300_453.t4 D.t1 a_216_453.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1744 pd=1.185 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 VPWR.t5 a_1829_398.t4 Q.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_846_74.t0 a_634_74.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.6426 ps=3.56 w=1.12 l=0.15
X18 a_1210_508.t0 a_634_74.t4 a_1044_100.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.084 pd=0.82 as=0.063 ps=0.72 w=0.42 l=0.15
X19 a_1592_424.t0 a_634_74.t5 a_1287_320.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.14715 pd=1.25 as=0.2226 ps=1.37 w=0.84 l=0.15
X20 a_216_453.t1 SCE.t2 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X21 a_1044_100.t2 a_846_74.t3 a_300_453.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X22 a_1287_320.t3 a_1044_100.t4 VPWR.t8 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2226 pd=1.37 as=0.16695 ps=1.37 w=0.84 l=0.15
X23 a_846_74.t1 a_634_74.t6 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X24 VGND.t2 a_1829_398.t5 Q.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2294 pd=2.1 as=0.12025 ps=1.065 w=0.74 l=0.15
X25 a_1829_398.t1 a_1592_424.t4 VPWR.t9 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.21335 ps=1.65 w=1 l=0.15
X26 a_442_74.t0 SCE.t3 a_300_453.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.11655 ps=0.975 w=0.42 l=0.15
X27 VPWR.t6 SCD.t1 a_439_453.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.28755 pd=1.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_1704_496.t1 a_846_74.t4 a_1592_424.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.14715 ps=1.25 w=0.42 l=0.15
X29 a_223_74.t1 a_27_74.t3 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
R0 CLK.n0 CLK.t0 226.809
R1 CLK.n0 CLK.t1 223.036
R2 CLK CLK.n0 179.667
R3 VPWR.n32 VPWR.t3 795.26
R4 VPWR.n25 VPWR.n8 614.697
R5 VPWR.n40 VPWR.n39 604.701
R6 VPWR.n12 VPWR.n11 585
R7 VPWR.n14 VPWR.n13 585
R8 VPWR.n47 VPWR.n1 317.094
R9 VPWR.n15 VPWR.t5 266.863
R10 VPWR.n13 VPWR.n12 164.167
R11 VPWR.n8 VPWR.t8 146.577
R12 VPWR.n39 VPWR.t6 104.656
R13 VPWR.n12 VPWR.t4 70.3576
R14 VPWR.n8 VPWR.t2 70.3576
R15 VPWR.n1 VPWR.t0 61.563
R16 VPWR.n39 VPWR.t7 46.3183
R17 VPWR.n1 VPWR.t1 46.1724
R18 VPWR.n41 VPWR.n2 36.1417
R19 VPWR.n45 VPWR.n2 36.1417
R20 VPWR.n46 VPWR.n45 36.1417
R21 VPWR.n26 VPWR.n6 36.1417
R22 VPWR.n30 VPWR.n6 36.1417
R23 VPWR.n31 VPWR.n30 36.1417
R24 VPWR.n33 VPWR.n31 36.1417
R25 VPWR.n19 VPWR.n18 36.1417
R26 VPWR.n19 VPWR.n9 36.1417
R27 VPWR.n23 VPWR.n9 36.1417
R28 VPWR.n24 VPWR.n23 36.1417
R29 VPWR.n38 VPWR.n37 35.3195
R30 VPWR.n13 VPWR.t9 33.6312
R31 VPWR.n18 VPWR.n17 32.256
R32 VPWR.n37 VPWR.n4 26.2751
R33 VPWR.n47 VPWR.n46 19.2005
R34 VPWR.n33 VPWR.n32 19.1192
R35 VPWR.n25 VPWR.n24 9.41227
R36 VPWR.n17 VPWR.n16 9.3005
R37 VPWR.n18 VPWR.n10 9.3005
R38 VPWR.n20 VPWR.n19 9.3005
R39 VPWR.n21 VPWR.n9 9.3005
R40 VPWR.n23 VPWR.n22 9.3005
R41 VPWR.n24 VPWR.n7 9.3005
R42 VPWR.n27 VPWR.n26 9.3005
R43 VPWR.n28 VPWR.n6 9.3005
R44 VPWR.n30 VPWR.n29 9.3005
R45 VPWR.n31 VPWR.n5 9.3005
R46 VPWR.n34 VPWR.n33 9.3005
R47 VPWR.n35 VPWR.n4 9.3005
R48 VPWR.n37 VPWR.n36 9.3005
R49 VPWR.n38 VPWR.n3 9.3005
R50 VPWR.n42 VPWR.n41 9.3005
R51 VPWR.n43 VPWR.n2 9.3005
R52 VPWR.n45 VPWR.n44 9.3005
R53 VPWR.n46 VPWR.n0 9.3005
R54 VPWR.n41 VPWR.n40 7.99674
R55 VPWR.n15 VPWR.n14 7.9067
R56 VPWR.n26 VPWR.n25 7.90638
R57 VPWR.n48 VPWR.n47 7.43488
R58 VPWR.n14 VPWR.n11 5.4308
R59 VPWR.n40 VPWR.n38 4.3013
R60 VPWR.n17 VPWR.n11 1.55202
R61 VPWR.n32 VPWR.n4 1.1269
R62 VPWR.n16 VPWR.n15 0.170963
R63 VPWR VPWR.n48 0.160103
R64 VPWR.n48 VPWR.n0 0.1477
R65 VPWR.n16 VPWR.n10 0.122949
R66 VPWR.n20 VPWR.n10 0.122949
R67 VPWR.n21 VPWR.n20 0.122949
R68 VPWR.n22 VPWR.n21 0.122949
R69 VPWR.n22 VPWR.n7 0.122949
R70 VPWR.n27 VPWR.n7 0.122949
R71 VPWR.n28 VPWR.n27 0.122949
R72 VPWR.n29 VPWR.n28 0.122949
R73 VPWR.n29 VPWR.n5 0.122949
R74 VPWR.n34 VPWR.n5 0.122949
R75 VPWR.n35 VPWR.n34 0.122949
R76 VPWR.n36 VPWR.n35 0.122949
R77 VPWR.n36 VPWR.n3 0.122949
R78 VPWR.n42 VPWR.n3 0.122949
R79 VPWR.n43 VPWR.n42 0.122949
R80 VPWR.n44 VPWR.n43 0.122949
R81 VPWR.n44 VPWR.n0 0.122949
R82 a_634_74.t0 a_634_74.n6 815.929
R83 a_634_74.n1 a_634_74.n0 580.299
R84 a_634_74.n2 a_634_74.n1 552.677
R85 a_634_74.n3 a_634_74.n2 402.046
R86 a_634_74.n4 a_634_74.t3 240.197
R87 a_634_74.n1 a_634_74.t5 213.954
R88 a_634_74.n6 a_634_74.t1 186.19
R89 a_634_74.n4 a_634_74.n3 184.101
R90 a_634_74.n6 a_634_74.n5 170.222
R91 a_634_74.n3 a_634_74.t2 163.881
R92 a_634_74.n2 a_634_74.t4 159.155
R93 a_634_74.n5 a_634_74.t6 154.24
R94 a_634_74.n5 a_634_74.n4 42.3225
R95 VPB.t15 VPB.t7 745.699
R96 VPB.t9 VPB.t3 630.78
R97 VPB.t3 VPB.t10 515.861
R98 VPB.t6 VPB.t15 408.603
R99 VPB.t11 VPB.t6 403.495
R100 VPB.t8 VPB.t9 377.957
R101 VPB.t12 VPB.t13 354.974
R102 VPB.t14 VPB.t1 347.312
R103 VPB.t5 VPB.t14 347.312
R104 VPB.t1 VPB.t11 286.022
R105 VPB.t2 VPB.t5 280.914
R106 VPB VPB.t0 257.93
R107 VPB.t0 VPB.t4 255.376
R108 VPB.t10 VPB.t2 229.839
R109 VPB.t13 VPB.t8 214.517
R110 VPB.t4 VPB.t12 214.517
R111 a_1829_398.t1 a_1829_398.n7 848.663
R112 a_1829_398.n5 a_1829_398.t3 341.818
R113 a_1829_398.n2 a_1829_398.t4 263.81
R114 a_1829_398.n3 a_1829_398.n1 261.62
R115 a_1829_398.n5 a_1829_398.t2 252.113
R116 a_1829_398.n6 a_1829_398.n5 196.505
R117 a_1829_398.n4 a_1829_398.n0 154.24
R118 a_1829_398.n2 a_1829_398.t5 154.24
R119 a_1829_398.n6 a_1829_398.t0 151.471
R120 a_1829_398.n7 a_1829_398.n4 112.749
R121 a_1829_398.n3 a_1829_398.n2 63.5369
R122 a_1829_398.n7 a_1829_398.n6 28.2358
R123 a_1829_398.n4 a_1829_398.n3 5.84292
R124 a_1704_496.t0 a_1704_496.t1 300.19
R125 a_1287_320.n3 a_1287_320.n2 661.801
R126 a_1287_320.n1 a_1287_320.t4 391.053
R127 a_1287_320.n2 a_1287_320.n0 206.425
R128 a_1287_320.n0 a_1287_320.t1 120.001
R129 a_1287_320.n2 a_1287_320.n1 116.638
R130 a_1287_320.n1 a_1287_320.t5 112.468
R131 a_1287_320.t0 a_1287_320.n3 89.1195
R132 a_1287_320.n3 a_1287_320.t3 35.1791
R133 a_1287_320.n0 a_1287_320.t2 30.546
R134 a_1210_508.t0 a_1210_508.t1 187.619
R135 VGND.n3 VGND.t3 242.133
R136 VGND.n34 VGND.n33 213.554
R137 VGND.n11 VGND.n10 207.498
R138 VGND.n42 VGND.n41 205.752
R139 VGND.n20 VGND.n8 199.934
R140 VGND.n12 VGND.t2 167.74
R141 VGND.n8 VGND.t9 120.001
R142 VGND.n33 VGND.t5 72.8576
R143 VGND.n41 VGND.t4 60.0005
R144 VGND.n8 VGND.t6 53.0654
R145 VGND.n10 VGND.t0 44.5565
R146 VGND.n10 VGND.t1 40.0005
R147 VGND.n41 VGND.t8 40.0005
R148 VGND.n15 VGND.n14 36.1417
R149 VGND.n16 VGND.n15 36.1417
R150 VGND.n16 VGND.n7 36.1417
R151 VGND.n22 VGND.n21 36.1417
R152 VGND.n22 VGND.n5 36.1417
R153 VGND.n26 VGND.n5 36.1417
R154 VGND.n27 VGND.n26 36.1417
R155 VGND.n28 VGND.n27 36.1417
R156 VGND.n32 VGND.n31 36.1417
R157 VGND.n35 VGND.n1 36.1417
R158 VGND.n39 VGND.n1 36.1417
R159 VGND.n40 VGND.n39 36.1417
R160 VGND.n14 VGND.n11 31.624
R161 VGND.n20 VGND.n7 29.3652
R162 VGND.n33 VGND.t7 29.2283
R163 VGND.n21 VGND.n20 18.0711
R164 VGND.n42 VGND.n40 15.8123
R165 VGND.n34 VGND.n32 10.9181
R166 VGND.n40 VGND.n0 9.3005
R167 VGND.n39 VGND.n38 9.3005
R168 VGND.n37 VGND.n1 9.3005
R169 VGND.n36 VGND.n35 9.3005
R170 VGND.n32 VGND.n2 9.3005
R171 VGND.n31 VGND.n30 9.3005
R172 VGND.n29 VGND.n28 9.3005
R173 VGND.n27 VGND.n4 9.3005
R174 VGND.n26 VGND.n25 9.3005
R175 VGND.n24 VGND.n5 9.3005
R176 VGND.n23 VGND.n22 9.3005
R177 VGND.n21 VGND.n6 9.3005
R178 VGND.n20 VGND.n19 9.3005
R179 VGND.n18 VGND.n7 9.3005
R180 VGND.n17 VGND.n16 9.3005
R181 VGND.n15 VGND.n9 9.3005
R182 VGND.n14 VGND.n13 9.3005
R183 VGND.n31 VGND.n3 7.90638
R184 VGND.n43 VGND.n42 7.56047
R185 VGND.n12 VGND.n11 6.62356
R186 VGND.n35 VGND.n34 5.64756
R187 VGND.n28 VGND.n3 3.38874
R188 VGND.n13 VGND.n12 0.171418
R189 VGND VGND.n43 0.161757
R190 VGND.n43 VGND.n0 0.146068
R191 VGND.n13 VGND.n9 0.122949
R192 VGND.n17 VGND.n9 0.122949
R193 VGND.n18 VGND.n17 0.122949
R194 VGND.n19 VGND.n18 0.122949
R195 VGND.n19 VGND.n6 0.122949
R196 VGND.n23 VGND.n6 0.122949
R197 VGND.n24 VGND.n23 0.122949
R198 VGND.n25 VGND.n24 0.122949
R199 VGND.n25 VGND.n4 0.122949
R200 VGND.n29 VGND.n4 0.122949
R201 VGND.n30 VGND.n29 0.122949
R202 VGND.n30 VGND.n2 0.122949
R203 VGND.n36 VGND.n2 0.122949
R204 VGND.n37 VGND.n36 0.122949
R205 VGND.n38 VGND.n37 0.122949
R206 VGND.n38 VGND.n0 0.122949
R207 VNB.t0 VNB.t1 3995.8
R208 VNB.t5 VNB.t9 3337.53
R209 VNB.t10 VNB.t4 2448.29
R210 VNB.t4 VNB.t5 2286.61
R211 VNB.t9 VNB.t13 2124.93
R212 VNB.t11 VNB.t2 2078.74
R213 VNB.t13 VNB.t11 1940.16
R214 VNB.t3 VNB.t6 1628.35
R215 VNB.t8 VNB.t10 1316.54
R216 VNB VNB.t7 1247.24
R217 VNB.t2 VNB.t0 1154.86
R218 VNB.t7 VNB.t12 1154.86
R219 VNB.t6 VNB.t8 900.788
R220 VNB.t12 VNB.t3 900.788
R221 a_300_453.n1 a_300_453.t3 721.707
R222 a_300_453.n2 a_300_453.n0 367.988
R223 a_300_453.n1 a_300_453.t1 362.486
R224 a_300_453.n3 a_300_453.n2 341.481
R225 a_300_453.n2 a_300_453.n1 100.483
R226 a_300_453.n3 a_300_453.t5 84.6489
R227 a_300_453.t4 a_300_453.n3 83.1099
R228 a_300_453.n0 a_300_453.t2 80.0005
R229 a_300_453.n0 a_300_453.t0 78.5719
R230 a_1044_100.n2 a_1044_100.n1 652.336
R231 a_1044_100.t1 a_1044_100.n2 350.479
R232 a_1044_100.n0 a_1044_100.t3 345.072
R233 a_1044_100.n2 a_1044_100.n0 267.447
R234 a_1044_100.n0 a_1044_100.t4 181.821
R235 a_1044_100.n1 a_1044_100.t0 70.3576
R236 a_1044_100.n1 a_1044_100.t2 70.3576
R237 a_1592_424.n2 a_1592_424.n1 661.066
R238 a_1592_424.n1 a_1592_424.t1 324.368
R239 a_1592_424.n1 a_1592_424.n0 234.927
R240 a_1592_424.n0 a_1592_424.t4 230.251
R241 a_1592_424.n0 a_1592_424.t3 218.737
R242 a_1592_424.n2 a_1592_424.t2 121.953
R243 a_1592_424.n3 a_1592_424.t0 28.9657
R244 a_1592_424.n4 a_1592_424.n3 24.8712
R245 a_1592_424.n3 a_1592_424.n2 6.44979
R246 a_846_74.t0 a_846_74.n4 832.554
R247 a_846_74.n0 a_846_74.t4 347.661
R248 a_846_74.n0 a_846_74.t2 299.813
R249 a_846_74.n2 a_846_74.n1 294.055
R250 a_846_74.n4 a_846_74.t3 279.875
R251 a_846_74.n2 a_846_74.n0 213.912
R252 a_846_74.n3 a_846_74.t1 206.231
R253 a_846_74.n4 a_846_74.n3 96.6149
R254 a_846_74.n3 a_846_74.n2 82.7328
R255 SCD.n1 SCD.t0 298.841
R256 SCD.n2 SCD.t1 173.788
R257 SCD.n1 SCD.n0 152
R258 SCD.n3 SCD.n2 152
R259 SCD.n2 SCD.n1 49.6611
R260 SCD.n3 SCD.n0 13.1884
R261 SCD.n0 SCD 0.776258
R262 SCD SCD.n3 0.388379
R263 a_442_74.t0 a_442_74.t1 68.5719
R264 SCE.n1 SCE.n0 398.745
R265 SCE SCE.t3 368.526
R266 SCE.n0 SCE.t2 287.594
R267 SCE SCE.n1 153.371
R268 SCE.n1 SCE.t1 126.927
R269 SCE.n0 SCE.t0 126.927
R270 a_27_74.n0 a_27_74.t3 480.344
R271 a_27_74.n0 a_27_74.t2 406.553
R272 a_27_74.t0 a_27_74.n1 362.017
R273 a_27_74.n1 a_27_74.t1 302.995
R274 a_27_74.n1 a_27_74.n0 8.68302
R275 a_439_453.t0 a_439_453.t1 83.1099
R276 D.n0 D.t1 260.738
R277 D.n0 D.t0 241.458
R278 D D.n0 72.8528
R279 a_223_74.t0 a_223_74.t1 68.5719
R280 a_216_453.t0 a_216_453.t1 83.1099
R281 Q.n1 Q 589.85
R282 Q.n1 Q.n0 585
R283 Q.n2 Q.n1 585
R284 Q Q.t1 204.582
R285 Q.n1 Q.t0 26.3844
R286 Q Q.n2 12.9944
R287 Q Q.n0 11.249
R288 Q Q.n0 3.10353
R289 Q.n2 Q 1.35808
C0 SCD VGND 0.009799f
C1 SCE SCD 0.038f
C2 VPWR CLK 0.016221f
C3 SCE VGND 0.076199f
C4 VPWR Q 0.216091f
C5 D VPWR 0.014061f
C6 VPB CLK 0.055255f
C7 VPWR SCD 0.012105f
C8 a_1219_100# VGND 0.003592f
C9 VPWR VGND 0.199731f
C10 VPB Q 0.006878f
C11 SCE VPWR 0.036298f
C12 D VPB 0.07144f
C13 VPB SCD 0.08297f
C14 VPB VGND 0.027791f
C15 SCE VPB 0.128469f
C16 a_1219_100# VPWR 4.73e-19
C17 SCD CLK 0.041841f
C18 CLK VGND 0.014465f
C19 D SCD 0.02092f
C20 VGND Q 0.161374f
C21 VPB VPWR 0.361172f
C22 D VGND 0.013582f
C23 SCE D 0.11554f
C24 Q VNB 0.031378f
C25 VGND VNB 1.43297f
C26 CLK VNB 0.137833f
C27 SCD VNB 0.138625f
C28 D VNB 0.142938f
C29 SCE VNB 0.341782f
C30 VPWR VNB 1.13056f
C31 VPB VNB 2.76322f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfxtp_4 VNB VPB VPWR VGND SCE CLK D SCD Q
X0 a_452_74.t1 SCE.t0 a_301_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.12705 ps=1.025 w=0.42 l=0.15
X1 VGND.t6 a_1814_48.t2 a_1766_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 VPWR.t9 SCE.t1 a_36_74.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.1888 ps=1.87 w=0.64 l=0.15
X3 a_630_74.t1 CLK.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1135 ps=1.09 w=0.74 l=0.15
X4 VPWR.t5 a_1814_48.t3 a_1764_476.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.195 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_828_74.t1 a_630_74.t2 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 Q.t5 a_1814_48.t4 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.13505 pd=1.105 as=0.12025 ps=1.065 w=0.74 l=0.15
X7 a_1764_476.t0 a_828_74.t2 a_1587_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1449 ps=1.23 w=0.42 l=0.15
X8 a_828_74.t0 a_630_74.t3 VPWR.t11 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.6216 ps=3.35 w=1.12 l=0.15
X9 VGND.t4 a_1814_48.t5 Q.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_412_464.t0 a_36_74.t2 a_301_74.t4 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1248 pd=1.03 as=0.096 ps=0.94 w=0.64 l=0.15
X11 a_301_74.t1 D.t0 a_238_464.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 a_301_74.t2 D.t1 a_223_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12705 pd=1.025 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 VGND.t3 SCD.t0 a_452_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1135 pd=1.09 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 a_1814_48.t0 a_1587_74.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1302 ps=1.195 w=0.84 l=0.15
X15 VPWR.t10 SCD.t1 a_412_464.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.2524 pd=1.71 as=0.1248 ps=1.03 w=0.64 l=0.15
X16 a_630_74.t0 CLK.t1 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2524 ps=1.71 w=1.12 l=0.15
X17 VGND.t8 SCE.t2 a_36_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X18 VPWR.t6 a_1814_48.t6 Q.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_1026_100.t0 a_630_74.t4 a_301_74.t5 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1197 ps=1.41 w=0.42 l=0.15
X20 a_1257_74.t1 a_1026_100.t4 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.74 as=0.185075 ps=1.52 w=0.84 l=0.15
X21 a_1766_74.t1 a_630_74.t5 a_1587_74.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.2 ps=1.295 w=0.42 l=0.15
X22 a_1214_506.t0 a_630_74.t6 a_1026_100.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.063 ps=0.72 w=0.42 l=0.15
X23 Q.t3 a_1814_48.t7 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_1026_100.t2 a_828_74.t3 a_301_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X25 a_1587_74.t2 a_630_74.t7 a_1257_74.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1449 pd=1.23 as=0.378 ps=1.74 w=0.84 l=0.15
X26 VPWR.t0 a_1257_74.t2 a_1214_506.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.185075 pd=1.52 as=0.0819 ps=0.81 w=0.42 l=0.15
X27 a_238_464.t1 SCE.t3 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X28 a_1162_100.t0 a_828_74.t4 a_1026_100.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.09975 pd=0.895 as=0.1113 ps=0.95 w=0.42 l=0.15
X29 VGND.t1 a_1587_74.t4 a_1814_48.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X30 VPWR.t4 a_1814_48.t8 Q.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X31 Q.t0 a_1814_48.t9 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1862 ps=1.475 w=1.12 l=0.15
X32 a_223_74.t1 a_36_74.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
R0 SCE.n1 SCE.n0 434.092
R1 SCE.n0 SCE.t3 287.594
R2 SCE SCE.t0 286.683
R3 SCE SCE.n1 190.627
R4 SCE.n1 SCE.t2 144.601
R5 SCE.n0 SCE.t1 126.927
R6 a_301_74.n1 a_301_74.t0 709.611
R7 a_301_74.n2 a_301_74.n0 379.906
R8 a_301_74.n3 a_301_74.n2 378.209
R9 a_301_74.n1 a_301_74.t5 340.878
R10 a_301_74.n2 a_301_74.n1 105.412
R11 a_301_74.n0 a_301_74.t3 87.1434
R12 a_301_74.n0 a_301_74.t2 85.7148
R13 a_301_74.n3 a_301_74.t4 46.1724
R14 a_301_74.t1 a_301_74.n3 46.1724
R15 a_452_74.t0 a_452_74.t1 68.5719
R16 VNB.t1 VNB.t12 6975.33
R17 VNB.t8 VNB.t2 2286.61
R18 VNB.t13 VNB.t14 2286.61
R19 VNB.t3 VNB.t13 2286.61
R20 VNB.t9 VNB.t11 2182.68
R21 VNB.t5 VNB.t7 1743.83
R22 VNB.t14 VNB.t1 1570.6
R23 VNB VNB.t6 1247.24
R24 VNB.t4 VNB.t3 1154.86
R25 VNB.t6 VNB.t0 1154.86
R26 VNB.t2 VNB.t9 1097.11
R27 VNB.t11 VNB.t10 993.177
R28 VNB.t12 VNB.t8 900.788
R29 VNB.t7 VNB.t4 900.788
R30 VNB.t0 VNB.t5 900.788
R31 a_1814_48.t0 a_1814_48.n15 412.577
R32 a_1814_48.n0 a_1814_48.t3 387.743
R33 a_1814_48.n5 a_1814_48.t6 240.197
R34 a_1814_48.n7 a_1814_48.n4 240.197
R35 a_1814_48.n10 a_1814_48.t8 240.197
R36 a_1814_48.n12 a_1814_48.t9 240.197
R37 a_1814_48.n1 a_1814_48.n0 223.22
R38 a_1814_48.n12 a_1814_48.t4 182.138
R39 a_1814_48.n5 a_1814_48.t5 181.407
R40 a_1814_48.n9 a_1814_48.n3 179.947
R41 a_1814_48.n6 a_1814_48.t7 179.947
R42 a_1814_48.n8 a_1814_48.n2 165.189
R43 a_1814_48.n1 a_1814_48.t1 160.28
R44 a_1814_48.n14 a_1814_48.n13 152
R45 a_1814_48.n11 a_1814_48.n2 152
R46 a_1814_48.n0 a_1814_48.t2 108.6
R47 a_1814_48.n6 a_1814_48.n5 61.346
R48 a_1814_48.n13 a_1814_48.n11 49.6611
R49 a_1814_48.n9 a_1814_48.n8 37.246
R50 a_1814_48.n15 a_1814_48.n14 25.2126
R51 a_1814_48.n8 a_1814_48.n7 21.1793
R52 a_1814_48.n14 a_1814_48.n2 13.1884
R53 a_1814_48.n13 a_1814_48.n12 10.955
R54 a_1814_48.n15 a_1814_48.n1 9.78874
R55 a_1814_48.n10 a_1814_48.n9 7.30353
R56 a_1814_48.n11 a_1814_48.n10 5.11262
R57 a_1814_48.n7 a_1814_48.n6 4.38232
R58 a_1766_74.t0 a_1766_74.t1 68.5719
R59 VGND.n11 VGND.t7 295.558
R60 VGND.n3 VGND.t9 286.334
R61 VGND.n12 VGND.t4 285.219
R62 VGND.n9 VGND.t6 245.946
R63 VGND.n41 VGND.n40 214.696
R64 VGND.n49 VGND.n48 206.916
R65 VGND.n16 VGND.n15 115.245
R66 VGND.n48 VGND.t8 60.0005
R67 VGND.n40 VGND.t2 44.5565
R68 VGND.n40 VGND.t3 40.0005
R69 VGND.n48 VGND.t0 40.0005
R70 VGND.n22 VGND.n21 36.1417
R71 VGND.n23 VGND.n22 36.1417
R72 VGND.n23 VGND.n7 36.1417
R73 VGND.n27 VGND.n7 36.1417
R74 VGND.n29 VGND.n28 36.1417
R75 VGND.n29 VGND.n5 36.1417
R76 VGND.n33 VGND.n5 36.1417
R77 VGND.n34 VGND.n33 36.1417
R78 VGND.n35 VGND.n34 36.1417
R79 VGND.n39 VGND.n38 36.1417
R80 VGND.n42 VGND.n1 36.1417
R81 VGND.n46 VGND.n1 36.1417
R82 VGND.n47 VGND.n46 36.1417
R83 VGND.n15 VGND.t5 30.0005
R84 VGND.n14 VGND.n11 28.2358
R85 VGND.n17 VGND.n16 25.977
R86 VGND.n17 VGND.n9 23.7181
R87 VGND.n21 VGND.n9 23.7181
R88 VGND.n15 VGND.t1 22.7032
R89 VGND.n16 VGND.n14 21.4593
R90 VGND.n49 VGND.n47 15.8123
R91 VGND.n41 VGND.n39 12.424
R92 VGND.n28 VGND.n27 11.2946
R93 VGND.n14 VGND.n13 9.3005
R94 VGND.n16 VGND.n10 9.3005
R95 VGND.n18 VGND.n17 9.3005
R96 VGND.n19 VGND.n9 9.3005
R97 VGND.n21 VGND.n20 9.3005
R98 VGND.n22 VGND.n8 9.3005
R99 VGND.n24 VGND.n23 9.3005
R100 VGND.n25 VGND.n7 9.3005
R101 VGND.n27 VGND.n26 9.3005
R102 VGND.n28 VGND.n6 9.3005
R103 VGND.n30 VGND.n29 9.3005
R104 VGND.n31 VGND.n5 9.3005
R105 VGND.n33 VGND.n32 9.3005
R106 VGND.n34 VGND.n4 9.3005
R107 VGND.n36 VGND.n35 9.3005
R108 VGND.n38 VGND.n37 9.3005
R109 VGND.n39 VGND.n2 9.3005
R110 VGND.n43 VGND.n42 9.3005
R111 VGND.n44 VGND.n1 9.3005
R112 VGND.n46 VGND.n45 9.3005
R113 VGND.n47 VGND.n0 9.3005
R114 VGND.n50 VGND.n49 7.56047
R115 VGND.n38 VGND.n3 6.4005
R116 VGND.n12 VGND.n11 6.26985
R117 VGND.n35 VGND.n3 4.89462
R118 VGND.n42 VGND.n41 4.89462
R119 VGND.n13 VGND.n12 0.733933
R120 VGND VGND.n50 0.161757
R121 VGND.n50 VGND.n0 0.146068
R122 VGND.n13 VGND.n10 0.122949
R123 VGND.n18 VGND.n10 0.122949
R124 VGND.n19 VGND.n18 0.122949
R125 VGND.n20 VGND.n19 0.122949
R126 VGND.n20 VGND.n8 0.122949
R127 VGND.n24 VGND.n8 0.122949
R128 VGND.n25 VGND.n24 0.122949
R129 VGND.n26 VGND.n25 0.122949
R130 VGND.n26 VGND.n6 0.122949
R131 VGND.n30 VGND.n6 0.122949
R132 VGND.n31 VGND.n30 0.122949
R133 VGND.n32 VGND.n31 0.122949
R134 VGND.n32 VGND.n4 0.122949
R135 VGND.n36 VGND.n4 0.122949
R136 VGND.n37 VGND.n36 0.122949
R137 VGND.n37 VGND.n2 0.122949
R138 VGND.n43 VGND.n2 0.122949
R139 VGND.n44 VGND.n43 0.122949
R140 VGND.n45 VGND.n44 0.122949
R141 VGND.n45 VGND.n0 0.122949
R142 a_36_74.n0 a_36_74.t3 498.019
R143 a_36_74.t0 a_36_74.n1 362.56
R144 a_36_74.n0 a_36_74.t2 345.736
R145 a_36_74.n1 a_36_74.t1 290.872
R146 a_36_74.n1 a_36_74.n0 9.17383
R147 VPWR.n37 VPWR.t11 732.307
R148 VPWR.n30 VPWR.n29 631.747
R149 VPWR.n21 VPWR.n11 613.703
R150 VPWR.n45 VPWR.n44 585
R151 VPWR.n15 VPWR.t3 401.68
R152 VPWR.n14 VPWR.t4 351.639
R153 VPWR.n13 VPWR.t6 350.642
R154 VPWR.n52 VPWR.n1 315.832
R155 VPWR.n29 VPWR.t0 131.333
R156 VPWR.n44 VPWR.t10 90.8052
R157 VPWR.n44 VPWR.t2 72.996
R158 VPWR.n11 VPWR.t5 70.3576
R159 VPWR.n11 VPWR.t1 64.4945
R160 VPWR.n1 VPWR.t9 61.563
R161 VPWR.n1 VPWR.t8 46.1724
R162 VPWR.n29 VPWR.t7 45.4667
R163 VPWR.n50 VPWR.n2 36.1417
R164 VPWR.n51 VPWR.n50 36.1417
R165 VPWR.n31 VPWR.n6 36.1417
R166 VPWR.n35 VPWR.n6 36.1417
R167 VPWR.n36 VPWR.n35 36.1417
R168 VPWR.n38 VPWR.n36 36.1417
R169 VPWR.n23 VPWR.n22 36.1417
R170 VPWR.n23 VPWR.n8 36.1417
R171 VPWR.n27 VPWR.n8 36.1417
R172 VPWR.n20 VPWR.n12 36.1417
R173 VPWR.n28 VPWR.n27 33.5198
R174 VPWR.n46 VPWR.n2 33.0282
R175 VPWR.n43 VPWR.n42 31.33
R176 VPWR.n16 VPWR.n14 31.2476
R177 VPWR.n16 VPWR.n15 30.8711
R178 VPWR.n22 VPWR.n21 25.977
R179 VPWR.n42 VPWR.n4 25.1031
R180 VPWR.n21 VPWR.n20 21.4593
R181 VPWR.n31 VPWR.n30 18.8308
R182 VPWR.n38 VPWR.n37 11.9129
R183 VPWR.n52 VPWR.n51 10.9181
R184 VPWR.n17 VPWR.n16 9.3005
R185 VPWR.n18 VPWR.n12 9.3005
R186 VPWR.n20 VPWR.n19 9.3005
R187 VPWR.n21 VPWR.n10 9.3005
R188 VPWR.n22 VPWR.n9 9.3005
R189 VPWR.n24 VPWR.n23 9.3005
R190 VPWR.n25 VPWR.n8 9.3005
R191 VPWR.n27 VPWR.n26 9.3005
R192 VPWR.n28 VPWR.n7 9.3005
R193 VPWR.n32 VPWR.n31 9.3005
R194 VPWR.n33 VPWR.n6 9.3005
R195 VPWR.n35 VPWR.n34 9.3005
R196 VPWR.n36 VPWR.n5 9.3005
R197 VPWR.n39 VPWR.n38 9.3005
R198 VPWR.n40 VPWR.n4 9.3005
R199 VPWR.n42 VPWR.n41 9.3005
R200 VPWR.n43 VPWR.n3 9.3005
R201 VPWR.n47 VPWR.n46 9.3005
R202 VPWR.n48 VPWR.n2 9.3005
R203 VPWR.n50 VPWR.n49 9.3005
R204 VPWR.n51 VPWR.n0 9.3005
R205 VPWR.n53 VPWR.n52 8.08026
R206 VPWR.n14 VPWR.n13 6.50549
R207 VPWR.n15 VPWR.n12 5.27109
R208 VPWR.n46 VPWR.n45 4.76546
R209 VPWR.n45 VPWR.n43 4.20488
R210 VPWR.n30 VPWR.n28 2.62907
R211 VPWR.n37 VPWR.n4 1.86911
R212 VPWR.n17 VPWR.n13 0.686474
R213 VPWR VPWR.n53 0.163644
R214 VPWR.n53 VPWR.n0 0.144205
R215 VPWR.n18 VPWR.n17 0.122949
R216 VPWR.n19 VPWR.n18 0.122949
R217 VPWR.n19 VPWR.n10 0.122949
R218 VPWR.n10 VPWR.n9 0.122949
R219 VPWR.n24 VPWR.n9 0.122949
R220 VPWR.n25 VPWR.n24 0.122949
R221 VPWR.n26 VPWR.n25 0.122949
R222 VPWR.n26 VPWR.n7 0.122949
R223 VPWR.n32 VPWR.n7 0.122949
R224 VPWR.n33 VPWR.n32 0.122949
R225 VPWR.n34 VPWR.n33 0.122949
R226 VPWR.n34 VPWR.n5 0.122949
R227 VPWR.n39 VPWR.n5 0.122949
R228 VPWR.n40 VPWR.n39 0.122949
R229 VPWR.n41 VPWR.n40 0.122949
R230 VPWR.n41 VPWR.n3 0.122949
R231 VPWR.n47 VPWR.n3 0.122949
R232 VPWR.n48 VPWR.n47 0.122949
R233 VPWR.n49 VPWR.n48 0.122949
R234 VPWR.n49 VPWR.n0 0.122949
R235 VPB.t5 VPB.t17 648.657
R236 VPB.t10 VPB.t15 536.29
R237 VPB.t17 VPB.t3 515.861
R238 VPB.t1 VPB.t6 487.769
R239 VPB.t7 VPB.t8 459.678
R240 VPB.t16 VPB.t5 377.957
R241 VPB.t0 VPB.t10 316.668
R242 VPB VPB.t13 314.113
R243 VPB.t15 VPB.t2 275.807
R244 VPB.t14 VPB.t0 275.807
R245 VPB.t11 VPB.t16 275.807
R246 VPB.t9 VPB.t1 257.93
R247 VPB.t13 VPB.t12 255.376
R248 VPB.t6 VPB.t7 229.839
R249 VPB.t3 VPB.t14 229.839
R250 VPB.t4 VPB.t11 229.839
R251 VPB.t2 VPB.t9 214.517
R252 VPB.t12 VPB.t4 214.517
R253 a_1587_74.n0 a_1587_74.n4 374.875
R254 a_1587_74.n4 a_1587_74.t1 318.3
R255 a_1587_74.n2 a_1587_74.t4 254.657
R256 a_1587_74.n2 a_1587_74.n1 250.105
R257 a_1587_74.n3 a_1587_74.t3 205.922
R258 a_1587_74.n4 a_1587_74.n3 172.559
R259 a_1587_74.n0 a_1587_74.t0 111.338
R260 a_1587_74.n3 a_1587_74.n2 88.6593
R261 a_1587_74.n5 a_1587_74.n0 49.2505
R262 a_1587_74.n0 a_1587_74.t2 34.8047
R263 CLK.n0 CLK.t1 261.62
R264 CLK.n0 CLK.t0 199.519
R265 CLK CLK.n0 183.024
R266 a_630_74.t0 a_630_74.n5 877.269
R267 a_630_74.n1 a_630_74.n0 538.976
R268 a_630_74.n0 a_630_74.t5 520.561
R269 a_630_74.n2 a_630_74.n1 341.783
R270 a_630_74.n3 a_630_74.t3 260.281
R271 a_630_74.n2 a_630_74.t4 247.428
R272 a_630_74.n0 a_630_74.t7 228.683
R273 a_630_74.n5 a_630_74.t1 204.321
R274 a_630_74.n4 a_630_74.t2 204.048
R275 a_630_74.n1 a_630_74.t6 162.542
R276 a_630_74.n5 a_630_74.n4 152
R277 a_630_74.n3 a_630_74.n2 138.173
R278 a_630_74.n4 a_630_74.n3 99.906
R279 a_1764_476.t0 a_1764_476.t1 126.644
R280 a_828_74.t0 a_828_74.n4 858.783
R281 a_828_74.n1 a_828_74.t2 468.896
R282 a_828_74.n4 a_828_74.t3 328.918
R283 a_828_74.n1 a_828_74.n0 316.5
R284 a_828_74.n2 a_828_74.t4 294.894
R285 a_828_74.n2 a_828_74.n1 215.341
R286 a_828_74.n3 a_828_74.t1 209.703
R287 a_828_74.n4 a_828_74.n3 121.6
R288 a_828_74.n3 a_828_74.n2 80.8036
R289 Q.n1 Q.n0 261.985
R290 Q.n1 Q.t2 235.286
R291 Q.n3 Q.t5 177.928
R292 Q.n3 Q.n2 98.2648
R293 Q Q.n1 30.4688
R294 Q.n0 Q.t1 26.3844
R295 Q.n0 Q.t0 26.3844
R296 Q.n2 Q.t4 22.7032
R297 Q.n2 Q.t3 22.7032
R298 Q Q.n3 16.3135
R299 a_412_464.t0 a_412_464.t1 120.047
R300 D.n0 D.t1 305.267
R301 D.n0 D.t0 274.204
R302 D D.n0 166.546
R303 a_238_464.t0 a_238_464.t1 83.1099
R304 a_223_74.t0 a_223_74.t1 68.5719
R305 SCD.n0 SCD.t0 355.074
R306 SCD.n0 SCD.t1 232.7
R307 SCD.n1 SCD.n0 152
R308 SCD.n1 SCD 7.56414
R309 SCD SCD.n1 6.78838
R310 a_1257_74.n2 a_1257_74.n1 831.38
R311 a_1257_74.n1 a_1257_74.t2 386.767
R312 a_1257_74.n1 a_1257_74.n0 151.924
R313 a_1257_74.t0 a_1257_74.n2 151.268
R314 a_1257_74.n2 a_1257_74.t1 59.8041
R315 a_1026_100.n3 a_1026_100.n0 648.144
R316 a_1026_100.n2 a_1026_100.n1 325.382
R317 a_1026_100.n4 a_1026_100.n3 259.166
R318 a_1026_100.n3 a_1026_100.n2 246.871
R319 a_1026_100.n2 a_1026_100.t4 201.132
R320 a_1026_100.t0 a_1026_100.n4 111.43
R321 a_1026_100.n0 a_1026_100.t1 70.3576
R322 a_1026_100.n0 a_1026_100.t2 70.3576
R323 a_1026_100.n4 a_1026_100.t3 40.0005
R324 a_1214_506.t0 a_1214_506.t1 182.929
C0 SCD SCE 0.038536f
C1 SCD VGND 0.011242f
C2 VGND SCE 0.079598f
C3 D SCD 0.003966f
C4 SCD VPWR 0.015363f
C5 D SCE 0.114536f
C6 VPWR SCE 0.042257f
C7 SCD VPB 0.084076f
C8 SCE VPB 0.140893f
C9 SCD CLK 0.037658f
C10 D VGND 0.012892f
C11 VGND VPWR 0.197546f
C12 D VPWR 0.014571f
C13 VGND VPB 0.025414f
C14 D VPB 0.064381f
C15 VPWR VPB 0.363956f
C16 VGND Q 0.281165f
C17 CLK VGND 0.015731f
C18 Q VPWR 0.410313f
C19 CLK VPWR 0.017394f
C20 Q VPB 0.015898f
C21 CLK VPB 0.047682f
C22 Q VNB 0.075286f
C23 VGND VNB 1.45547f
C24 CLK VNB 0.14426f
C25 SCD VNB 0.132222f
C26 D VNB 0.12578f
C27 SCE VNB 0.352582f
C28 VPWR VNB 1.14893f
C29 VPB VNB 2.87035f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdlclkp_4 VNB VPB VPWR VGND SCE GATE CLK GCLK
X0 a_1289_368.t1 a_792_48.t2 a_1292_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 GCLK.t7 a_1289_368.t3 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t1 a_792_48.t3 a_785_455.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.18725 pd=1.52 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_634_74.t3 a_324_79.t2 a_119_143.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.105125 pd=0.95 as=0.38225 ps=2.49 w=0.55 l=0.15
X4 a_116_395.t1 SCE.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_354_105.t0 a_324_79.t3 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4033 pd=3.02 as=0.4872 ps=2.84 w=0.84 l=0.15
X6 a_785_455.t1 a_324_79.t4 a_634_74.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1428 ps=1.225 w=0.42 l=0.15
X7 VPWR.t2 a_792_48.t4 a_1289_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2772 ps=1.615 w=1.12 l=0.15
X8 a_119_143.t4 SCE.t1 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.089375 pd=0.875 as=0.1705 ps=1.72 w=0.55 l=0.15
X9 a_634_74.t1 a_354_105.t2 a_119_143.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X10 GCLK.t0 a_1289_368.t4 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.196 ps=1.47 w=1.12 l=0.15
X11 a_792_48.t0 a_634_74.t4 VGND.t10 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1891 ps=1.45 w=0.74 l=0.15
X12 a_792_48.t1 a_634_74.t5 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.18725 ps=1.52 w=1.12 l=0.15
X13 a_1289_368.t2 CLK.t0 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2772 pd=1.615 as=0.203 ps=1.505 w=1.12 l=0.15
X14 VGND.t1 a_792_48.t5 a_744_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1891 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X15 a_354_105.t1 a_324_79.t5 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.274375 ps=1.68 w=0.74 l=0.15
X16 VPWR.t9 CLK.t1 a_324_79.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.252 ps=2.28 w=0.84 l=0.15
X17 a_1292_74.t0 CLK.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 a_119_143.t0 GATE.t0 a_116_395.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1134 ps=1.11 w=0.84 l=0.15
X19 GCLK.t6 a_1289_368.t5 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t7 a_1289_368.t6 GCLK.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2408 ps=1.55 w=1.12 l=0.15
X21 VGND.t3 GATE.t1 a_119_143.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.274375 pd=1.68 as=0.089375 ps=0.875 w=0.55 l=0.15
X22 VGND.t2 CLK.t3 a_324_79.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X23 VGND.t7 a_1289_368.t7 GCLK.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VPWR.t6 a_1289_368.t8 GCLK.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.1932 ps=1.465 w=1.12 l=0.15
X25 GCLK.t1 a_1289_368.t9 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2408 pd=1.55 as=0.196 ps=1.47 w=1.12 l=0.15
X26 VGND.t6 a_1289_368.t10 GCLK.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X27 a_744_74.t1 a_354_105.t3 a_634_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.105125 ps=0.95 w=0.42 l=0.15
R0 a_792_48.n0 a_792_48.t5 339.61
R1 a_792_48.n3 a_792_48.n2 304.676
R2 a_792_48.n1 a_792_48.t0 270.055
R3 a_792_48.n2 a_792_48.t4 259.834
R4 a_792_48.t1 a_792_48.n3 219.778
R5 a_792_48.n1 a_792_48.n0 202.825
R6 a_792_48.n2 a_792_48.t2 199.584
R7 a_792_48.n0 a_792_48.t3 190.458
R8 a_792_48.n3 a_792_48.n1 11.641
R9 a_1292_74.t0 a_1292_74.t1 38.9194
R10 a_1289_368.n12 a_1289_368.n11 257.671
R11 a_1289_368.n9 a_1289_368.t9 251.151
R12 a_1289_368.n1 a_1289_368.t8 240.197
R13 a_1289_368.n3 a_1289_368.t4 240.197
R14 a_1289_368.n6 a_1289_368.t6 240.197
R15 a_1289_368.n11 a_1289_368.t1 182.216
R16 a_1289_368.n1 a_1289_368.t7 182.138
R17 a_1289_368.n8 a_1289_368.t3 179.947
R18 a_1289_368.n5 a_1289_368.t10 179.947
R19 a_1289_368.n2 a_1289_368.t5 179.947
R20 a_1289_368.n4 a_1289_368.n0 165.189
R21 a_1289_368.n10 a_1289_368.n9 152
R22 a_1289_368.n7 a_1289_368.n0 152
R23 a_1289_368.n12 a_1289_368.t2 60.6835
R24 a_1289_368.n2 a_1289_368.n1 60.6157
R25 a_1289_368.n4 a_1289_368.n3 47.4702
R26 a_1289_368.t0 a_1289_368.n12 26.3844
R27 a_1289_368.n9 a_1289_368.n8 25.5611
R28 a_1289_368.n7 a_1289_368.n6 24.1005
R29 a_1289_368.n8 a_1289_368.n7 24.1005
R30 a_1289_368.n6 a_1289_368.n5 21.9096
R31 a_1289_368.n10 a_1289_368.n0 13.1884
R32 a_1289_368.n3 a_1289_368.n2 11.6853
R33 a_1289_368.n11 a_1289_368.n10 5.4308
R34 a_1289_368.n5 a_1289_368.n4 3.65202
R35 VNB.n0 VNB 12403.2
R36 VNB VNB.n1 10323.1
R37 VNB.t7 VNB.t6 3250.66
R38 VNB.t3 VNB.t12 2286.61
R39 VNB.t6 VNB.t5 1625.33
R40 VNB.n1 VNB.t13 1510.99
R41 VNB.t0 VNB.t7 1277.04
R42 VNB.t8 VNB 1207.39
R43 VNB.n0 VNB.t4 1189.5
R44 VNB.t4 VNB.t1 1154.86
R45 VNB.t13 VNB.n0 1148.35
R46 VNB.t12 VNB.t9 1108.66
R47 VNB.t5 VNB.t8 1102.9
R48 VNB.t11 VNB.t10 993.177
R49 VNB.t9 VNB.t11 993.177
R50 VNB.t2 VNB.t0 905.542
R51 VNB.t1 VNB.t3 900.788
R52 VNB.n1 VNB.t2 545.646
R53 VGND.n14 VGND.t9 285.764
R54 VGND.n2 VGND.n1 280.606
R55 VGND.n41 VGND.t5 259.401
R56 VGND.n12 VGND.n11 214.185
R57 VGND.n28 VGND.n27 205.752
R58 VGND.n10 VGND.t7 178.81
R59 VGND.n27 VGND.t10 141.7
R60 VGND.n20 VGND.n19 116.288
R61 VGND.n1 VGND.t3 67.6369
R62 VGND.n27 VGND.t1 45.7148
R63 VGND.n1 VGND.t4 38.9194
R64 VGND.n18 VGND.n8 36.1417
R65 VGND.n22 VGND.n21 36.1417
R66 VGND.n22 VGND.n6 36.1417
R67 VGND.n26 VGND.n6 36.1417
R68 VGND.n30 VGND.n29 36.1417
R69 VGND.n30 VGND.n4 36.1417
R70 VGND.n34 VGND.n4 36.1417
R71 VGND.n35 VGND.n34 36.1417
R72 VGND.n36 VGND.n35 36.1417
R73 VGND.n19 VGND.t2 34.0546
R74 VGND.n40 VGND.n39 32.3059
R75 VGND.n14 VGND.n8 32.0005
R76 VGND.n13 VGND.n12 28.2358
R77 VGND.n11 VGND.t8 22.7032
R78 VGND.n11 VGND.t6 22.7032
R79 VGND.n19 VGND.t0 22.7032
R80 VGND.n14 VGND.n13 21.4593
R81 VGND.n41 VGND.n40 20.7064
R82 VGND.n36 VGND.n2 13.9725
R83 VGND.n20 VGND.n18 10.9181
R84 VGND.n28 VGND.n26 9.41227
R85 VGND.n42 VGND.n41 9.3005
R86 VGND.n13 VGND.n9 9.3005
R87 VGND.n15 VGND.n14 9.3005
R88 VGND.n16 VGND.n8 9.3005
R89 VGND.n18 VGND.n17 9.3005
R90 VGND.n21 VGND.n7 9.3005
R91 VGND.n23 VGND.n22 9.3005
R92 VGND.n24 VGND.n6 9.3005
R93 VGND.n26 VGND.n25 9.3005
R94 VGND.n29 VGND.n5 9.3005
R95 VGND.n31 VGND.n30 9.3005
R96 VGND.n32 VGND.n4 9.3005
R97 VGND.n34 VGND.n33 9.3005
R98 VGND.n35 VGND.n3 9.3005
R99 VGND.n37 VGND.n36 9.3005
R100 VGND.n39 VGND.n38 9.3005
R101 VGND.n40 VGND.n0 9.3005
R102 VGND.n12 VGND.n10 6.79022
R103 VGND.n39 VGND.n2 3.50239
R104 VGND.n29 VGND.n28 1.88285
R105 VGND.n10 VGND.n9 0.5771
R106 VGND.n21 VGND.n20 0.376971
R107 VGND.n15 VGND.n9 0.122949
R108 VGND.n16 VGND.n15 0.122949
R109 VGND.n17 VGND.n16 0.122949
R110 VGND.n17 VGND.n7 0.122949
R111 VGND.n23 VGND.n7 0.122949
R112 VGND.n24 VGND.n23 0.122949
R113 VGND.n25 VGND.n24 0.122949
R114 VGND.n25 VGND.n5 0.122949
R115 VGND.n31 VGND.n5 0.122949
R116 VGND.n32 VGND.n31 0.122949
R117 VGND.n33 VGND.n32 0.122949
R118 VGND.n33 VGND.n3 0.122949
R119 VGND.n37 VGND.n3 0.122949
R120 VGND.n38 VGND.n37 0.122949
R121 VGND.n38 VGND.n0 0.122949
R122 VGND.n42 VGND.n0 0.122949
R123 VGND VGND.n42 0.0617245
R124 GCLK.n2 GCLK.n0 254.282
R125 GCLK.n2 GCLK.n1 207.6
R126 GCLK.n5 GCLK.n3 147.95
R127 GCLK.n5 GCLK.n4 99.7716
R128 GCLK.n0 GCLK.t1 49.2505
R129 GCLK.n1 GCLK.t2 34.2996
R130 GCLK.n3 GCLK.t7 30.8113
R131 GCLK GCLK.n2 30.255
R132 GCLK.n1 GCLK.t0 26.3844
R133 GCLK.n0 GCLK.t3 26.3844
R134 GCLK.n4 GCLK.t5 22.7032
R135 GCLK.n4 GCLK.t6 22.7032
R136 GCLK.n3 GCLK.t4 22.7032
R137 GCLK GCLK.n5 6.4005
R138 a_785_455.t0 a_785_455.t1 126.644
R139 VPWR.n3 VPWR.t3 664.819
R140 VPWR.n21 VPWR.n9 651.098
R141 VPWR.n39 VPWR.t0 415.183
R142 VPWR.n26 VPWR.n6 335.337
R143 VPWR.n14 VPWR.n13 325.255
R144 VPWR.n11 VPWR.n10 317.341
R145 VPWR.n12 VPWR.t6 257.664
R146 VPWR.n6 VPWR.t1 117.263
R147 VPWR.n9 VPWR.t9 55.1136
R148 VPWR.n38 VPWR.n37 36.1417
R149 VPWR.n27 VPWR.n4 36.1417
R150 VPWR.n31 VPWR.n4 36.1417
R151 VPWR.n32 VPWR.n31 36.1417
R152 VPWR.n33 VPWR.n32 36.1417
R153 VPWR.n25 VPWR.n7 36.1417
R154 VPWR.n20 VPWR.n19 36.1417
R155 VPWR.n10 VPWR.t2 35.1791
R156 VPWR.n13 VPWR.t8 35.1791
R157 VPWR.n15 VPWR.n11 35.0123
R158 VPWR.n21 VPWR.n7 34.6358
R159 VPWR.n9 VPWR.t4 29.6087
R160 VPWR.n37 VPWR.n1 28.2358
R161 VPWR.n6 VPWR.t10 27.9716
R162 VPWR.n26 VPWR.n25 27.1064
R163 VPWR.n10 VPWR.t5 26.3844
R164 VPWR.n13 VPWR.t7 26.3844
R165 VPWR.n27 VPWR.n26 26.3534
R166 VPWR.n15 VPWR.n14 23.7181
R167 VPWR.n39 VPWR.n38 20.7064
R168 VPWR.n21 VPWR.n20 12.8005
R169 VPWR.n19 VPWR.n11 12.424
R170 VPWR.n16 VPWR.n15 9.3005
R171 VPWR.n17 VPWR.n11 9.3005
R172 VPWR.n19 VPWR.n18 9.3005
R173 VPWR.n20 VPWR.n8 9.3005
R174 VPWR.n22 VPWR.n21 9.3005
R175 VPWR.n23 VPWR.n7 9.3005
R176 VPWR.n25 VPWR.n24 9.3005
R177 VPWR.n26 VPWR.n5 9.3005
R178 VPWR.n28 VPWR.n27 9.3005
R179 VPWR.n29 VPWR.n4 9.3005
R180 VPWR.n31 VPWR.n30 9.3005
R181 VPWR.n32 VPWR.n2 9.3005
R182 VPWR.n34 VPWR.n33 9.3005
R183 VPWR.n35 VPWR.n1 9.3005
R184 VPWR.n37 VPWR.n36 9.3005
R185 VPWR.n38 VPWR.n0 9.3005
R186 VPWR.n40 VPWR.n39 9.3005
R187 VPWR.n14 VPWR.n12 6.96039
R188 VPWR.n3 VPWR.n1 5.18743
R189 VPWR.n33 VPWR.n3 2.84494
R190 VPWR.n16 VPWR.n12 0.594857
R191 VPWR.n17 VPWR.n16 0.122949
R192 VPWR.n18 VPWR.n17 0.122949
R193 VPWR.n18 VPWR.n8 0.122949
R194 VPWR.n22 VPWR.n8 0.122949
R195 VPWR.n23 VPWR.n22 0.122949
R196 VPWR.n24 VPWR.n23 0.122949
R197 VPWR.n24 VPWR.n5 0.122949
R198 VPWR.n28 VPWR.n5 0.122949
R199 VPWR.n29 VPWR.n28 0.122949
R200 VPWR.n30 VPWR.n29 0.122949
R201 VPWR.n30 VPWR.n2 0.122949
R202 VPWR.n34 VPWR.n2 0.122949
R203 VPWR.n35 VPWR.n34 0.122949
R204 VPWR.n36 VPWR.n35 0.122949
R205 VPWR.n36 VPWR.n0 0.122949
R206 VPWR.n40 VPWR.n0 0.122949
R207 VPWR VPWR.n40 0.0617245
R208 VPB.n0 VPB 2742.74
R209 VPB VPB.n1 703.611
R210 VPB.t5 VPB.t4 556.284
R211 VPB.n1 VPB.t5 424.199
R212 VPB.t7 VPB.t2 329.435
R213 VPB.t8 VPB.t10 296.238
R214 VPB.t13 VPB.n0 279.413
R215 VPB.t3 VPB.t13 279.413
R216 VPB.t12 VPB.t7 273.253
R217 VPB.t4 VPB.t6 271.791
R218 VPB.t0 VPB 257.93
R219 VPB.t10 VPB.t11 255.376
R220 VPB.t2 VPB.t8 255.376
R221 VPB.t11 VPB.t9 252.823
R222 VPB.n0 VPB.t12 237.5
R223 VPB.n1 VPB.t1 234.946
R224 VPB.t1 VPB.t0 214.517
R225 VPB.t6 VPB.t3 213.369
R226 a_324_79.t3 a_324_79.t4 849.124
R227 a_324_79.t1 a_324_79.n2 842.029
R228 a_324_79.n2 a_324_79.n1 503.714
R229 a_324_79.n1 a_324_79.t2 313.5
R230 a_324_79.n0 a_324_79.t3 307.678
R231 a_324_79.n0 a_324_79.t5 292.522
R232 a_324_79.n2 a_324_79.t0 132.249
R233 a_324_79.n1 a_324_79.n0 20.5803
R234 a_119_143.t0 a_119_143.n0 777.639
R235 a_119_143.t0 a_119_143.n3 768.644
R236 a_119_143.n0 a_119_143.t1 479.945
R237 a_119_143.n2 a_119_143.t3 353.509
R238 a_119_143.n2 a_119_143.n1 243.308
R239 a_119_143.n3 a_119_143.n2 91.2469
R240 a_119_143.n1 a_119_143.t4 40.3641
R241 a_119_143.n1 a_119_143.t2 30.546
R242 a_119_143.n3 a_119_143.n0 5.25423
R243 a_634_74.n0 a_634_74.n3 332.699
R244 a_634_74.n1 a_634_74.t5 256.337
R245 a_634_74.n3 a_634_74.n1 225.788
R246 a_634_74.n3 a_634_74.n2 218.079
R247 a_634_74.n1 a_634_74.t4 180.555
R248 a_634_74.n0 a_634_74.t2 111.418
R249 a_634_74.n2 a_634_74.t0 68.5719
R250 a_634_74.n2 a_634_74.t3 34.9096
R251 a_634_74.n0 a_634_74.t1 31.3024
R252 a_634_74.n4 a_634_74.n0 14.5065
R253 SCE.n0 SCE.t0 211.062
R254 SCE.n0 SCE.t1 170.629
R255 SCE SCE.n0 160.922
R256 a_116_395.t0 a_116_395.t1 63.3219
R257 a_354_105.t0 a_354_105.n1 901.237
R258 a_354_105.n0 a_354_105.t3 355.365
R259 a_354_105.n1 a_354_105.t1 332.382
R260 a_354_105.n1 a_354_105.n0 212.255
R261 a_354_105.n0 a_354_105.t2 181.821
R262 CLK.n0 CLK.t0 261.62
R263 CLK.n1 CLK.t1 223.935
R264 CLK CLK.n2 158.788
R265 CLK.n0 CLK.t2 156.431
R266 CLK.n1 CLK.t3 154.24
R267 CLK.n2 CLK.n0 61.346
R268 CLK.n2 CLK.n1 9.49444
R269 a_744_74.t0 a_744_74.t1 68.5719
R270 GATE.n0 GATE.t0 213.954
R271 GATE.n0 GATE.t1 173.52
R272 GATE GATE.n0 156.462
C0 GCLK VGND 0.2748f
C1 CLK GCLK 1.31e-19
C2 VPWR VGND 0.168397f
C3 SCE VGND 0.047123f
C4 GATE GCLK 1.17e-20
C5 VPB GCLK 0.013106f
C6 VPWR CLK 0.02632f
C7 VPWR GATE 0.017602f
C8 VPB VPWR 0.313936f
C9 SCE GATE 0.07811f
C10 VPB SCE 0.049638f
C11 VPWR GCLK 0.408978f
C12 VPWR SCE 0.052078f
C13 CLK VGND 0.05091f
C14 GATE VGND 0.008219f
C15 VPB VGND 0.023484f
C16 VPB CLK 0.080982f
C17 VPB GATE 0.053055f
C18 VGND VNB 1.21174f
C19 GCLK VNB 0.038649f
C20 CLK VNB 0.211976f
C21 VPWR VNB 0.955987f
C22 GATE VNB 0.103409f
C23 SCE VNB 0.139194f
C24 VPB VNB 2.24222f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sedfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sedfxbp_1 VNB VPB VPWR VGND Q_N CLK Q SCD SCE DE D
X0 a_1348_368.t0 CLK.t0 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_1549_74.t0 a_1348_368.t1 VPWR.t2 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_556_464.t1 DE.t0 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1696 ps=1.17 w=0.64 l=0.15
X3 a_2391_74.t0 a_1972_92.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1824 ps=1.85 w=0.64 l=0.15
X4 a_1068_462.t1 SCD.t0 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1488 ps=1.105 w=0.64 l=0.15
X5 VGND.t2 DE.t1 a_157_90.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6 a_697_113.t2 a_667_87.t2 a_27_90.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR.t3 a_2463_74.t4 Q.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X8 a_2463_74.t1 a_1549_74.t2 a_2391_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.10695 pd=1 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 VPWR.t0 SCE.t0 a_667_87.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1488 pd=1.105 as=0.2304 ps=2 w=0.64 l=0.15
X10 a_533_113.t0 a_161_394.t2 VGND.t9 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 a_2345_392.t0 a_1972_92.t3 VPWR.t12 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.4125 pd=1.825 as=0.4032 ps=2.92 w=1 l=0.15
X12 VGND.t6 a_575_305.t2 a_2565_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.20915 pd=1.505 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 a_1972_92.t0 a_1747_118# VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.149975 ps=1.365 w=0.84 l=0.15
X14 a_116_464.t0 D.t0 a_27_90.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1888 ps=1.87 w=0.64 l=0.15
X15 VGND.t3 SCE.t1 a_667_87.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.1197 ps=1.41 w=0.42 l=0.15
X16 a_697_113.t3 SCE.t2 a_1075_125.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X17 VPWR.t13 a_1972_92.t4 a_1931_508.t0 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.149975 pd=1.365 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 Q_N.t0 a_575_305.t3 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1961 ps=1.27 w=0.74 l=0.15
X19 a_1075_125.t0 SCD.t1 VGND.t8 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X20 VGND.t1 DE.t2 a_161_394.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X21 a_157_90.t1 D.t1 a_27_90.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21 ps=1.84 w=0.42 l=0.15
X22 a_1549_74.t1 a_1348_368.t2 VGND.t10 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X23 a_575_305.t1 a_2463_74.t5 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.19445 ps=1.56 w=1 l=0.15
X24 a_575_305.t0 a_2463_74.t6 VGND.t11 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.20915 ps=1.505 w=0.64 l=0.15
X25 VPWR.t7 DE.t3 a_161_394.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X26 a_2463_74.t3 a_1348_368.t3 a_2345_392.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.4125 ps=1.825 w=1 l=0.15
X27 VPWR.t9 a_575_305.t4 a_2647_508.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.19445 pd=1.56 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 Q_N.t1 a_575_305.t5 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X29 VPWR.t5 a_161_394.t3 a_116_464.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0768 ps=0.88 w=0.64 l=0.15
X30 a_27_90.t4 a_575_305.t6 a_533_113.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X31 a_1972_92.t1 a_1747_118# VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.192 pd=1.88 as=0.20615 ps=1.31 w=0.64 l=0.15
X32 a_2565_74.t1 a_1348_368.t4 a_2463_74.t2 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.10695 ps=1 w=0.42 l=0.15
X33 a_697_113.t0 SCE.t3 a_27_90.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.096 ps=0.94 w=0.64 l=0.15
X34 VGND.t4 a_1972_92.t5 a_1895_118.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.20615 pd=1.31 as=0.08085 ps=0.805 w=0.42 l=0.15
X35 VGND.t12 a_2463_74.t7 Q.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=1.27 as=0.2109 ps=2.05 w=0.74 l=0.15
X36 a_697_113.t1 a_667_87.t3 a_1068_462.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0768 ps=0.88 w=0.64 l=0.15
X37 a_2647_508.t1 a_1549_74.t3 a_2463_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1664 ps=1.385 w=0.42 l=0.15
X38 a_27_90.t0 a_575_305.t7 a_556_464.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
R0 CLK.n1 CLK.t0 285.719
R1 CLK.n1 CLK.n0 178.34
R2 CLK CLK.n1 156.481
R3 VPWR.n44 VPWR.t6 882.111
R4 VPWR.n10 VPWR.t2 882.111
R5 VPWR.n30 VPWR.t12 827.386
R6 VPWR.n0 VPWR.t5 722.067
R7 VPWR.n49 VPWR.n7 612.136
R8 VPWR.n56 VPWR.n3 611.369
R9 VPWR.n32 VPWR.n14 604.976
R10 VPWR.n19 VPWR.n18 585
R11 VPWR.n21 VPWR.n20 239.088
R12 VPWR.n18 VPWR.t9 131.333
R13 VPWR.n3 VPWR.t7 116.969
R14 VPWR.n14 VPWR.t1 99.5923
R15 VPWR.n7 VPWR.t0 96.9614
R16 VPWR.n18 VPWR.t4 94.6074
R17 VPWR.n14 VPWR.t13 77.1507
R18 VPWR.n3 VPWR.t11 46.1724
R19 VPWR.n7 VPWR.t8 46.1724
R20 VPWR.n58 VPWR.n57 36.1417
R21 VPWR.n51 VPWR.n50 36.1417
R22 VPWR.n51 VPWR.n4 36.1417
R23 VPWR.n55 VPWR.n4 36.1417
R24 VPWR.n48 VPWR.n8 36.1417
R25 VPWR.n43 VPWR.n42 36.1417
R26 VPWR.n36 VPWR.n12 36.1417
R27 VPWR.n37 VPWR.n36 36.1417
R28 VPWR.n38 VPWR.n37 36.1417
R29 VPWR.n25 VPWR.n24 36.1417
R30 VPWR.n25 VPWR.n16 36.1417
R31 VPWR.n29 VPWR.n16 36.1417
R32 VPWR.n58 VPWR.n0 35.7652
R33 VPWR.n56 VPWR.n55 35.7652
R34 VPWR.n20 VPWR.t10 35.1791
R35 VPWR.n24 VPWR.n23 33.7992
R36 VPWR.n38 VPWR.n10 30.4946
R37 VPWR.n50 VPWR.n49 29.7417
R38 VPWR.n32 VPWR.n31 29.3652
R39 VPWR.n31 VPWR.n30 28.2358
R40 VPWR.n44 VPWR.n43 26.7299
R41 VPWR.n20 VPWR.t3 26.3844
R42 VPWR.n49 VPWR.n48 23.7181
R43 VPWR.n44 VPWR.n8 20.7064
R44 VPWR.n30 VPWR.n29 19.2005
R45 VPWR.n32 VPWR.n12 18.0711
R46 VPWR.n57 VPWR.n56 17.6946
R47 VPWR.n42 VPWR.n10 16.9417
R48 VPWR.n21 VPWR.n19 11.2201
R49 VPWR.n23 VPWR.n22 9.3005
R50 VPWR.n24 VPWR.n17 9.3005
R51 VPWR.n26 VPWR.n25 9.3005
R52 VPWR.n27 VPWR.n16 9.3005
R53 VPWR.n29 VPWR.n28 9.3005
R54 VPWR.n30 VPWR.n15 9.3005
R55 VPWR.n31 VPWR.n13 9.3005
R56 VPWR.n33 VPWR.n32 9.3005
R57 VPWR.n34 VPWR.n12 9.3005
R58 VPWR.n36 VPWR.n35 9.3005
R59 VPWR.n37 VPWR.n11 9.3005
R60 VPWR.n39 VPWR.n38 9.3005
R61 VPWR.n40 VPWR.n10 9.3005
R62 VPWR.n42 VPWR.n41 9.3005
R63 VPWR.n43 VPWR.n9 9.3005
R64 VPWR.n45 VPWR.n44 9.3005
R65 VPWR.n46 VPWR.n8 9.3005
R66 VPWR.n48 VPWR.n47 9.3005
R67 VPWR.n49 VPWR.n6 9.3005
R68 VPWR.n50 VPWR.n5 9.3005
R69 VPWR.n52 VPWR.n51 9.3005
R70 VPWR.n53 VPWR.n4 9.3005
R71 VPWR.n55 VPWR.n54 9.3005
R72 VPWR.n56 VPWR.n2 9.3005
R73 VPWR.n57 VPWR.n1 9.3005
R74 VPWR.n59 VPWR.n58 9.3005
R75 VPWR.n60 VPWR.n0 6.78023
R76 VPWR.n23 VPWR.n19 4.26717
R77 VPWR VPWR.n60 0.268898
R78 VPWR.n22 VPWR.n21 0.208513
R79 VPWR.n60 VPWR.n59 0.161808
R80 VPWR.n22 VPWR.n17 0.122949
R81 VPWR.n26 VPWR.n17 0.122949
R82 VPWR.n27 VPWR.n26 0.122949
R83 VPWR.n28 VPWR.n27 0.122949
R84 VPWR.n28 VPWR.n15 0.122949
R85 VPWR.n15 VPWR.n13 0.122949
R86 VPWR.n33 VPWR.n13 0.122949
R87 VPWR.n34 VPWR.n33 0.122949
R88 VPWR.n35 VPWR.n34 0.122949
R89 VPWR.n35 VPWR.n11 0.122949
R90 VPWR.n39 VPWR.n11 0.122949
R91 VPWR.n40 VPWR.n39 0.122949
R92 VPWR.n41 VPWR.n40 0.122949
R93 VPWR.n41 VPWR.n9 0.122949
R94 VPWR.n45 VPWR.n9 0.122949
R95 VPWR.n46 VPWR.n45 0.122949
R96 VPWR.n47 VPWR.n46 0.122949
R97 VPWR.n47 VPWR.n6 0.122949
R98 VPWR.n6 VPWR.n5 0.122949
R99 VPWR.n52 VPWR.n5 0.122949
R100 VPWR.n53 VPWR.n52 0.122949
R101 VPWR.n54 VPWR.n53 0.122949
R102 VPWR.n54 VPWR.n2 0.122949
R103 VPWR.n2 VPWR.n1 0.122949
R104 VPWR.n59 VPWR.n1 0.122949
R105 a_1348_368.t0 a_1348_368.n6 1097.41
R106 a_1348_368.n2 a_1348_368.n1 585.458
R107 a_1348_368.n1 a_1348_368.t4 310.087
R108 a_1348_368.n4 a_1348_368.n2 306.873
R109 a_1348_368.n4 a_1348_368.n3 285.988
R110 a_1348_368.n6 a_1348_368.t2 281.168
R111 a_1348_368.n1 a_1348_368.t3 231.629
R112 a_1348_368.n5 a_1348_368.t1 204.048
R113 a_1348_368.n2 a_1348_368.n0 171.913
R114 a_1348_368.n5 a_1348_368.n4 170.308
R115 a_1348_368.n6 a_1348_368.n5 123.713
R116 VPB.t17 VPB.t19 998.521
R117 VPB.t9 VPB.t17 709.947
R118 VPB.t7 VPB.t10 577.152
R119 VPB.t2 VPB.t18 559.274
R120 VPB.t8 VPB.t1 549.059
R121 VPB.t5 VPB.t4 515.861
R122 VPB.t6 VPB.t9 515.861
R123 VPB.t18 VPB.t16 497.985
R124 VPB.t12 VPB.t5 362.635
R125 VPB.t10 VPB.t14 347.312
R126 VPB.t1 VPB.t11 314.113
R127 VPB.t19 VPB.t2 278.361
R128 VPB.t16 VPB.t0 273.253
R129 VPB VPB.t15 257.93
R130 VPB.t4 VPB.t13 255.376
R131 VPB.t3 VPB.t8 229.839
R132 VPB.t0 VPB.t12 214.517
R133 VPB.t14 VPB.t3 214.517
R134 VPB.t11 VPB.t6 199.195
R135 VPB.t15 VPB.t7 199.195
R136 a_1549_74.t0 a_1549_74.n5 856.563
R137 a_1549_74.n1 a_1549_74.t3 605.109
R138 a_1549_74.n1 a_1549_74.t2 442.055
R139 a_1549_74.n5 a_1549_74.n0 337.993
R140 a_1549_74.n3 a_1549_74.n2 297.58
R141 a_1549_74.n3 a_1549_74.n1 252.415
R142 a_1549_74.n4 a_1549_74.t1 209.703
R143 a_1549_74.n5 a_1549_74.n4 107.436
R144 a_1549_74.n4 a_1549_74.n3 91.1629
R145 DE.n1 DE.t1 363.108
R146 DE.n0 DE.t0 345.433
R147 DE.n1 DE.t2 175.127
R148 DE DE.n2 164.607
R149 DE.n2 DE.n0 130.141
R150 DE.n0 DE.t3 126.927
R151 DE.n2 DE.n1 101.221
R152 a_556_464.t0 a_556_464.t1 83.1099
R153 a_1972_92.t0 a_1972_92.n2 823.986
R154 a_1972_92.n1 a_1972_92.t4 378.103
R155 a_1972_92.n0 a_1972_92.t3 282.507
R156 a_1972_92.n2 a_1972_92.t1 242.674
R157 a_1972_92.n2 a_1972_92.n1 216.88
R158 a_1972_92.n0 a_1972_92.t2 190.528
R159 a_1972_92.n1 a_1972_92.t5 138.173
R160 a_1972_92.n2 a_1972_92.n0 107.302
R161 VGND.n42 VGND.t10 286.334
R162 VGND.n12 VGND.t5 285.053
R163 VGND.n62 VGND.t2 250.601
R164 VGND.n50 VGND.n49 216.225
R165 VGND.n2 VGND.n1 215.061
R166 VGND.n32 VGND.n31 205.284
R167 VGND.n17 VGND.n14 185
R168 VGND.n19 VGND.n18 185
R169 VGND.n18 VGND.n17 147.143
R170 VGND.n16 VGND.n15 141.496
R171 VGND.n31 VGND.t0 77.813
R172 VGND.n15 VGND.t12 63.2437
R173 VGND.n49 VGND.t3 60.0005
R174 VGND.n1 VGND.t1 60.0005
R175 VGND.n31 VGND.t4 55.1791
R176 VGND.n18 VGND.t11 47.7237
R177 VGND.n49 VGND.t8 42.8576
R178 VGND.n17 VGND.t6 40.0005
R179 VGND.n1 VGND.t9 40.0005
R180 VGND.n25 VGND.n24 36.1417
R181 VGND.n30 VGND.n29 36.1417
R182 VGND.n36 VGND.n10 36.1417
R183 VGND.n37 VGND.n36 36.1417
R184 VGND.n38 VGND.n37 36.1417
R185 VGND.n38 VGND.n8 36.1417
R186 VGND.n44 VGND.n43 36.1417
R187 VGND.n44 VGND.n6 36.1417
R188 VGND.n48 VGND.n6 36.1417
R189 VGND.n51 VGND.n4 36.1417
R190 VGND.n55 VGND.n4 36.1417
R191 VGND.n56 VGND.n55 36.1417
R192 VGND.n57 VGND.n56 36.1417
R193 VGND.n61 VGND.n60 36.1417
R194 VGND.n24 VGND.n23 35.5756
R195 VGND.n25 VGND.n12 30.8711
R196 VGND.n32 VGND.n30 30.8711
R197 VGND.n51 VGND.n50 26.3534
R198 VGND.n43 VGND.n42 24.8476
R199 VGND.n15 VGND.t7 22.7032
R200 VGND.n29 VGND.n12 22.5887
R201 VGND.n42 VGND.n8 22.5887
R202 VGND.n50 VGND.n48 21.0829
R203 VGND.n19 VGND.n16 20.1051
R204 VGND.n32 VGND.n10 16.9417
R205 VGND.n62 VGND.n61 15.0593
R206 VGND.n21 VGND.n20 9.3005
R207 VGND.n23 VGND.n22 9.3005
R208 VGND.n24 VGND.n13 9.3005
R209 VGND.n26 VGND.n25 9.3005
R210 VGND.n27 VGND.n12 9.3005
R211 VGND.n29 VGND.n28 9.3005
R212 VGND.n30 VGND.n11 9.3005
R213 VGND.n33 VGND.n32 9.3005
R214 VGND.n34 VGND.n10 9.3005
R215 VGND.n36 VGND.n35 9.3005
R216 VGND.n37 VGND.n9 9.3005
R217 VGND.n39 VGND.n38 9.3005
R218 VGND.n40 VGND.n8 9.3005
R219 VGND.n42 VGND.n41 9.3005
R220 VGND.n43 VGND.n7 9.3005
R221 VGND.n45 VGND.n44 9.3005
R222 VGND.n46 VGND.n6 9.3005
R223 VGND.n48 VGND.n47 9.3005
R224 VGND.n50 VGND.n5 9.3005
R225 VGND.n52 VGND.n51 9.3005
R226 VGND.n53 VGND.n4 9.3005
R227 VGND.n55 VGND.n54 9.3005
R228 VGND.n56 VGND.n3 9.3005
R229 VGND.n58 VGND.n57 9.3005
R230 VGND.n60 VGND.n59 9.3005
R231 VGND.n61 VGND.n0 9.3005
R232 VGND.n57 VGND.n2 7.52991
R233 VGND.n63 VGND.n62 7.52757
R234 VGND.n20 VGND.n14 6.07349
R235 VGND.n60 VGND.n2 3.76521
R236 VGND.n20 VGND.n19 3.55086
R237 VGND.n23 VGND.n14 2.89685
R238 VGND VGND.n63 0.280446
R239 VGND.n21 VGND.n16 0.189781
R240 VGND.n63 VGND.n0 0.150435
R241 VGND.n22 VGND.n21 0.122949
R242 VGND.n22 VGND.n13 0.122949
R243 VGND.n26 VGND.n13 0.122949
R244 VGND.n27 VGND.n26 0.122949
R245 VGND.n28 VGND.n27 0.122949
R246 VGND.n28 VGND.n11 0.122949
R247 VGND.n33 VGND.n11 0.122949
R248 VGND.n34 VGND.n33 0.122949
R249 VGND.n35 VGND.n34 0.122949
R250 VGND.n35 VGND.n9 0.122949
R251 VGND.n39 VGND.n9 0.122949
R252 VGND.n40 VGND.n39 0.122949
R253 VGND.n41 VGND.n40 0.122949
R254 VGND.n41 VGND.n7 0.122949
R255 VGND.n45 VGND.n7 0.122949
R256 VGND.n46 VGND.n45 0.122949
R257 VGND.n47 VGND.n46 0.122949
R258 VGND.n47 VGND.n5 0.122949
R259 VGND.n52 VGND.n5 0.122949
R260 VGND.n53 VGND.n52 0.122949
R261 VGND.n54 VGND.n53 0.122949
R262 VGND.n54 VGND.n3 0.122949
R263 VGND.n58 VGND.n3 0.122949
R264 VGND.n59 VGND.n58 0.122949
R265 VGND.n59 VGND.n0 0.122949
R266 a_2391_74.t0 a_2391_74.t1 39.3755
R267 VNB.t15 VNB.t4 5231.5
R268 VNB.t18 VNB.t15 4573.23
R269 VNB.t6 VNB.t3 3187.4
R270 VNB.t0 VNB.t5 2598.43
R271 VNB.t7 VNB.t16 2344.36
R272 VNB.t16 VNB.t17 2286.61
R273 VNB.t2 VNB.t1 2286.61
R274 VNB.t4 VNB.t0 1893.96
R275 VNB VNB.t12 1639.9
R276 VNB.t17 VNB.t8 1570.6
R277 VNB.t10 VNB.t14 1177.95
R278 VNB.t3 VNB.t9 1177.95
R279 VNB.t1 VNB.t11 1154.86
R280 VNB.t13 VNB.t6 993.177
R281 VNB.t14 VNB.t7 900.788
R282 VNB.t9 VNB.t18 900.788
R283 VNB.t11 VNB.t13 900.788
R284 VNB.t12 VNB.t2 900.788
R285 VNB.t5 VNB.t10 831.496
R286 SCD.n0 SCD.t0 345.166
R287 SCD SCD.n0 159.565
R288 SCD.n0 SCD.t1 134.96
R289 a_1068_462.t0 a_1068_462.t1 73.8755
R290 a_157_90.t0 a_157_90.t1 68.5719
R291 a_667_87.t0 a_667_87.n1 677.417
R292 a_667_87.n1 a_667_87.t3 435.092
R293 a_667_87.n0 a_667_87.t2 321.384
R294 a_667_87.n0 a_667_87.t1 239.126
R295 a_667_87.n1 a_667_87.n0 34.2658
R296 a_27_90.n0 a_27_90.t5 357.786
R297 a_27_90.n0 a_27_90.t2 351.175
R298 a_27_90.n3 a_27_90.n2 298.337
R299 a_27_90.n2 a_27_90.n1 287.024
R300 a_27_90.n2 a_27_90.n0 271.812
R301 a_27_90.n3 a_27_90.t1 46.1724
R302 a_27_90.t0 a_27_90.n3 46.1724
R303 a_27_90.n1 a_27_90.t3 40.0005
R304 a_27_90.n1 a_27_90.t4 40.0005
R305 a_697_113.t0 a_697_113.n1 701.865
R306 a_697_113.t0 a_697_113.n2 701.865
R307 a_697_113.n2 a_697_113.t2 359.248
R308 a_697_113.n0 a_697_113.t1 354.058
R309 a_697_113.n0 a_697_113.t3 344.836
R310 a_697_113.n1 a_697_113.n0 185.346
R311 a_697_113.n2 a_697_113.n1 17.9205
R312 a_2463_74.n5 a_2463_74.n4 705.177
R313 a_2463_74.n1 a_2463_74.t4 363.642
R314 a_2463_74.n3 a_2463_74.t5 298.993
R315 a_2463_74.n2 a_2463_74.n1 245.821
R316 a_2463_74.n4 a_2463_74.n0 203.356
R317 a_2463_74.n2 a_2463_74.t6 173.218
R318 a_2463_74.n4 a_2463_74.n3 165.189
R319 a_2463_74.n1 a_2463_74.t7 142.994
R320 a_2463_74.n5 a_2463_74.t0 110.227
R321 a_2463_74.n0 a_2463_74.t2 62.8576
R322 a_2463_74.t3 a_2463_74.n5 30.9107
R323 a_2463_74.n0 a_2463_74.t1 26.2505
R324 a_2463_74.n3 a_2463_74.n2 9.87279
R325 Q.n1 Q 589.052
R326 Q.n1 Q.n0 585
R327 Q.n2 Q.n1 585
R328 Q Q.t0 283.445
R329 Q.n1 Q.t1 26.3844
R330 Q Q.n2 10.8562
R331 Q Q.n0 9.39797
R332 Q Q.n0 2.59291
R333 Q.n2 Q 1.13468
R334 SCE.t1 SCE.t2 661.947
R335 SCE.t0 SCE.t3 597.48
R336 SCE.n0 SCE.t0 272.866
R337 SCE.n0 SCE.t1 221.72
R338 SCE SCE.n0 160.727
R339 a_161_394.t1 a_161_394.n1 660.913
R340 a_161_394.n1 a_161_394.t2 470.764
R341 a_161_394.n0 a_161_394.t0 291.562
R342 a_161_394.n0 a_161_394.t3 290.038
R343 a_161_394.n1 a_161_394.n0 42.0742
R344 a_533_113.t0 a_533_113.t1 68.5719
R345 a_2345_392.t0 a_2345_392.t1 162.525
R346 a_575_305.n2 a_575_305.t2 621.78
R347 a_575_305.n1 a_575_305.n0 300.257
R348 a_575_305.n3 a_575_305.t6 264.392
R349 a_575_305.n0 a_575_305.t5 258.942
R350 a_575_305.n3 a_575_305.t7 254.751
R351 a_575_305.t1 a_575_305.n5 230.054
R352 a_575_305.n0 a_575_305.t3 204.048
R353 a_575_305.n4 a_575_305.n3 193.738
R354 a_575_305.n4 a_575_305.n2 171.743
R355 a_575_305.n2 a_575_305.t4 138.441
R356 a_575_305.n1 a_575_305.t0 126.569
R357 a_575_305.n5 a_575_305.n1 77.9088
R358 a_575_305.n5 a_575_305.n4 9.87876
R359 a_2565_74.t0 a_2565_74.t1 68.5719
R360 D.n2 D.t0 286.327
R361 D.n1 D.n0 152
R362 D.n3 D.n2 152
R363 D.n1 D.t1 150.029
R364 D.n2 D.n1 44.2924
R365 D.n3 D.n0 11.4531
R366 D D.n3 0.505763
R367 D.n0 D 0.505763
R368 a_116_464.t0 a_116_464.t1 73.8755
R369 a_1075_125.t0 a_1075_125.t1 68.5719
R370 Q_N.n1 Q_N 589.268
R371 Q_N.n1 Q_N.n0 585
R372 Q_N.n2 Q_N.n1 585
R373 Q_N Q_N.t0 204.51
R374 Q_N.n1 Q_N.t1 26.3844
R375 Q_N Q_N.n2 11.4352
R376 Q_N Q_N.n0 9.89917
R377 Q_N Q_N.n0 2.73117
R378 Q_N.n2 Q_N 1.19517
R379 a_2647_508.t0 a_2647_508.t1 126.644
C0 DE SCE 4.07e-19
C1 VPWR SCE 0.031438f
C2 DE VGND 0.035278f
C3 SCE CLK 0.003801f
C4 Q Q_N 0.003643f
C5 VPWR Q_N 0.13858f
C6 VPWR SCD 0.012773f
C7 Q VGND 0.007393f
C8 SCD CLK 0.008701f
C9 VPWR VGND 0.080634f
C10 CLK VGND 0.020717f
C11 VPB a_1747_118# 0.090814f
C12 VPB D 0.073439f
C13 VPWR DE 0.021954f
C14 VPWR Q 0.133524f
C15 a_1747_118# SCE 9.98e-22
C16 VPWR CLK 0.013809f
C17 Q_N a_1747_118# 1.4e-20
C18 a_1747_118# VGND 0.014343f
C19 D VGND 0.015574f
C20 Q a_1747_118# 2.21e-20
C21 VPWR a_1747_118# 0.063786f
C22 VPB SCE 0.186924f
C23 D DE 0.036698f
C24 VPB Q_N 0.015803f
C25 SCD VPB 0.062204f
C26 VPWR D 0.012707f
C27 VPB VGND 0.029529f
C28 SCD SCE 0.115495f
C29 SCE VGND 0.071931f
C30 Q_N VGND 0.101602f
C31 SCD VGND 0.037665f
C32 VPB DE 0.155192f
C33 VPB Q 0.014561f
C34 VPWR VPB 0.453226f
C35 VPB CLK 0.039915f
C36 Q_N VNB 0.111572f
C37 Q VNB 0.008841f
C38 VGND VNB 1.92844f
C39 CLK VNB 0.136106f
C40 SCD VNB 0.119804f
C41 VPWR VNB 1.42615f
C42 SCE VNB 0.368347f
C43 DE VNB 0.293709f
C44 D VNB 0.184881f
C45 VPB VNB 3.72744f
C46 a_1747_118# VNB 0.147827f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sedfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sedfxbp_2 VNB VPB VPWR VGND Q Q_N D CLK SCD SCE DE
X0 a_575_87.t1 a_2489_74.t3 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.21035 ps=1.68 w=1.12 l=0.15
X1 a_132_464.t0 D.t0 a_32_74.t4 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1888 ps=1.87 w=0.64 l=0.15
X2 a_691_113.t0 SCE.t0 a_32_74.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.096 ps=0.94 w=0.64 l=0.15
X3 a_1920_97# a_1586_74.t2 a_1784_97.t2 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.09765 pd=0.885 as=0.1113 ps=0.95 w=0.42 l=0.15
X4 a_32_74.t1 a_575_87.t2 a_578_462.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0768 ps=0.88 w=0.64 l=0.15
X5 a_691_113.t3 a_661_87.t2 a_1088_453.t0 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 a_691_113.t4 a_661_87.t3 a_32_74.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND.t5 SCE.t1 a_661_87.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 a_2489_74.t2 a_1374_368.t2 a_2374_392.t1 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.4025 ps=1.805 w=1 l=0.15
X9 VGND.t2 a_575_87.t3 Q_N.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_1088_453.t1 SCD.t0 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1728 ps=1.18 w=0.64 l=0.15
X11 VPWR.t5 a_575_87.t4 a_2672_508.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.21035 pd=1.68 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_2417_74.t0 a_2013_71.t2 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1824 ps=1.85 w=0.64 l=0.15
X13 VPWR.t4 DE.t0 a_183_290.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X14 a_578_462.t1 DE.t1 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1696 ps=1.17 w=0.64 l=0.15
X15 a_691_113.t1 SCE.t2 a_1091_125.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X16 VGND.t4 DE.t2 a_183_290.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X17 VGND.t10 a_2489_74.t4 Q.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_1091_125.t1 SCD.t1 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_2489_74.t1 a_1586_74.t3 a_2417_74.t1 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.10695 pd=1 as=0.0672 ps=0.85 w=0.64 l=0.15
X20 a_2374_392.t0 a_2013_71.t3 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4025 pd=1.805 as=0.4032 ps=2.92 w=1 l=0.15
X21 VPWR.t6 a_575_87.t5 Q_N.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_2013_71.t0 a_1784_97.t4 VGND.t11 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.171975 ps=1.25 w=0.64 l=0.15
X23 VPWR.t8 a_2489_74.t5 Q.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_1784_97.t1 a_1374_368.t3 a_691_113.t5 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1197 ps=1.41 w=0.42 l=0.15
X25 VGND.t3 a_575_87.t6 a_2591_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.27575 pd=1.775 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 a_1586_74.t1 a_1374_368.t4 VGND.t12 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X27 Q.t1 a_2489_74.t6 VPWR.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X28 Q_N.t0 a_575_87.t7 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 a_1374_368.t1 CLK.t0 VPWR.t14 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X30 VPWR.t2 a_2013_71.t4 a_1944_508.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.149975 pd=1.365 as=0.0756 ps=0.78 w=0.42 l=0.15
X31 a_2591_74.t1 a_1374_368.t5 a_2489_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.10695 ps=1 w=0.42 l=0.15
X32 VGND.t13 DE.t3 a_141_74.t0 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X33 a_141_74.t1 D.t1 a_32_74.t5 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1659 ps=1.63 w=0.42 l=0.15
X34 a_2013_71.t1 a_1784_97.t5 VPWR.t12 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.149975 ps=1.365 w=0.84 l=0.15
X35 VPWR.t13 a_183_290.t2 a_132_464.t1 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0864 ps=0.91 w=0.64 l=0.15
X36 a_1944_508.t1 a_1374_368.t6 a_1784_97.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0756 pd=0.78 as=0.063 ps=0.72 w=0.42 l=0.15
X37 VPWR.t3 SCE.t3 a_661_87.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1728 pd=1.18 as=0.1952 ps=1.89 w=0.64 l=0.15
X38 a_575_87.t0 a_2489_74.t7 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.27575 ps=1.775 w=0.74 l=0.15
X39 a_1586_74.t0 a_1374_368.t7 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X40 a_1784_97.t3 a_1586_74.t4 a_691_113.t2 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X41 a_32_74.t0 a_575_87.t8 a_527_113.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X42 a_1374_368.t0 CLK.t1 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X43 a_527_113.t1 a_183_290.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
R0 a_2489_74.n8 a_2489_74.n7 687.245
R1 a_2489_74.n2 a_2489_74.t5 240.197
R2 a_2489_74.n4 a_2489_74.t6 240.197
R3 a_2489_74.n6 a_2489_74.t3 240.197
R4 a_2489_74.n7 a_2489_74.n0 200.344
R5 a_2489_74.n7 a_2489_74.n6 185.749
R6 a_2489_74.n2 a_2489_74.t4 179.947
R7 a_2489_74.n5 a_2489_74.t7 179.947
R8 a_2489_74.n3 a_2489_74.n1 179.947
R9 a_2489_74.n5 a_2489_74.n4 141.679
R10 a_2489_74.n8 a_2489_74.t2 129.81
R11 a_2489_74.n0 a_2489_74.t0 62.8576
R12 a_2489_74.n3 a_2489_74.n2 62.8066
R13 a_2489_74.n0 a_2489_74.t1 26.2505
R14 a_2489_74.n6 a_2489_74.n5 5.84292
R15 a_2489_74.n4 a_2489_74.n3 2.92171
R16 VPWR.n53 VPWR.t14 888.505
R17 VPWR.n10 VPWR.t0 882.111
R18 VPWR.n19 VPWR.t9 860.096
R19 VPWR.n21 VPWR.t8 855.867
R20 VPWR.n15 VPWR.t1 827.386
R21 VPWR.n0 VPWR.t13 722.067
R22 VPWR.n66 VPWR.n3 612.136
R23 VPWR.n59 VPWR.n7 612.023
R24 VPWR.n41 VPWR.n14 604.976
R25 VPWR.n29 VPWR.n28 585
R26 VPWR.n20 VPWR.t6 351.858
R27 VPWR.n28 VPWR.t5 119.608
R28 VPWR.n28 VPWR.t7 119.108
R29 VPWR.n3 VPWR.t4 116.969
R30 VPWR.n7 VPWR.t3 116.969
R31 VPWR.n14 VPWR.t12 99.5923
R32 VPWR.n14 VPWR.t2 77.1507
R33 VPWR.n7 VPWR.t11 49.2505
R34 VPWR.n3 VPWR.t10 46.1724
R35 VPWR.n68 VPWR.n67 36.1417
R36 VPWR.n61 VPWR.n60 36.1417
R37 VPWR.n61 VPWR.n4 36.1417
R38 VPWR.n65 VPWR.n4 36.1417
R39 VPWR.n54 VPWR.n8 36.1417
R40 VPWR.n58 VPWR.n8 36.1417
R41 VPWR.n52 VPWR.n51 36.1417
R42 VPWR.n45 VPWR.n12 36.1417
R43 VPWR.n46 VPWR.n45 36.1417
R44 VPWR.n47 VPWR.n46 36.1417
R45 VPWR.n40 VPWR.n39 36.1417
R46 VPWR.n30 VPWR.n17 36.1417
R47 VPWR.n34 VPWR.n17 36.1417
R48 VPWR.n35 VPWR.n34 36.1417
R49 VPWR.n36 VPWR.n35 36.1417
R50 VPWR.n60 VPWR.n59 35.7652
R51 VPWR.n26 VPWR.n19 29.7417
R52 VPWR.n41 VPWR.n12 28.9887
R53 VPWR.n27 VPWR.n26 27.6502
R54 VPWR.n68 VPWR.n0 27.4829
R55 VPWR.n66 VPWR.n65 27.4829
R56 VPWR.n51 VPWR.n10 26.7299
R57 VPWR.n67 VPWR.n66 25.977
R58 VPWR.n22 VPWR.n21 25.224
R59 VPWR.n47 VPWR.n10 20.7064
R60 VPWR.n41 VPWR.n40 18.4476
R61 VPWR.n22 VPWR.n19 17.6946
R62 VPWR.n53 VPWR.n52 16.9417
R63 VPWR.n59 VPWR.n58 16.1887
R64 VPWR.n30 VPWR.n29 10.9181
R65 VPWR.n23 VPWR.n22 9.3005
R66 VPWR.n24 VPWR.n19 9.3005
R67 VPWR.n26 VPWR.n25 9.3005
R68 VPWR.n27 VPWR.n18 9.3005
R69 VPWR.n31 VPWR.n30 9.3005
R70 VPWR.n32 VPWR.n17 9.3005
R71 VPWR.n34 VPWR.n33 9.3005
R72 VPWR.n35 VPWR.n16 9.3005
R73 VPWR.n37 VPWR.n36 9.3005
R74 VPWR.n39 VPWR.n38 9.3005
R75 VPWR.n40 VPWR.n13 9.3005
R76 VPWR.n42 VPWR.n41 9.3005
R77 VPWR.n43 VPWR.n12 9.3005
R78 VPWR.n45 VPWR.n44 9.3005
R79 VPWR.n46 VPWR.n11 9.3005
R80 VPWR.n48 VPWR.n47 9.3005
R81 VPWR.n49 VPWR.n10 9.3005
R82 VPWR.n51 VPWR.n50 9.3005
R83 VPWR.n52 VPWR.n9 9.3005
R84 VPWR.n55 VPWR.n54 9.3005
R85 VPWR.n56 VPWR.n8 9.3005
R86 VPWR.n58 VPWR.n57 9.3005
R87 VPWR.n59 VPWR.n6 9.3005
R88 VPWR.n60 VPWR.n5 9.3005
R89 VPWR.n62 VPWR.n61 9.3005
R90 VPWR.n63 VPWR.n4 9.3005
R91 VPWR.n65 VPWR.n64 9.3005
R92 VPWR.n66 VPWR.n2 9.3005
R93 VPWR.n67 VPWR.n1 9.3005
R94 VPWR.n69 VPWR.n68 9.3005
R95 VPWR.n36 VPWR.n15 8.28285
R96 VPWR.n70 VPWR.n0 7.26437
R97 VPWR.n21 VPWR.n20 6.50549
R98 VPWR.n39 VPWR.n15 3.01226
R99 VPWR.n29 VPWR.n27 2.092
R100 VPWR.n23 VPWR.n20 0.686474
R101 VPWR.n54 VPWR.n53 0.376971
R102 VPWR VPWR.n70 0.276379
R103 VPWR.n70 VPWR.n69 0.15444
R104 VPWR.n24 VPWR.n23 0.122949
R105 VPWR.n25 VPWR.n24 0.122949
R106 VPWR.n25 VPWR.n18 0.122949
R107 VPWR.n31 VPWR.n18 0.122949
R108 VPWR.n32 VPWR.n31 0.122949
R109 VPWR.n33 VPWR.n32 0.122949
R110 VPWR.n33 VPWR.n16 0.122949
R111 VPWR.n37 VPWR.n16 0.122949
R112 VPWR.n38 VPWR.n37 0.122949
R113 VPWR.n38 VPWR.n13 0.122949
R114 VPWR.n42 VPWR.n13 0.122949
R115 VPWR.n43 VPWR.n42 0.122949
R116 VPWR.n44 VPWR.n43 0.122949
R117 VPWR.n44 VPWR.n11 0.122949
R118 VPWR.n48 VPWR.n11 0.122949
R119 VPWR.n49 VPWR.n48 0.122949
R120 VPWR.n50 VPWR.n49 0.122949
R121 VPWR.n50 VPWR.n9 0.122949
R122 VPWR.n55 VPWR.n9 0.122949
R123 VPWR.n56 VPWR.n55 0.122949
R124 VPWR.n57 VPWR.n56 0.122949
R125 VPWR.n57 VPWR.n6 0.122949
R126 VPWR.n6 VPWR.n5 0.122949
R127 VPWR.n62 VPWR.n5 0.122949
R128 VPWR.n63 VPWR.n62 0.122949
R129 VPWR.n64 VPWR.n63 0.122949
R130 VPWR.n64 VPWR.n2 0.122949
R131 VPWR.n2 VPWR.n1 0.122949
R132 VPWR.n69 VPWR.n1 0.122949
R133 a_575_87.n0 a_575_87.t6 631.42
R134 a_575_87.n4 a_575_87.n3 287.058
R135 a_575_87.n6 a_575_87.n5 278.038
R136 a_575_87.n1 a_575_87.t8 256.723
R137 a_575_87.n1 a_575_87.t2 250.297
R138 a_575_87.n2 a_575_87.t5 246.04
R139 a_575_87.t1 a_575_87.n7 222.59
R140 a_575_87.n6 a_575_87.n1 193.02
R141 a_575_87.n6 a_575_87.t0 192.365
R142 a_575_87.n7 a_575_87.n0 183.708
R143 a_575_87.n4 a_575_87.t7 182.138
R144 a_575_87.n2 a_575_87.t3 179.947
R145 a_575_87.n0 a_575_87.t4 138.441
R146 a_575_87.n5 a_575_87.n2 49.6611
R147 a_575_87.n5 a_575_87.n4 10.955
R148 a_575_87.n7 a_575_87.n6 5.66079
R149 VPB.t21 VPB.t1 709.947
R150 VPB.t19 VPB.t8 577.152
R151 VPB.t18 VPB.t5 559.274
R152 VPB.t9 VPB.t7 520.968
R153 VPB.t12 VPB.t10 515.861
R154 VPB.t1 VPB.t14 515.861
R155 VPB.t17 VPB.t21 515.861
R156 VPB.t20 VPB.t3 487.769
R157 VPB.t5 VPB.t20 487.769
R158 VPB.t11 VPB.t2 459.678
R159 VPB.t3 VPB.t12 362.635
R160 VPB.t7 VPB.t16 352.42
R161 VPB.t8 VPB.t13 347.312
R162 VPB VPB.t15 298.791
R163 VPB.t6 VPB.t18 278.361
R164 VPB.t0 VPB.t6 260.485
R165 VPB.t10 VPB.t11 229.839
R166 VPB.t14 VPB.t0 229.839
R167 VPB.t4 VPB.t9 229.839
R168 VPB.t16 VPB.t17 214.517
R169 VPB.t15 VPB.t19 214.517
R170 VPB.t13 VPB.t4 199.195
R171 D.n0 D.t0 219.31
R172 D D.n0 159.649
R173 D.n1 D 154.03
R174 D.n1 D.t1 152.633
R175 D.n3 D.n2 152
R176 D.n2 D.n0 49.6611
R177 D.n2 D.n1 49.6611
R178 D.n3 D 8.58587
R179 D D.n3 2.96635
R180 a_32_74.n0 a_32_74.t4 356.079
R181 a_32_74.n0 a_32_74.t5 355.048
R182 a_32_74.n3 a_32_74.n2 300.103
R183 a_32_74.n2 a_32_74.n1 288.639
R184 a_32_74.n2 a_32_74.n0 273.318
R185 a_32_74.n3 a_32_74.t2 46.1724
R186 a_32_74.t1 a_32_74.n3 46.1724
R187 a_32_74.n1 a_32_74.t3 40.0005
R188 a_32_74.n1 a_32_74.t0 40.0005
R189 a_132_464.t0 a_132_464.t1 83.1099
R190 SCE.t1 SCE.t2 671.587
R191 SCE.t3 SCE.t0 584.827
R192 SCE.n0 SCE.t3 333.116
R193 SCE SCE.n0 162.667
R194 SCE.n0 SCE.t1 134.96
R195 a_691_113.n0 a_691_113.t2 726.194
R196 a_691_113.t0 a_691_113.n3 701.865
R197 a_691_113.t0 a_691_113.n4 701.865
R198 a_691_113.n4 a_691_113.t4 357.849
R199 a_691_113.n0 a_691_113.t5 351.675
R200 a_691_113.n2 a_691_113.t3 349.257
R201 a_691_113.n1 a_691_113.t1 339.459
R202 a_691_113.n3 a_691_113.n2 190.319
R203 a_691_113.n1 a_691_113.n0 116.329
R204 a_691_113.n4 a_691_113.n3 17.9205
R205 a_691_113.n2 a_691_113.n1 5.63632
R206 a_1586_74.t0 a_1586_74.n4 851.364
R207 a_1586_74.n1 a_1586_74.n0 579.51
R208 a_1586_74.n1 a_1586_74.t3 443.284
R209 a_1586_74.n4 a_1586_74.t4 352.88
R210 a_1586_74.n2 a_1586_74.t2 289.74
R211 a_1586_74.n2 a_1586_74.n1 249.839
R212 a_1586_74.n3 a_1586_74.t1 206.231
R213 a_1586_74.n4 a_1586_74.n3 111.242
R214 a_1586_74.n3 a_1586_74.n2 86.9522
R215 a_1784_97.n2 a_1784_97.n0 643.447
R216 a_1784_97.n1 a_1784_97.t4 282.07
R217 a_1784_97.n2 a_1784_97.n1 256.283
R218 a_1784_97.n3 a_1784_97.n2 255.024
R219 a_1784_97.n1 a_1784_97.t5 203.611
R220 a_1784_97.t1 a_1784_97.n3 111.43
R221 a_1784_97.n0 a_1784_97.t0 70.3576
R222 a_1784_97.n0 a_1784_97.t3 70.3576
R223 a_1784_97.n3 a_1784_97.t2 40.0005
R224 VNB.t14 VNB.t8 3372.18
R225 VNB.t12 VNB.t13 3279.79
R226 VNB.t21 VNB.t16 3175.85
R227 VNB.t4 VNB.t12 2737.01
R228 VNB.t16 VNB.t11 2563.78
R229 VNB.t7 VNB.t9 2529.13
R230 VNB.t19 VNB.t6 2402.1
R231 VNB.t18 VNB.t17 2286.61
R232 VNB.t9 VNB.t18 2286.61
R233 VNB.t17 VNB.t21 1570.6
R234 VNB VNB.t15 1455.12
R235 VNB.t8 VNB.t10 1247.24
R236 VNB.t20 VNB.t0 1177.95
R237 VNB.t6 VNB.t1 1154.86
R238 VNB.t3 VNB.t5 993.177
R239 VNB.t13 VNB.t3 993.177
R240 VNB.t2 VNB.t14 993.177
R241 VNB.t0 VNB.t4 900.788
R242 VNB.t10 VNB.t7 900.788
R243 VNB.t1 VNB.t2 900.788
R244 VNB.t15 VNB.t19 900.788
R245 VNB.t11 VNB.t20 831.496
R246 a_578_462.t0 a_578_462.t1 73.8755
R247 a_661_87.t0 a_661_87.n7 665.045
R248 a_661_87.n0 a_661_87.t2 373.628
R249 a_661_87.n2 a_661_87.t3 295.627
R250 a_661_87.n3 a_661_87.t1 237.049
R251 a_661_87.n7 a_661_87.n6 201.661
R252 a_661_87.n6 a_661_87.n5 152
R253 a_661_87.n4 a_661_87.n1 152
R254 a_661_87.n3 a_661_87.n2 127.081
R255 a_661_87.n6 a_661_87.n1 49.6611
R256 a_661_87.n4 a_661_87.n3 18.7722
R257 a_661_87.n5 a_661_87.n4 17.4085
R258 a_661_87.n5 a_661_87.n0 11.0085
R259 a_661_87.n2 a_661_87.n1 10.955
R260 a_661_87.n7 a_661_87.n0 6.4005
R261 a_1088_453.t0 a_1088_453.t1 83.1099
R262 VGND.n48 VGND.t11 292.856
R263 VGND.n43 VGND.t8 285.053
R264 VGND.n78 VGND.t13 247.498
R265 VGND.n21 VGND.t2 243.585
R266 VGND.n66 VGND.n65 216.225
R267 VGND.n2 VGND.n1 215.061
R268 VGND.n32 VGND.n31 201.831
R269 VGND.n36 VGND.n35 185
R270 VGND.n34 VGND.n16 185
R271 VGND.n29 VGND.n17 185
R272 VGND.n8 VGND.t12 180.233
R273 VGND.n60 VGND.t6 148.939
R274 VGND.n22 VGND.n20 132.637
R275 VGND.n35 VGND.n34 102.858
R276 VGND.n34 VGND.n33 100.001
R277 VGND.n65 VGND.t5 60.0005
R278 VGND.n1 VGND.t4 60.0005
R279 VGND.n32 VGND.t9 52.5005
R280 VGND.n65 VGND.t7 51.4291
R281 VGND.n22 VGND.n21 40.4356
R282 VGND.t9 VGND.n17 40.0005
R283 VGND.n35 VGND.t3 40.0005
R284 VGND.n1 VGND.t0 40.0005
R285 VGND.n24 VGND.n23 36.1417
R286 VGND.n41 VGND.n14 36.1417
R287 VGND.n42 VGND.n41 36.1417
R288 VGND.n47 VGND.n12 36.1417
R289 VGND.n49 VGND.n10 36.1417
R290 VGND.n53 VGND.n10 36.1417
R291 VGND.n54 VGND.n53 36.1417
R292 VGND.n55 VGND.n54 36.1417
R293 VGND.n59 VGND.n58 36.1417
R294 VGND.n64 VGND.n6 36.1417
R295 VGND.n67 VGND.n4 36.1417
R296 VGND.n71 VGND.n4 36.1417
R297 VGND.n72 VGND.n71 36.1417
R298 VGND.n73 VGND.n72 36.1417
R299 VGND.n77 VGND.n76 36.1417
R300 VGND.n43 VGND.n12 32.377
R301 VGND.n49 VGND.n48 32.377
R302 VGND.n28 VGND.n18 32.0005
R303 VGND.n60 VGND.n6 31.2476
R304 VGND.n67 VGND.n66 30.1181
R305 VGND.n29 VGND.n28 24.7404
R306 VGND.n20 VGND.t1 22.7032
R307 VGND.n20 VGND.t10 22.7032
R308 VGND.n24 VGND.n18 21.4593
R309 VGND.n43 VGND.n42 21.0829
R310 VGND.n48 VGND.n47 21.0829
R311 VGND.n55 VGND.n8 21.0829
R312 VGND.n78 VGND.n77 21.0829
R313 VGND.n66 VGND.n64 17.3181
R314 VGND.n33 VGND.n32 16.8755
R315 VGND.n60 VGND.n59 16.1887
R316 VGND.n58 VGND.n8 15.0593
R317 VGND.n33 VGND.n17 12.8576
R318 VGND.n36 VGND.n14 12.119
R319 VGND.n73 VGND.n2 9.78874
R320 VGND.n77 VGND.n0 9.3005
R321 VGND.n76 VGND.n75 9.3005
R322 VGND.n74 VGND.n73 9.3005
R323 VGND.n72 VGND.n3 9.3005
R324 VGND.n71 VGND.n70 9.3005
R325 VGND.n69 VGND.n4 9.3005
R326 VGND.n68 VGND.n67 9.3005
R327 VGND.n66 VGND.n5 9.3005
R328 VGND.n64 VGND.n63 9.3005
R329 VGND.n62 VGND.n6 9.3005
R330 VGND.n61 VGND.n60 9.3005
R331 VGND.n59 VGND.n7 9.3005
R332 VGND.n58 VGND.n57 9.3005
R333 VGND.n56 VGND.n55 9.3005
R334 VGND.n54 VGND.n9 9.3005
R335 VGND.n53 VGND.n52 9.3005
R336 VGND.n51 VGND.n10 9.3005
R337 VGND.n50 VGND.n49 9.3005
R338 VGND.n48 VGND.n11 9.3005
R339 VGND.n47 VGND.n46 9.3005
R340 VGND.n45 VGND.n12 9.3005
R341 VGND.n44 VGND.n43 9.3005
R342 VGND.n42 VGND.n13 9.3005
R343 VGND.n41 VGND.n40 9.3005
R344 VGND.n39 VGND.n14 9.3005
R345 VGND.n38 VGND.n37 9.3005
R346 VGND.n30 VGND.n15 9.3005
R347 VGND.n23 VGND.n19 9.3005
R348 VGND.n25 VGND.n24 9.3005
R349 VGND.n26 VGND.n18 9.3005
R350 VGND.n28 VGND.n27 9.3005
R351 VGND.n79 VGND.n78 7.282
R352 VGND.n30 VGND.n16 5.88663
R353 VGND.n37 VGND.n36 3.6443
R354 VGND.n37 VGND.n16 3.08371
R355 VGND.n21 VGND.n19 2.26417
R356 VGND.n76 VGND.n2 1.50638
R357 VGND.n23 VGND.n22 0.753441
R358 VGND.n31 VGND.n29 0.747945
R359 VGND.n31 VGND.n30 0.747945
R360 VGND VGND.n79 0.276651
R361 VGND.n79 VGND.n0 0.154172
R362 VGND.n25 VGND.n19 0.122949
R363 VGND.n26 VGND.n25 0.122949
R364 VGND.n27 VGND.n26 0.122949
R365 VGND.n27 VGND.n15 0.122949
R366 VGND.n38 VGND.n15 0.122949
R367 VGND.n39 VGND.n38 0.122949
R368 VGND.n40 VGND.n39 0.122949
R369 VGND.n40 VGND.n13 0.122949
R370 VGND.n44 VGND.n13 0.122949
R371 VGND.n45 VGND.n44 0.122949
R372 VGND.n46 VGND.n45 0.122949
R373 VGND.n46 VGND.n11 0.122949
R374 VGND.n50 VGND.n11 0.122949
R375 VGND.n51 VGND.n50 0.122949
R376 VGND.n52 VGND.n51 0.122949
R377 VGND.n52 VGND.n9 0.122949
R378 VGND.n56 VGND.n9 0.122949
R379 VGND.n57 VGND.n56 0.122949
R380 VGND.n57 VGND.n7 0.122949
R381 VGND.n61 VGND.n7 0.122949
R382 VGND.n62 VGND.n61 0.122949
R383 VGND.n63 VGND.n62 0.122949
R384 VGND.n63 VGND.n5 0.122949
R385 VGND.n68 VGND.n5 0.122949
R386 VGND.n69 VGND.n68 0.122949
R387 VGND.n70 VGND.n69 0.122949
R388 VGND.n70 VGND.n3 0.122949
R389 VGND.n74 VGND.n3 0.122949
R390 VGND.n75 VGND.n74 0.122949
R391 VGND.n75 VGND.n0 0.122949
R392 a_1374_368.t1 a_1374_368.n5 852.196
R393 a_1374_368.n1 a_1374_368.n0 574.173
R394 a_1374_368.n2 a_1374_368.n1 361.5
R395 a_1374_368.n0 a_1374_368.t5 310.087
R396 a_1374_368.n2 a_1374_368.t3 285.988
R397 a_1374_368.n4 a_1374_368.t4 234.573
R398 a_1374_368.n0 a_1374_368.t2 231.629
R399 a_1374_368.n3 a_1374_368.n2 207.261
R400 a_1374_368.n3 a_1374_368.t7 204.048
R401 a_1374_368.n5 a_1374_368.t0 183.982
R402 a_1374_368.n1 a_1374_368.t6 143.798
R403 a_1374_368.n5 a_1374_368.n4 125.805
R404 a_1374_368.n4 a_1374_368.n3 90.762
R405 a_2374_392.t0 a_2374_392.t1 158.585
R406 Q_N.n0 Q_N.t2 857.518
R407 Q_N.n2 Q_N.n1 185
R408 Q_N.n3 Q_N.n2 185
R409 Q_N.n1 Q_N 33.4676
R410 Q_N.n2 Q_N.t1 22.7032
R411 Q_N.n2 Q_N.t0 22.7032
R412 Q_N.n0 Q_N 18.644
R413 Q_N.n3 Q_N 12.6066
R414 Q_N.n1 Q_N 4.84898
R415 Q_N Q_N.n0 1.94833
R416 Q_N Q_N.n3 1.74595
R417 SCD.n0 SCD.t0 333.116
R418 SCD SCD.n0 157.625
R419 SCD.n0 SCD.t1 134.96
R420 a_2013_71.t1 a_2013_71.n4 836.785
R421 a_2013_71.n2 a_2013_71.t4 368.731
R422 a_2013_71.n0 a_2013_71.t3 282.507
R423 a_2013_71.n3 a_2013_71.t0 240.238
R424 a_2013_71.n3 a_2013_71.n2 212.613
R425 a_2013_71.n0 a_2013_71.t2 185.708
R426 a_2013_71.n2 a_2013_71.n1 183.161
R427 a_2013_71.n4 a_2013_71.n0 100.709
R428 a_2013_71.n4 a_2013_71.n3 10.8269
R429 a_2417_74.t0 a_2417_74.t1 39.3755
R430 DE.n1 DE.t3 356.68
R431 DE.n0 DE.t1 345.433
R432 DE.n1 DE.t2 223.327
R433 DE.n2 DE.n0 220.113
R434 DE DE.n2 157.625
R435 DE.n0 DE.t0 126.927
R436 DE.n2 DE.n1 101.221
R437 a_183_290.t1 a_183_290.n1 660.538
R438 a_183_290.n1 a_183_290.t3 457.399
R439 a_183_290.n0 a_183_290.t0 290.632
R440 a_183_290.n0 a_183_290.t2 260.846
R441 a_183_290.n1 a_183_290.n0 52.0257
R442 a_1091_125.t0 a_1091_125.t1 68.5719
R443 Q Q.n0 586.318
R444 Q.n2 Q.t0 281.43
R445 Q.t0 Q.n1 281.43
R446 Q.n0 Q.t2 26.3844
R447 Q.n0 Q.t1 26.3844
R448 Q.n1 Q 12.2358
R449 Q Q.n2 9.22403
R450 Q.n2 Q 4.70638
R451 Q.n1 Q 1.69462
R452 a_2591_74.t0 a_2591_74.t1 68.5719
R453 CLK.n0 CLK.t0 285.719
R454 CLK.n0 CLK.t1 178.34
R455 CLK CLK.n0 158.589
R456 a_1944_508.t0 a_1944_508.t1 168.857
R457 a_141_74.t0 a_141_74.t1 68.5719
R458 a_527_113.t0 a_527_113.t1 68.5719
C0 VPB Q 0.002363f
C1 Q_N VPWR 0.172756f
C2 Q_N VGND 0.174054f
C3 VPB SCE 0.181116f
C4 SCD VPWR 0.012929f
C5 SCE DE 5.45e-19
C6 Q Q_N 0.005181f
C7 VPB CLK 0.038251f
C8 VGND VPWR 0.081381f
C9 VGND SCD 0.035734f
C10 Q VPWR 0.014738f
C11 Q VGND 0.167833f
C12 VPB D 0.07453f
C13 SCE VPWR 0.03159f
C14 SCE SCD 0.119016f
C15 D DE 0.044518f
C16 CLK VPWR 0.01427f
C17 VGND SCE 0.073709f
C18 CLK SCD 0.003268f
C19 VGND a_1920_97# 0.005048f
C20 CLK VGND 0.022857f
C21 VPB DE 0.174038f
C22 D VPWR 0.012868f
C23 CLK SCE 0.003752f
C24 D VGND 0.021194f
C25 VPB Q_N 0.009481f
C26 VPB VPWR 0.498678f
C27 VPB SCD 0.058535f
C28 VPWR DE 0.023964f
C29 VPB VGND 0.014147f
C30 VGND DE 0.03635f
C31 Q_N VNB 0.063207f
C32 Q VNB 0.007595f
C33 VGND VNB 2.05886f
C34 CLK VNB 0.127916f
C35 SCD VNB 0.112144f
C36 SCE VNB 0.371815f
C37 DE VNB 0.311198f
C38 VPWR VNB 1.52506f
C39 D VNB 0.189882f
C40 VPB VNB 3.94171f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sedfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sedfxtp_1 VNB VPB VPWR VGND CLK Q SCD SCE DE D
X0 a_114_464.t1 D.t0 a_27_74.t4 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X1 a_1890_508.t0 a_1295_74.t1 a_1688_97.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2 VGND.t10 DE.t0 a_143_74.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 a_1492_74# a_1295_74.t2 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 a_547_301.t0 a_2385_74.t3 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.20475 ps=1.395 w=0.42 l=0.15
X5 VGND.t5 a_2385_74.t4 Q.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VPWR.t9 DE.t1 a_159_404.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X7 a_1824_97.t0 a_1492_74# a_1688_97.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0903 pd=0.85 as=0.1113 ps=0.95 w=0.42 l=0.15
X8 a_27_74.t2 a_547_301.t2 a_554_463.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0768 ps=0.88 w=0.64 l=0.15
X9 VGND.t9 DE.t2 a_159_404.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X10 a_27_74.t1 a_547_301.t3 a_505_111.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X11 a_1910_71.t1 a_1688_97.t4 VPWR.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.231 pd=2.23 as=0.144725 ps=1.34 w=0.84 l=0.15
X12 VPWR.t11 a_1910_71.t2 a_1890_508.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.144725 pd=1.34 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 a_554_463.t1 DE.t3 VPWR.t8 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1696 ps=1.17 w=0.64 l=0.15
X14 a_1295_74.t0 CLK.t0 VPWR.t4 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X15 a_1688_97.t2 a_1492_74# a_669_111.t4 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1176 ps=1.4 w=0.42 l=0.15
X16 VGND.t11 a_1910_71.t3 a_1824_97.t1 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.17065 pd=1.245 as=0.0903 ps=0.85 w=0.42 l=0.15
X17 a_2487_74.t0 a_1295_74.t3 a_2385_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.10695 ps=1 w=0.42 l=0.15
X18 VPWR.t7 SCE.t0 a_639_85.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1792 ps=1.84 w=0.64 l=0.15
X19 a_505_111.t1 a_159_404.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 VPWR.t10 a_159_404.t3 a_114_464.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0768 ps=0.88 w=0.64 l=0.15
X21 a_143_74.t0 D.t1 a_27_74.t5 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1806 ps=1.7 w=0.42 l=0.15
X22 a_1688_97.t0 a_1295_74.t4 a_669_111.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1176 ps=1.4 w=0.42 l=0.15
X23 a_669_111.t2 a_639_85.t2 a_27_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 a_669_111.t1 SCE.t1 a_1026_125.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 a_2313_74.t1 a_1910_71.t4 VGND.t6 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1824 ps=1.85 w=0.64 l=0.15
X26 VGND.t2 SCE.t2 a_639_85.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X27 a_2274_392.t1 a_1910_71.t5 VPWR.t5 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3925 pd=1.785 as=0.275 ps=2.55 w=1 l=0.15
X28 a_1026_125.t1 SCD.t0 VGND.t7 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 a_2385_74.t2 a_1492_74# a_2313_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.10695 pd=1 as=0.0672 ps=0.85 w=0.64 l=0.15
X30 a_1053_455.t0 SCD.t1 VPWR.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1696 ps=1.17 w=0.64 l=0.15
X31 a_2385_74.t1 a_1295_74.t5 a_2274_392.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.3925 ps=1.785 w=1 l=0.15
X32 VPWR.t0 a_547_301.t4 a_2568_508.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.14675 pd=1.2 as=0.0567 ps=0.69 w=0.42 l=0.15
X33 a_1910_71.t0 a_1688_97.t5 VGND.t8 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.17065 ps=1.245 w=0.64 l=0.15
X34 VGND.t3 a_547_301.t5 a_2487_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.20475 pd=1.395 as=0.0504 ps=0.66 w=0.42 l=0.15
X35 a_669_111.t3 SCE.t3 a_27_74.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.83 as=0.096 ps=0.94 w=0.64 l=0.15
X36 a_547_301.t1 a_2385_74.t5 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.83 as=0.14675 ps=1.2 w=0.64 l=0.15
X37 VPWR.t2 a_2385_74.t6 Q.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.308 ps=2.79 w=1.12 l=0.15
R0 D.n0 D.t0 274.836
R1 D.n1 D.t1 193.698
R2 D D.n0 153.179
R3 D.n2 D.n1 152
R4 D.n1 D.n0 48.2005
R5 D D.n2 10.2742
R6 D.n2 D 2.18997
R7 a_27_74.n0 a_27_74.t5 367.954
R8 a_27_74.n0 a_27_74.t4 359.447
R9 a_27_74.n3 a_27_74.n2 301.264
R10 a_27_74.n2 a_27_74.n1 286.846
R11 a_27_74.n2 a_27_74.n0 271.06
R12 a_27_74.n3 a_27_74.t3 46.1724
R13 a_27_74.t2 a_27_74.n3 46.1724
R14 a_27_74.n1 a_27_74.t0 40.0005
R15 a_27_74.n1 a_27_74.t1 40.0005
R16 a_114_464.t0 a_114_464.t1 73.8755
R17 VPB.t10 VPB.t13 1187.5
R18 VPB.t9 VPB.t10 694.625
R19 VPB.t4 VPB.t12 577.152
R20 VPB.t11 VPB.t16 497.985
R21 VPB.t3 VPB.t0 495.43
R22 VPB.t2 VPB.t14 495.43
R23 VPB.t8 VPB.t1 487.769
R24 VPB.t14 VPB.t8 477.555
R25 VPB.t1 VPB.t3 362.635
R26 VPB.t16 VPB.t9 347.312
R27 VPB.t12 VPB.t5 347.312
R28 VPB.t17 VPB.t2 265.591
R29 VPB.t13 VPB.t6 255.376
R30 VPB VPB.t15 252.823
R31 VPB.t7 VPB.t11 229.839
R32 VPB.t6 VPB.t17 219.625
R33 VPB.t5 VPB.t7 199.195
R34 VPB.t15 VPB.t4 199.195
R35 a_1295_74.t0 a_1295_74.n5 1104.1
R36 a_1295_74.n2 a_1295_74.n1 577.374
R37 a_1295_74.n3 a_1295_74.n2 359.894
R38 a_1295_74.n1 a_1295_74.t3 295.627
R39 a_1295_74.n3 a_1295_74.t4 295.627
R40 a_1295_74.n5 a_1295_74.t2 281.168
R41 a_1295_74.n1 a_1295_74.t5 243.679
R42 a_1295_74.n4 a_1295_74.n0 204.048
R43 a_1295_74.n2 a_1295_74.t1 171.913
R44 a_1295_74.n5 a_1295_74.n4 165.488
R45 a_1295_74.n4 a_1295_74.n3 149.421
R46 a_1688_97.n2 a_1688_97.n0 654.865
R47 a_1688_97.n1 a_1688_97.t5 284.38
R48 a_1688_97.n3 a_1688_97.n2 256.529
R49 a_1688_97.n2 a_1688_97.n1 251.606
R50 a_1688_97.n1 a_1688_97.t4 205.922
R51 a_1688_97.t0 a_1688_97.n3 111.43
R52 a_1688_97.n0 a_1688_97.t2 93.81
R53 a_1688_97.n0 a_1688_97.t1 70.3576
R54 a_1688_97.n3 a_1688_97.t3 40.0005
R55 a_1890_508.t0 a_1890_508.t1 131.333
R56 DE.n0 DE.t3 345.433
R57 DE.n1 DE.t0 306.873
R58 DE.n2 DE.n0 253.853
R59 DE DE.n2 155.685
R60 DE.n1 DE.t2 147.814
R61 DE.n0 DE.t1 126.927
R62 DE.n2 DE.n1 52.5823
R63 a_143_74.t0 a_143_74.t1 68.5719
R64 VGND.n39 VGND.t1 286.334
R65 VGND.n26 VGND.t6 285.053
R66 VGND.n60 VGND.t10 247.498
R67 VGND.n47 VGND.n46 226.216
R68 VGND.n58 VGND.n2 214.673
R69 VGND.n31 VGND.n11 211.369
R70 VGND.n20 VGND.n19 185
R71 VGND.n18 VGND.n17 185
R72 VGND.n16 VGND.t5 179.31
R73 VGND.n19 VGND.n18 178.571
R74 VGND.n11 VGND.t8 81.4873
R75 VGND.n18 VGND.t4 60.0005
R76 VGND.n11 VGND.t11 52.8309
R77 VGND.n19 VGND.t3 40.0005
R78 VGND.n46 VGND.t7 40.0005
R79 VGND.n46 VGND.t2 40.0005
R80 VGND.n2 VGND.t0 40.0005
R81 VGND.n2 VGND.t9 40.0005
R82 VGND.n21 VGND.n13 36.1417
R83 VGND.n25 VGND.n13 36.1417
R84 VGND.n27 VGND.n10 36.1417
R85 VGND.n33 VGND.n32 36.1417
R86 VGND.n33 VGND.n8 36.1417
R87 VGND.n37 VGND.n8 36.1417
R88 VGND.n38 VGND.n37 36.1417
R89 VGND.n40 VGND.n6 36.1417
R90 VGND.n45 VGND.n44 36.1417
R91 VGND.n48 VGND.n45 36.1417
R92 VGND.n52 VGND.n4 36.1417
R93 VGND.n53 VGND.n52 36.1417
R94 VGND.n54 VGND.n53 36.1417
R95 VGND.n54 VGND.n1 36.1417
R96 VGND.n27 VGND.n26 29.3652
R97 VGND.n32 VGND.n31 29.3652
R98 VGND.n59 VGND.n58 29.3652
R99 VGND.n26 VGND.n25 24.0946
R100 VGND.n31 VGND.n10 24.0946
R101 VGND.n60 VGND.n59 20.3299
R102 VGND.n58 VGND.n1 18.0711
R103 VGND.n44 VGND.n6 16.5652
R104 VGND.n47 VGND.n4 14.6829
R105 VGND.n59 VGND.n0 9.3005
R106 VGND.n58 VGND.n57 9.3005
R107 VGND.n56 VGND.n1 9.3005
R108 VGND.n55 VGND.n54 9.3005
R109 VGND.n53 VGND.n3 9.3005
R110 VGND.n52 VGND.n51 9.3005
R111 VGND.n50 VGND.n4 9.3005
R112 VGND.n49 VGND.n48 9.3005
R113 VGND.n45 VGND.n5 9.3005
R114 VGND.n44 VGND.n43 9.3005
R115 VGND.n42 VGND.n6 9.3005
R116 VGND.n41 VGND.n40 9.3005
R117 VGND.n38 VGND.n7 9.3005
R118 VGND.n37 VGND.n36 9.3005
R119 VGND.n35 VGND.n8 9.3005
R120 VGND.n34 VGND.n33 9.3005
R121 VGND.n32 VGND.n9 9.3005
R122 VGND.n31 VGND.n30 9.3005
R123 VGND.n29 VGND.n10 9.3005
R124 VGND.n28 VGND.n27 9.3005
R125 VGND.n26 VGND.n12 9.3005
R126 VGND.n25 VGND.n24 9.3005
R127 VGND.n23 VGND.n13 9.3005
R128 VGND.n22 VGND.n21 9.3005
R129 VGND.n15 VGND.n14 9.3005
R130 VGND.n17 VGND.n16 9.12543
R131 VGND.n21 VGND.n20 9.10724
R132 VGND.n39 VGND.n38 7.90638
R133 VGND.n61 VGND.n60 7.31635
R134 VGND.n17 VGND.n15 7.28809
R135 VGND.n20 VGND.n15 4.39174
R136 VGND.n40 VGND.n39 3.38874
R137 VGND.n48 VGND.n47 2.63579
R138 VGND VGND.n61 0.277182
R139 VGND.n16 VGND.n14 0.215162
R140 VGND.n61 VGND.n0 0.15365
R141 VGND.n22 VGND.n14 0.122949
R142 VGND.n23 VGND.n22 0.122949
R143 VGND.n24 VGND.n23 0.122949
R144 VGND.n24 VGND.n12 0.122949
R145 VGND.n28 VGND.n12 0.122949
R146 VGND.n29 VGND.n28 0.122949
R147 VGND.n30 VGND.n29 0.122949
R148 VGND.n30 VGND.n9 0.122949
R149 VGND.n34 VGND.n9 0.122949
R150 VGND.n35 VGND.n34 0.122949
R151 VGND.n36 VGND.n35 0.122949
R152 VGND.n36 VGND.n7 0.122949
R153 VGND.n41 VGND.n7 0.122949
R154 VGND.n42 VGND.n41 0.122949
R155 VGND.n43 VGND.n42 0.122949
R156 VGND.n43 VGND.n5 0.122949
R157 VGND.n49 VGND.n5 0.122949
R158 VGND.n50 VGND.n49 0.122949
R159 VGND.n51 VGND.n50 0.122949
R160 VGND.n51 VGND.n3 0.122949
R161 VGND.n55 VGND.n3 0.122949
R162 VGND.n56 VGND.n55 0.122949
R163 VGND.n57 VGND.n56 0.122949
R164 VGND.n57 VGND.n0 0.122949
R165 VNB.n0 VNB 16352.8
R166 VNB VNB.n1 14356.6
R167 VNB.t4 VNB.t7 3129.66
R168 VNB.t5 VNB.t8 2598.43
R169 VNB.t16 VNB.t13 2563.78
R170 VNB.n1 VNB.n0 2527.91
R171 VNB.t8 VNB.t9 2286.61
R172 VNB.t17 VNB.t18 2286.61
R173 VNB.t3 VNB.t1 2263.52
R174 VNB.t19 VNB.t16 1743.83
R175 VNB.t1 VNB.t12 1570.6
R176 VNB.t15 VNB 1478.22
R177 VNB.n1 VNB.t6 1397.38
R178 VNB.t12 VNB.t19 1339.63
R179 VNB.t11 VNB.t2 1177.95
R180 VNB.t14 VNB.t4 993.177
R181 VNB.t7 VNB.t10 993.177
R182 VNB.t0 VNB.t17 993.177
R183 VNB.t2 VNB.t5 900.788
R184 VNB.t10 VNB.t0 900.788
R185 VNB.t18 VNB.t15 900.788
R186 VNB.t13 VNB.t11 831.496
R187 VNB.t6 VNB.t14 831.496
R188 VNB.n0 VNB.t3 704.462
R189 a_2385_74.n7 a_2385_74.n5 633.659
R190 a_2385_74.n2 a_2385_74.t5 294.288
R191 a_2385_74.n6 a_2385_74.n5 291.502
R192 a_2385_74.n1 a_2385_74.t6 242.875
R193 a_2385_74.n4 a_2385_74.n0 233.096
R194 a_2385_74.n4 a_2385_74.n3 225.889
R195 a_2385_74.n3 a_2385_74.t3 184.403
R196 a_2385_74.n1 a_2385_74.t4 157.453
R197 a_2385_74.n2 a_2385_74.n1 119.882
R198 a_2385_74.n7 a_2385_74.n6 107.456
R199 a_2385_74.n0 a_2385_74.t0 62.8576
R200 a_2385_74.n5 a_2385_74.n4 53.5438
R201 a_2385_74.n0 a_2385_74.t2 26.2505
R202 a_2385_74.n6 a_2385_74.t1 22.3551
R203 a_2385_74.n3 a_2385_74.n2 13.4525
R204 a_547_301.n0 a_547_301.t5 621.78
R205 a_547_301.t1 a_547_301.n3 367.854
R206 a_547_301.n2 a_547_301.t0 295.029
R207 a_547_301.n1 a_547_301.t3 255.863
R208 a_547_301.n1 a_547_301.t2 253.452
R209 a_547_301.n2 a_547_301.n1 190.869
R210 a_547_301.n3 a_547_301.n0 182.427
R211 a_547_301.n0 a_547_301.t4 138.441
R212 a_547_301.n3 a_547_301.n2 27.6853
R213 Q.n3 Q 589.707
R214 Q.n3 Q.n0 585
R215 Q.n4 Q.n3 585
R216 Q.n2 Q.t0 279.738
R217 Q.t0 Q.n1 279.738
R218 Q.n3 Q.t1 26.3844
R219 Q Q.n4 12.6123
R220 Q.n1 Q 12.2358
R221 Q Q.n0 10.9181
R222 Q Q.n2 9.22403
R223 Q.n2 Q 4.70638
R224 Q Q.n0 3.01226
R225 Q.n1 Q 1.69462
R226 Q.n4 Q 1.31815
R227 a_159_404.t1 a_159_404.n1 660.913
R228 a_159_404.n1 a_159_404.t2 461.729
R229 a_159_404.n0 a_159_404.t0 301.007
R230 a_159_404.n0 a_159_404.t3 271.57
R231 a_159_404.n1 a_159_404.n0 45.4738
R232 VPWR.n41 VPWR.t4 904.595
R233 VPWR.n25 VPWR.t5 859.285
R234 VPWR.n61 VPWR.t10 722.067
R235 VPWR.n46 VPWR.n5 613.928
R236 VPWR.n54 VPWR.n53 612.136
R237 VPWR.n28 VPWR.n27 604.976
R238 VPWR.n15 VPWR.n14 599.489
R239 VPWR.n16 VPWR.t2 266.74
R240 VPWR.n14 VPWR.t0 138.369
R241 VPWR.n53 VPWR.t9 116.969
R242 VPWR.n5 VPWR.t7 116.969
R243 VPWR.n14 VPWR.t1 102.531
R244 VPWR.n27 VPWR.t6 89.4026
R245 VPWR.n27 VPWR.t11 72.4603
R246 VPWR.n53 VPWR.t8 46.1724
R247 VPWR.n5 VPWR.t3 46.1724
R248 VPWR.n59 VPWR.n1 36.1417
R249 VPWR.n60 VPWR.n59 36.1417
R250 VPWR.n47 VPWR.n3 36.1417
R251 VPWR.n51 VPWR.n3 36.1417
R252 VPWR.n52 VPWR.n51 36.1417
R253 VPWR.n55 VPWR.n52 36.1417
R254 VPWR.n45 VPWR.n6 36.1417
R255 VPWR.n40 VPWR.n39 36.1417
R256 VPWR.n33 VPWR.n10 36.1417
R257 VPWR.n34 VPWR.n33 36.1417
R258 VPWR.n35 VPWR.n34 36.1417
R259 VPWR.n35 VPWR.n8 36.1417
R260 VPWR.n29 VPWR.n26 36.1417
R261 VPWR.n19 VPWR.n18 36.1417
R262 VPWR.n20 VPWR.n19 36.1417
R263 VPWR.n20 VPWR.n12 36.1417
R264 VPWR.n24 VPWR.n12 36.1417
R265 VPWR.n41 VPWR.n40 35.3887
R266 VPWR.n46 VPWR.n45 29.3652
R267 VPWR.n62 VPWR.n61 24.645
R268 VPWR.n47 VPWR.n46 24.0946
R269 VPWR.n54 VPWR.n1 16.9417
R270 VPWR.n41 VPWR.n6 12.0476
R271 VPWR.n39 VPWR.n8 11.2946
R272 VPWR.n18 VPWR.n15 9.78874
R273 VPWR.n29 VPWR.n28 9.41227
R274 VPWR.n18 VPWR.n17 9.3005
R275 VPWR.n19 VPWR.n13 9.3005
R276 VPWR.n21 VPWR.n20 9.3005
R277 VPWR.n22 VPWR.n12 9.3005
R278 VPWR.n24 VPWR.n23 9.3005
R279 VPWR.n26 VPWR.n11 9.3005
R280 VPWR.n30 VPWR.n29 9.3005
R281 VPWR.n31 VPWR.n10 9.3005
R282 VPWR.n33 VPWR.n32 9.3005
R283 VPWR.n34 VPWR.n9 9.3005
R284 VPWR.n36 VPWR.n35 9.3005
R285 VPWR.n37 VPWR.n8 9.3005
R286 VPWR.n39 VPWR.n38 9.3005
R287 VPWR.n40 VPWR.n7 9.3005
R288 VPWR.n42 VPWR.n41 9.3005
R289 VPWR.n43 VPWR.n6 9.3005
R290 VPWR.n45 VPWR.n44 9.3005
R291 VPWR.n46 VPWR.n4 9.3005
R292 VPWR.n48 VPWR.n47 9.3005
R293 VPWR.n49 VPWR.n3 9.3005
R294 VPWR.n51 VPWR.n50 9.3005
R295 VPWR.n52 VPWR.n2 9.3005
R296 VPWR.n56 VPWR.n55 9.3005
R297 VPWR.n57 VPWR.n1 9.3005
R298 VPWR.n59 VPWR.n58 9.3005
R299 VPWR.n60 VPWR.n0 9.3005
R300 VPWR.n26 VPWR.n25 7.90638
R301 VPWR.n16 VPWR.n15 7.29491
R302 VPWR.n25 VPWR.n24 3.38874
R303 VPWR.n28 VPWR.n10 1.88285
R304 VPWR.n61 VPWR.n60 0.376971
R305 VPWR.n55 VPWR.n54 0.376971
R306 VPWR.n17 VPWR.n16 0.221392
R307 VPWR VPWR.n62 0.163644
R308 VPWR.n62 VPWR.n0 0.144205
R309 VPWR.n17 VPWR.n13 0.122949
R310 VPWR.n21 VPWR.n13 0.122949
R311 VPWR.n22 VPWR.n21 0.122949
R312 VPWR.n23 VPWR.n22 0.122949
R313 VPWR.n23 VPWR.n11 0.122949
R314 VPWR.n30 VPWR.n11 0.122949
R315 VPWR.n31 VPWR.n30 0.122949
R316 VPWR.n32 VPWR.n31 0.122949
R317 VPWR.n32 VPWR.n9 0.122949
R318 VPWR.n36 VPWR.n9 0.122949
R319 VPWR.n37 VPWR.n36 0.122949
R320 VPWR.n38 VPWR.n37 0.122949
R321 VPWR.n38 VPWR.n7 0.122949
R322 VPWR.n42 VPWR.n7 0.122949
R323 VPWR.n43 VPWR.n42 0.122949
R324 VPWR.n44 VPWR.n43 0.122949
R325 VPWR.n44 VPWR.n4 0.122949
R326 VPWR.n48 VPWR.n4 0.122949
R327 VPWR.n49 VPWR.n48 0.122949
R328 VPWR.n50 VPWR.n49 0.122949
R329 VPWR.n50 VPWR.n2 0.122949
R330 VPWR.n56 VPWR.n2 0.122949
R331 VPWR.n57 VPWR.n56 0.122949
R332 VPWR.n58 VPWR.n57 0.122949
R333 VPWR.n58 VPWR.n0 0.122949
R334 a_1824_97.t0 a_1824_97.t1 122.858
R335 a_554_463.t0 a_554_463.t1 73.8755
R336 a_505_111.t0 a_505_111.t1 68.5719
R337 a_1910_71.t1 a_1910_71.n3 851.861
R338 a_1910_71.n1 a_1910_71.t2 377.055
R339 a_1910_71.n0 a_1910_71.t5 281.168
R340 a_1910_71.n2 a_1910_71.t0 240.238
R341 a_1910_71.n2 a_1910_71.n1 212.829
R342 a_1910_71.n0 a_1910_71.t4 179.154
R343 a_1910_71.n1 a_1910_71.t3 170.865
R344 a_1910_71.n3 a_1910_71.n0 95.7752
R345 a_1910_71.n3 a_1910_71.n2 26.5381
R346 CLK.n1 CLK.t0 269.293
R347 CLK.n1 CLK.n0 177.981
R348 CLK CLK.n1 158.788
R349 a_669_111.n0 a_669_111.t4 730.457
R350 a_669_111.t3 a_669_111.n2 710.365
R351 a_669_111.t3 a_669_111.n3 710.365
R352 a_669_111.n3 a_669_111.t2 358.959
R353 a_669_111.n1 a_669_111.t1 343.772
R354 a_669_111.n0 a_669_111.t0 338.498
R355 a_669_111.n2 a_669_111.n1 180.804
R356 a_669_111.n1 a_669_111.n0 119.341
R357 a_669_111.n3 a_669_111.n2 16.0005
R358 a_2487_74.t0 a_2487_74.t1 68.5719
R359 SCE.t2 SCE.t1 626.601
R360 SCE.t0 SCE.t3 569.029
R361 SCE.n0 SCE.t0 335.793
R362 SCE SCE.n0 157.237
R363 SCE.n0 SCE.t2 134.96
R364 a_639_85.t1 a_639_85.n2 656.511
R365 a_639_85.n2 a_639_85.n0 372.204
R366 a_639_85.n1 a_639_85.t2 313.983
R367 a_639_85.n1 a_639_85.t0 246.389
R368 a_639_85.n2 a_639_85.n1 32.1576
R369 a_1026_125.t0 a_1026_125.t1 60.0005
R370 a_2313_74.t0 a_2313_74.t1 39.3755
R371 a_2274_392.t0 a_2274_392.t1 154.645
R372 SCD.n0 SCD.t1 272.866
R373 SCD.n0 SCD.t0 210.474
R374 SCD SCD.n0 165.341
C0 VGND DE 0.037318f
C1 SCE CLK 0.003737f
C2 VPWR D 0.012559f
C3 DE VPB 0.165139f
C4 VGND a_1492_74# 0.54695f
C5 Q VPWR 0.130719f
C6 VGND VPWR 0.068739f
C7 a_1492_74# VPB 0.225504f
C8 VGND D 0.017722f
C9 VPWR VPB 0.453221f
C10 SCD VPWR 0.013229f
C11 SCE DE 6.97e-20
C12 Q VGND 0.102271f
C13 CLK VPWR 0.013331f
C14 VPB D 0.071654f
C15 Q VPB 0.01206f
C16 SCE a_1492_74# 3.61e-19
C17 VGND VPB 0.016741f
C18 SCD VGND 0.0231f
C19 SCE VPWR 0.031355f
C20 CLK VGND 0.017315f
C21 SCD VPB 0.061524f
C22 VPWR DE 0.022365f
C23 CLK VPB 0.039424f
C24 SCE VGND 0.063484f
C25 SCD CLK 0.003409f
C26 DE D 0.04224f
C27 a_1492_74# VPWR 0.017509f
C28 SCE VPB 0.182669f
C29 SCE SCD 0.129102f
C30 Q VNB 0.032549f
C31 VGND VNB 1.85704f
C32 CLK VNB 0.122603f
C33 SCD VNB 0.10684f
C34 SCE VNB 0.347229f
C35 DE VNB 0.294181f
C36 VPWR VNB 1.39402f
C37 D VNB 0.186413f
C38 VPB VNB 3.5208f
C39 a_1492_74# VNB 0.362449f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sedfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sedfxtp_2 VNB VPB VPWR VGND SCE CLK D DE SCD Q
X0 a_575_463.t0 DE.t0 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1696 ps=1.17 w=0.64 l=0.15
X1 VPWR.t5 DE.t1 a_180_290.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X2 a_1872_97.t0 a_1538_74.t2 a_1736_97.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.11235 pd=0.955 as=0.1113 ps=0.95 w=0.42 l=0.15
X3 VGND.t0 a_1979_71.t2 a_1872_97.t1 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.176 pd=1.265 as=0.11235 ps=0.955 w=0.42 l=0.15
X4 a_40_464.t4 a_548_87.t2 a_500_113.t0 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.08925 pd=0.845 as=0.0504 ps=0.66 w=0.42 l=0.15
X5 a_693_113.t3 SCE.t0 a_1068_125.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR.t1 a_180_290.t2 a_129_464.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0864 ps=0.91 w=0.64 l=0.15
X7 VGND.t12 a_548_87.t3 a_2569_74.t0 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.20055 pd=1.375 as=0.0504 ps=0.66 w=0.42 l=0.15
X8 a_138_74.t0 D.t0 a_40_464.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 a_2402_74.t0 a_1979_71.t3 VGND.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1824 ps=1.85 w=0.64 l=0.15
X10 VPWR.t9 SCE.t1 a_663_87.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1856 ps=1.86 w=0.64 l=0.15
X11 a_500_113.t1 a_180_290.t3 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 a_1079_455.t0 SCD.t0 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1696 ps=1.17 w=0.64 l=0.15
X13 a_1979_71.t0 a_1736_97.t4 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.147875 ps=1.355 w=0.84 l=0.15
X14 a_2474_74.t1 a_1538_74.t3 a_2402_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.09575 pd=0.965 as=0.0672 ps=0.85 w=0.64 l=0.15
X15 a_1936_508.t1 a_1340_74.t2 a_1736_97.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.084 pd=0.82 as=0.063 ps=0.72 w=0.42 l=0.15
X16 a_1068_125.t0 SCD.t1 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X17 VPWR.t8 a_2474_74.t4 Q.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X18 a_1736_97.t2 a_1538_74.t4 a_693_113.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X19 a_2357_392.t0 a_1979_71.t4 VPWR.t12 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.405 pd=1.81 as=0.305 ps=2.61 w=1 l=0.15
X20 a_1538_74.t1 a_1340_74.t3 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X21 a_693_113.t0 a_663_87.t2 a_40_464.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.08925 ps=0.845 w=0.42 l=0.15
X22 a_2474_74.t3 a_1340_74.t4 a_2357_392.t1 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.15875 pd=1.39 as=0.405 ps=1.81 w=1 l=0.15
X23 a_1340_74.t1 CLK.t0 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2183 ps=2.07 w=0.74 l=0.15
X24 a_1736_97.t0 a_1340_74.t5 a_693_113.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1197 ps=1.41 w=0.42 l=0.15
X25 a_1538_74.t0 a_1340_74.t6 VGND.t10 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X26 VPWR.t4 a_1979_71.t5 a_1936_508.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.147875 pd=1.355 as=0.084 ps=0.82 w=0.42 l=0.15
X27 VGND.t11 a_2474_74.t5 Q.t0 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VGND.t4 SCE.t2 a_663_87.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X29 VPWR.t13 a_548_87.t4 a_2657_508.t0 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.14675 pd=1.2 as=0.0567 ps=0.69 w=0.42 l=0.15
X30 a_129_464.t1 D.t1 a_40_464.t5 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1888 ps=1.87 w=0.64 l=0.15
X31 a_2657_508.t1 a_1538_74.t5 a_2474_74.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.15875 ps=1.39 w=0.42 l=0.15
X32 VGND.t9 DE.t2 a_138_74.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X33 a_548_87.t0 a_2474_74.t6 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.14675 ps=1.2 w=0.64 l=0.15
X34 a_2569_74.t1 a_1340_74.t7 a_2474_74.t2 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.09575 ps=0.965 w=0.42 l=0.15
X35 a_1340_74.t0 CLK.t1 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.336 ps=2.84 w=1.12 l=0.15
X36 a_693_113.t4 SCE.t3 a_40_464.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1856 pd=1.86 as=0.096 ps=0.94 w=0.64 l=0.15
X37 a_40_464.t3 a_548_87.t5 a_575_463.t1 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0768 ps=0.88 w=0.64 l=0.15
X38 Q.t1 a_2474_74.t7 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.3304 ps=2.83 w=1.12 l=0.15
X39 a_1979_71.t1 a_1736_97.t5 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.176 ps=1.265 w=0.64 l=0.15
X40 VGND.t8 DE.t3 a_180_290.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X41 a_548_87.t1 a_2474_74.t8 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.20055 ps=1.375 w=0.42 l=0.15
R0 DE.n0 DE.t0 345.433
R1 DE.n1 DE.t2 318.12
R2 DE.n2 DE.n0 287.594
R3 DE DE.n2 155.685
R4 DE.n1 DE.t3 139.78
R5 DE.n0 DE.t1 126.927
R6 DE.n2 DE.n1 51.1217
R7 VPWR.n49 VPWR.t0 877.958
R8 VPWR.n10 VPWR.t11 875.822
R9 VPWR.n15 VPWR.t12 833.683
R10 VPWR.n0 VPWR.t1 722.067
R11 VPWR.n54 VPWR.n7 613.928
R12 VPWR.n61 VPWR.n3 612.136
R13 VPWR.n37 VPWR.n14 604.976
R14 VPWR.n25 VPWR.n24 585
R15 VPWR.n20 VPWR.t8 349.394
R16 VPWR.n19 VPWR.t3 249.631
R17 VPWR.n24 VPWR.t2 121.293
R18 VPWR.n24 VPWR.t13 119.608
R19 VPWR.n3 VPWR.t5 116.969
R20 VPWR.n7 VPWR.t9 116.969
R21 VPWR.n14 VPWR.t10 99.5923
R22 VPWR.n14 VPWR.t4 71.409
R23 VPWR.n3 VPWR.t6 46.1724
R24 VPWR.n7 VPWR.t7 46.1724
R25 VPWR.n63 VPWR.n62 36.1417
R26 VPWR.n56 VPWR.n55 36.1417
R27 VPWR.n56 VPWR.n4 36.1417
R28 VPWR.n60 VPWR.n4 36.1417
R29 VPWR.n53 VPWR.n8 36.1417
R30 VPWR.n48 VPWR.n47 36.1417
R31 VPWR.n41 VPWR.n12 36.1417
R32 VPWR.n42 VPWR.n41 36.1417
R33 VPWR.n43 VPWR.n42 36.1417
R34 VPWR.n36 VPWR.n35 36.1417
R35 VPWR.n26 VPWR.n17 36.1417
R36 VPWR.n30 VPWR.n17 36.1417
R37 VPWR.n31 VPWR.n30 36.1417
R38 VPWR.n32 VPWR.n31 36.1417
R39 VPWR.n55 VPWR.n54 33.8829
R40 VPWR.n23 VPWR.n22 32.0423
R41 VPWR.n63 VPWR.n0 28.6123
R42 VPWR.n61 VPWR.n60 28.6123
R43 VPWR.n37 VPWR.n12 28.2358
R44 VPWR.n49 VPWR.n8 27.1064
R45 VPWR.n62 VPWR.n61 24.8476
R46 VPWR.n22 VPWR.n19 24.0946
R47 VPWR.n47 VPWR.n10 23.7181
R48 VPWR.n43 VPWR.n10 23.7181
R49 VPWR.n49 VPWR.n48 19.9534
R50 VPWR.n54 VPWR.n53 19.577
R51 VPWR.n37 VPWR.n36 19.2005
R52 VPWR.n22 VPWR.n21 9.3005
R53 VPWR.n23 VPWR.n18 9.3005
R54 VPWR.n27 VPWR.n26 9.3005
R55 VPWR.n28 VPWR.n17 9.3005
R56 VPWR.n30 VPWR.n29 9.3005
R57 VPWR.n31 VPWR.n16 9.3005
R58 VPWR.n33 VPWR.n32 9.3005
R59 VPWR.n35 VPWR.n34 9.3005
R60 VPWR.n36 VPWR.n13 9.3005
R61 VPWR.n38 VPWR.n37 9.3005
R62 VPWR.n39 VPWR.n12 9.3005
R63 VPWR.n41 VPWR.n40 9.3005
R64 VPWR.n42 VPWR.n11 9.3005
R65 VPWR.n44 VPWR.n43 9.3005
R66 VPWR.n45 VPWR.n10 9.3005
R67 VPWR.n47 VPWR.n46 9.3005
R68 VPWR.n48 VPWR.n9 9.3005
R69 VPWR.n50 VPWR.n49 9.3005
R70 VPWR.n51 VPWR.n8 9.3005
R71 VPWR.n53 VPWR.n52 9.3005
R72 VPWR.n54 VPWR.n6 9.3005
R73 VPWR.n55 VPWR.n5 9.3005
R74 VPWR.n57 VPWR.n56 9.3005
R75 VPWR.n58 VPWR.n4 9.3005
R76 VPWR.n60 VPWR.n59 9.3005
R77 VPWR.n61 VPWR.n2 9.3005
R78 VPWR.n62 VPWR.n1 9.3005
R79 VPWR.n64 VPWR.n63 9.3005
R80 VPWR.n32 VPWR.n15 8.28285
R81 VPWR.n65 VPWR.n0 7.2096
R82 VPWR.n20 VPWR.n19 6.58468
R83 VPWR.n26 VPWR.n25 5.27109
R84 VPWR.n25 VPWR.n23 3.34691
R85 VPWR.n35 VPWR.n15 2.25932
R86 VPWR.n21 VPWR.n20 0.670526
R87 VPWR VPWR.n65 0.275532
R88 VPWR.n65 VPWR.n64 0.155274
R89 VPWR.n21 VPWR.n18 0.122949
R90 VPWR.n27 VPWR.n18 0.122949
R91 VPWR.n28 VPWR.n27 0.122949
R92 VPWR.n29 VPWR.n28 0.122949
R93 VPWR.n29 VPWR.n16 0.122949
R94 VPWR.n33 VPWR.n16 0.122949
R95 VPWR.n34 VPWR.n33 0.122949
R96 VPWR.n34 VPWR.n13 0.122949
R97 VPWR.n38 VPWR.n13 0.122949
R98 VPWR.n39 VPWR.n38 0.122949
R99 VPWR.n40 VPWR.n39 0.122949
R100 VPWR.n40 VPWR.n11 0.122949
R101 VPWR.n44 VPWR.n11 0.122949
R102 VPWR.n45 VPWR.n44 0.122949
R103 VPWR.n46 VPWR.n45 0.122949
R104 VPWR.n46 VPWR.n9 0.122949
R105 VPWR.n50 VPWR.n9 0.122949
R106 VPWR.n51 VPWR.n50 0.122949
R107 VPWR.n52 VPWR.n51 0.122949
R108 VPWR.n52 VPWR.n6 0.122949
R109 VPWR.n6 VPWR.n5 0.122949
R110 VPWR.n57 VPWR.n5 0.122949
R111 VPWR.n58 VPWR.n57 0.122949
R112 VPWR.n59 VPWR.n58 0.122949
R113 VPWR.n59 VPWR.n2 0.122949
R114 VPWR.n2 VPWR.n1 0.122949
R115 VPWR.n64 VPWR.n1 0.122949
R116 a_575_463.t0 a_575_463.t1 73.8755
R117 VPB.t10 VPB.t2 732.931
R118 VPB.t2 VPB.t15 709.947
R119 VPB.t3 VPB.t8 577.152
R120 VPB.t14 VPB.t17 520.968
R121 VPB.t4 VPB.t5 515.861
R122 VPB.t15 VPB.t13 515.861
R123 VPB.t0 VPB.t12 510.753
R124 VPB.t17 VPB.t18 490.324
R125 VPB.t19 VPB.t4 362.635
R126 VPB.t12 VPB.t10 347.312
R127 VPB.t8 VPB.t9 347.312
R128 VPB VPB.t16 291.13
R129 VPB.t7 VPB.t6 280.914
R130 VPB.t18 VPB.t1 275.807
R131 VPB.t6 VPB.t14 273.253
R132 VPB.t5 VPB.t11 237.5
R133 VPB.t13 VPB.t7 229.839
R134 VPB.t20 VPB.t0 229.839
R135 VPB.t1 VPB.t19 214.517
R136 VPB.t16 VPB.t3 214.517
R137 VPB.t9 VPB.t20 199.195
R138 a_180_290.t0 a_180_290.n1 660.913
R139 a_180_290.n1 a_180_290.t3 446.959
R140 a_180_290.n0 a_180_290.t1 291.62
R141 a_180_290.n0 a_180_290.t2 261.834
R142 a_180_290.n1 a_180_290.n0 53.1323
R143 a_1538_74.t1 a_1538_74.n3 857.567
R144 a_1538_74.n0 a_1538_74.t5 565.143
R145 a_1538_74.n0 a_1538_74.t3 440.704
R146 a_1538_74.n3 a_1538_74.t4 342.803
R147 a_1538_74.n1 a_1538_74.t2 294.272
R148 a_1538_74.n1 a_1538_74.n0 266.074
R149 a_1538_74.n2 a_1538_74.t0 206.231
R150 a_1538_74.n3 a_1538_74.n2 105.035
R151 a_1538_74.n2 a_1538_74.n1 86.4975
R152 a_1736_97.n2 a_1736_97.n0 645.131
R153 a_1736_97.n1 a_1736_97.t5 282.07
R154 a_1736_97.n3 a_1736_97.n2 267.825
R155 a_1736_97.n2 a_1736_97.n1 248.264
R156 a_1736_97.n1 a_1736_97.t4 203.611
R157 a_1736_97.t0 a_1736_97.n3 111.43
R158 a_1736_97.n0 a_1736_97.t3 70.3576
R159 a_1736_97.n0 a_1736_97.t2 70.3576
R160 a_1736_97.n3 a_1736_97.t1 40.0005
R161 a_1872_97.t0 a_1872_97.t1 152.857
R162 VNB.n0 VNB 16872.4
R163 VNB VNB.n1 14472.1
R164 VNB.t7 VNB.t16 3441.47
R165 VNB.t8 VNB.t0 3175.85
R166 VNB.t9 VNB.t18 2748.56
R167 VNB.t20 VNB.t7 2552.23
R168 VNB.t15 VNB.t1 2286.61
R169 VNB.t13 VNB.t14 2286.61
R170 VNB.t17 VNB.t9 1790.03
R171 VNB.t10 VNB.n0 1587.27
R172 VNB.t5 VNB.t17 1582.15
R173 VNB.t1 VNB.t5 1570.6
R174 VNB.t2 VNB 1420.47
R175 VNB.n1 VNB.t3 1328.08
R176 VNB.t0 VNB.t19 1328.08
R177 VNB.t12 VNB.t8 1154.86
R178 VNB.t4 VNB.t11 1097.11
R179 VNB.t6 VNB.t13 993.177
R180 VNB.n1 VNB.t10 992.043
R181 VNB.t11 VNB.t20 900.788
R182 VNB.t19 VNB.t6 900.788
R183 VNB.t14 VNB.t2 900.788
R184 VNB.t18 VNB.t4 831.496
R185 VNB.t3 VNB.t12 831.496
R186 VNB.n0 VNB.t15 716.01
R187 a_1979_71.t0 a_1979_71.n0 817.962
R188 a_1979_71.n2 a_1979_71.t5 371.37
R189 a_1979_71.n1 a_1979_71.t4 282.507
R190 a_1979_71.n0 a_1979_71.t1 233.179
R191 a_1979_71.n0 a_1979_71.n2 208.798
R192 a_1979_71.n1 a_1979_71.t3 188.921
R193 a_1979_71.n2 a_1979_71.t2 176.964
R194 a_1979_71.n0 a_1979_71.n1 108.347
R195 VGND.n6 VGND.t6 301.88
R196 VGND.n27 VGND.t1 285.053
R197 VGND.n60 VGND.t9 247.498
R198 VGND.n48 VGND.n47 216.225
R199 VGND.n58 VGND.n2 215.061
R200 VGND.n11 VGND.n10 209.875
R201 VGND.n21 VGND.n20 185
R202 VGND.n19 VGND.n18 185
R203 VGND.n20 VGND.n19 172.857
R204 VGND.n40 VGND.t10 171.77
R205 VGND.n17 VGND.t11 162.089
R206 VGND.n10 VGND.t5 83.7303
R207 VGND.n19 VGND.t3 60.0005
R208 VGND.n47 VGND.t4 60.0005
R209 VGND.n10 VGND.t0 55.0739
R210 VGND.n20 VGND.t12 40.0005
R211 VGND.n47 VGND.t7 40.0005
R212 VGND.n2 VGND.t2 40.0005
R213 VGND.n2 VGND.t8 40.0005
R214 VGND.n23 VGND.n22 36.1417
R215 VGND.n23 VGND.n13 36.1417
R216 VGND.n29 VGND.n28 36.1417
R217 VGND.n34 VGND.n33 36.1417
R218 VGND.n35 VGND.n34 36.1417
R219 VGND.n35 VGND.n8 36.1417
R220 VGND.n39 VGND.n8 36.1417
R221 VGND.n46 VGND.n45 36.1417
R222 VGND.n52 VGND.n4 36.1417
R223 VGND.n53 VGND.n52 36.1417
R224 VGND.n54 VGND.n53 36.1417
R225 VGND.n54 VGND.n1 36.1417
R226 VGND.n41 VGND.n6 35.0123
R227 VGND.n29 VGND.n11 32.7534
R228 VGND.n40 VGND.n39 32.7534
R229 VGND.n59 VGND.n58 27.4829
R230 VGND.n27 VGND.n13 26.7299
R231 VGND.n28 VGND.n27 26.7299
R232 VGND.n48 VGND.n4 24.4711
R233 VGND.n48 VGND.n46 22.9652
R234 VGND.n60 VGND.n59 22.2123
R235 VGND.n41 VGND.n40 20.7064
R236 VGND.n58 VGND.n1 19.9534
R237 VGND.n33 VGND.n11 19.577
R238 VGND.n45 VGND.n6 17.6946
R239 VGND.n18 VGND.n17 11.4891
R240 VGND.n59 VGND.n0 9.3005
R241 VGND.n58 VGND.n57 9.3005
R242 VGND.n56 VGND.n1 9.3005
R243 VGND.n55 VGND.n54 9.3005
R244 VGND.n53 VGND.n3 9.3005
R245 VGND.n52 VGND.n51 9.3005
R246 VGND.n50 VGND.n4 9.3005
R247 VGND.n49 VGND.n48 9.3005
R248 VGND.n46 VGND.n5 9.3005
R249 VGND.n45 VGND.n44 9.3005
R250 VGND.n43 VGND.n6 9.3005
R251 VGND.n42 VGND.n41 9.3005
R252 VGND.n16 VGND.n15 9.3005
R253 VGND.n22 VGND.n14 9.3005
R254 VGND.n24 VGND.n23 9.3005
R255 VGND.n25 VGND.n13 9.3005
R256 VGND.n27 VGND.n26 9.3005
R257 VGND.n28 VGND.n12 9.3005
R258 VGND.n30 VGND.n29 9.3005
R259 VGND.n31 VGND.n11 9.3005
R260 VGND.n33 VGND.n32 9.3005
R261 VGND.n34 VGND.n9 9.3005
R262 VGND.n36 VGND.n35 9.3005
R263 VGND.n37 VGND.n8 9.3005
R264 VGND.n39 VGND.n38 9.3005
R265 VGND.n40 VGND.n7 9.3005
R266 VGND.n61 VGND.n60 7.22818
R267 VGND.n21 VGND.n15 5.10377
R268 VGND.n18 VGND.n15 5.02011
R269 VGND.n22 VGND.n21 3.51423
R270 VGND VGND.n61 0.27582
R271 VGND.n17 VGND.n16 0.173703
R272 VGND.n61 VGND.n0 0.154991
R273 VGND.n16 VGND.n14 0.122949
R274 VGND.n24 VGND.n14 0.122949
R275 VGND.n25 VGND.n24 0.122949
R276 VGND.n26 VGND.n25 0.122949
R277 VGND.n26 VGND.n12 0.122949
R278 VGND.n30 VGND.n12 0.122949
R279 VGND.n31 VGND.n30 0.122949
R280 VGND.n32 VGND.n31 0.122949
R281 VGND.n32 VGND.n9 0.122949
R282 VGND.n36 VGND.n9 0.122949
R283 VGND.n37 VGND.n36 0.122949
R284 VGND.n38 VGND.n37 0.122949
R285 VGND.n38 VGND.n7 0.122949
R286 VGND.n42 VGND.n7 0.122949
R287 VGND.n43 VGND.n42 0.122949
R288 VGND.n44 VGND.n43 0.122949
R289 VGND.n44 VGND.n5 0.122949
R290 VGND.n49 VGND.n5 0.122949
R291 VGND.n50 VGND.n49 0.122949
R292 VGND.n51 VGND.n50 0.122949
R293 VGND.n51 VGND.n3 0.122949
R294 VGND.n55 VGND.n3 0.122949
R295 VGND.n56 VGND.n55 0.122949
R296 VGND.n57 VGND.n56 0.122949
R297 VGND.n57 VGND.n0 0.122949
R298 a_548_87.n0 a_548_87.t3 642.668
R299 a_548_87.t0 a_548_87.n3 357.031
R300 a_548_87.n2 a_548_87.t1 279.452
R301 a_548_87.n1 a_548_87.t5 274.327
R302 a_548_87.n1 a_548_87.t2 250.933
R303 a_548_87.n2 a_548_87.n1 217.243
R304 a_548_87.n3 a_548_87.n0 200.76
R305 a_548_87.n0 a_548_87.t4 138.441
R306 a_548_87.n3 a_548_87.n2 42.262
R307 a_500_113.t0 a_500_113.t1 68.5719
R308 a_40_464.n0 a_40_464.t5 356.26
R309 a_40_464.n0 a_40_464.t2 345.396
R310 a_40_464.n3 a_40_464.n2 301.264
R311 a_40_464.n2 a_40_464.n1 284.346
R312 a_40_464.n2 a_40_464.n0 273.318
R313 a_40_464.n1 a_40_464.t0 61.4291
R314 a_40_464.n1 a_40_464.t4 60.0005
R315 a_40_464.t1 a_40_464.n3 46.1724
R316 a_40_464.n3 a_40_464.t3 46.1724
R317 SCE.t2 SCE.t0 649.093
R318 SCE.t1 SCE.t3 577.062
R319 SCE.n0 SCE.t1 335.435
R320 SCE SCE.n0 159.565
R321 SCE.n0 SCE.t2 134.601
R322 a_1068_125.t0 a_1068_125.t1 60.0005
R323 a_693_113.n0 a_693_113.t2 715.313
R324 a_693_113.t4 a_693_113.n2 703.88
R325 a_693_113.t4 a_693_113.n3 703.88
R326 a_693_113.n3 a_693_113.t0 358.594
R327 a_693_113.n0 a_693_113.t1 341.135
R328 a_693_113.n1 a_693_113.t3 329.356
R329 a_693_113.n2 a_693_113.n1 198.935
R330 a_693_113.n1 a_693_113.n0 133.701
R331 a_693_113.n3 a_693_113.n2 16.0005
R332 a_129_464.t0 a_129_464.t1 83.1099
R333 a_2569_74.t0 a_2569_74.t1 68.5719
R334 a_663_87.t1 a_663_87.n2 655.981
R335 a_663_87.n2 a_663_87.n0 375.022
R336 a_663_87.n1 a_663_87.t2 319.199
R337 a_663_87.n1 a_663_87.t0 247.482
R338 a_663_87.n2 a_663_87.n1 31.4839
R339 D.n0 D.t1 219.31
R340 D D.n0 160.254
R341 D.n1 D 154.19
R342 D.n1 D.t0 152.633
R343 D.n3 D.n2 152
R344 D.n2 D.n0 49.6611
R345 D.n2 D.n1 49.6611
R346 D.n3 D 9.26366
R347 D D.n3 3.2005
R348 a_138_74.t0 a_138_74.t1 68.5719
R349 a_2402_74.t0 a_2402_74.t1 39.3755
R350 SCD.n0 SCD.t0 272.866
R351 SCD.n0 SCD.t1 210.474
R352 SCD SCD.n0 162.41
R353 a_2474_74.n8 a_2474_74.n7 655.831
R354 a_2474_74.n7 a_2474_74.n0 328.276
R355 a_2474_74.n5 a_2474_74.t8 275.745
R356 a_2474_74.n2 a_2474_74.t4 255.382
R357 a_2474_74.n3 a_2474_74.t7 245.553
R358 a_2474_74.n6 a_2474_74.t6 218.644
R359 a_2474_74.n4 a_2474_74.n1 199.227
R360 a_2474_74.n2 a_2474_74.t5 199.227
R361 a_2474_74.n5 a_2474_74.n4 172.556
R362 a_2474_74.n7 a_2474_74.n6 93.4785
R363 a_2474_74.n3 a_2474_74.n2 78.0845
R364 a_2474_74.t3 a_2474_74.n8 77.2057
R365 a_2474_74.n8 a_2474_74.t0 70.3576
R366 a_2474_74.n6 a_2474_74.n5 56.5206
R367 a_2474_74.n0 a_2474_74.t1 40.5809
R368 a_2474_74.n0 a_2474_74.t2 40.0005
R369 a_2474_74.n4 a_2474_74.n3 4.8205
R370 a_1340_74.t0 a_1340_74.n5 841.75
R371 a_1340_74.n1 a_1340_74.n0 579.292
R372 a_1340_74.n2 a_1340_74.n1 410.296
R373 a_1340_74.n0 a_1340_74.t7 310.087
R374 a_1340_74.n2 a_1340_74.t5 273.134
R375 a_1340_74.n4 a_1340_74.t6 268.731
R376 a_1340_74.n0 a_1340_74.t4 231.629
R377 a_1340_74.n3 a_1340_74.t3 204.048
R378 a_1340_74.n5 a_1340_74.t1 185.839
R379 a_1340_74.n1 a_1340_74.t2 145.097
R380 a_1340_74.n3 a_1340_74.n2 100.782
R381 a_1340_74.n4 a_1340_74.n3 99.6869
R382 a_1340_74.n5 a_1340_74.n4 88.4945
R383 a_1936_508.t0 a_1936_508.t1 187.619
R384 Q Q.n0 211.446
R385 Q Q.t0 173.814
R386 Q.n0 Q.t2 28.1434
R387 Q.n0 Q.t1 27.2639
R388 a_2357_392.t0 a_2357_392.t1 159.571
R389 CLK.n0 CLK.t1 273.938
R390 CLK.n0 CLK.t0 171.913
R391 CLK CLK.n0 158.788
R392 a_2657_508.t0 a_2657_508.t1 126.644
C0 SCE VPB 0.183867f
C1 VPB CLK 0.044277f
C2 DE D 0.0429f
C3 D VPWR 0.013131f
C4 VGND DE 0.037274f
C5 VGND VPWR 0.058423f
C6 VGND SCD 0.03952f
C7 VGND Q 0.173866f
C8 DE VPB 0.173309f
C9 VPB VPWR 0.482128f
C10 VPB SCD 0.062614f
C11 Q VPB 0.010794f
C12 SCE CLK 0.003876f
C13 VGND D 0.020729f
C14 VPB D 0.073858f
C15 DE SCE 6.65e-20
C16 SCE VPWR 0.030224f
C17 VGND VPB 0.012547f
C18 SCE SCD 0.126583f
C19 CLK VPWR 0.01713f
C20 SCD CLK 0.003688f
C21 DE VPWR 0.024856f
C22 SCD VPWR 0.013215f
C23 VGND SCE 0.069415f
C24 Q VPWR 0.214153f
C25 VGND CLK 0.025559f
C26 Q VNB 0.054009f
C27 VGND VNB 1.96012f
C28 CLK VNB 0.137413f
C29 SCD VNB 0.110095f
C30 SCE VNB 0.358133f
C31 DE VNB 0.296334f
C32 VPWR VNB 1.43942f
C33 D VNB 0.188586f
C34 VPB VNB 3.73009f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xnor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor2_4 VNB VPB VPWR VGND Y B A
X0 a_116_368.t5 A.t0 VPWR.t4 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 a_950_368.t3 B.t0 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t3 B.t1 a_950_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t7 a_116_368.t6 a_511_74.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.16465 ps=1.185 w=0.74 l=0.15
X4 a_950_368.t1 B.t2 Y.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 Y.t2 B.t3 a_950_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_27_74.t1 B.t4 a_116_368.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.112 ps=0.99 w=0.64 l=0.15
X7 Y.t6 a_116_368.t7 a_511_74.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 a_950_368.t7 A.t1 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.297275 ps=1.825 w=1.12 l=0.15
X9 VGND.t4 A.t2 a_27_74.t2 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X10 VGND.t2 B.t5 a_511_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1889 pd=1.36 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t7 A.t3 a_950_368.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.30065 pd=1.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X12 VPWR.t6 A.t4 a_950_368.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.297275 pd=1.825 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_950_368.t4 A.t5 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.30065 ps=1.83 w=1.12 l=0.15
X14 a_511_74.t0 B.t6 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1889 ps=1.36 w=0.74 l=0.15
X15 a_116_368.t0 B.t7 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 VPWR.t2 B.t8 a_116_368.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.29145 pd=1.835 as=0.126 ps=1.14 w=0.84 l=0.15
X17 VGND.t7 A.t6 a_511_74.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1889 pd=1.36 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 a_511_74.t2 B.t9 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.205 ps=1.395 w=0.74 l=0.15
X19 a_116_368.t2 B.t10 VPWR.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X20 VPWR.t5 A.t7 a_116_368.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X21 a_511_74.t8 A.t8 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1889 ps=1.36 w=0.74 l=0.15
X22 VPWR.t1 a_116_368.t8 Y.t9 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.49375 pd=3.47 as=0.168 ps=1.42 w=1.12 l=0.15
X23 Y.t8 a_116_368.t9 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.29145 ps=1.835 w=1.12 l=0.15
X24 a_27_74.t3 A.t9 VGND.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
X25 a_511_74.t4 a_116_368.t10 Y.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 a_511_74.t3 a_116_368.t11 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.16465 pd=1.185 as=0.1295 ps=1.09 w=0.74 l=0.15
X27 a_511_74.t7 A.t10 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1889 ps=1.36 w=0.74 l=0.15
R0 A.n2 A.t1 279.024
R1 A.n5 A.t5 226.809
R2 A.n9 A.t3 226.809
R3 A.n2 A.t10 220.113
R4 A.n3 A.t4 214.758
R5 A.n12 A.t9 209.087
R6 A.n13 A.t2 203.901
R7 A.n10 A.t6 203.316
R8 A.n4 A.n1 196.013
R9 A.n7 A.t8 196.013
R10 A.n15 A.n14 193.34
R11 A.n12 A.t7 189.855
R12 A.n13 A.t0 189.855
R13 A.n6 A.n0 162.24
R14 A.n11 A.n10 152
R15 A.n8 A.n0 152
R16 A.n3 A.n2 57.0372
R17 A.n4 A.n3 53.0205
R18 A.n5 A.n4 39.9237
R19 A.n14 A.n12 35.7853
R20 A.n9 A.n8 30.6732
R21 A.n14 A.n13 29.9429
R22 A.n8 A.n7 29.2126
R23 A.n7 A.n6 20.449
R24 A.n10 A.n9 18.9884
R25 A.n15 A.n11 12.9511
R26 A.n6 A.n5 10.955
R27 A.n11 A.n0 10.2405
R28 A A.n15 2.5605
R29 VPWR.n4 VPWR.t1 936.455
R30 VPWR.n21 VPWR.n20 785.537
R31 VPWR.n10 VPWR.n9 652.628
R32 VPWR.n8 VPWR.n7 645.102
R33 VPWR.n27 VPWR.n1 641.471
R34 VPWR.n29 VPWR.t4 431.94
R35 VPWR.n20 VPWR.t2 66.8398
R36 VPWR.n7 VPWR.t9 42.2148
R37 VPWR.n9 VPWR.t8 41.3353
R38 VPWR.n9 VPWR.t6 41.3353
R39 VPWR.n7 VPWR.t7 41.3353
R40 VPWR.n26 VPWR.n2 36.1417
R41 VPWR.n13 VPWR.n6 36.1417
R42 VPWR.n14 VPWR.n13 36.1417
R43 VPWR.n15 VPWR.n14 36.1417
R44 VPWR.n1 VPWR.t3 35.1791
R45 VPWR.n1 VPWR.t5 35.1791
R46 VPWR.n28 VPWR.n27 34.6358
R47 VPWR.n20 VPWR.t0 34.5586
R48 VPWR.n19 VPWR.n18 34.2677
R49 VPWR.n22 VPWR.n2 28.6457
R50 VPWR.n21 VPWR.n19 27.4243
R51 VPWR.n29 VPWR.n28 26.7299
R52 VPWR.n8 VPWR.n6 21.635
R53 VPWR.n15 VPWR.n4 18.9997
R54 VPWR.n10 VPWR.n8 9.80424
R55 VPWR.n11 VPWR.n6 9.3005
R56 VPWR.n13 VPWR.n12 9.3005
R57 VPWR.n14 VPWR.n5 9.3005
R58 VPWR.n16 VPWR.n15 9.3005
R59 VPWR.n18 VPWR.n17 9.3005
R60 VPWR.n19 VPWR.n3 9.3005
R61 VPWR.n23 VPWR.n22 9.3005
R62 VPWR.n24 VPWR.n2 9.3005
R63 VPWR.n26 VPWR.n25 9.3005
R64 VPWR.n28 VPWR.n0 9.3005
R65 VPWR.n30 VPWR.n29 9.3005
R66 VPWR.n18 VPWR.n4 3.55606
R67 VPWR.n27 VPWR.n26 1.50638
R68 VPWR.n11 VPWR.n10 0.424093
R69 VPWR.n22 VPWR.n21 0.284944
R70 VPWR.n12 VPWR.n11 0.122949
R71 VPWR.n12 VPWR.n5 0.122949
R72 VPWR.n16 VPWR.n5 0.122949
R73 VPWR.n17 VPWR.n16 0.122949
R74 VPWR.n17 VPWR.n3 0.122949
R75 VPWR.n23 VPWR.n3 0.122949
R76 VPWR.n24 VPWR.n23 0.122949
R77 VPWR.n25 VPWR.n24 0.122949
R78 VPWR.n25 VPWR.n0 0.122949
R79 VPWR.n30 VPWR.n0 0.122949
R80 VPWR VPWR.n30 0.0617245
R81 a_116_368.n13 a_116_368.n11 530.303
R82 a_116_368.n14 a_116_368.n13 351.825
R83 a_116_368.n11 a_116_368.t10 321.041
R84 a_116_368.n13 a_116_368.n12 288.485
R85 a_116_368.n3 a_116_368.n2 255.571
R86 a_116_368.n4 a_116_368.t9 237.762
R87 a_116_368.n7 a_116_368.t8 226.809
R88 a_116_368.n11 a_116_368.t6 196.013
R89 a_116_368.n6 a_116_368.t7 196.013
R90 a_116_368.n0 a_116_368.t11 196.013
R91 a_116_368.n4 a_116_368.n3 152
R92 a_116_368.n5 a_116_368.n1 152
R93 a_116_368.n9 a_116_368.n8 152
R94 a_116_368.n10 a_116_368.n9 81.6328
R95 a_116_368.n5 a_116_368.n4 49.6611
R96 a_116_368.n10 a_116_368.n0 44.6774
R97 a_116_368.n8 a_116_368.n7 44.549
R98 a_116_368.n2 a_116_368.t0 39.3755
R99 a_116_368.n11 a_116_368.n10 35.5081
R100 a_116_368.n12 a_116_368.t1 35.1791
R101 a_116_368.n12 a_116_368.t2 35.1791
R102 a_116_368.n14 a_116_368.t4 35.1791
R103 a_116_368.t5 a_116_368.n14 35.1791
R104 a_116_368.n2 a_116_368.t3 26.2505
R105 a_116_368.n8 a_116_368.n0 25.5611
R106 a_116_368.n9 a_116_368.n1 13.1884
R107 a_116_368.n3 a_116_368.n1 13.1884
R108 a_116_368.n7 a_116_368.n6 2.92171
R109 a_116_368.n6 a_116_368.n5 2.19141
R110 VPB.t5 VPB.t11 1115.99
R111 VPB.t0 VPB.t4 321.774
R112 VPB.t11 VPB.t9 319.221
R113 VPB.t10 VPB.t12 316.668
R114 VPB VPB.t13 257.93
R115 VPB.t6 VPB.t3 229.839
R116 VPB.t7 VPB.t6 229.839
R117 VPB.t2 VPB.t7 229.839
R118 VPB.t12 VPB.t2 229.839
R119 VPB.t9 VPB.t10 229.839
R120 VPB.t4 VPB.t5 229.839
R121 VPB.t1 VPB.t0 229.839
R122 VPB.t8 VPB.t1 229.839
R123 VPB.t13 VPB.t8 229.839
R124 B.n12 B.n11 366.397
R125 B.n0 B.t0 295.091
R126 B.n6 B.n5 231.506
R127 B.n1 B.t1 226.809
R128 B.n4 B.t2 226.809
R129 B.n6 B.t3 226.809
R130 B.n0 B.t6 216.097
R131 B.n7 B.t7 212.081
R132 B.n10 B.t4 212.081
R133 B.n15 B.t9 196.013
R134 B.n2 B.t5 196.013
R135 B.n7 B.t10 184.743
R136 B.n9 B.t8 181.821
R137 B.n11 B.n8 165.189
R138 B.n11 B.n10 161.494
R139 B B.n3 156.781
R140 B.n14 B.n13 152
R141 B.n17 B.n16 152
R142 B.n1 B.n0 99.906
R143 B.n15 B.n14 43.0884
R144 B.n4 B.n3 40.1672
R145 B.n8 B.n7 32.8641
R146 B.n9 B.n8 29.9429
R147 B.n2 B.n1 18.9884
R148 B.n13 B 13.4174
R149 B B.n12 13.1089
R150 B.n10 B.n9 10.2247
R151 B.n16 B.n4 9.49444
R152 B.n17 B 9.09929
R153 B.n3 B.n2 6.57323
R154 B.n16 B.n15 6.57323
R155 B.n14 B.n6 6.57323
R156 B B.n17 5.70652
R157 B.n12 B 1.69689
R158 B.n13 B 1.38845
R159 Y.n7 Y.n5 937.707
R160 Y.n4 Y.n3 366.438
R161 Y.n4 Y.n0 300.091
R162 Y.n7 Y.n6 291.832
R163 Y.n3 Y.n1 250.055
R164 Y.n3 Y.n2 185
R165 Y.n8 Y.n4 42.9181
R166 Y.n1 Y.t6 34.0546
R167 Y.n6 Y.t0 26.3844
R168 Y.n6 Y.t2 26.3844
R169 Y.n5 Y.t9 26.3844
R170 Y.n5 Y.t8 26.3844
R171 Y.n0 Y.t1 26.3844
R172 Y.n0 Y.t3 26.3844
R173 Y.n2 Y.t5 22.7032
R174 Y.n2 Y.t7 22.7032
R175 Y.n1 Y.t4 22.7032
R176 Y.n8 Y.n7 8.26006
R177 Y Y.n8 2.71565
R178 a_950_368.n2 a_950_368.t6 920.111
R179 a_950_368.n2 a_950_368.n1 585
R180 a_950_368.n4 a_950_368.n3 585
R181 a_950_368.n5 a_950_368.n0 306.171
R182 a_950_368.t3 a_950_368.n5 301.632
R183 a_950_368.n5 a_950_368.n4 71.0932
R184 a_950_368.n4 a_950_368.n2 66.2754
R185 a_950_368.n3 a_950_368.t0 26.3844
R186 a_950_368.n3 a_950_368.t7 26.3844
R187 a_950_368.n1 a_950_368.t5 26.3844
R188 a_950_368.n1 a_950_368.t4 26.3844
R189 a_950_368.n0 a_950_368.t2 26.3844
R190 a_950_368.n0 a_950_368.t1 26.3844
R191 a_511_74.n6 a_511_74.t5 310.002
R192 a_511_74.n3 a_511_74.t8 247.143
R193 a_511_74.n2 a_511_74.t7 247.143
R194 a_511_74.n1 a_511_74.t0 200.496
R195 a_511_74.n1 a_511_74.n0 185
R196 a_511_74.n5 a_511_74.n4 185
R197 a_511_74.n7 a_511_74.n6 185
R198 a_511_74.n6 a_511_74.n5 65.8311
R199 a_511_74.n2 a_511_74.n1 63.2091
R200 a_511_74.n5 a_511_74.n3 62.4697
R201 a_511_74.n3 a_511_74.n2 60.5738
R202 a_511_74.t6 a_511_74.n7 38.1086
R203 a_511_74.n4 a_511_74.t4 34.0546
R204 a_511_74.n7 a_511_74.t3 34.0546
R205 a_511_74.n4 a_511_74.t9 22.7032
R206 a_511_74.n0 a_511_74.t1 22.7032
R207 a_511_74.n0 a_511_74.t2 22.7032
R208 VNB.t9 VNB.t0 2436.75
R209 VNB.t11 VNB.t9 2355.91
R210 VNB.t4 VNB.t7 2286.61
R211 VNB.t5 VNB.t8 1374.28
R212 VNB.t3 VNB.t2 1362.73
R213 VNB.t12 VNB.t11 1362.73
R214 VNB.t6 VNB.t12 1154.86
R215 VNB.t7 VNB.t5 1154.86
R216 VNB.t1 VNB.t4 1154.86
R217 VNB.t13 VNB.t10 1154.86
R218 VNB VNB.t13 1143.31
R219 VNB.t0 VNB.t3 993.177
R220 VNB.t8 VNB.t6 993.177
R221 VNB.t10 VNB.t1 993.177
R222 a_27_74.t1 a_27_74.n1 305.952
R223 a_27_74.n1 a_27_74.t2 209.419
R224 a_27_74.n1 a_27_74.n0 89.2272
R225 a_27_74.n0 a_27_74.t0 26.2505
R226 a_27_74.n0 a_27_74.t3 26.2505
R227 VGND.n11 VGND.t5 313.387
R228 VGND.n9 VGND.t0 291.397
R229 VGND.n8 VGND.n7 218.093
R230 VGND.n18 VGND.n17 212.477
R231 VGND.n33 VGND.n32 207.498
R232 VGND.n32 VGND.t3 39.3755
R233 VGND.n12 VGND.n10 36.1417
R234 VGND.n16 VGND.n5 36.1417
R235 VGND.n20 VGND.n19 36.1417
R236 VGND.n20 VGND.n3 36.1417
R237 VGND.n24 VGND.n3 36.1417
R238 VGND.n25 VGND.n24 36.1417
R239 VGND.n26 VGND.n25 36.1417
R240 VGND.n26 VGND.n1 36.1417
R241 VGND.n30 VGND.n1 36.1417
R242 VGND.n31 VGND.n30 36.1417
R243 VGND.n7 VGND.t1 35.6762
R244 VGND.n7 VGND.t2 35.6762
R245 VGND.n17 VGND.t6 35.6762
R246 VGND.n17 VGND.t7 35.6762
R247 VGND.n32 VGND.t4 26.2505
R248 VGND.n33 VGND.n31 24.4711
R249 VGND.n10 VGND.n9 15.2331
R250 VGND.n9 VGND.n8 10.4812
R251 VGND.n10 VGND.n6 9.3005
R252 VGND.n13 VGND.n12 9.3005
R253 VGND.n14 VGND.n5 9.3005
R254 VGND.n16 VGND.n15 9.3005
R255 VGND.n19 VGND.n4 9.3005
R256 VGND.n21 VGND.n20 9.3005
R257 VGND.n22 VGND.n3 9.3005
R258 VGND.n24 VGND.n23 9.3005
R259 VGND.n25 VGND.n2 9.3005
R260 VGND.n27 VGND.n26 9.3005
R261 VGND.n28 VGND.n1 9.3005
R262 VGND.n30 VGND.n29 9.3005
R263 VGND.n31 VGND.n0 9.3005
R264 VGND.n18 VGND.n16 9.03579
R265 VGND.n34 VGND.n33 7.19894
R266 VGND.n11 VGND.n5 6.77697
R267 VGND.n12 VGND.n11 4.51815
R268 VGND.n19 VGND.n18 2.25932
R269 VGND.n8 VGND.n6 0.514322
R270 VGND VGND.n34 0.156997
R271 VGND.n34 VGND.n0 0.150766
R272 VGND.n13 VGND.n6 0.122949
R273 VGND.n14 VGND.n13 0.122949
R274 VGND.n15 VGND.n14 0.122949
R275 VGND.n15 VGND.n4 0.122949
R276 VGND.n21 VGND.n4 0.122949
R277 VGND.n22 VGND.n21 0.122949
R278 VGND.n23 VGND.n22 0.122949
R279 VGND.n23 VGND.n2 0.122949
R280 VGND.n27 VGND.n2 0.122949
R281 VGND.n28 VGND.n27 0.122949
R282 VGND.n29 VGND.n28 0.122949
R283 VGND.n29 VGND.n0 0.122949
C0 B VGND 0.064816f
C1 VPWR A 0.182592f
C2 VPWR VPB 0.260777f
C3 VPWR VGND 0.090347f
C4 B VPWR 0.090532f
C5 Y A 0.218993f
C6 Y VPB 0.028178f
C7 Y VGND 0.055833f
C8 B Y 0.771074f
C9 A VPB 0.268659f
C10 A VGND 0.1773f
C11 VGND VPB 0.008713f
C12 Y VPWR 0.085056f
C13 B A 0.431882f
C14 B VPB 0.251116f
C15 VGND VNB 1.02929f
C16 Y VNB 0.060315f
C17 B VNB 0.7033f
C18 A VNB 0.733779f
C19 VPWR VNB 0.85745f
C20 VPB VNB 2.1204f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xnor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor2_2 VNB VPB VPWR VGND Y B A
X0 VGND.t1 B.t0 a_340_107.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1958 pd=1.375 as=0.111 ps=1.04 w=0.74 l=0.15
X1 a_340_107.t4 A.t0 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.20355 pd=2.05 as=0.1958 ps=1.375 w=0.74 l=0.15
X2 VPWR.t5 a_133_368.t3 Y.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.27625 pd=1.68 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t4 a_133_368.t4 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.451225 ps=1.94 w=1.12 l=0.15
X4 VPWR.t1 A.t1 a_638_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X5 a_638_368.t0 A.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2823 pd=1.69 as=0.27625 ps=1.68 w=1.12 l=0.15
X6 Y.t3 a_133_368.t5 a_340_107.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2004 pd=1.335 as=0.197775 ps=2.05 w=0.74 l=0.15
X7 VGND.t3 A.t3 a_340_107.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1912 pd=1.365 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t3 B.t1 a_133_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.451225 pd=1.94 as=0.1725 ps=1.345 w=1 l=0.15
X9 a_340_107.t2 B.t2 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1912 ps=1.365 w=0.74 l=0.15
X10 a_638_368.t3 B.t3 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t0 B.t4 a_638_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2823 ps=1.69 w=1.12 l=0.15
X12 a_340_107.t1 a_133_368.t6 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2004 ps=1.335 w=0.74 l=0.15
X13 a_133_368.t1 B.t5 a_151_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.206875 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X14 a_151_74.t0 A.t4 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.25 ps=2.44 w=0.74 l=0.15
X15 a_133_368.t0 A.t5 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.4177 ps=3.02 w=1 l=0.15
R0 B B.n3 631.856
R1 B.n0 B.t3 261.62
R2 B.n1 B.t4 261.62
R3 B.n3 B.t1 207.529
R4 B.n3 B.t5 198.204
R5 B B.n2 158.788
R6 B.n1 B.t2 156.431
R7 B.n0 B.t0 154.24
R8 B.n2 B.n1 50.3914
R9 B.n2 B.n0 13.146
R10 a_340_107.n1 a_340_107.t4 275.735
R11 a_340_107.n4 a_340_107.n3 254.647
R12 a_340_107.n1 a_340_107.n0 185
R13 a_340_107.n3 a_340_107.n2 95.7792
R14 a_340_107.n3 a_340_107.n1 58.3642
R15 a_340_107.n5 a_340_107.n4 40.8005
R16 a_340_107.n0 a_340_107.t3 25.9464
R17 a_340_107.n0 a_340_107.t2 22.7032
R18 a_340_107.n2 a_340_107.t5 22.7032
R19 a_340_107.n2 a_340_107.t1 22.7032
R20 a_340_107.n4 a_340_107.t0 21.0457
R21 VGND.n16 VGND.t4 286.567
R22 VGND.n6 VGND.n5 205.578
R23 VGND.n4 VGND.n3 199.238
R24 VGND.n5 VGND.t2 37.2978
R25 VGND.n3 VGND.t0 36.487
R26 VGND.n5 VGND.t1 36.487
R27 VGND.n9 VGND.n8 36.1417
R28 VGND.n10 VGND.n9 36.1417
R29 VGND.n10 VGND.n1 36.1417
R30 VGND.n14 VGND.n1 36.1417
R31 VGND.n15 VGND.n14 36.1417
R32 VGND.n3 VGND.t3 35.6762
R33 VGND.n16 VGND.n15 16.9417
R34 VGND.n8 VGND.n4 14.5284
R35 VGND.n6 VGND.n4 10.968
R36 VGND.n17 VGND.n16 9.3005
R37 VGND.n8 VGND.n7 9.3005
R38 VGND.n9 VGND.n2 9.3005
R39 VGND.n11 VGND.n10 9.3005
R40 VGND.n12 VGND.n1 9.3005
R41 VGND.n14 VGND.n13 9.3005
R42 VGND.n15 VGND.n0 9.3005
R43 VGND.n7 VGND.n6 0.534576
R44 VGND.n7 VGND.n2 0.122949
R45 VGND.n11 VGND.n2 0.122949
R46 VGND.n12 VGND.n11 0.122949
R47 VGND.n13 VGND.n12 0.122949
R48 VGND.n13 VGND.n0 0.122949
R49 VGND.n17 VGND.n0 0.122949
R50 VGND VGND.n17 0.0617245
R51 VNB.t2 VNB.t0 2286.61
R52 VNB VNB.t7 1570.6
R53 VNB.t0 VNB.t1 1489.76
R54 VNB.t4 VNB.t5 1397.38
R55 VNB.t6 VNB.t3 1374.28
R56 VNB.t3 VNB.t4 1039.37
R57 VNB.t1 VNB.t6 993.177
R58 VNB.t7 VNB.t2 900.788
R59 A.n1 A.t2 285.719
R60 A.n0 A.t5 266.44
R61 A.n3 A.t1 250.548
R62 A.n3 A.t0 219.755
R63 A.n2 A.n0 180.43
R64 A.n1 A.t3 178.34
R65 A.n0 A.t4 178.34
R66 A.n4 A.n3 157.042
R67 A.n2 A.n1 152
R68 A.n4 A.n2 104.953
R69 A A.n4 5.56572
R70 A.n4 A 3.29747
R71 a_133_368.n4 a_133_368.n3 645.524
R72 a_133_368.n1 a_133_368.t4 263.81
R73 a_133_368.n0 a_133_368.t3 261.62
R74 a_133_368.n3 a_133_368.t1 216.431
R75 a_133_368.n0 a_133_368.t6 205.946
R76 a_133_368.n1 a_133_368.t5 154.24
R77 a_133_368.n3 a_133_368.n2 106.183
R78 a_133_368.n4 a_133_368.t2 34.4755
R79 a_133_368.t0 a_133_368.n4 33.4905
R80 a_133_368.n2 a_133_368.n0 32.9301
R81 a_133_368.n2 a_133_368.n1 23.7903
R82 Y.n4 Y.n1 694.457
R83 Y.n3 Y.n2 618.081
R84 Y Y.n0 590.745
R85 Y Y.n0 589.432
R86 Y.n4 Y.n0 585
R87 Y.n2 Y.t2 40.541
R88 Y.n2 Y.t3 39.7302
R89 Y.n0 Y.t5 26.3844
R90 Y.n0 Y.t4 26.3844
R91 Y.n1 Y.t1 26.3844
R92 Y.n1 Y.t0 26.3844
R93 Y Y.n4 6.72871
R94 Y.n3 Y 2.79024
R95 Y.n4 Y.n3 2.62614
R96 VPWR.n15 VPWR.t2 856.023
R97 VPWR.n5 VPWR.n4 601.486
R98 VPWR.n9 VPWR.n8 591.573
R99 VPWR.n7 VPWR.n1 585
R100 VPWR.n3 VPWR.t1 357.878
R101 VPWR.n8 VPWR.n7 68.6106
R102 VPWR.n7 VPWR.t3 42.3555
R103 VPWR.n4 VPWR.t0 41.3353
R104 VPWR.n4 VPWR.t5 41.3353
R105 VPWR.n14 VPWR.n13 36.1417
R106 VPWR.n6 VPWR.n5 36.1417
R107 VPWR.n9 VPWR.n6 22.9004
R108 VPWR.n8 VPWR.t4 22.3156
R109 VPWR.n15 VPWR.n14 20.7064
R110 VPWR.n6 VPWR.n2 9.3005
R111 VPWR.n11 VPWR.n10 9.3005
R112 VPWR.n13 VPWR.n12 9.3005
R113 VPWR.n14 VPWR.n0 9.3005
R114 VPWR.n16 VPWR.n15 9.3005
R115 VPWR.n5 VPWR.n3 6.2019
R116 VPWR.n10 VPWR.n1 5.17136
R117 VPWR.n13 VPWR.n1 4.7176
R118 VPWR.n10 VPWR.n9 1.8654
R119 VPWR.n3 VPWR.n2 0.176375
R120 VPWR.n11 VPWR.n2 0.122949
R121 VPWR.n12 VPWR.n11 0.122949
R122 VPWR.n12 VPWR.n0 0.122949
R123 VPWR.n16 VPWR.n0 0.122949
R124 VPWR VPWR.n16 0.0617245
R125 VPB.t5 VPB.t6 490.324
R126 VPB.t1 VPB.t3 321.774
R127 VPB.t7 VPB.t1 316.668
R128 VPB VPB.t0 301.344
R129 VPB.t4 VPB.t2 255.376
R130 VPB.t0 VPB.t5 252.823
R131 VPB.t3 VPB.t4 229.839
R132 VPB.t6 VPB.t7 229.839
R133 a_638_368.n1 a_638_368.n0 946.74
R134 a_638_368.n0 a_638_368.t2 42.2148
R135 a_638_368.n0 a_638_368.t0 42.2148
R136 a_638_368.n1 a_638_368.t3 35.1791
R137 a_638_368.t1 a_638_368.n1 26.3844
R138 a_151_74.t0 a_151_74.t1 38.9194
C0 Y VPB 0.020106f
C1 Y A 0.144761f
C2 A VPB 0.118077f
C3 Y VGND 0.296934f
C4 B Y 0.255241f
C5 VPB VGND 0.004518f
C6 B VPB 0.132105f
C7 B A 0.542907f
C8 Y VPWR 0.333466f
C9 A VGND 0.130403f
C10 VPWR VPB 0.146428f
C11 VPWR A 0.115726f
C12 B VGND 0.041313f
C13 VPWR VGND 0.044519f
C14 B VPWR 0.103643f
C15 VGND VNB 0.647649f
C16 Y VNB 0.106875f
C17 B VNB 0.408088f
C18 A VNB 0.419458f
C19 VPWR VNB 0.534116f
C20 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xnor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor2_1 VNB VPB VPWR VGND A Y B
X0 a_138_385.t1 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2898 ps=2.37 w=0.84 l=0.15
X1 a_138_385.t0 B.t0 a_112_119.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.176 pd=1.83 as=0.0672 ps=0.85 w=0.64 l=0.15
X2 VGND.t1 A.t1 a_293_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.182 pd=1.345 as=0.2035 ps=2.03 w=0.74 l=0.15
X3 a_293_74.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.182 ps=1.345 w=0.74 l=0.15
X4 Y.t0 B.t2 a_376_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X5 a_376_368.t1 A.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.287825 ps=1.71 w=1.12 l=0.15
X6 VPWR.t3 B.t3 a_138_385.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.287825 pd=1.71 as=0.126 ps=1.14 w=0.84 l=0.15
X7 VPWR.t0 a_138_385.t3 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X8 Y.t1 a_138_385.t4 a_293_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2294 pd=2.1 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_112_119.t1 A.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.176 ps=1.83 w=0.64 l=0.15
R0 A.t1 A.t3 795.301
R1 A.t3 A.t0 435.815
R2 A.n0 A.t2 247.738
R3 A.n0 A.t1 216.942
R4 A A.n0 154.53
R5 VPWR.n7 VPWR.t2 375.342
R6 VPWR.n3 VPWR.t0 350.644
R7 VPWR.n2 VPWR.n1 324.637
R8 VPWR.n1 VPWR.t3 103.191
R9 VPWR.n6 VPWR.n5 36.1417
R10 VPWR.n1 VPWR.t1 28.734
R11 VPWR.n5 VPWR.n2 16.1887
R12 VPWR.n7 VPWR.n6 16.1887
R13 VPWR.n5 VPWR.n4 9.3005
R14 VPWR.n6 VPWR.n0 9.3005
R15 VPWR.n8 VPWR.n7 9.3005
R16 VPWR.n3 VPWR.n2 7.39741
R17 VPWR.n4 VPWR.n3 0.237078
R18 VPWR.n4 VPWR.n0 0.122949
R19 VPWR.n8 VPWR.n0 0.122949
R20 VPWR VPWR.n8 0.0617245
R21 a_138_385.n2 a_138_385.n1 373.262
R22 a_138_385.n1 a_138_385.n0 280.64
R23 a_138_385.n0 a_138_385.t3 264.298
R24 a_138_385.n0 a_138_385.t4 204.048
R25 a_138_385.n1 a_138_385.t0 134.185
R26 a_138_385.n2 a_138_385.t2 35.1791
R27 a_138_385.t1 a_138_385.n2 35.1791
R28 VPB.t4 VPB.t1 377.957
R29 VPB VPB.t2 314.113
R30 VPB.t3 VPB.t0 291.13
R31 VPB.t2 VPB.t4 229.839
R32 VPB.t1 VPB.t3 214.517
R33 B.n2 B.n0 261.894
R34 B.n0 B.t2 250.909
R35 B.n0 B.t1 220.113
R36 B.n1 B.t3 205.922
R37 B.n1 B.t0 190.464
R38 B.n2 B.n1 152
R39 B B.n2 0.6405
R40 a_112_119.t0 a_112_119.t1 39.3755
R41 VNB.t1 VNB.t4 2240.42
R42 VNB.t4 VNB.t0 1328.08
R43 VNB VNB.t3 1120.21
R44 VNB.t0 VNB.t2 993.177
R45 VNB.t3 VNB.t1 831.496
R46 a_293_74.n0 a_293_74.t2 456.327
R47 a_293_74.n0 a_293_74.t1 22.7032
R48 a_293_74.t0 a_293_74.n0 22.7032
R49 VGND.n1 VGND.n0 205.534
R50 VGND.n1 VGND.t2 169.702
R51 VGND.n0 VGND.t0 34.8654
R52 VGND.n0 VGND.t1 34.0546
R53 VGND VGND.n1 0.112484
R54 a_376_368.t0 a_376_368.t1 47.4916
R55 Y.n1 Y.n0 585
R56 Y Y.n0 296.387
R57 Y.n1 Y.t1 243.065
R58 Y.n0 Y.t0 38.6969
R59 Y.n0 Y.t2 35.1791
R60 Y Y.n1 11.2672
C0 VPB A 0.081856f
C1 B A 0.267566f
C2 VPWR VPB 0.127789f
C3 Y A 0.005772f
C4 VGND VPB 0.010821f
C5 B VPWR 0.078694f
C6 VPWR Y 0.216144f
C7 B VGND 0.023037f
C8 Y VGND 0.042936f
C9 Y VPB 0.014546f
C10 B VPB 0.093824f
C11 B Y 0.077205f
C12 VGND A 0.076551f
C13 VPWR A 0.039376f
C14 VPWR VGND 0.067723f
C15 VGND VNB 0.474927f
C16 Y VNB 0.08802f
C17 VPWR VNB 0.414375f
C18 B VNB 0.21418f
C19 A VNB 0.401644f
C20 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__tapvpwrvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tapvpwrvgnd_1 VPWR VGND
C0 VPWR VGND 0.378723f
.ends

* NGSPICE file created from sky130_fd_sc_hs__tapvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tapvgnd_1 VPB VPWR VGND
C0 VPB VPWR 0.08054f
C1 VPWR VGND 0.0962f
C2 VPB VGND 0.317545f
.ends

* NGSPICE file created from sky130_fd_sc_hs__tapvgnd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tapvgnd2_1 VPB VPWR VGND
C0 VPB VPWR 0.0712f
C1 VPWR VGND 0.0962f
C2 VPB VGND 0.319242f
.ends

* NGSPICE file created from sky130_fd_sc_hs__tapmet1_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tapmet1_2 VNB VPB VPWR VGND
C0 VPWR VGND 0.006005f
C1 VPB VPWR 0.152242f
C2 VPB VGND 0.011046f
C3 VGND VNB 0.28126f
C4 VPWR VNB 0.140162f
C5 VPB VNB 0.403384f
.ends

* NGSPICE file created from sky130_fd_sc_hs__tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tap_2 VNB VPB VPWR VGND
R0 VPB.n3 VPB.n2 337.661
R1 VPB.n4 VPB.n0 185
R2 VPB.n4 VPB.n3 185
R3 VPB.n2 VPB 122.582
R4 VPB.n2 VPB.n0 92.5005
R5 VPB.n1 VPB 79.9256
R6 VPB.n1 VPB.n0 28.9261
R7 VPB.n3 VPB.n1 28.9261
R8 VPB.n4 VPB 5.16973
R9 VPB VPB.n4 0.903064
R10 VNB.n2 VNB 1826.2
R11 VNB.n3 VNB.n1 585
R12 VNB.n1 VNB.n0 585
R13 VNB.n2 VNB.n0 292.502
R14 VNB.n3 VNB.n2 292.5
R15 VNB.n5 VNB.n4 266.404
R16 VNB.n4 VNB.n3 52.1968
R17 VNB.n4 VNB.n0 52.1968
R18 VNB.n1 VNB 5.16973
R19 VNB VNB.n5 4.43127
R20 VNB.n5 VNB 1.64153
R21 VNB.n1 VNB 0.903064
C0 VPWR VGND 0.015118f
C1 VPB VGND 0.007684f
C2 VPB VPWR 0.130375f
C3 VGND VNB 0.259442f
C4 VPWR VNB 0.13675f
C5 VPB VNB 0.422331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__tap_1 VNB VPB VPWR VGND
R0 VPB.n0 VPB 555.936
R1 VPB VPB.n0 10.2452
R2 VPB.n0 VPB 5.2481
R3 VNB.n1 VNB 3105.83
R4 VNB.n1 VNB.n0 930.092
R5 VNB.n2 VNB.n1 659.543
R6 VNB.n2 VNB 13.4405
R7 VNB.n0 VNB 11.5205
R8 VNB.n0 VNB 4.26717
R9 VNB VNB.n2 2.34717
C0 VPB VGND 0.004807f
C1 VPB VPWR 0.058009f
C2 VPWR VGND 0.008283f
C3 VGND VNB 0.14762f
C4 VPWR VNB 0.094419f
C5 VPB VNB 0.290558f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sedfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sedfxtp_4 VNB VPB VPWR VGND SCE CLK D DE SCD Q
X0 a_2586_508.t1 a_1510_74# a_2403_74.t2 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.15245 ps=1.36 w=0.42 l=0.15
X1 a_545_87.t1 a_2403_74.t4 VGND.t8 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.21 ps=1.42 w=0.42 l=0.15
X2 Q.t3 a_2403_74.t5 VGND.t10 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 a_545_87.t0 a_2403_74.t6 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.83 as=0.14675 ps=1.2 w=0.64 l=0.15
X4 VGND.t11 a_1943_53.t2 a_1858_79.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1388 pd=1.17 as=0.08925 ps=0.845 w=0.42 l=0.15
X5 a_126_464.t1 D.t0 a_37_464.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1888 ps=1.87 w=0.64 l=0.15
X6 a_1313_74.t0 CLK.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.3136 ps=2.8 w=1.12 l=0.15
X7 Q.t6 a_2403_74.t7 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X8 a_1044_125.t0 SCD.t0 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 a_2403_74.t3 a_1510_74# a_2331_74.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.09575 pd=0.965 as=0.0672 ps=0.85 w=0.64 l=0.15
X10 a_661_113.t3 SCE.t0 a_37_464.t3 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.83 as=0.096 ps=0.94 w=0.64 l=0.15
X11 a_135_74.t1 D.t1 a_37_464.t4 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X12 Q.t2 a_2403_74.t8 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 VGND.t7 a_2403_74.t9 Q.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_37_464.t1 a_545_87.t2 a_572_463.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0768 ps=0.88 w=0.64 l=0.15
X15 a_1943_53.t0 a_1756_97.t3 VGND.t13 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1388 ps=1.17 w=0.64 l=0.15
X16 VGND.t4 DE.t0 a_177_290.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X17 a_572_463.t0 DE.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1696 ps=1.17 w=0.64 l=0.15
X18 a_1510_74# a_1313_74.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.2109 ps=2.05 w=0.74 l=0.15
X19 a_1943_53.t1 a_1756_97.t4 VPWR.t11 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.231 pd=2.23 as=0.143675 ps=1.335 w=0.84 l=0.15
X20 VPWR.t4 DE.t2 a_177_290.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X21 a_2498_74.t0 a_1313_74.t3 a_2403_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.09575 ps=0.965 w=0.42 l=0.15
X22 a_37_464.t2 a_545_87.t3 a_497_113.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 VPWR.t9 a_177_290.t2 a_126_464.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1756_97.t0 a_1510_74# a_661_113.t4 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1155 ps=1.39 w=0.42 l=0.15
X25 a_661_113.t2 SCE.t1 a_1044_125.t1 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 VPWR.t6 a_2403_74.t10 Q.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X27 a_497_113.t1 a_177_290.t3 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 a_2292_392.t0 a_1943_53.t3 VPWR.t10 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.405 pd=1.81 as=0.275 ps=2.55 w=1 l=0.15
X29 Q.t4 a_2403_74.t11 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_661_113.t0 a_631_87.t2 a_1071_455.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.84 as=0.0768 ps=0.88 w=0.64 l=0.15
X31 VGND.t2 DE.t3 a_135_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X32 a_2403_74.t1 a_1313_74.t4 a_2292_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15245 pd=1.36 as=0.405 ps=1.81 w=1 l=0.15
X33 a_1858_79.t1 a_1510_74# a_1756_97.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.08925 pd=0.845 as=0.083475 ps=0.87 w=0.42 l=0.15
X34 VPWR.t12 SCE.t2 a_631_87.t0 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.1696 pd=1.17 as=0.1792 ps=1.84 w=0.64 l=0.15
X35 a_661_113.t1 a_631_87.t3 a_37_464.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.21 pd=1.84 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 VGND.t14 SCE.t3 a_631_87.t1 VNB.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X37 a_1756_97.t2 a_1313_74.t5 a_661_113.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.083475 pd=0.87 as=0.2226 ps=1.9 w=0.42 l=0.15
X38 VGND.t6 a_2403_74.t12 Q.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.10915 ps=1.035 w=0.74 l=0.15
X39 a_1071_455.t0 SCD.t1 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.1696 ps=1.17 w=0.64 l=0.15
X40 a_1313_74.t1 CLK.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.2109 ps=2.05 w=0.74 l=0.15
X41 VPWR.t2 a_545_87.t4 a_2586_508.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.14675 pd=1.2 as=0.0567 ps=0.69 w=0.42 l=0.15
X42 a_2331_74.t0 a_1943_53.t4 VGND.t12 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1824 ps=1.85 w=0.64 l=0.15
R0 a_2403_74.n13 a_2403_74.n0 672.806
R1 a_2403_74.n0 a_2403_74.n12 305.688
R2 a_2403_74.n3 a_2403_74.t10 226.809
R3 a_2403_74.n5 a_2403_74.t11 226.809
R4 a_2403_74.n6 a_2403_74.n2 226.809
R5 a_2403_74.n8 a_2403_74.t7 226.809
R6 a_2403_74.n10 a_2403_74.t6 217.934
R7 a_2403_74.n10 a_2403_74.n0 159.019
R8 a_2403_74.n0 a_2403_74.n1 67.5585
R9 a_2403_74.n11 a_2403_74.n9 147.137
R10 a_2403_74.n3 a_2403_74.t12 145.53
R11 a_2403_74.n9 a_2403_74.t8 142.994
R12 a_2403_74.n7 a_2403_74.t9 142.994
R13 a_2403_74.n4 a_2403_74.t5 142.994
R14 a_2403_74.n6 a_2403_74.n5 76.1058
R15 a_2403_74.n4 a_2403_74.n3 72.7233
R16 a_2403_74.n8 a_2403_74.n7 71.0321
R17 a_2403_74.n13 a_2403_74.t2 70.3576
R18 a_2403_74.t1 a_2403_74.n13 63.1343
R19 a_2403_74.t4 a_2403_74.n1 171.983
R20 a_2403_74.n12 a_2403_74.t3 40.5809
R21 a_2403_74.n12 a_2403_74.t0 40.0005
R22 a_2403_74.n11 a_2403_74.n10 39.9376
R23 a_2403_74.n1 a_2403_74.n11 26.8566
R24 a_2403_74.n7 a_2403_74.n6 5.07418
R25 a_2403_74.n5 a_2403_74.n4 3.38296
R26 a_2403_74.n9 a_2403_74.n8 1.69173
R27 a_2586_508.t0 a_2586_508.t1 126.644
R28 VPB.t3 VPB.t14 1184.95
R29 VPB.t14 VPB.t17 738.038
R30 VPB.t13 VPB.t7 577.152
R31 VPB.t2 VPB.t3 500.538
R32 VPB.t18 VPB.t19 497.985
R33 VPB.t11 VPB.t10 495.43
R34 VPB.t17 VPB.t16 495.43
R35 VPB.t16 VPB.t4 490.324
R36 VPB.t10 VPB.t8 459.678
R37 VPB.t5 VPB.t11 362.635
R38 VPB.t19 VPB.t6 347.312
R39 VPB.t7 VPB.t0 347.312
R40 VPB VPB.t1 283.469
R41 VPB.t4 VPB.t15 260.485
R42 VPB.t8 VPB.t9 229.839
R43 VPB.t12 VPB.t18 229.839
R44 VPB.t15 VPB.t5 214.517
R45 VPB.t1 VPB.t13 214.517
R46 VPB.t6 VPB.t2 199.195
R47 VPB.t0 VPB.t12 199.195
R48 a_545_87.n1 a_545_87.n0 642.668
R49 a_545_87.t0 a_545_87.n4 365.67
R50 a_545_87.n3 a_545_87.t1 288.267
R51 a_545_87.n2 a_545_87.t2 272.988
R52 a_545_87.n2 a_545_87.t3 252.54
R53 a_545_87.n3 a_545_87.n2 209.275
R54 a_545_87.n4 a_545_87.n1 202.447
R55 a_545_87.n1 a_545_87.t4 138.441
R56 a_545_87.n4 a_545_87.n3 33.2267
R57 VGND.n30 VGND.n29 370.714
R58 VGND.n18 VGND.t6 313.656
R59 VGND.n49 VGND.t1 286.334
R60 VGND.n36 VGND.t12 283.204
R61 VGND.n69 VGND.t2 247.498
R62 VGND.n6 VGND.t0 239.447
R63 VGND.n57 VGND.n56 216.225
R64 VGND.n67 VGND.n2 215.061
R65 VGND.n20 VGND.n19 213.703
R66 VGND.n11 VGND.n10 211.881
R67 VGND.n29 VGND.n28 185
R68 VGND.n22 VGND.t9 172.222
R69 VGND.n10 VGND.t13 99.1523
R70 VGND.n29 VGND.t8 60.0005
R71 VGND.n10 VGND.t11 40.0005
R72 VGND.n56 VGND.t5 40.0005
R73 VGND.n56 VGND.t14 40.0005
R74 VGND.n2 VGND.t3 40.0005
R75 VGND.n2 VGND.t4 40.0005
R76 VGND.n32 VGND.n31 36.1417
R77 VGND.n32 VGND.n13 36.1417
R78 VGND.n37 VGND.n36 36.1417
R79 VGND.n38 VGND.n37 36.1417
R80 VGND.n42 VGND.n11 36.1417
R81 VGND.n43 VGND.n42 36.1417
R82 VGND.n44 VGND.n43 36.1417
R83 VGND.n44 VGND.n8 36.1417
R84 VGND.n48 VGND.n8 36.1417
R85 VGND.n51 VGND.n50 36.1417
R86 VGND.n55 VGND.n54 36.1417
R87 VGND.n61 VGND.n4 36.1417
R88 VGND.n62 VGND.n61 36.1417
R89 VGND.n63 VGND.n62 36.1417
R90 VGND.n63 VGND.n1 36.1417
R91 VGND.n19 VGND.t7 34.0546
R92 VGND.n57 VGND.n55 32.0005
R93 VGND.n22 VGND.n16 30.4946
R94 VGND.n21 VGND.n20 28.2358
R95 VGND.n27 VGND.n16 27.0646
R96 VGND.n68 VGND.n67 26.3534
R97 VGND.n69 VGND.n68 23.3417
R98 VGND.n19 VGND.t10 22.7032
R99 VGND.n67 VGND.n1 21.0829
R100 VGND.n36 VGND.n13 17.3181
R101 VGND.n38 VGND.n11 17.3181
R102 VGND.n22 VGND.n21 16.9417
R103 VGND.n57 VGND.n4 15.4358
R104 VGND.n31 VGND.n30 12.926
R105 VGND.n50 VGND.n49 10.1652
R106 VGND.n68 VGND.n0 9.3005
R107 VGND.n67 VGND.n66 9.3005
R108 VGND.n65 VGND.n1 9.3005
R109 VGND.n64 VGND.n63 9.3005
R110 VGND.n62 VGND.n3 9.3005
R111 VGND.n61 VGND.n60 9.3005
R112 VGND.n59 VGND.n4 9.3005
R113 VGND.n58 VGND.n57 9.3005
R114 VGND.n55 VGND.n5 9.3005
R115 VGND.n54 VGND.n53 9.3005
R116 VGND.n52 VGND.n51 9.3005
R117 VGND.n50 VGND.n7 9.3005
R118 VGND.n48 VGND.n47 9.3005
R119 VGND.n46 VGND.n8 9.3005
R120 VGND.n45 VGND.n44 9.3005
R121 VGND.n43 VGND.n9 9.3005
R122 VGND.n42 VGND.n41 9.3005
R123 VGND.n40 VGND.n11 9.3005
R124 VGND.n39 VGND.n38 9.3005
R125 VGND.n37 VGND.n12 9.3005
R126 VGND.n36 VGND.n35 9.3005
R127 VGND.n34 VGND.n13 9.3005
R128 VGND.n33 VGND.n32 9.3005
R129 VGND.n31 VGND.n14 9.3005
R130 VGND.n25 VGND.n15 9.3005
R131 VGND.n27 VGND.n26 9.3005
R132 VGND.n24 VGND.n16 9.3005
R133 VGND.n23 VGND.n22 9.3005
R134 VGND.n21 VGND.n17 9.3005
R135 VGND.n51 VGND.n6 9.03579
R136 VGND.n54 VGND.n6 8.28285
R137 VGND.n28 VGND.n15 7.86455
R138 VGND.n70 VGND.n69 7.17141
R139 VGND.n20 VGND.n18 6.29111
R140 VGND.n30 VGND.n15 3.01226
R141 VGND.n49 VGND.n48 1.12991
R142 VGND.n18 VGND.n17 0.71681
R143 VGND VGND.n70 0.274942
R144 VGND.n28 VGND.n27 0.16782
R145 VGND.n70 VGND.n0 0.155855
R146 VGND.n23 VGND.n17 0.122949
R147 VGND.n24 VGND.n23 0.122949
R148 VGND.n26 VGND.n24 0.122949
R149 VGND.n26 VGND.n25 0.122949
R150 VGND.n25 VGND.n14 0.122949
R151 VGND.n33 VGND.n14 0.122949
R152 VGND.n34 VGND.n33 0.122949
R153 VGND.n35 VGND.n34 0.122949
R154 VGND.n35 VGND.n12 0.122949
R155 VGND.n39 VGND.n12 0.122949
R156 VGND.n40 VGND.n39 0.122949
R157 VGND.n41 VGND.n40 0.122949
R158 VGND.n41 VGND.n9 0.122949
R159 VGND.n45 VGND.n9 0.122949
R160 VGND.n46 VGND.n45 0.122949
R161 VGND.n47 VGND.n46 0.122949
R162 VGND.n47 VGND.n7 0.122949
R163 VGND.n52 VGND.n7 0.122949
R164 VGND.n53 VGND.n52 0.122949
R165 VGND.n53 VGND.n5 0.122949
R166 VGND.n58 VGND.n5 0.122949
R167 VGND.n59 VGND.n58 0.122949
R168 VGND.n60 VGND.n59 0.122949
R169 VGND.n60 VGND.n3 0.122949
R170 VGND.n64 VGND.n3 0.122949
R171 VGND.n65 VGND.n64 0.122949
R172 VGND.n66 VGND.n65 0.122949
R173 VGND.n66 VGND.n0 0.122949
R174 VNB.n0 VNB 16583.7
R175 VNB VNB.n1 14388.2
R176 VNB.t3 VNB.t14 3556.96
R177 VNB.t22 VNB.t0 3429.92
R178 VNB.t2 VNB.t4 2840.95
R179 VNB.t19 VNB.t18 2563.78
R180 VNB.t14 VNB.t12 2286.61
R181 VNB.t8 VNB.t6 2286.61
R182 VNB.t1 VNB.n0 1623.53
R183 VNB.t17 VNB.t19 1570.6
R184 VNB.n1 VNB.t20 1408.92
R185 VNB.t21 VNB 1385.83
R186 VNB.t15 VNB.t17 1328.08
R187 VNB.t4 VNB.t15 1177.95
R188 VNB.t11 VNB.t13 1154.86
R189 VNB.t16 VNB.t3 1097.11
R190 VNB.t13 VNB.t10 1027.82
R191 VNB.t12 VNB.t11 993.177
R192 VNB.t9 VNB.t22 993.177
R193 VNB.t0 VNB.t5 993.177
R194 VNB.t7 VNB.t8 993.177
R195 VNB.t5 VNB.t7 900.788
R196 VNB.t6 VNB.t21 900.788
R197 VNB.n1 VNB.t1 882.354
R198 VNB.t18 VNB.t16 831.496
R199 VNB.t20 VNB.t9 831.496
R200 VNB.n0 VNB.t2 681.365
R201 Q.n6 Q.n5 585
R202 Q.n5 Q.n3 295.854
R203 Q.n10 Q.n9 204.935
R204 Q.n11 Q.n0 97.6592
R205 Q.n2 Q.n1 84.9229
R206 Q.n4 Q.n3 80.7144
R207 Q.n8 Q.n2 44.0509
R208 Q.n7 Q.n3 37.6588
R209 Q.n4 Q.n2 26.9085
R210 Q.n9 Q.t5 26.3844
R211 Q.n9 Q.t4 26.3844
R212 Q.n5 Q.t6 26.3844
R213 Q.n0 Q.t0 24.3248
R214 Q.n0 Q.t3 23.514
R215 Q.n1 Q.t1 22.7032
R216 Q.n1 Q.t2 22.7032
R217 Q.n10 Q.n8 10.0448
R218 Q Q.n11 4.58918
R219 Q.n7 Q.n6 0.543896
R220 Q.n8 Q.n7 0.242009
R221 Q.n11 Q.n10 0.221354
R222 Q.n6 Q.n4 0.181632
R223 VPWR.n50 VPWR.t1 891.668
R224 VPWR.n35 VPWR.t10 859.285
R225 VPWR.n0 VPWR.t9 722.067
R226 VPWR.n37 VPWR.t11 690.981
R227 VPWR.n55 VPWR.n7 613.928
R228 VPWR.n62 VPWR.n3 612.136
R229 VPWR.n28 VPWR.n27 585
R230 VPWR.n19 VPWR.t6 349.418
R231 VPWR.n20 VPWR.t5 342.784
R232 VPWR.n22 VPWR.t7 249.317
R233 VPWR.n27 VPWR.t8 121.293
R234 VPWR.n27 VPWR.t2 119.608
R235 VPWR.n3 VPWR.t4 116.969
R236 VPWR.n7 VPWR.t12 116.969
R237 VPWR.n3 VPWR.t0 46.1724
R238 VPWR.n7 VPWR.t3 46.1724
R239 VPWR.n64 VPWR.n63 36.1417
R240 VPWR.n57 VPWR.n56 36.1417
R241 VPWR.n57 VPWR.n4 36.1417
R242 VPWR.n61 VPWR.n4 36.1417
R243 VPWR.n54 VPWR.n8 36.1417
R244 VPWR.n49 VPWR.n48 36.1417
R245 VPWR.n42 VPWR.n12 36.1417
R246 VPWR.n43 VPWR.n42 36.1417
R247 VPWR.n44 VPWR.n43 36.1417
R248 VPWR.n38 VPWR.n36 36.1417
R249 VPWR.n30 VPWR.n29 36.1417
R250 VPWR.n30 VPWR.n15 36.1417
R251 VPWR.n34 VPWR.n15 36.1417
R252 VPWR.n44 VPWR.n10 34.6358
R253 VPWR.n35 VPWR.n34 32.7534
R254 VPWR.n56 VPWR.n55 30.8711
R255 VPWR.n22 VPWR.n17 30.4946
R256 VPWR.n64 VPWR.n0 29.7417
R257 VPWR.n62 VPWR.n61 29.7417
R258 VPWR.n50 VPWR.n49 27.8593
R259 VPWR.n21 VPWR.n20 25.977
R260 VPWR.n26 VPWR.n17 24.7221
R261 VPWR.n63 VPWR.n62 23.7181
R262 VPWR.n55 VPWR.n54 22.5887
R263 VPWR.n50 VPWR.n8 19.577
R264 VPWR.n22 VPWR.n21 16.9417
R265 VPWR.n29 VPWR.n28 14.6829
R266 VPWR.n36 VPWR.n35 14.6829
R267 VPWR.n48 VPWR.n10 12.8005
R268 VPWR.n21 VPWR.n18 9.3005
R269 VPWR.n23 VPWR.n22 9.3005
R270 VPWR.n24 VPWR.n17 9.3005
R271 VPWR.n26 VPWR.n25 9.3005
R272 VPWR.n29 VPWR.n16 9.3005
R273 VPWR.n31 VPWR.n30 9.3005
R274 VPWR.n32 VPWR.n15 9.3005
R275 VPWR.n34 VPWR.n33 9.3005
R276 VPWR.n35 VPWR.n14 9.3005
R277 VPWR.n36 VPWR.n13 9.3005
R278 VPWR.n39 VPWR.n38 9.3005
R279 VPWR.n40 VPWR.n12 9.3005
R280 VPWR.n42 VPWR.n41 9.3005
R281 VPWR.n43 VPWR.n11 9.3005
R282 VPWR.n45 VPWR.n44 9.3005
R283 VPWR.n46 VPWR.n10 9.3005
R284 VPWR.n48 VPWR.n47 9.3005
R285 VPWR.n49 VPWR.n9 9.3005
R286 VPWR.n51 VPWR.n50 9.3005
R287 VPWR.n52 VPWR.n8 9.3005
R288 VPWR.n54 VPWR.n53 9.3005
R289 VPWR.n55 VPWR.n6 9.3005
R290 VPWR.n56 VPWR.n5 9.3005
R291 VPWR.n58 VPWR.n57 9.3005
R292 VPWR.n59 VPWR.n4 9.3005
R293 VPWR.n61 VPWR.n60 9.3005
R294 VPWR.n62 VPWR.n2 9.3005
R295 VPWR.n63 VPWR.n1 9.3005
R296 VPWR.n65 VPWR.n64 9.3005
R297 VPWR.n37 VPWR.n12 9.03579
R298 VPWR.n66 VPWR.n0 7.1518
R299 VPWR.n20 VPWR.n19 6.46335
R300 VPWR.n38 VPWR.n37 2.25932
R301 VPWR.n28 VPWR.n26 1.2554
R302 VPWR.n19 VPWR.n18 0.686829
R303 VPWR VPWR.n66 0.274639
R304 VPWR.n66 VPWR.n65 0.156154
R305 VPWR.n23 VPWR.n18 0.122949
R306 VPWR.n24 VPWR.n23 0.122949
R307 VPWR.n25 VPWR.n24 0.122949
R308 VPWR.n25 VPWR.n16 0.122949
R309 VPWR.n31 VPWR.n16 0.122949
R310 VPWR.n32 VPWR.n31 0.122949
R311 VPWR.n33 VPWR.n32 0.122949
R312 VPWR.n33 VPWR.n14 0.122949
R313 VPWR.n14 VPWR.n13 0.122949
R314 VPWR.n39 VPWR.n13 0.122949
R315 VPWR.n40 VPWR.n39 0.122949
R316 VPWR.n41 VPWR.n40 0.122949
R317 VPWR.n41 VPWR.n11 0.122949
R318 VPWR.n45 VPWR.n11 0.122949
R319 VPWR.n46 VPWR.n45 0.122949
R320 VPWR.n47 VPWR.n46 0.122949
R321 VPWR.n47 VPWR.n9 0.122949
R322 VPWR.n51 VPWR.n9 0.122949
R323 VPWR.n52 VPWR.n51 0.122949
R324 VPWR.n53 VPWR.n52 0.122949
R325 VPWR.n53 VPWR.n6 0.122949
R326 VPWR.n6 VPWR.n5 0.122949
R327 VPWR.n58 VPWR.n5 0.122949
R328 VPWR.n59 VPWR.n58 0.122949
R329 VPWR.n60 VPWR.n59 0.122949
R330 VPWR.n60 VPWR.n2 0.122949
R331 VPWR.n2 VPWR.n1 0.122949
R332 VPWR.n65 VPWR.n1 0.122949
R333 a_1943_53.t1 a_1943_53.n4 847.37
R334 a_1943_53.n2 a_1943_53.n1 379.442
R335 a_1943_53.n0 a_1943_53.t3 303.928
R336 a_1943_53.n3 a_1943_53.t0 239.486
R337 a_1943_53.n3 a_1943_53.n2 210.492
R338 a_1943_53.n2 a_1943_53.t2 199.227
R339 a_1943_53.n0 a_1943_53.t4 194.992
R340 a_1943_53.n4 a_1943_53.n0 166.683
R341 a_1943_53.n4 a_1943_53.n3 32.377
R342 a_1858_79.t0 a_1858_79.t1 121.43
R343 D.n0 D.t0 219.31
R344 D D.n0 159.84
R345 D.n1 D 154.081
R346 D.n1 D.t1 152.633
R347 D.n3 D.n2 152
R348 D.n2 D.n0 49.6611
R349 D.n2 D.n1 49.6611
R350 D.n3 D 8.8005
R351 D D.n3 3.0405
R352 a_37_464.n0 a_37_464.t5 356.454
R353 a_37_464.n0 a_37_464.t4 345.558
R354 a_37_464.n3 a_37_464.n2 301.264
R355 a_37_464.n2 a_37_464.n1 295.882
R356 a_37_464.n2 a_37_464.n0 273.318
R357 a_37_464.n3 a_37_464.t3 46.1724
R358 a_37_464.t1 a_37_464.n3 46.1724
R359 a_37_464.n1 a_37_464.t0 40.0005
R360 a_37_464.n1 a_37_464.t2 40.0005
R361 a_126_464.t0 a_126_464.t1 83.1099
R362 CLK.n0 CLK.t0 276.348
R363 CLK.n0 CLK.t1 178.34
R364 CLK CLK.n0 162.206
R365 a_1313_74.t0 a_1313_74.n7 879.54
R366 a_1313_74.n3 a_1313_74.n2 568.939
R367 a_1313_74.n2 a_1313_74.t3 310.087
R368 a_1313_74.n4 a_1313_74.n3 305.267
R369 a_1313_74.n4 a_1313_74.t5 295.627
R370 a_1313_74.n6 a_1313_74.t2 290.437
R371 a_1313_74.n7 a_1313_74.t1 233.076
R372 a_1313_74.n2 a_1313_74.t4 231.629
R373 a_1313_74.n5 a_1313_74.n4 226.541
R374 a_1313_74.n5 a_1313_74.n0 204.048
R375 a_1313_74.n7 a_1313_74.n6 184.133
R376 a_1313_74.n3 a_1313_74.n1 151.831
R377 a_1313_74.n6 a_1313_74.n5 144.601
R378 SCD.n0 SCD.t1 272.866
R379 SCD.n0 SCD.t0 210.474
R380 SCD SCD.n0 163.412
R381 a_1044_125.t0 a_1044_125.t1 60.0005
R382 a_2331_74.t0 a_2331_74.t1 39.3755
R383 SCE.t3 SCE.t1 626.601
R384 SCE.t2 SCE.t0 569.029
R385 SCE.n0 SCE.t2 335.435
R386 SCE SCE.n0 157.625
R387 SCE.n0 SCE.t3 134.601
R388 a_661_113.t0 a_661_113.n3 718.404
R389 a_661_113.t0 a_661_113.n3 708.125
R390 a_661_113.n0 a_661_113.t4 701.72
R391 a_661_113.n0 a_661_113.t5 409.55
R392 a_661_113.n2 a_661_113.t1 382.031
R393 a_661_113.n2 a_661_113.t3 351.228
R394 a_661_113.n1 a_661_113.t2 330.971
R395 a_661_113.n3 a_661_113.n2 195.882
R396 a_661_113.n1 a_661_113.n0 125.2
R397 a_661_113.n3 a_661_113.n1 11.2645
R398 a_135_74.t0 a_135_74.t1 68.5719
R399 a_572_463.t0 a_572_463.t1 73.8755
R400 a_1756_97.n1 a_1756_97.t0 717.747
R401 a_1756_97.n0 a_1756_97.t3 273.134
R402 a_1756_97.n2 a_1756_97.n1 262.93
R403 a_1756_97.n1 a_1756_97.n0 248.218
R404 a_1756_97.n0 a_1756_97.t4 208.6
R405 a_1756_97.n2 a_1756_97.t2 40.0005
R406 a_1756_97.n3 a_1756_97.n2 34.546
R407 a_1756_97.n3 a_1756_97.t1 25.4063
R408 a_1756_97.n4 a_1756_97.n3 21.6005
R409 DE.n0 DE.t1 345.433
R410 DE.n1 DE.t3 329.368
R411 DE.n2 DE.n0 276.348
R412 DE DE.n2 154.923
R413 DE.n1 DE.t0 128.534
R414 DE.n0 DE.t2 126.927
R415 DE.n2 DE.n1 51.1217
R416 a_177_290.t0 a_177_290.n1 660.913
R417 a_177_290.n1 a_177_290.t3 451.839
R418 a_177_290.n0 a_177_290.t1 288.93
R419 a_177_290.n0 a_177_290.t2 259.634
R420 a_177_290.n1 a_177_290.n0 50.5479
R421 a_497_113.t0 a_497_113.t1 68.5719
R422 a_2292_392.t0 a_2292_392.t1 159.571
R423 a_631_87.t0 a_631_87.n1 656.511
R424 a_631_87.n1 a_631_87.t2 373.161
R425 a_631_87.n0 a_631_87.t3 354.491
R426 a_631_87.n0 a_631_87.t1 246.544
R427 a_631_87.n1 a_631_87.n0 32.0025
R428 a_1071_455.t0 a_1071_455.t1 73.8755
C0 VGND Q 0.279523f
C1 SCD VGND 0.029929f
C2 SCE VGND 0.069248f
C3 VGND VPWR 0.080094f
C4 DE SCE 6.71e-20
C5 DE VPWR 0.024746f
C6 VGND VPB 0.013134f
C7 D VPWR 0.013628f
C8 DE VPB 0.170447f
C9 D VPB 0.073462f
C10 VGND a_1510_74# 0.567892f
C11 DE VGND 0.03786f
C12 VGND D 0.022407f
C13 DE D 0.043496f
C14 SCD CLK 0.003409f
C15 CLK SCE 0.003821f
C16 CLK VPWR 0.014837f
C17 CLK VPB 0.039516f
C18 CLK VGND 0.014686f
C19 SCD SCE 0.129969f
C20 Q VPWR 0.39346f
C21 SCD VPWR 0.01323f
C22 SCE VPWR 0.029698f
C23 Q VPB 0.015904f
C24 SCD VPB 0.061824f
C25 SCE VPB 0.18306f
C26 VPWR VPB 0.486569f
C27 a_1899_508# VPWR 0.006969f
C28 SCE a_1510_74# 4.03e-19
C29 VPWR a_1510_74# 0.020773f
C30 a_1510_74# VPB 0.224642f
C31 Q VNB 0.065249f
C32 VGND VNB 2.00461f
C33 CLK VNB 0.130454f
C34 SCD VNB 0.108168f
C35 SCE VNB 0.348104f
C36 DE VNB 0.295705f
C37 VPWR VNB 1.47927f
C38 D VNB 0.190752f
C39 VPB VNB 3.83905f
C40 a_1510_74# VNB 0.364478f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xnor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor3_1 VNB VPB VPWR VGND X B C A
X0 a_1113_383.t0 a_897_54.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1376 ps=1.07 w=0.64 l=0.15
X1 a_81_268.t1 C.t0 a_363_394.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.208975 pd=1.425 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 VGND.t3 a_81_268.t4 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.19575 pd=1.49 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_232_162.t0 C.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1575 pd=1.59 as=0.19575 ps=1.49 w=0.42 l=0.15
X4 a_786_100.t0 B.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.36 ps=2.83 w=0.74 l=0.15
X5 a_363_394.t0 a_786_100.t2 a_897_54.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1527 pd=1.225 as=0.36585 ps=2.87 w=0.84 l=0.15
X6 a_371_74.t0 a_786_100.t3 a_897_54.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1328 pd=1.055 as=0.374625 ps=2.77 w=0.64 l=0.15
X7 a_371_74.t4 a_232_162.t2 a_81_268.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=2.26 as=0.208975 ps=1.425 w=0.84 l=0.15
X8 a_1113_383.t2 B.t1 a_371_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1136 pd=1.05 as=0.1328 ps=1.055 w=0.64 l=0.15
X9 VGND.t4 A.t0 a_897_54.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.07 as=0.1104 ps=0.985 w=0.64 l=0.15
X10 a_232_162.t1 C.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.2404 ps=1.65 w=0.64 l=0.15
X11 a_786_100.t1 B.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.4194 ps=3.08 w=1.12 l=0.15
X12 a_897_54.t3 B.t3 a_371_74.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1858 pd=1.39 as=0.1852 ps=1.325 w=0.84 l=0.15
X13 a_363_394.t2 a_232_162.t3 a_81_268.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.112 ps=0.99 w=0.64 l=0.15
X14 a_1113_383.t1 a_897_54.t7 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.1925 ps=1.385 w=1 l=0.15
X15 a_363_394.t3 a_786_100.t4 a_1113_383.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.09995 pd=0.985 as=0.1136 ps=1.05 w=0.42 l=0.15
X16 VPWR.t1 A.t1 a_897_54.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1925 pd=1.385 as=0.1858 ps=1.39 w=1 l=0.15
X17 VPWR.t0 a_81_268.t5 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2404 pd=1.65 as=0.3192 ps=2.81 w=1.12 l=0.15
X18 a_81_268.t0 C.t3 a_371_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X19 a_1113_383.t4 B.t4 a_363_394.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1527 ps=1.225 w=0.64 l=0.15
X20 a_897_54.t5 B.t5 a_363_394.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1104 pd=0.985 as=0.09995 ps=0.985 w=0.64 l=0.15
R0 a_897_54.n4 a_897_54.t1 1058.32
R1 a_897_54.n1 a_897_54.t4 519.34
R2 a_897_54.n5 a_897_54.n4 287.779
R3 a_897_54.n2 a_897_54.t7 231.629
R4 a_897_54.n2 a_897_54.t6 184.768
R5 a_897_54.n3 a_897_54.n2 152
R6 a_897_54.n1 a_897_54.n0 89.3175
R7 a_897_54.n4 a_897_54.n3 62.9506
R8 a_897_54.n3 a_897_54.n1 62.4528
R9 a_897_54.n5 a_897_54.t3 55.1136
R10 a_897_54.n0 a_897_54.t5 38.438
R11 a_897_54.t0 a_897_54.n5 32.4514
R12 a_897_54.n0 a_897_54.t2 26.2505
R13 VGND.n6 VGND.t0 387.914
R14 VGND.n1 VGND.n0 268.276
R15 VGND.n5 VGND.n4 214.97
R16 VGND.n0 VGND.t1 74.2862
R17 VGND.n4 VGND.t4 46.8755
R18 VGND.n7 VGND.n3 36.1417
R19 VGND.n11 VGND.n3 36.1417
R20 VGND.n12 VGND.n11 36.1417
R21 VGND.n13 VGND.n12 36.1417
R22 VGND.n4 VGND.t2 33.7505
R23 VGND.n0 VGND.t3 29.1897
R24 VGND.n13 VGND.n1 22.1206
R25 VGND.n7 VGND.n6 20.7064
R26 VGND.n14 VGND.n13 9.3005
R27 VGND.n12 VGND.n2 9.3005
R28 VGND.n11 VGND.n10 9.3005
R29 VGND.n9 VGND.n3 9.3005
R30 VGND.n8 VGND.n7 9.3005
R31 VGND.n15 VGND.n1 9.10055
R32 VGND.n6 VGND.n5 7.296
R33 VGND VGND.n15 0.161517
R34 VGND.n8 VGND.n5 0.155071
R35 VGND.n15 VGND.n14 0.146304
R36 VGND.n9 VGND.n8 0.122949
R37 VGND.n10 VGND.n9 0.122949
R38 VGND.n10 VGND.n2 0.122949
R39 VGND.n14 VGND.n2 0.122949
R40 a_1113_383.n1 a_1113_383.t4 806.506
R41 a_1113_383.t1 a_1113_383.n2 381.726
R42 a_1113_383.n1 a_1113_383.n0 193.053
R43 a_1113_383.n2 a_1113_383.t0 141.668
R44 a_1113_383.n0 a_1113_383.t2 59.1523
R45 a_1113_383.n0 a_1113_383.t3 45.7148
R46 a_1113_383.n2 a_1113_383.n1 20.2135
R47 VNB.t7 VNB.t1 2633.07
R48 VNB.t2 VNB.t0 2609.97
R49 VNB.t1 VNB.t9 2575.33
R50 VNB.t4 VNB.t2 1362.73
R51 VNB.t6 VNB.t3 1339.63
R52 VNB.t9 VNB.t5 1304.99
R53 VNB.t5 VNB.t8 1293.44
R54 VNB.t0 VNB.t7 1154.86
R55 VNB.t10 VNB.t6 1143.31
R56 VNB.t8 VNB.t10 1143.31
R57 VNB VNB.t4 1143.31
R58 C.n1 C.n0 271.527
R59 C.n0 C.t0 264.832
R60 C.n0 C.t3 200.958
R61 C.n2 C.t2 173.788
R62 C C.n2 154.522
R63 C.n1 C.t1 116.996
R64 C.n2 C.n1 13.146
R65 a_363_394.n3 a_363_394.t1 472.361
R66 a_363_394.n0 a_363_394.n3 418.301
R67 a_363_394.n2 a_363_394.n1 406.947
R68 a_363_394.n2 a_363_394.t2 136.167
R69 a_363_394.n3 a_363_394.n2 105.412
R70 a_363_394.n0 a_363_394.t4 72.3364
R71 a_363_394.n1 a_363_394.t3 58.5719
R72 a_363_394.n4 a_363_394.n0 50.0852
R73 a_363_394.n0 a_363_394.t0 32.7911
R74 a_363_394.n1 a_363_394.t5 27.7237
R75 a_81_268.n3 a_81_268.n2 800.971
R76 a_81_268.n2 a_81_268.n0 288.702
R77 a_81_268.n1 a_81_268.t5 252.208
R78 a_81_268.n1 a_81_268.t4 176.964
R79 a_81_268.n2 a_81_268.n1 152
R80 a_81_268.t1 a_81_268.n3 53.941
R81 a_81_268.n3 a_81_268.t2 52.7684
R82 a_81_268.n0 a_81_268.t0 39.3755
R83 a_81_268.n0 a_81_268.t3 26.2505
R84 VPB.t6 VPB.t2 559.274
R85 VPB.t9 VPB.t7 554.168
R86 VPB.t8 VPB.t6 546.505
R87 VPB.t3 VPB.t4 515.861
R88 VPB.t1 VPB.t3 347.312
R89 VPB.t4 VPB.t8 309.005
R90 VPB.t7 VPB.t0 275.807
R91 VPB.t0 VPB.t5 273.253
R92 VPB.t2 VPB.t9 273.253
R93 VPB VPB.t1 252.823
R94 X.n0 X.t1 295.872
R95 X.n1 X.t0 279.738
R96 X.t0 X.n0 246.054
R97 X X.n1 7.28939
R98 X X.n0 5.86717
R99 X.n1 X 5.86717
R100 a_232_162.t1 a_232_162.n1 656.288
R101 a_232_162.n1 a_232_162.t0 276.954
R102 a_232_162.n0 a_232_162.t3 275.642
R103 a_232_162.n1 a_232_162.n0 228.8
R104 a_232_162.n0 a_232_162.t2 203.611
R105 B.n2 B.n0 824.227
R106 B.n0 B.t3 535.557
R107 B.t3 B.t5 445.048
R108 B.t4 B.t1 407.175
R109 B.n0 B.t4 266.171
R110 B.n1 B.t2 226.809
R111 B.n1 B.t0 154.97
R112 B B.n2 67.806
R113 B.n2 B.n1 22.7194
R114 a_786_100.t1 a_786_100.n2 834.082
R115 a_786_100.t3 a_786_100.t4 821.008
R116 a_786_100.t4 a_786_100.n0 367.392
R117 a_786_100.n2 a_786_100.t0 339.303
R118 a_786_100.n1 a_786_100.t2 211.278
R119 a_786_100.n1 a_786_100.t3 162.274
R120 a_786_100.n2 a_786_100.n1 152
R121 a_371_74.n1 a_371_74.t4 899.992
R122 a_371_74.n3 a_371_74.n2 701.194
R123 a_371_74.n1 a_371_74.t1 231.636
R124 a_371_74.n2 a_371_74.n0 192.376
R125 a_371_74.n3 a_371_74.t3 40.6191
R126 a_371_74.n0 a_371_74.t2 39.3755
R127 a_371_74.n0 a_371_74.t0 38.438
R128 a_371_74.n2 a_371_74.n1 21.4992
R129 A.n0 A.t1 231.629
R130 A.n0 A.t0 184.768
R131 A A.n0 157.95
R132 VPWR.n6 VPWR.t4 862.58
R133 VPWR.n5 VPWR.n4 325.087
R134 VPWR.n14 VPWR.n1 323.55
R135 VPWR.n1 VPWR.t2 117.749
R136 VPWR.n4 VPWR.t1 46.2955
R137 VPWR.n8 VPWR.n7 36.1417
R138 VPWR.n8 VPWR.n2 36.1417
R139 VPWR.n12 VPWR.n2 36.1417
R140 VPWR.n13 VPWR.n12 36.1417
R141 VPWR.n14 VPWR.n13 29.7417
R142 VPWR.n4 VPWR.t3 29.5505
R143 VPWR.n1 VPWR.t0 26.2634
R144 VPWR.n7 VPWR.n6 20.7064
R145 VPWR.n7 VPWR.n3 9.3005
R146 VPWR.n9 VPWR.n8 9.3005
R147 VPWR.n10 VPWR.n2 9.3005
R148 VPWR.n12 VPWR.n11 9.3005
R149 VPWR.n13 VPWR.n0 9.3005
R150 VPWR.n6 VPWR.n5 7.296
R151 VPWR.n15 VPWR.n14 7.23624
R152 VPWR VPWR.n15 0.157488
R153 VPWR.n5 VPWR.n3 0.15507
R154 VPWR.n15 VPWR.n0 0.150282
R155 VPWR.n9 VPWR.n3 0.122949
R156 VPWR.n10 VPWR.n9 0.122949
R157 VPWR.n11 VPWR.n10 0.122949
R158 VPWR.n11 VPWR.n0 0.122949
C0 VPWR VGND 0.038062f
C1 VPB VPWR 0.195167f
C2 B X 1.02e-19
C3 A B 0.053708f
C4 C X 0.001082f
C5 VPB VGND 0.007415f
C6 VPWR X 0.088853f
C7 VPWR A 0.012661f
C8 C B 6.83e-19
C9 VGND X 0.039597f
C10 A VGND 0.008997f
C11 VPB X 0.013215f
C12 VPWR B 0.083707f
C13 VPB A 0.038862f
C14 VPWR C 0.010249f
C15 VGND B 0.013742f
C16 C VGND 0.010226f
C17 VPB B 0.490007f
C18 VPB C 0.116963f
C19 VGND VNB 0.952735f
C20 A VNB 0.094939f
C21 C VNB 0.288269f
C22 X VNB 0.110441f
C23 B VNB 0.401745f
C24 VPWR VNB 0.744927f
C25 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xnor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor3_2 VNB VPB VPWR VGND X B C A
X0 VPWR.t1 a_83_247.t6 a_27_373.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.295 ps=2.59 w=1 l=0.15
X1 VPWR.t0 C.t0 a_1027_48.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2404 pd=1.65 as=0.1856 ps=1.86 w=0.64 l=0.15
X2 a_329_81.t0 C.t1 a_1057_74.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=2.26 as=0.213825 ps=1.435 w=0.84 l=0.15
X3 a_332_373.t3 B.t0 a_83_247.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1742 pd=1.3 as=0.1866 ps=1.39 w=0.84 l=0.15
X4 VGND.t5 B.t1 a_397_21.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.3368 pd=2.67 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_329_81.t4 B.t2 a_83_247.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1198 pd=1.2 as=0.12 ps=1.015 w=0.64 l=0.15
X6 a_1057_74.t2 a_1027_48.t2 a_329_81.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X7 VGND.t1 a_83_247.t7 a_27_373.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1152 pd=1 as=0.1824 ps=1.85 w=0.64 l=0.15
X8 X.t2 a_1057_74.t4 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2404 ps=1.65 w=1.12 l=0.15
X9 a_329_81.t2 B.t3 a_27_373.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1543 pd=1.23 as=0.1024 ps=0.96 w=0.64 l=0.15
X10 VGND.t3 a_1057_74.t5 X.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_1057_74.t3 a_1027_48.t3 a_332_373.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.213825 pd=1.435 as=0.2436 ps=2.26 w=0.84 l=0.15
X12 a_83_247.t3 a_397_21.t2 a_332_373.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.3525 pd=2.83 as=0.112 ps=0.99 w=0.64 l=0.15
X13 VGND.t0 C.t2 a_1027_48.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.382125 pd=1.845 as=0.1197 ps=1.41 w=0.42 l=0.15
X14 a_83_247.t1 a_397_21.t3 a_329_81.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3766 pd=2.89 as=0.1543 ps=1.23 w=0.84 l=0.15
X15 a_83_247.t2 A.t0 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12 pd=1.015 as=0.1152 ps=1 w=0.64 l=0.15
X16 X.t0 a_1057_74.t6 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.382125 ps=1.845 w=0.74 l=0.15
X17 a_27_373.t0 a_397_21.t4 a_332_373.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1024 pd=0.96 as=0.1742 ps=1.3 w=0.64 l=0.15
X18 VPWR.t2 B.t4 a_397_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4382 pd=3.15 as=0.3248 ps=2.82 w=1.12 l=0.15
X19 a_332_373.t4 B.t5 a_27_373.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1031 ps=1 w=0.64 l=0.15
X20 a_83_247.t4 A.t1 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1866 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X21 a_27_373.t5 a_397_21.t5 a_329_81.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1031 pd=1 as=0.1198 ps=1.2 w=0.42 l=0.15
X22 a_332_373.t0 C.t3 a_1057_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.112 ps=0.99 w=0.64 l=0.15
R0 a_83_247.n7 a_83_247.t1 1040.18
R1 a_83_247.n6 a_83_247.n5 585
R2 a_83_247.n8 a_83_247.n7 585
R3 a_83_247.n2 a_83_247.t3 569.947
R4 a_83_247.n3 a_83_247.t6 269.118
R5 a_83_247.n3 a_83_247.t7 187.981
R6 a_83_247.n4 a_83_247.n3 152
R7 a_83_247.n2 a_83_247.n1 88.228
R8 a_83_247.n4 a_83_247.n2 63.2709
R9 a_83_247.n6 a_83_247.n4 62.5226
R10 a_83_247.n5 a_83_247.t0 53.941
R11 a_83_247.n9 a_83_247.n8 44.9303
R12 a_83_247.n1 a_83_247.t5 44.063
R13 a_83_247.n0 a_83_247.t4 28.8091
R14 a_83_247.n7 a_83_247.n6 27.6576
R15 a_83_247.n1 a_83_247.t2 26.2505
R16 a_83_247.n8 a_83_247.n0 10.3689
R17 a_83_247.n5 a_83_247.n0 4.69098
R18 a_27_373.n2 a_27_373.n1 447.87
R19 a_27_373.t2 a_27_373.n3 381.175
R20 a_27_373.n2 a_27_373.n0 220.28
R21 a_27_373.n3 a_27_373.t1 151.619
R22 a_27_373.n1 a_27_373.t0 52.3286
R23 a_27_373.n0 a_27_373.t3 50.5809
R24 a_27_373.n1 a_27_373.t4 46.1724
R25 a_27_373.n0 a_27_373.t5 40.0005
R26 a_27_373.n3 a_27_373.n2 19.7849
R27 VPWR.n5 VPWR.t2 867.895
R28 VPWR.n18 VPWR.n1 622.029
R29 VPWR.n7 VPWR.n6 389.217
R30 VPWR.n6 VPWR.t0 116.969
R31 VPWR.n1 VPWR.t4 44.3255
R32 VPWR.n10 VPWR.n4 36.1417
R33 VPWR.n11 VPWR.n10 36.1417
R34 VPWR.n12 VPWR.n11 36.1417
R35 VPWR.n12 VPWR.n2 36.1417
R36 VPWR.n16 VPWR.n2 36.1417
R37 VPWR.n17 VPWR.n16 36.1417
R38 VPWR.n1 VPWR.t1 32.5055
R39 VPWR.n5 VPWR.n4 28.2358
R40 VPWR.n6 VPWR.t3 24.7674
R41 VPWR.n18 VPWR.n17 20.7064
R42 VPWR.n8 VPWR.n4 9.3005
R43 VPWR.n10 VPWR.n9 9.3005
R44 VPWR.n11 VPWR.n3 9.3005
R45 VPWR.n13 VPWR.n12 9.3005
R46 VPWR.n14 VPWR.n2 9.3005
R47 VPWR.n16 VPWR.n15 9.3005
R48 VPWR.n17 VPWR.n0 9.3005
R49 VPWR.n19 VPWR.n18 7.52053
R50 VPWR.n7 VPWR.n5 6.87981
R51 VPWR.n8 VPWR.n7 0.161921
R52 VPWR VPWR.n19 0.161231
R53 VPWR.n19 VPWR.n0 0.146587
R54 VPWR.n9 VPWR.n8 0.122949
R55 VPWR.n9 VPWR.n3 0.122949
R56 VPWR.n13 VPWR.n3 0.122949
R57 VPWR.n14 VPWR.n13 0.122949
R58 VPWR.n15 VPWR.n14 0.122949
R59 VPWR.n15 VPWR.n0 0.122949
R60 VPB.t2 VPB.t5 566.936
R61 VPB.t5 VPB.t10 551.614
R62 VPB.t7 VPB.t1 510.753
R63 VPB.t1 VPB.t6 347.312
R64 VPB.t10 VPB.t7 314.113
R65 VPB.t0 VPB.t3 311.56
R66 VPB.t8 VPB.t2 275.807
R67 VPB.t9 VPB.t0 275.807
R68 VPB.t4 VPB.t9 275.807
R69 VPB VPB.t4 257.93
R70 VPB.t3 VPB.t8 240.054
R71 C.n0 C.t1 271.527
R72 C.n0 C.t3 265.101
R73 C.n1 C.n0 215.293
R74 C.n2 C.t0 166.257
R75 C C.n2 156.019
R76 C.n1 C.t2 113.572
R77 C.n2 C.n1 9.038
R78 a_1027_48.t1 a_1027_48.n1 654.062
R79 a_1027_48.n0 a_1027_48.t2 267.541
R80 a_1027_48.n1 a_1027_48.t0 242.517
R81 a_1027_48.n0 a_1027_48.t3 205.149
R82 a_1027_48.n1 a_1027_48.n0 192.339
R83 a_1057_74.n6 a_1057_74.n5 800.634
R84 a_1057_74.n5 a_1057_74.n0 289.682
R85 a_1057_74.n4 a_1057_74.t4 251.275
R86 a_1057_74.n2 a_1057_74.n1 246.892
R87 a_1057_74.n3 a_1057_74.t6 171.407
R88 a_1057_74.n2 a_1057_74.t5 155.149
R89 a_1057_74.n5 a_1057_74.n4 152
R90 a_1057_74.n3 a_1057_74.n2 63.6609
R91 a_1057_74.t0 a_1057_74.n6 55.1136
R92 a_1057_74.n6 a_1057_74.t3 53.941
R93 a_1057_74.n0 a_1057_74.t2 39.3755
R94 a_1057_74.n0 a_1057_74.t1 26.2505
R95 a_1057_74.n4 a_1057_74.n3 4.62242
R96 a_329_81.t0 a_329_81.n3 470.428
R97 a_329_81.n3 a_329_81.n0 405.147
R98 a_329_81.n2 a_329_81.n1 392.952
R99 a_329_81.n2 a_329_81.t3 143.775
R100 a_329_81.n3 a_329_81.n2 112.189
R101 a_329_81.n1 a_329_81.t5 86.7148
R102 a_329_81.n0 a_329_81.t2 73.8755
R103 a_329_81.n0 a_329_81.t1 35.1315
R104 a_329_81.n1 a_329_81.t4 24.3755
R105 B.n3 B.n2 798.659
R106 B.n2 B.t0 547.338
R107 B.t0 B.t2 486.017
R108 B.t3 B.t5 370.832
R109 B.n2 B.t3 279.56
R110 B.n0 B.t4 237.762
R111 B.n1 B.t1 171.913
R112 B B.n0 159.293
R113 B B.n3 154.828
R114 B.n3 B.n1 35.055
R115 B.n1 B.n0 14.6066
R116 a_332_373.n1 a_332_373.t5 814.806
R117 a_332_373.n3 a_332_373.n2 668.861
R118 a_332_373.n1 a_332_373.t0 295.276
R119 a_332_373.n2 a_332_373.n0 190.553
R120 a_332_373.n5 a_332_373.n4 72.9635
R121 a_332_373.n4 a_332_373.n3 53.8677
R122 a_332_373.n3 a_332_373.t1 46.1724
R123 a_332_373.n0 a_332_373.t2 36.563
R124 a_332_373.n4 a_332_373.t3 33.0098
R125 a_332_373.n0 a_332_373.t4 29.063
R126 a_332_373.n2 a_332_373.n1 20.642
R127 a_397_21.t1 a_397_21.n1 833.434
R128 a_397_21.t2 a_397_21.t5 803.333
R129 a_397_21.n1 a_397_21.t0 337.217
R130 a_397_21.t5 a_397_21.t4 322.94
R131 a_397_21.n0 a_397_21.t3 198.053
R132 a_397_21.n0 a_397_21.t2 154.405
R133 a_397_21.n1 a_397_21.n0 152
R134 VGND.n20 VGND.t5 355.781
R135 VGND.n11 VGND.n9 254.678
R136 VGND.n12 VGND.n11 252.743
R137 VGND.n33 VGND.n32 215.256
R138 VGND.n10 VGND.n7 194.555
R139 VGND.n8 VGND.t3 184.993
R140 VGND.n11 VGND.t0 73.321
R141 VGND.n32 VGND.t2 41.2505
R142 VGND.n10 VGND.t4 39.7302
R143 VGND.n14 VGND.n5 36.1417
R144 VGND.n18 VGND.n5 36.1417
R145 VGND.n19 VGND.n18 36.1417
R146 VGND.n24 VGND.n3 36.1417
R147 VGND.n25 VGND.n24 36.1417
R148 VGND.n26 VGND.n25 36.1417
R149 VGND.n26 VGND.n1 36.1417
R150 VGND.n30 VGND.n1 36.1417
R151 VGND.n31 VGND.n30 36.1417
R152 VGND.n20 VGND.n19 33.1299
R153 VGND.n14 VGND.n13 32.9597
R154 VGND.n32 VGND.t1 26.2505
R155 VGND.n11 VGND.n10 25.1356
R156 VGND.n33 VGND.n31 21.4593
R157 VGND.n20 VGND.n3 14.3064
R158 VGND.n31 VGND.n0 9.3005
R159 VGND.n30 VGND.n29 9.3005
R160 VGND.n28 VGND.n1 9.3005
R161 VGND.n27 VGND.n26 9.3005
R162 VGND.n25 VGND.n2 9.3005
R163 VGND.n24 VGND.n23 9.3005
R164 VGND.n22 VGND.n3 9.3005
R165 VGND.n21 VGND.n20 9.3005
R166 VGND.n19 VGND.n4 9.3005
R167 VGND.n18 VGND.n17 9.3005
R168 VGND.n16 VGND.n5 9.3005
R169 VGND.n15 VGND.n14 9.3005
R170 VGND.n13 VGND.n6 9.3005
R171 VGND.n12 VGND.n7 7.5692
R172 VGND.n9 VGND.n8 7.41446
R173 VGND.n34 VGND.n33 7.34058
R174 VGND.n13 VGND.n12 2.33789
R175 VGND.n8 VGND.n6 0.544755
R176 VGND.n9 VGND.n7 0.334413
R177 VGND VGND.n34 0.158861
R178 VGND.n34 VGND.n0 0.148926
R179 VGND.n15 VGND.n6 0.122949
R180 VGND.n16 VGND.n15 0.122949
R181 VGND.n17 VGND.n16 0.122949
R182 VGND.n17 VGND.n4 0.122949
R183 VGND.n21 VGND.n4 0.122949
R184 VGND.n22 VGND.n21 0.122949
R185 VGND.n23 VGND.n22 0.122949
R186 VGND.n23 VGND.n2 0.122949
R187 VGND.n27 VGND.n2 0.122949
R188 VGND.n28 VGND.n27 0.122949
R189 VGND.n29 VGND.n28 0.122949
R190 VGND.n29 VGND.n0 0.122949
R191 VNB.t10 VNB.t11 2471.39
R192 VNB.t3 VNB.t10 2471.39
R193 VNB.t0 VNB.t1 2448.29
R194 VNB.t1 VNB.t6 2182.68
R195 VNB VNB.t4 1235.7
R196 VNB.t5 VNB.t9 1212.6
R197 VNB.t2 VNB.t8 1177.95
R198 VNB.t4 VNB.t5 1177.95
R199 VNB.t11 VNB.t0 1154.86
R200 VNB.t8 VNB.t3 1154.86
R201 VNB.t9 VNB.t2 1131.76
R202 VNB.t6 VNB.t7 993.177
R203 X.n0 X.t2 292.507
R204 X.n1 X.n0 185
R205 X.n2 X.n1 185
R206 X.n1 X.t1 22.7032
R207 X.n1 X.t0 22.7032
R208 X X.n2 7.95202
R209 X X.n0 6.4005
R210 X.n2 X 6.4005
R211 A.n0 A.t0 232.968
R212 A.n0 A.t1 231.629
R213 A A.n0 153.423
C0 C VGND 0.014653f
C1 VPB VGND 0.010733f
C2 VPB C 0.126647f
C3 X VGND 0.13172f
C4 C X 0.001007f
C5 VPWR VGND 0.079504f
C6 VGND A 0.011946f
C7 VPB X 0.006028f
C8 VPWR C 0.011021f
C9 VPB VPWR 0.218891f
C10 VPB A 0.036484f
C11 VPWR X 0.187104f
C12 VGND B 0.014164f
C13 VPWR A 0.01389f
C14 C B 3.4e-19
C15 VPB B 0.49008f
C16 X B 1.48e-19
C17 VPWR B 0.082232f
C18 B A 0.058852f
C19 VGND VNB 1.02596f
C20 X VNB 0.02506f
C21 C VNB 0.314947f
C22 VPWR VNB 0.830907f
C23 A VNB 0.106911f
C24 B VNB 0.418322f
C25 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xnor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor3_4 VNB VPB VPWR VGND X B C A
X0 VPWR.t3 a_1057_74.t3 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t4 a_75_227.t6 a_27_373.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X2 a_75_227.t4 a_386_23.t2 a_324_373.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.3467 pd=2.79 as=0.096 ps=0.94 w=0.64 l=0.15
X3 a_1057_74.t1 a_1024_300# a_324_373.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.22785 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X4 a_324_373.t2 C.t0 a_1057_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.192 pd=1.88 as=0.1296 ps=1.045 w=0.64 l=0.15
X5 VPWR.t0 B.t0 a_386_23.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 VGND.t0 B.t1 a_386_23.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.3368 pd=2.67 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 a_1057_74.t2 a_1024_300# a_321_77.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1296 pd=1.045 as=0.1824 ps=1.85 w=0.64 l=0.15
X8 a_321_77.t2 B.t2 a_27_373.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1417 pd=1.2 as=0.096 ps=0.94 w=0.64 l=0.15
X9 a_27_373.t4 a_386_23.t3 a_321_77.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14055 pd=1.105 as=0.09575 ps=0.965 w=0.42 l=0.15
X10 a_324_373.t4 B.t3 a_27_373.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.096 pd=0.94 as=0.14055 ps=1.105 w=0.64 l=0.15
X11 a_75_227.t1 A.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1874 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X12 VGND.t7 C.t1 a_1024_300# VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.686625 pd=2.425 as=0.1197 ps=1.41 w=0.42 l=0.15
X13 a_27_373.t5 a_386_23.t4 a_324_373.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.2025 ps=1.39 w=0.64 l=0.15
X14 a_75_227.t5 a_386_23.t5 a_321_77.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.38735 pd=2.91 as=0.1417 ps=1.2 w=0.84 l=0.15
X15 VPWR C a_1024_300# VPB sky130_fd_pr__pfet_01v8 ad=0.5316 pd=2.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X16 VGND.t5 a_1057_74.t4 X.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_324_373.t5 B.t4 a_75_227.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2025 pd=1.39 as=0.1874 ps=1.39 w=0.84 l=0.15
X18 VGND.t6 a_75_227.t7 a_27_373.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X19 VGND.t4 a_1057_74.t5 X.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t2 a_1057_74.t6 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X21 X.t3 a_1057_74.t7 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_321_77.t3 B.t5 a_75_227.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.09575 pd=0.965 as=0.1072 ps=0.975 w=0.64 l=0.15
X23 X.t2 a_1057_74.t8 VGND.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.686625 ps=2.425 w=0.74 l=0.15
X24 a_75_227.t2 A.t1 VGND.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1072 pd=0.975 as=0.112 ps=0.99 w=0.64 l=0.15
R0 a_1057_74.t1 a_1057_74.n10 1004.27
R1 a_1057_74.n10 a_1057_74.n0 277.154
R2 a_1057_74.n3 a_1057_74.t6 230.825
R3 a_1057_74.n5 a_1057_74.n2 229.487
R4 a_1057_74.n7 a_1057_74.t3 229.487
R5 a_1057_74.n9 a_1057_74.n1 229.487
R6 a_1057_74.n3 a_1057_74.t4 156.465
R7 a_1057_74.n8 a_1057_74.t8 154.24
R8 a_1057_74.n6 a_1057_74.t5 154.24
R9 a_1057_74.n4 a_1057_74.t7 153.058
R10 a_1057_74.n10 a_1057_74.n9 93.2014
R11 a_1057_74.n4 a_1057_74.n3 60.785
R12 a_1057_74.n6 a_1057_74.n5 57.6944
R13 a_1057_74.n8 a_1057_74.n7 54.7732
R14 a_1057_74.n0 a_1057_74.t2 39.3755
R15 a_1057_74.n0 a_1057_74.t0 36.563
R16 a_1057_74.n9 a_1057_74.n8 10.955
R17 a_1057_74.n7 a_1057_74.n6 8.03383
R18 a_1057_74.n5 a_1057_74.n4 5.01811
R19 X.n8 X.n7 585
R20 X.n7 X.n0 291.033
R21 X.n2 X.t1 252.197
R22 X.n5 X.n4 185
R23 X.n4 X.n3 185
R24 X.n2 X.n1 117.966
R25 X.n6 X.n2 38.0883
R26 X.n7 X.t0 26.3844
R27 X.n1 X.t4 22.7032
R28 X.n1 X.t2 22.7032
R29 X.n4 X.t5 22.7032
R30 X.n4 X.t3 22.7032
R31 X X.n8 12.0794
R32 X.n6 X 11.7516
R33 X.n5 X 9.50353
R34 X X.n0 8.04766
R35 X.n3 X 7.95202
R36 X.n3 X 6.4005
R37 X.n0 X 5.20292
R38 X X.n5 4.84898
R39 X X.n6 2.16388
R40 X.n8 X 1.26247
R41 VPWR.n25 VPWR.t0 882.111
R42 VPWR.n37 VPWR.n1 319.615
R43 VPWR.n11 VPWR.t3 270.3
R44 VPWR.n10 VPWR.t2 264.682
R45 VPWR.n11 VPWR.n10 40.4499
R46 VPWR.n1 VPWR.t1 39.4005
R47 VPWR.n29 VPWR.n4 36.1417
R48 VPWR.n30 VPWR.n29 36.1417
R49 VPWR.n31 VPWR.n30 36.1417
R50 VPWR.n31 VPWR.n2 36.1417
R51 VPWR.n35 VPWR.n2 36.1417
R52 VPWR.n36 VPWR.n35 36.1417
R53 VPWR.n18 VPWR.n17 36.1417
R54 VPWR.n19 VPWR.n18 36.1417
R55 VPWR.n19 VPWR.n6 36.1417
R56 VPWR.n23 VPWR.n6 36.1417
R57 VPWR.n24 VPWR.n23 36.1417
R58 VPWR.n13 VPWR.n12 36.1417
R59 VPWR.n1 VPWR.t4 29.5505
R60 VPWR.n25 VPWR.n24 24.0946
R61 VPWR.n25 VPWR.n4 23.3417
R62 VPWR.n37 VPWR.n36 22.9652
R63 VPWR.n13 VPWR.n8 21.8358
R64 VPWR.n12 VPWR.n9 9.3005
R65 VPWR.n14 VPWR.n13 9.3005
R66 VPWR.n15 VPWR.n8 9.3005
R67 VPWR.n17 VPWR.n16 9.3005
R68 VPWR.n18 VPWR.n7 9.3005
R69 VPWR.n20 VPWR.n19 9.3005
R70 VPWR.n21 VPWR.n6 9.3005
R71 VPWR.n23 VPWR.n22 9.3005
R72 VPWR.n24 VPWR.n5 9.3005
R73 VPWR.n26 VPWR.n25 9.3005
R74 VPWR.n27 VPWR.n4 9.3005
R75 VPWR.n29 VPWR.n28 9.3005
R76 VPWR.n30 VPWR.n3 9.3005
R77 VPWR.n32 VPWR.n31 9.3005
R78 VPWR.n33 VPWR.n2 9.3005
R79 VPWR.n35 VPWR.n34 9.3005
R80 VPWR.n36 VPWR.n0 9.3005
R81 VPWR.n38 VPWR.n37 7.27223
R82 VPWR.n17 VPWR.n8 3.38874
R83 VPWR.n10 VPWR.n9 2.0675
R84 VPWR.n12 VPWR.n11 1.12991
R85 VPWR VPWR.n38 0.157962
R86 VPWR.n38 VPWR.n0 0.149814
R87 VPWR.n14 VPWR.n9 0.122949
R88 VPWR.n15 VPWR.n14 0.122949
R89 VPWR.n16 VPWR.n15 0.122949
R90 VPWR.n16 VPWR.n7 0.122949
R91 VPWR.n20 VPWR.n7 0.122949
R92 VPWR.n21 VPWR.n20 0.122949
R93 VPWR.n22 VPWR.n21 0.122949
R94 VPWR.n22 VPWR.n5 0.122949
R95 VPWR.n26 VPWR.n5 0.122949
R96 VPWR.n27 VPWR.n26 0.122949
R97 VPWR.n28 VPWR.n27 0.122949
R98 VPWR.n28 VPWR.n3 0.122949
R99 VPWR.n32 VPWR.n3 0.122949
R100 VPWR.n33 VPWR.n32 0.122949
R101 VPWR.n34 VPWR.n33 0.122949
R102 VPWR.n34 VPWR.n0 0.122949
R103 VPB.t3 VPB.t5 1700.81
R104 VPB.t9 VPB.t0 574.597
R105 VPB.t0 VPB.t3 515.861
R106 VPB.t5 VPB.t4 459.678
R107 VPB.t6 VPB.t8 357.527
R108 VPB.t2 VPB.t6 275.807
R109 VPB.t1 VPB.t9 260.485
R110 VPB VPB.t7 257.93
R111 VPB.t7 VPB.t2 255.376
R112 VPB.t8 VPB.t1 229.839
R113 a_75_227.n6 a_75_227.t5 1029.11
R114 a_75_227.n7 a_75_227.n6 585
R115 a_75_227.n2 a_75_227.t4 554.622
R116 a_75_227.n3 a_75_227.t6 295.894
R117 a_75_227.n5 a_75_227.n0 289.24
R118 a_75_227.n3 a_75_227.t7 162.274
R119 a_75_227.n4 a_75_227.n3 152
R120 a_75_227.n2 a_75_227.n1 88.228
R121 a_75_227.n5 a_75_227.n4 84.993
R122 a_75_227.n4 a_75_227.n2 65.4393
R123 a_75_227.n0 a_75_227.t3 56.2862
R124 a_75_227.n8 a_75_227.n7 43.4073
R125 a_75_227.n1 a_75_227.t0 36.563
R126 a_75_227.n0 a_75_227.t1 29.5767
R127 a_75_227.n1 a_75_227.t2 26.2505
R128 a_75_227.n6 a_75_227.n5 19.9033
R129 a_75_227.n7 a_75_227.n0 11.1901
R130 a_27_373.n2 a_27_373.n0 673.247
R131 a_27_373.n2 a_27_373.n1 297.063
R132 a_27_373.n3 a_27_373.t3 290.063
R133 a_27_373.t2 a_27_373.n3 232.595
R134 a_27_373.n1 a_27_373.t4 77.1434
R135 a_27_373.n0 a_27_373.t0 46.1724
R136 a_27_373.n0 a_27_373.t5 46.1724
R137 a_27_373.n1 a_27_373.t1 36.563
R138 a_27_373.n3 a_27_373.n2 20.1821
R139 a_386_23.t0 a_386_23.n1 815.274
R140 a_386_23.t2 a_386_23.t3 731.034
R141 a_386_23.t3 a_386_23.t4 443.173
R142 a_386_23.n1 a_386_23.t1 316.632
R143 a_386_23.n0 a_386_23.t5 205.922
R144 a_386_23.n1 a_386_23.n0 172.364
R145 a_386_23.n0 a_386_23.t2 168.701
R146 a_324_373.t3 a_324_373.n3 772.201
R147 a_324_373.n2 a_324_373.n1 585
R148 a_324_373.n3 a_324_373.t2 351.366
R149 a_324_373.n2 a_324_373.n0 259.226
R150 a_324_373.n1 a_324_373.t5 115.26
R151 a_324_373.n1 a_324_373.t0 46.1724
R152 a_324_373.n0 a_324_373.t1 28.1255
R153 a_324_373.n0 a_324_373.t4 28.1255
R154 a_324_373.n3 a_324_373.n2 22.9287
R155 VNB.t3 VNB.t8 3522.31
R156 VNB.t5 VNB.t6 2471.39
R157 VNB.t1 VNB.t5 2471.39
R158 VNB.t2 VNB.t3 2321.26
R159 VNB.t0 VNB.t12 1420.47
R160 VNB.t6 VNB.t2 1281.89
R161 VNB VNB.t13 1258.79
R162 VNB.t13 VNB.t7 1154.86
R163 VNB.t7 VNB.t4 1120.21
R164 VNB.t4 VNB.t0 1097.11
R165 VNB.t12 VNB.t1 1039.37
R166 VNB.t9 VNB.t11 993.177
R167 VNB.t10 VNB.t9 993.177
R168 VNB.t8 VNB.t10 993.177
R169 C.n2 C.n1 290.272
R170 C.n2 C.t0 245.821
R171 C.n3 C.n2 207.261
R172 C.n4 C.n0 168.852
R173 C C.n4 154.084
R174 C.n3 C.t1 114.751
R175 C.n4 C.n3 10.4535
R176 B.n2 B.n1 843.5
R177 B.n1 B.t4 569.832
R178 B.t4 B.t5 499.673
R179 B.t2 B.t3 386.805
R180 B.n1 B.t2 279.56
R181 B.n0 B.t0 254.56
R182 B.n0 B.t1 171.913
R183 B B.n2 155.274
R184 B.n2 B.n0 5.11262
R185 VGND.n37 VGND.t0 355.781
R186 VGND.n50 VGND.n49 208.856
R187 VGND.n27 VGND.n7 185
R188 VGND.n9 VGND.n8 185
R189 VGND.n26 VGND.n25 185
R190 VGND.n20 VGND.n19 185
R191 VGND.n29 VGND.n28 185
R192 VGND.n13 VGND.t5 183.456
R193 VGND.n12 VGND.n11 141.673
R194 VGND.n18 VGND.n17 94.4277
R195 VGND.n49 VGND.t6 39.3755
R196 VGND.n28 VGND.t7 38.0005
R197 VGND.n13 VGND.n12 37.0937
R198 VGND.n16 VGND.n15 36.1417
R199 VGND.n31 VGND.n5 36.1417
R200 VGND.n35 VGND.n5 36.1417
R201 VGND.n36 VGND.n35 36.1417
R202 VGND.n41 VGND.n3 36.1417
R203 VGND.n42 VGND.n41 36.1417
R204 VGND.n43 VGND.n42 36.1417
R205 VGND.n43 VGND.n1 36.1417
R206 VGND.n47 VGND.n1 36.1417
R207 VGND.n48 VGND.n47 36.1417
R208 VGND.n19 VGND.n8 33.7148
R209 VGND.n37 VGND.n36 33.1299
R210 VGND.n31 VGND.n30 32.9597
R211 VGND.n28 VGND.n27 28.5719
R212 VGND.n49 VGND.t1 26.2505
R213 VGND.n27 VGND.n26 24.5719
R214 VGND.n11 VGND.t3 22.7032
R215 VGND.n11 VGND.t4 22.7032
R216 VGND.n26 VGND.n8 20.0005
R217 VGND.n18 VGND.t2 19.5912
R218 VGND.n17 VGND.n16 19.1415
R219 VGND.n50 VGND.n48 15.4358
R220 VGND.n37 VGND.n3 14.3064
R221 VGND.n48 VGND.n0 9.3005
R222 VGND.n47 VGND.n46 9.3005
R223 VGND.n45 VGND.n1 9.3005
R224 VGND.n44 VGND.n43 9.3005
R225 VGND.n42 VGND.n2 9.3005
R226 VGND.n41 VGND.n40 9.3005
R227 VGND.n39 VGND.n3 9.3005
R228 VGND.n38 VGND.n37 9.3005
R229 VGND.n36 VGND.n4 9.3005
R230 VGND.n35 VGND.n34 9.3005
R231 VGND.n33 VGND.n5 9.3005
R232 VGND.n32 VGND.n31 9.3005
R233 VGND.n30 VGND.n6 9.3005
R234 VGND.n24 VGND.n23 9.3005
R235 VGND.n22 VGND.n21 9.3005
R236 VGND.n16 VGND.n10 9.3005
R237 VGND.n15 VGND.n14 9.3005
R238 VGND.n19 VGND.n18 9.14336
R239 VGND.n51 VGND.n50 7.57339
R240 VGND.n29 VGND.n7 4.84976
R241 VGND.n15 VGND.n12 4.51815
R242 VGND.n21 VGND.n9 2.97564
R243 VGND.n25 VGND.n9 2.42212
R244 VGND.n30 VGND.n29 2.33789
R245 VGND.n14 VGND.n13 2.0514
R246 VGND.n24 VGND.n7 1.73023
R247 VGND.n25 VGND.n24 1.24591
R248 VGND.n21 VGND.n20 1.10753
R249 VGND.n20 VGND.n17 0.837035
R250 VGND VGND.n51 0.161927
R251 VGND.n51 VGND.n0 0.1459
R252 VGND.n14 VGND.n10 0.122949
R253 VGND.n22 VGND.n10 0.122949
R254 VGND.n23 VGND.n22 0.122949
R255 VGND.n23 VGND.n6 0.122949
R256 VGND.n32 VGND.n6 0.122949
R257 VGND.n33 VGND.n32 0.122949
R258 VGND.n34 VGND.n33 0.122949
R259 VGND.n34 VGND.n4 0.122949
R260 VGND.n38 VGND.n4 0.122949
R261 VGND.n39 VGND.n38 0.122949
R262 VGND.n40 VGND.n39 0.122949
R263 VGND.n40 VGND.n2 0.122949
R264 VGND.n44 VGND.n2 0.122949
R265 VGND.n45 VGND.n44 0.122949
R266 VGND.n46 VGND.n45 0.122949
R267 VGND.n46 VGND.n0 0.122949
R268 a_321_77.n2 a_321_77.n1 505.428
R269 a_321_77.n1 a_321_77.n0 378.661
R270 a_321_77.n1 a_321_77.t4 144.803
R271 a_321_77.n2 a_321_77.t2 64.6411
R272 a_321_77.n0 a_321_77.t3 40.5809
R273 a_321_77.n0 a_321_77.t0 40.0005
R274 a_321_77.t1 a_321_77.n2 37.7532
R275 A.n0 A.t1 239.393
R276 A.n0 A.t0 231.629
R277 A A.n0 153.28
C0 C VGND 0.015559f
C1 VGND A 0.016524f
C2 VPB VGND 0.015567f
C3 a_1024_300# VGND 0.017724f
C4 VPB C 0.129699f
C5 VPB A 0.036002f
C6 a_1024_300# C 0.154435f
C7 a_1024_300# VPB 0.080675f
C8 X VGND 0.33712f
C9 C X 7.74e-19
C10 VPWR VGND 0.100395f
C11 VGND B 0.017405f
C12 VPB X 0.014365f
C13 VPWR C 0.012452f
C14 C B 3.4e-19
C15 VPWR A 0.013641f
C16 B A 0.063939f
C17 VPB VPWR 0.251605f
C18 VPB B 0.49412f
C19 a_1024_300# VPWR 0.018343f
C20 a_1024_300# B 0.017938f
C21 VPWR X 0.480563f
C22 X B 2.05e-19
C23 VPWR B 0.080509f
C24 VGND VNB 1.18496f
C25 X VNB 0.032001f
C26 C VNB 0.300353f
C27 VPWR VNB 0.94483f
C28 A VNB 0.107742f
C29 B VNB 0.411557f
C30 VPB VNB 2.33467f
C31 a_1024_300# VNB 0.140682f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor2_1 VNB VPB VPWR VGND A B X
X0 X.t1 B.t0 a_455_87.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 X.t0 a_194_125.t3 a_355_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_194_125.t1 B.t1 a_158_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t1 A.t0 a_355_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X4 a_158_392.t1 A.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5 a_355_368.t2 B.t2 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X6 a_194_125.t2 A.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.177375 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X7 a_455_87.t0 A.t3 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.126075 ps=1.1 w=0.74 l=0.15
X8 VGND.t1 B.t3 a_194_125.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.177375 ps=1.195 w=0.55 l=0.15
X9 VGND.t0 a_194_125.t4 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
R0 B.n0 B.t1 272.087
R1 B.n1 B.t2 250.909
R2 B.n1 B.t0 199.227
R3 B B.n0 194.862
R4 B.n0 B.t3 184.476
R5 B.n2 B.n1 152
R6 B B.n2 18.824
R7 B.n2 B 4.84898
R8 a_455_87.t0 a_455_87.t1 38.9194
R9 X.n0 X.t0 348.457
R10 X.n1 X.n0 185
R11 X.n2 X.n1 185
R12 X.n1 X.t2 45.4059
R13 X.n1 X.t1 22.7032
R14 X X.n2 7.47915
R15 X X.n0 4.17129
R16 X.n2 X 3.16454
R17 VNB VNB.t4 2067.19
R18 VNB.t4 VNB.t1 1836.22
R19 VNB.t2 VNB.t3 1316.54
R20 VNB.t1 VNB.t0 1177.95
R21 VNB.t0 VNB.t2 900.788
R22 a_194_125.n2 a_194_125.n0 299.346
R23 a_194_125.n0 a_194_125.t3 258.942
R24 a_194_125.t1 a_194_125.n2 230.556
R25 a_194_125.n0 a_194_125.t4 189.588
R26 a_194_125.n2 a_194_125.n1 152.939
R27 a_194_125.n1 a_194_125.t0 64.7431
R28 a_194_125.n1 a_194_125.t2 62.3121
R29 a_355_368.t0 a_355_368.n0 690.256
R30 a_355_368.n0 a_355_368.t2 35.1791
R31 a_355_368.n0 a_355_368.t1 26.3844
R32 VPB.t3 VPB.t0 536.29
R33 VPB VPB.t4 365.188
R34 VPB.t0 VPB.t2 291.13
R35 VPB.t2 VPB.t1 255.376
R36 VPB.t4 VPB.t3 214.517
R37 a_158_392.t0 a_158_392.t1 53.1905
R38 A.t2 A.t3 803.333
R39 A.t3 A.t0 484.947
R40 A.n0 A.t1 260.281
R41 A.n0 A.t2 173.228
R42 A A.n0 106.367
R43 VPWR.n1 VPWR.n0 605.418
R44 VPWR.n1 VPWR.t2 258.94
R45 VPWR.n0 VPWR.t1 37.8175
R46 VPWR.n0 VPWR.t0 36.0585
R47 VPWR VPWR.n1 0.153593
R48 VGND.n3 VGND.t0 281.322
R49 VGND.n7 VGND.t3 156.095
R50 VGND.n2 VGND.n1 123.984
R51 VGND.n1 VGND.t1 47.2956
R52 VGND.n6 VGND.n5 36.1417
R53 VGND.n7 VGND.n6 32.0005
R54 VGND.n1 VGND.t2 21.9347
R55 VGND.n5 VGND.n2 10.5417
R56 VGND.n6 VGND.n0 9.3005
R57 VGND.n5 VGND.n4 9.3005
R58 VGND.n3 VGND.n2 8.2678
R59 VGND.n8 VGND.n7 4.62059
R60 VGND.n4 VGND.n3 0.283861
R61 VGND.n8 VGND.n0 0.184273
R62 VGND VGND.n8 0.123049
R63 VGND.n4 VGND.n0 0.122949
C0 A VGND 0.148411f
C1 A VPWR 0.059856f
C2 A B 0.16657f
C3 VPB X 0.016429f
C4 VPWR X 0.047071f
C5 VGND X 0.152626f
C6 B X 0.040653f
C7 VGND VPB 0.010925f
C8 VPB VPWR 0.124002f
C9 B VPB 0.106329f
C10 VGND VPWR 0.064893f
C11 A X 0.004787f
C12 B VGND 0.059011f
C13 B VPWR 0.023003f
C14 A VPB 0.102444f
C15 VGND VNB 0.55128f
C16 X VNB 0.101097f
C17 VPWR VNB 0.425233f
C18 B VNB 0.236191f
C19 A VNB 0.480314f
C20 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor2_2 VNB VPB VPWR VGND A B X
X0 a_313_368.t5 A.t0 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1 a_399_74.t1 B.t0 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1794 pd=1.285 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_116_392.t1 A.t1 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X3 X.t1 B.t1 a_399_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1794 ps=1.285 w=0.74 l=0.15
X4 a_183_74.t2 A.t2 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.5031 ps=2.9 w=0.64 l=0.15
X5 VPWR.t3 A.t3 a_313_368.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 VGND.t4 A.t4 a_399_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.3156 pd=1.7 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VGND.t0 B.t2 a_183_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1725 pd=1.24 as=0.0896 ps=0.92 w=0.64 l=0.15
X8 a_183_74.t0 B.t3 a_116_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X9 a_313_368.t1 B.t4 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3416 pd=2.85 as=0.196 ps=1.47 w=1.12 l=0.15
X10 a_399_74.t2 A.t5 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1725 ps=1.24 w=0.74 l=0.15
X11 VPWR.t1 B.t5 a_313_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X12 X.t4 a_183_74.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3156 ps=1.7 w=0.74 l=0.15
X13 a_313_368.t0 a_183_74.t4 X.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 X.t3 a_183_74.t5 a_313_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n3 A.t1 324.986
R1 A.n1 A.t0 239.224
R2 A.n0 A.t3 226.809
R3 A.n0 A.t5 198.204
R4 A.n1 A.t4 196.013
R5 A.n3 A.t2 165.78
R6 A A.n3 161.697
R7 A A.n2 147.359
R8 A.n2 A.n0 31.7185
R9 A.n2 A.n1 22.1151
R10 VPWR.n5 VPWR.n2 617.774
R11 VPWR.n4 VPWR.n3 605.17
R12 VPWR.n10 VPWR.t2 345.382
R13 VPWR.n8 VPWR.n1 36.1417
R14 VPWR.n9 VPWR.n8 36.1417
R15 VPWR.n3 VPWR.t4 35.1791
R16 VPWR.n2 VPWR.t0 35.1791
R17 VPWR.n3 VPWR.t3 26.3844
R18 VPWR.n2 VPWR.t1 26.3844
R19 VPWR.n4 VPWR.n1 23.7181
R20 VPWR.n10 VPWR.n9 20.7064
R21 VPWR.n6 VPWR.n1 9.3005
R22 VPWR.n8 VPWR.n7 9.3005
R23 VPWR.n9 VPWR.n0 9.3005
R24 VPWR.n11 VPWR.n10 9.3005
R25 VPWR.n5 VPWR.n4 7.13405
R26 VPWR.n6 VPWR.n5 0.171369
R27 VPWR.n7 VPWR.n6 0.122949
R28 VPWR.n7 VPWR.n0 0.122949
R29 VPWR.n11 VPWR.n0 0.122949
R30 VPWR VPWR.n11 0.0617245
R31 a_313_368.t4 a_313_368.n3 389.913
R32 a_313_368.n1 a_313_368.t1 387.295
R33 a_313_368.n3 a_313_368.n2 289.146
R34 a_313_368.n1 a_313_368.n0 286.457
R35 a_313_368.n3 a_313_368.n1 76.5049
R36 a_313_368.n2 a_313_368.t3 26.3844
R37 a_313_368.n2 a_313_368.t5 26.3844
R38 a_313_368.n0 a_313_368.t2 26.3844
R39 a_313_368.n0 a_313_368.t0 26.3844
R40 VPB.t1 VPB.t5 515.861
R41 VPB VPB.t6 257.93
R42 VPB.t3 VPB.t2 255.376
R43 VPB.t5 VPB.t7 255.376
R44 VPB.t0 VPB.t3 229.839
R45 VPB.t4 VPB.t0 229.839
R46 VPB.t7 VPB.t4 229.839
R47 VPB.t6 VPB.t1 214.517
R48 B.n3 B.t3 398.454
R49 B B.n3 310.67
R50 B.n0 B.t4 261.62
R51 B.n1 B.t5 261.62
R52 B.n1 B.t0 165.196
R53 B B.n2 163.023
R54 B.n3 B.t2 162.274
R55 B.n0 B.t1 156.781
R56 B.n2 B.n0 44.549
R57 B.n2 B.n1 28.4823
R58 X X.n0 410.01
R59 X.n4 X.t1 279.738
R60 X.t1 X.n3 279.738
R61 X.n2 X.n1 245.951
R62 X.n0 X.t2 26.3844
R63 X.n0 X.t3 26.3844
R64 X.n1 X.t0 22.7032
R65 X.n1 X.t4 22.7032
R66 X X.n4 9.50353
R67 X.n3 X.n2 9.30959
R68 X.n4 X 4.84898
R69 X.n2 X 3.29747
R70 X.n3 X 1.74595
R71 a_399_74.n1 a_399_74.n0 517.332
R72 a_399_74.n1 a_399_74.t0 36.487
R73 a_399_74.t1 a_399_74.n1 35.6762
R74 a_399_74.n0 a_399_74.t3 22.7032
R75 a_399_74.n0 a_399_74.t2 22.7032
R76 VNB.t5 VNB.t3 2148.03
R77 VNB VNB.t6 1940.16
R78 VNB.t0 VNB.t4 1501.31
R79 VNB.t2 VNB.t1 1374.28
R80 VNB.t3 VNB.t2 993.177
R81 VNB.t4 VNB.t5 993.177
R82 VNB.t6 VNB.t0 993.177
R83 a_116_392.t0 a_116_392.t1 53.1905
R84 VGND.n8 VGND.t2 259.13
R85 VGND.n2 VGND.n1 208.079
R86 VGND.n4 VGND.n3 205.089
R87 VGND.n3 VGND.t1 90.0005
R88 VGND.n1 VGND.t3 50.7861
R89 VGND.n1 VGND.t0 39.3755
R90 VGND.n3 VGND.t4 36.487
R91 VGND.n7 VGND.n6 36.1417
R92 VGND.n6 VGND.n2 14.3064
R93 VGND.n9 VGND.n8 13.0202
R94 VGND.n7 VGND.n0 9.3005
R95 VGND.n6 VGND.n5 9.3005
R96 VGND.n8 VGND.n7 7.31754
R97 VGND.n4 VGND.n2 7.25585
R98 VGND.n5 VGND.n4 0.4354
R99 VGND.n5 VGND.n0 0.122949
R100 VGND.n9 VGND.n0 0.122949
R101 VGND VGND.n9 0.0617245
R102 a_183_74.n3 a_183_74.n0 371.147
R103 a_183_74.n3 a_183_74.n2 290.005
R104 a_183_74.t0 a_183_74.n3 238.192
R105 a_183_74.n2 a_183_74.t5 237.762
R106 a_183_74.n1 a_183_74.t4 234.841
R107 a_183_74.n1 a_183_74.t3 196.013
R108 a_183_74.n2 a_183_74.n1 46.7399
R109 a_183_74.n0 a_183_74.t1 26.2505
R110 a_183_74.n0 a_183_74.t2 26.2505
C0 B X 0.221546f
C1 X VPB 0.010158f
C2 B VPB 0.131453f
C3 VPWR VGND 0.081126f
C4 VGND A 0.044536f
C5 VPWR A 0.051815f
C6 X VGND 0.0573f
C7 VPWR X 0.019053f
C8 B VGND 0.093076f
C9 X A 0.001228f
C10 B VPWR 0.049427f
C11 VGND VPB 0.009237f
C12 VPWR VPB 0.135999f
C13 B A 0.267476f
C14 VPB A 0.118962f
C15 VGND VNB 0.575244f
C16 X VNB 0.085376f
C17 VPWR VNB 0.489772f
C18 B VNB 0.399817f
C19 A VNB 0.384715f
C20 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor2_4 VNB VPB VPWR VGND A B X
X0 VGND.t5 A.t0 a_877_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1889 pd=1.36 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VPWR.t3 A.t1 a_514_368.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.270175 pd=1.785 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_160_98.t3 B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.20775 ps=1.49 w=0.74 l=0.15
X3 VGND.t8 B.t1 a_160_98.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.20775 pd=1.49 as=0.1443 ps=1.13 w=0.74 l=0.15
X4 a_877_74.t5 B.t2 X.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_514_368.t5 A.t2 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.27695 ps=1.795 w=1.12 l=0.15
X6 VPWR.t1 A.t3 a_514_368.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.27695 pd=1.795 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_514_368.t0 a_160_98.t6 X.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_877_74.t3 A.t4 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1889 ps=1.36 w=0.74 l=0.15
X9 X.t5 a_160_98.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.20905 pd=1.305 as=0.20775 ps=1.49 w=0.74 l=0.15
X10 X.t2 a_160_98.t8 a_514_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_514_368.t2 a_160_98.t9 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 X.t0 a_160_98.t10 a_514_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X13 a_514_368.t8 B.t3 VPWR.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR.t7 B.t4 a_514_368.t9 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_514_368.t10 B.t5 VPWR.t8 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VPWR.t9 B.t6 a_514_368.t11 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_514_368.t7 A.t5 VPWR.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.270175 ps=1.785 w=1.12 l=0.15
X18 VGND.t9 a_160_98.t11 X.t4 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.44175 pd=2.96 as=0.20905 ps=1.305 w=0.74 l=0.15
X19 a_877_74.t6 B.t7 X.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t5 A.t6 a_36_392.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X21 a_160_98.t1 A.t7 VGND.t7 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3811 ps=2.51 w=0.74 l=0.15
X22 VGND.t3 A.t8 a_877_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1889 pd=1.36 as=0.2109 ps=2.05 w=0.74 l=0.15
X23 X.t7 B.t8 a_877_74.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X24 a_877_74.t1 A.t9 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1889 ps=1.36 w=0.74 l=0.15
X25 a_36_392.t3 B.t9 a_160_98.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X26 a_160_98.t4 B.t10 a_36_392.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X27 VGND.t6 A.t10 a_160_98.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.20775 pd=1.49 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 X.t6 B.t11 a_877_74.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 a_36_392.t0 A.t11 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
R0 A A.n10 334.433
R1 A.n0 A.t5 242.875
R2 A.n5 A.t3 229.73
R3 A.n9 A.t6 228.951
R4 A.n1 A.t1 226.809
R5 A.n4 A.t2 226.809
R6 A.n6 A.t11 220.917
R7 A.n6 A.t10 200.589
R8 A.n0 A.t4 197.799
R9 A.n1 A.t0 196.013
R10 A.n5 A.t8 196.013
R11 A.n3 A.t9 196.013
R12 A.n8 A.t7 179.947
R13 A.n10 A.n7 165.189
R14 A A.n2 152.452
R15 A.n10 A.n9 152
R16 A.n12 A.n11 152
R17 A.n14 A.n13 152
R18 A.n1 A.n0 100.621
R19 A.n13 A.n12 49.6611
R20 A.n2 A.n1 46.0096
R21 A.n8 A.n7 32.1338
R22 A.n13 A.n4 29.9429
R23 A.n9 A.n8 17.5278
R24 A.n3 A.n2 16.7975
R25 A.n7 A.n6 15.3369
R26 A A.n14 9.78874
R27 A.n11 A 8.88521
R28 A.n11 A 5.57226
R29 A.n14 A 4.66874
R30 A.n12 A.n5 3.65202
R31 A.n4 A.n3 2.92171
R32 a_877_74.n4 a_877_74.t2 268.276
R33 a_877_74.n1 a_877_74.t6 260.603
R34 a_877_74.n1 a_877_74.n0 197.994
R35 a_877_74.n3 a_877_74.n2 185
R36 a_877_74.n5 a_877_74.n4 185
R37 a_877_74.n3 a_877_74.n1 68.3525
R38 a_877_74.n4 a_877_74.n3 60.3596
R39 a_877_74.n0 a_877_74.t5 34.0546
R40 a_877_74.n2 a_877_74.t4 22.7032
R41 a_877_74.n2 a_877_74.t3 22.7032
R42 a_877_74.n0 a_877_74.t7 22.7032
R43 a_877_74.t0 a_877_74.n5 22.7032
R44 a_877_74.n5 a_877_74.t1 22.7032
R45 VGND.n14 VGND.t9 330.067
R46 VGND.n19 VGND.n5 262.132
R47 VGND.n2 VGND.n1 253.276
R48 VGND.n10 VGND.n9 218.101
R49 VGND.n8 VGND.n7 212.477
R50 VGND.n26 VGND.t7 193.679
R51 VGND.n15 VGND.n4 36.1417
R52 VGND.n21 VGND.n20 36.1417
R53 VGND.n25 VGND.n24 36.1417
R54 VGND.n1 VGND.t1 35.6762
R55 VGND.n1 VGND.t6 35.6762
R56 VGND.n9 VGND.t4 35.6762
R57 VGND.n9 VGND.t5 35.6762
R58 VGND.n7 VGND.t2 35.6762
R59 VGND.n7 VGND.t3 35.6762
R60 VGND.n5 VGND.t0 35.6762
R61 VGND.n5 VGND.t8 35.6762
R62 VGND.n13 VGND.n12 33.1837
R63 VGND.n19 VGND.n4 28.2358
R64 VGND.n26 VGND.n25 28.2358
R65 VGND.n12 VGND.n8 23.7181
R66 VGND.n20 VGND.n19 19.2005
R67 VGND.n15 VGND.n14 13.4459
R68 VGND.n24 VGND.n2 10.6672
R69 VGND.n27 VGND.n26 9.3005
R70 VGND.n12 VGND.n11 9.3005
R71 VGND.n13 VGND.n6 9.3005
R72 VGND.n16 VGND.n15 9.3005
R73 VGND.n17 VGND.n4 9.3005
R74 VGND.n19 VGND.n18 9.3005
R75 VGND.n20 VGND.n3 9.3005
R76 VGND.n22 VGND.n21 9.3005
R77 VGND.n24 VGND.n23 9.3005
R78 VGND.n25 VGND.n0 9.3005
R79 VGND.n21 VGND.n2 9.16128
R80 VGND.n10 VGND.n8 6.79999
R81 VGND.n14 VGND.n13 3.33495
R82 VGND.n11 VGND.n10 0.48894
R83 VGND.n11 VGND.n6 0.122949
R84 VGND.n16 VGND.n6 0.122949
R85 VGND.n17 VGND.n16 0.122949
R86 VGND.n18 VGND.n17 0.122949
R87 VGND.n18 VGND.n3 0.122949
R88 VGND.n22 VGND.n3 0.122949
R89 VGND.n23 VGND.n22 0.122949
R90 VGND.n23 VGND.n0 0.122949
R91 VGND.n27 VGND.n0 0.122949
R92 VGND VGND.n27 0.0617245
R93 VNB.t13 VNB.t4 2667.72
R94 VNB VNB.t5 1674.54
R95 VNB.t0 VNB.t13 1651.44
R96 VNB.t7 VNB.t6 1362.73
R97 VNB.t4 VNB.t3 1362.73
R98 VNB.t10 VNB.t0 1362.73
R99 VNB.t2 VNB.t1 1362.73
R100 VNB.t1 VNB.t10 1247.24
R101 VNB.t9 VNB.t12 1154.86
R102 VNB.t12 VNB.t11 993.177
R103 VNB.t8 VNB.t9 993.177
R104 VNB.t6 VNB.t8 993.177
R105 VNB.t3 VNB.t7 993.177
R106 VNB.t5 VNB.t2 993.177
R107 a_514_368.n1 a_514_368.n0 592.907
R108 a_514_368.n7 a_514_368.n6 585
R109 a_514_368.n9 a_514_368.n8 585
R110 a_514_368.n1 a_514_368.t3 394.981
R111 a_514_368.n4 a_514_368.t8 368.354
R112 a_514_368.n4 a_514_368.n3 299.053
R113 a_514_368.n5 a_514_368.n2 289.803
R114 a_514_368.n7 a_514_368.n5 77.2342
R115 a_514_368.n8 a_514_368.n1 71.0932
R116 a_514_368.n8 a_514_368.n7 64.0166
R117 a_514_368.n5 a_514_368.n4 61.4809
R118 a_514_368.n0 a_514_368.t1 26.3844
R119 a_514_368.n0 a_514_368.t2 26.3844
R120 a_514_368.n6 a_514_368.t6 26.3844
R121 a_514_368.n6 a_514_368.t5 26.3844
R122 a_514_368.n3 a_514_368.t9 26.3844
R123 a_514_368.n3 a_514_368.t10 26.3844
R124 a_514_368.n2 a_514_368.t11 26.3844
R125 a_514_368.n2 a_514_368.t7 26.3844
R126 a_514_368.n9 a_514_368.t4 26.3844
R127 a_514_368.t0 a_514_368.n9 26.3844
R128 VPWR.n12 VPWR.n11 655.92
R129 VPWR.n20 VPWR.n19 653.192
R130 VPWR.n8 VPWR.n7 624.564
R131 VPWR.n10 VPWR.n9 611.88
R132 VPWR.n33 VPWR.n1 323.777
R133 VPWR.n1 VPWR.t4 39.4005
R134 VPWR.n19 VPWR.t2 38.6969
R135 VPWR.n19 VPWR.t1 38.6969
R136 VPWR.n11 VPWR.t0 37.8175
R137 VPWR.n11 VPWR.t3 37.8175
R138 VPWR.n21 VPWR.n4 36.1417
R139 VPWR.n25 VPWR.n4 36.1417
R140 VPWR.n26 VPWR.n25 36.1417
R141 VPWR.n27 VPWR.n26 36.1417
R142 VPWR.n27 VPWR.n2 36.1417
R143 VPWR.n31 VPWR.n2 36.1417
R144 VPWR.n32 VPWR.n31 36.1417
R145 VPWR.n17 VPWR.n6 30.9882
R146 VPWR.n1 VPWR.t5 29.5505
R147 VPWR.n18 VPWR.n17 29.3485
R148 VPWR.n13 VPWR.n10 28.2358
R149 VPWR.n21 VPWR.n20 26.9056
R150 VPWR.n7 VPWR.t6 26.3844
R151 VPWR.n7 VPWR.t7 26.3844
R152 VPWR.n9 VPWR.t8 26.3844
R153 VPWR.n9 VPWR.t9 26.3844
R154 VPWR.n13 VPWR.n12 24.2703
R155 VPWR.n33 VPWR.n32 19.577
R156 VPWR.n14 VPWR.n13 9.3005
R157 VPWR.n15 VPWR.n6 9.3005
R158 VPWR.n17 VPWR.n16 9.3005
R159 VPWR.n18 VPWR.n5 9.3005
R160 VPWR.n22 VPWR.n21 9.3005
R161 VPWR.n23 VPWR.n4 9.3005
R162 VPWR.n25 VPWR.n24 9.3005
R163 VPWR.n26 VPWR.n3 9.3005
R164 VPWR.n28 VPWR.n27 9.3005
R165 VPWR.n29 VPWR.n2 9.3005
R166 VPWR.n31 VPWR.n30 9.3005
R167 VPWR.n32 VPWR.n0 9.3005
R168 VPWR.n34 VPWR.n33 7.63521
R169 VPWR.n10 VPWR.n8 6.92957
R170 VPWR.n12 VPWR.n6 1.56494
R171 VPWR.n20 VPWR.n18 0.569389
R172 VPWR.n14 VPWR.n8 0.451354
R173 VPWR VPWR.n34 0.162741
R174 VPWR.n34 VPWR.n0 0.145097
R175 VPWR.n15 VPWR.n14 0.122949
R176 VPWR.n16 VPWR.n15 0.122949
R177 VPWR.n16 VPWR.n5 0.122949
R178 VPWR.n22 VPWR.n5 0.122949
R179 VPWR.n23 VPWR.n22 0.122949
R180 VPWR.n24 VPWR.n23 0.122949
R181 VPWR.n24 VPWR.n3 0.122949
R182 VPWR.n28 VPWR.n3 0.122949
R183 VPWR.n29 VPWR.n28 0.122949
R184 VPWR.n30 VPWR.n29 0.122949
R185 VPWR.n30 VPWR.n0 0.122949
R186 VPB.t10 VPB.t3 497.985
R187 VPB.t7 VPB.t8 301.344
R188 VPB.t9 VPB.t6 296.238
R189 VPB VPB.t5 280.914
R190 VPB.t5 VPB.t4 255.376
R191 VPB.t13 VPB.t12 229.839
R192 VPB.t14 VPB.t13 229.839
R193 VPB.t15 VPB.t14 229.839
R194 VPB.t6 VPB.t15 229.839
R195 VPB.t8 VPB.t9 229.839
R196 VPB.t0 VPB.t7 229.839
R197 VPB.t1 VPB.t0 229.839
R198 VPB.t2 VPB.t1 229.839
R199 VPB.t3 VPB.t2 229.839
R200 VPB.t11 VPB.t10 229.839
R201 VPB.t4 VPB.t11 229.839
R202 B.t11 B.t6 502.351
R203 B.n8 B.n7 438.829
R204 B.t2 B.t11 424.161
R205 B.n5 B.t10 247.746
R206 B.n0 B.t3 226.809
R207 B.n3 B.t4 226.809
R208 B.n4 B.t5 226.809
R209 B.n7 B.t1 207.582
R210 B.n0 B.t7 196.013
R211 B.n2 B.t8 196.013
R212 B.n5 B.t0 196.013
R213 B.n6 B.t9 195.478
R214 B.n4 B.t2 193.822
R215 B B.n1 156.912
R216 B.n12 B.n11 152
R217 B.n10 B.n9 152
R218 B.n11 B.n10 49.6611
R219 B.n2 B.n1 41.6278
R220 B.n7 B.n6 31.4912
R221 B.n6 B.n5 28.8904
R222 B.n1 B.n0 21.1793
R223 B B.n8 13.9585
R224 B.n9 B 13.247
R225 B.n10 B.n4 10.955
R226 B.n12 B 9.07957
R227 B B.n12 5.2098
R228 B.n11 B.n3 5.11262
R229 B.n3 B.n2 2.92171
R230 B.n9 B 1.04236
R231 B.n8 B 0.327293
R232 a_160_98.n2 a_160_98.t6 352.111
R233 a_160_98.n12 a_160_98.n0 345.183
R234 a_160_98.n5 a_160_98.t9 226.809
R235 a_160_98.n7 a_160_98.t10 226.809
R236 a_160_98.n13 a_160_98.n12 223.144
R237 a_160_98.n2 a_160_98.t8 204.048
R238 a_160_98.n11 a_160_98.n10 185
R239 a_160_98.n9 a_160_98.n8 170.258
R240 a_160_98.n4 a_160_98.n1 165.601
R241 a_160_98.n8 a_160_98.t7 157.453
R242 a_160_98.n3 a_160_98.t11 157.453
R243 a_160_98.n6 a_160_98.n1 152
R244 a_160_98.n3 a_160_98.n2 51.908
R245 a_160_98.n11 a_160_98.n9 48.9205
R246 a_160_98.n6 a_160_98.n5 41.6278
R247 a_160_98.n10 a_160_98.t2 31.6221
R248 a_160_98.n10 a_160_98.t3 31.6221
R249 a_160_98.n0 a_160_98.t5 29.5505
R250 a_160_98.n0 a_160_98.t4 29.5505
R251 a_160_98.n7 a_160_98.n6 24.1005
R252 a_160_98.n4 a_160_98.n3 23.3702
R253 a_160_98.n13 a_160_98.t0 22.7032
R254 a_160_98.t1 a_160_98.n13 22.7032
R255 a_160_98.n12 a_160_98.n11 16.8965
R256 a_160_98.n9 a_160_98.n1 13.6005
R257 a_160_98.n5 a_160_98.n4 8.03383
R258 a_160_98.n8 a_160_98.n7 7.30353
R259 X.n6 X.n5 585
R260 X.n3 X.n1 450.7
R261 X.n6 X.n4 428.599
R262 X X.n7 342.173
R263 X.n4 X.n0 200.435
R264 X.n3 X.n2 197.994
R265 X.n1 X.t5 68.9194
R266 X.n4 X.n3 57.6005
R267 X.n5 X.t3 26.3844
R268 X.n5 X.t2 26.3844
R269 X.n7 X.t1 26.3844
R270 X.n7 X.t0 26.3844
R271 X.n1 X.t4 22.7032
R272 X.n2 X.t9 22.7032
R273 X.n2 X.t6 22.7032
R274 X.n0 X.t8 22.7032
R275 X.n0 X.t7 22.7032
R276 X X.n6 1.56494
R277 a_36_392.n1 a_36_392.t3 408.764
R278 a_36_392.t1 a_36_392.n1 305.349
R279 a_36_392.n1 a_36_392.n0 187.186
R280 a_36_392.n0 a_36_392.t2 29.5505
R281 a_36_392.n0 a_36_392.t0 29.5505
C0 VGND VPWR 0.13974f
C1 VGND B 0.056654f
C2 X VGND 0.147364f
C3 B VPWR 0.099205f
C4 VGND VPB 0.013448f
C5 X VPWR 0.0772f
C6 VPB VPWR 0.207848f
C7 VGND A 0.329884f
C8 X B 0.768863f
C9 B VPB 0.245369f
C10 A VPWR 0.079829f
C11 X VPB 0.008048f
C12 A B 0.370069f
C13 X A 0.322025f
C14 A VPB 0.244733f
C15 VGND VNB 1.03463f
C16 X VNB 0.09172f
C17 B VNB 0.671421f
C18 A VNB 0.717643f
C19 VPWR VNB 0.782249f
C20 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor3_1 VNB VPB VPWR VGND B C A X
X0 a_84_108.t0 A.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1702 pd=1.41 as=0.34745 ps=1.81 w=0.64 l=0.15
X1 X.t1 a_1215_396# VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2436 ps=1.66 w=1.12 l=0.15
X2 a_27_134.t5 a_452_288.t2 a_384_392.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1024 pd=0.96 as=0.1401 ps=1.195 w=0.64 l=0.15
X3 a_84_108.t2 a_452_288.t3 a_384_392.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2848 pd=2.17 as=0.169075 ps=1.275 w=0.64 l=0.15
X4 X.t0 a_1215_396# VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1212 ps=1.1 w=0.74 l=0.15
X5 a_384_392.t5 B.t0 a_84_108.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1401 pd=1.195 as=0.1837 ps=1.385 w=0.84 l=0.15
X6 a_84_108.t1 A.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1837 pd=1.385 as=0.25 ps=1.5 w=1 l=0.15
X7 VPWR.t1 a_84_108.t6 a_27_134.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.295 ps=2.59 w=1 l=0.15
X8 a_27_134.t4 a_452_288.t4 a_416_86# VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.15815 pd=1.16 as=0.10375 ps=0.99 w=0.42 l=0.15
X9 VPWR.t2 C.t0 a_1157_298.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=1.66 as=0.2528 ps=2.07 w=0.64 l=0.15
X10 a_416_86# C.t1 a_1215_396# VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.24 pd=2.03 as=0.1696 ps=1.17 w=0.64 l=0.15
X11 a_384_392.t4 C.t2 a_1215_396# VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2982 pd=2.39 as=0.2541 ps=1.445 w=0.84 l=0.15
X12 a_416_86# B.t1 a_84_108.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.10375 pd=0.99 as=0.1702 ps=1.41 w=0.64 l=0.15
X13 a_1215_396# a_1157_298.t2 a_384_392.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.17 as=0.176 ps=1.83 w=0.64 l=0.15
X14 VGND.t0 B.t2 a_452_288.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3885 pd=2.53 as=0.2035 ps=2.03 w=0.74 l=0.15
X15 a_84_108.t3 a_452_288.t5 a_416_86# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.5082 pd=2.89 as=0.150675 ps=1.225 w=0.84 l=0.15
X16 a_416_86# B.t3 a_27_134.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.150675 pd=1.225 as=0.1024 ps=0.96 w=0.64 l=0.15
X17 a_384_392.t1 B.t4 a_27_134.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.169075 pd=1.275 as=0.15815 ps=1.16 w=0.64 l=0.15
X18 VGND.t4 C.t3 a_1157_298.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.1197 ps=1.41 w=0.42 l=0.15
X19 VGND.t2 a_84_108.t7 a_27_134.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.34745 pd=1.81 as=0.1824 ps=1.85 w=0.64 l=0.15
X20 VPWR.t4 B.t5 a_452_288.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 A.n0 A.t1 238.993
R1 A A.n0 166.769
R2 A.n0 A.t0 156.249
R3 VGND.n11 VGND.t0 274.611
R4 VGND.n1 VGND.n0 263.113
R5 VGND.n9 VGND.n6 202.456
R6 VGND.n9 VGND.n8 185
R7 VGND.n0 VGND.t1 63.7505
R8 VGND.n0 VGND.t2 63.7505
R9 VGND.n7 VGND.t4 61.4291
R10 VGND.t3 VGND.n6 52.5005
R11 VGND.n8 VGND.t3 40.0005
R12 VGND.n12 VGND.n5 36.1417
R13 VGND.n16 VGND.n5 36.1417
R14 VGND.n17 VGND.n16 36.1417
R15 VGND.n18 VGND.n17 36.1417
R16 VGND.n18 VGND.n3 36.1417
R17 VGND.n22 VGND.n3 36.1417
R18 VGND.n23 VGND.n22 36.1417
R19 VGND.n24 VGND.n23 36.1417
R20 VGND.n10 VGND.n9 28.475
R21 VGND.n12 VGND.n11 20.7064
R22 VGND.n26 VGND.n1 11.7718
R23 VGND.n25 VGND.n24 9.3005
R24 VGND.n23 VGND.n2 9.3005
R25 VGND.n22 VGND.n21 9.3005
R26 VGND.n20 VGND.n3 9.3005
R27 VGND.n19 VGND.n18 9.3005
R28 VGND.n17 VGND.n4 9.3005
R29 VGND.n16 VGND.n15 9.3005
R30 VGND.n14 VGND.n5 9.3005
R31 VGND.n13 VGND.n12 9.3005
R32 VGND.n11 VGND.n10 7.53798
R33 VGND.n24 VGND.n1 6.72132
R34 VGND.n7 VGND.n6 1.8755
R35 VGND.n8 VGND.n7 1.42907
R36 VGND VGND.n26 0.161517
R37 VGND.n13 VGND.n10 0.151527
R38 VGND.n26 VGND.n25 0.146304
R39 VGND.n14 VGND.n13 0.122949
R40 VGND.n15 VGND.n14 0.122949
R41 VGND.n15 VGND.n4 0.122949
R42 VGND.n19 VGND.n4 0.122949
R43 VGND.n20 VGND.n19 0.122949
R44 VGND.n21 VGND.n20 0.122949
R45 VGND.n21 VGND.n2 0.122949
R46 VGND.n25 VGND.n2 0.122949
R47 a_84_108.n8 a_84_108.n7 600.562
R48 a_84_108.n1 a_84_108.t3 379.158
R49 a_84_108.n1 a_84_108.t2 305.791
R50 a_84_108.n6 a_84_108.n5 288.053
R51 a_84_108.n7 a_84_108.n1 261.017
R52 a_84_108.n4 a_84_108.n3 246.114
R53 a_84_108.n2 a_84_108.t6 231.629
R54 a_84_108.n4 a_84_108.n2 213.256
R55 a_84_108.n2 a_84_108.t7 178.34
R56 a_84_108.n3 a_84_108.t5 102.939
R57 a_84_108.n5 a_84_108.t4 55.1136
R58 a_84_108.n9 a_84_108.n8 46.5641
R59 a_84_108.n0 a_84_108.t1 28.0191
R60 a_84_108.n3 a_84_108.t0 26.2505
R61 a_84_108.n6 a_84_108.n4 13.9185
R62 a_84_108.n7 a_84_108.n6 10.9067
R63 a_84_108.n8 a_84_108.n0 10.746
R64 a_84_108.n5 a_84_108.n0 3.51836
R65 VNB.t1 VNB.t10 2956.43
R66 VNB.t2 VNB.t0 2817.85
R67 VNB.t5 VNB.t2 2702.36
R68 VNB.t4 VNB.t3 1917.06
R69 VNB.t0 VNB.t1 1570.6
R70 VNB.t3 VNB.t9 1570.6
R71 VNB.t6 VNB.t7 1547.51
R72 VNB.t7 VNB.t5 1362.73
R73 VNB.t10 VNB.t8 1177.95
R74 VNB.t9 VNB.t6 1154.86
R75 VNB VNB.t4 1143.31
R76 VPWR.n20 VPWR.n1 316.209
R77 VPWR.n7 VPWR.t4 257.433
R78 VPWR.n6 VPWR.n5 249.149
R79 VPWR.n5 VPWR.t2 120.047
R80 VPWR.n1 VPWR.t0 59.1005
R81 VPWR.n1 VPWR.t1 39.4005
R82 VPWR.n8 VPWR.n4 36.1417
R83 VPWR.n12 VPWR.n4 36.1417
R84 VPWR.n13 VPWR.n12 36.1417
R85 VPWR.n14 VPWR.n13 36.1417
R86 VPWR.n14 VPWR.n2 36.1417
R87 VPWR.n18 VPWR.n2 36.1417
R88 VPWR.n19 VPWR.n18 36.1417
R89 VPWR.n8 VPWR.n7 29.3652
R90 VPWR.n5 VPWR.t3 25.8278
R91 VPWR.n21 VPWR.n20 11.4685
R92 VPWR.n9 VPWR.n8 9.3005
R93 VPWR.n10 VPWR.n4 9.3005
R94 VPWR.n12 VPWR.n11 9.3005
R95 VPWR.n13 VPWR.n3 9.3005
R96 VPWR.n15 VPWR.n14 9.3005
R97 VPWR.n16 VPWR.n2 9.3005
R98 VPWR.n18 VPWR.n17 9.3005
R99 VPWR.n19 VPWR.n0 9.3005
R100 VPWR.n20 VPWR.n19 7.52991
R101 VPWR.n7 VPWR.n6 7.16768
R102 VPWR VPWR.n21 0.163644
R103 VPWR.n9 VPWR.n6 0.157145
R104 VPWR.n21 VPWR.n0 0.144205
R105 VPWR.n10 VPWR.n9 0.122949
R106 VPWR.n11 VPWR.n10 0.122949
R107 VPWR.n11 VPWR.n3 0.122949
R108 VPWR.n15 VPWR.n3 0.122949
R109 VPWR.n16 VPWR.n15 0.122949
R110 VPWR.n17 VPWR.n16 0.122949
R111 VPWR.n17 VPWR.n0 0.122949
R112 X.n3 X 591.4
R113 X.n3 X.n0 585
R114 X.n4 X.n3 585
R115 X.n2 X.t0 279.738
R116 X.t0 X.n1 279.738
R117 X.n3 X.t1 26.3844
R118 X X.n4 17.1525
R119 X X.n0 14.8485
R120 X.n1 X 14.0805
R121 X X.n2 9.9845
R122 X.n2 X 8.9605
R123 X.n1 X 4.8645
R124 X X.n0 4.0965
R125 X.n4 X 1.7925
R126 VPB.t9 VPB.t7 952.554
R127 VPB.t5 VPB.t9 784.005
R128 VPB.t7 VPB.t3 597.582
R129 VPB.t3 VPB.t6 352.42
R130 VPB VPB.t2 337.098
R131 VPB.t2 VPB.t1 331.99
R132 VPB.t0 VPB.t5 273.253
R133 VPB.t1 VPB.t8 273.253
R134 VPB.t8 VPB.t4 257.93
R135 VPB.t4 VPB.t0 240.054
R136 a_452_288.t1 a_452_288.n3 317.659
R137 a_452_288.n3 a_452_288.n2 294.158
R138 a_452_288.n0 a_452_288.t2 255.728
R139 a_452_288.n1 a_452_288.n0 244.214
R140 a_452_288.n1 a_452_288.t5 240.732
R141 a_452_288.n3 a_452_288.t0 207.703
R142 a_452_288.n0 a_452_288.t4 186.374
R143 a_452_288.n2 a_452_288.t3 147.814
R144 a_452_288.n2 a_452_288.n1 89.6817
R145 a_384_392.t4 a_384_392.n5 626.707
R146 a_384_392.n1 a_384_392.n0 503.325
R147 a_384_392.n5 a_384_392.n4 223.76
R148 a_384_392.n5 a_384_392.t0 211.25
R149 a_384_392.n4 a_384_392.n3 209.615
R150 a_384_392.n2 a_384_392.n1 206.538
R151 a_384_392.n0 a_384_392.t3 55.4067
R152 a_384_392.n0 a_384_392.t5 46.0016
R153 a_384_392.n4 a_384_392.n1 41.0358
R154 a_384_392.n2 a_384_392.t2 34.688
R155 a_384_392.n3 a_384_392.t1 33.7505
R156 a_384_392.n3 a_384_392.n2 20.2252
R157 a_27_134.n2 a_27_134.n0 618.359
R158 a_27_134.t2 a_27_134.n3 411.851
R159 a_27_134.n2 a_27_134.n1 212.421
R160 a_27_134.n3 a_27_134.n2 190.279
R161 a_27_134.n3 a_27_134.t1 125.329
R162 a_27_134.n1 a_27_134.t3 62.813
R163 a_27_134.n0 a_27_134.t5 52.3286
R164 a_27_134.n0 a_27_134.t0 46.1724
R165 a_27_134.n1 a_27_134.t4 42.0541
R166 B.n2 B.n1 996.134
R167 B.n2 B.n0 756.74
R168 B.n0 B.t1 535.02
R169 B.n1 B.t0 488.159
R170 B.n1 B.t3 254.121
R171 B.n4 B.t5 244.482
R172 B.n3 B.t2 204.048
R173 B.n0 B.t4 159.06
R174 B B.n4 155.87
R175 B.n3 B.n2 117.287
R176 B.n4 B.n3 9.6405
R177 C.n1 C.t2 290.272
R178 C.n2 C.n0 270.724
R179 C.n0 C.t3 250.641
R180 C.n0 C.t0 203.244
R181 C.n1 C.t1 177.001
R182 C C.n2 164.024
R183 C.n2 C.n1 16.0672
R184 a_1157_298.t1 a_1157_298.n2 646.562
R185 a_1157_298.n2 a_1157_298.n1 378.928
R186 a_1157_298.n2 a_1157_298.t0 346.991
R187 a_1157_298.n1 a_1157_298.n0 199.694
R188 a_1157_298.n1 a_1157_298.t2 199.425
C0 VPWR VPB 0.224347f
C1 B A 0.011285f
C2 a_416_86# VPB 0.036474f
C3 a_416_86# VPWR 0.195269f
C4 a_1215_396# B 0.001263f
C5 B VGND 0.078836f
C6 a_1215_396# X 0.056611f
C7 VGND X 0.091329f
C8 B VPB 0.506832f
C9 X VPB 0.012381f
C10 B VPWR 0.126187f
C11 VPWR X 0.111185f
C12 a_416_86# B 0.123484f
C13 a_1215_396# C 0.133084f
C14 VGND C 0.025182f
C15 C VPB 0.130819f
C16 VGND A 0.013726f
C17 B X 1.51e-19
C18 VPWR C 0.00904f
C19 VPB A 0.052079f
C20 a_1215_396# VGND 0.124016f
C21 a_416_86# C 0.039963f
C22 VPWR A 0.017364f
C23 a_1215_396# VPB 0.066707f
C24 a_416_86# A 8.23e-19
C25 VGND VPB 0.010188f
C26 a_1215_396# VPWR 0.138223f
C27 VPWR VGND 0.070329f
C28 B C 0.003039f
C29 C X 0.001363f
C30 a_416_86# a_1215_396# 0.096382f
C31 a_416_86# VGND 0.216545f
C32 X VNB 0.109996f
C33 C VNB 0.336344f
C34 VGND VNB 1.04461f
C35 VPWR VNB 0.83043f
C36 B VNB 0.820474f
C37 A VNB 0.11454f
C38 VPB VNB 2.1204f
C39 a_1215_396# VNB 0.168542f
C40 a_416_86# VNB 0.062961f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor3_2 VNB VPB VPWR VGND B C A X
X0 a_83_289.t3 A.t0 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.16985 pd=1.275 as=0.34745 ps=1.81 w=0.64 l=0.15
X1 VPWR.t1 a_1195_424# X.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 X.t0 a_1195_424# VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3956 ps=1.865 w=1.12 l=0.15
X3 a_27_134.t0 a_440_315.t2 a_416_113.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.15815 pd=1.16 as=0.10375 ps=0.99 w=0.42 l=0.15
X4 a_83_289.t1 a_440_315.t3 a_372_419# VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2848 pd=2.17 as=0.1495 ps=1.14 w=0.64 l=0.15
X5 a_1195_424# a_1162_379.t2 a_372_419# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.169775 pd=1.24 as=0.176 ps=1.83 w=0.64 l=0.15
X6 VPWR.t4 a_83_289.t6 a_27_134.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2225 pd=1.445 as=0.295 ps=2.59 w=1 l=0.15
X7 a_83_289.t4 A.t1 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2225 ps=1.445 w=1 l=0.15
X8 VGND.t1 a_1195_424# X.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_416_113.t0 B.t0 a_83_289.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10375 pd=0.99 as=0.16985 ps=1.275 w=0.64 l=0.15
X10 VPWR.t3 C.t0 a_1162_379.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3956 pd=1.865 as=0.24 ps=2.03 w=0.64 l=0.15
X11 a_372_419# C a_1195_424# VPB sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2562 ps=1.45 w=0.84 l=0.15
X12 a_416_113.t3 B.t1 a_27_134.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1527 pd=1.225 as=0.096 ps=0.94 w=0.64 l=0.15
X13 a_416_113.t4 C.t1 a_1195_424# VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2144 pd=1.95 as=0.169775 ps=1.24 w=0.64 l=0.15
X14 a_27_134.t1 a_440_315.t4 a_372_419# VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1401 ps=1.195 w=0.64 l=0.15
X15 VGND.t4 B.t2 a_440_315.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.46725 pd=2.88 as=0.2035 ps=2.03 w=0.74 l=0.15
X16 X.t1 a_1195_424# VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1471 ps=1.17 w=0.74 l=0.15
X17 a_372_419# B.t3 a_83_289.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1401 pd=1.195 as=0.1853 ps=1.385 w=0.84 l=0.15
X18 a_83_289.t2 a_440_315.t5 a_416_113.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.5544 pd=3 as=0.1527 ps=1.225 w=0.84 l=0.15
X19 VGND.t2 C.t2 a_1162_379.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1471 pd=1.17 as=0.1197 ps=1.41 w=0.42 l=0.15
X20 a_372_419# B.t4 a_27_134.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1495 pd=1.14 as=0.15815 ps=1.16 w=0.64 l=0.15
X21 VGND.t3 a_83_289.t7 a_27_134.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.34745 pd=1.81 as=0.1824 ps=1.85 w=0.64 l=0.15
X22 VPWR.t2 B.t5 a_440_315.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 A.n0 A.t1 232.095
R1 A A.n0 166.546
R2 A.n0 A.t0 156.046
R3 VGND.n20 VGND.t4 348.695
R4 VGND.n1 VGND.n0 263.113
R5 VGND.n11 VGND.t1 179.755
R6 VGND.n10 VGND.n9 117.826
R7 VGND.n9 VGND.t2 66.7516
R8 VGND.n0 VGND.t5 63.7505
R9 VGND.n0 VGND.t3 63.7505
R10 VGND.n14 VGND.n13 36.1417
R11 VGND.n15 VGND.n14 36.1417
R12 VGND.n15 VGND.n7 36.1417
R13 VGND.n19 VGND.n7 36.1417
R14 VGND.n21 VGND.n5 36.1417
R15 VGND.n25 VGND.n5 36.1417
R16 VGND.n26 VGND.n25 36.1417
R17 VGND.n27 VGND.n26 36.1417
R18 VGND.n27 VGND.n3 36.1417
R19 VGND.n31 VGND.n3 36.1417
R20 VGND.n32 VGND.n31 36.1417
R21 VGND.n33 VGND.n32 36.1417
R22 VGND.n9 VGND.t0 33.6878
R23 VGND.n20 VGND.n19 32.7534
R24 VGND.n13 VGND.n10 21.4593
R25 VGND.n21 VGND.n20 20.7064
R26 VGND.n35 VGND.n1 11.7718
R27 VGND.n34 VGND.n33 9.3005
R28 VGND.n32 VGND.n2 9.3005
R29 VGND.n31 VGND.n30 9.3005
R30 VGND.n29 VGND.n3 9.3005
R31 VGND.n28 VGND.n27 9.3005
R32 VGND.n26 VGND.n4 9.3005
R33 VGND.n25 VGND.n24 9.3005
R34 VGND.n23 VGND.n5 9.3005
R35 VGND.n22 VGND.n21 9.3005
R36 VGND.n20 VGND.n6 9.3005
R37 VGND.n19 VGND.n18 9.3005
R38 VGND.n17 VGND.n7 9.3005
R39 VGND.n16 VGND.n15 9.3005
R40 VGND.n14 VGND.n8 9.3005
R41 VGND.n13 VGND.n12 9.3005
R42 VGND.n11 VGND.n10 6.81625
R43 VGND.n33 VGND.n1 6.72132
R44 VGND.n12 VGND.n11 0.584177
R45 VGND VGND.n35 0.161517
R46 VGND.n35 VGND.n34 0.146304
R47 VGND.n12 VGND.n8 0.122949
R48 VGND.n16 VGND.n8 0.122949
R49 VGND.n17 VGND.n16 0.122949
R50 VGND.n18 VGND.n17 0.122949
R51 VGND.n18 VGND.n6 0.122949
R52 VGND.n22 VGND.n6 0.122949
R53 VGND.n23 VGND.n22 0.122949
R54 VGND.n24 VGND.n23 0.122949
R55 VGND.n24 VGND.n4 0.122949
R56 VGND.n28 VGND.n4 0.122949
R57 VGND.n29 VGND.n28 0.122949
R58 VGND.n30 VGND.n29 0.122949
R59 VGND.n30 VGND.n2 0.122949
R60 VGND.n34 VGND.n2 0.122949
R61 a_83_289.n4 a_83_289.n3 543.673
R62 a_83_289.n3 a_83_289.t2 397.92
R63 a_83_289.n3 a_83_289.t1 305.791
R64 a_83_289.n5 a_83_289.n4 291.305
R65 a_83_289.n2 a_83_289.n1 245.302
R66 a_83_289.n0 a_83_289.t6 231.629
R67 a_83_289.n2 a_83_289.n0 210.341
R68 a_83_289.n0 a_83_289.t7 170.308
R69 a_83_289.n1 a_83_289.t0 81.4873
R70 a_83_289.n5 a_83_289.t5 55.1136
R71 a_83_289.t4 a_83_289.n5 30.7494
R72 a_83_289.n1 a_83_289.t3 23.315
R73 a_83_289.n4 a_83_289.n2 16.229
R74 VNB.t10 VNB.t4 2864.04
R75 VNB.t9 VNB.t7 2817.85
R76 VNB.t6 VNB.t9 2702.36
R77 VNB.t8 VNB.t11 1917.06
R78 VNB.t7 VNB.t10 1570.6
R79 VNB.t11 VNB.t2 1570.6
R80 VNB.t5 VNB.t3 1547.51
R81 VNB.t3 VNB.t6 1362.73
R82 VNB.t4 VNB.t0 1339.63
R83 VNB.t2 VNB.t5 1154.86
R84 VNB VNB.t8 1143.31
R85 VNB.t0 VNB.t1 993.177
R86 X.n4 X 589.85
R87 X.n4 X.n0 585
R88 X.n5 X.n4 585
R89 X.n3 X.n2 185
R90 X.n2 X.n1 185
R91 X.n4 X.t3 26.3844
R92 X.n4 X.t0 26.3844
R93 X.n2 X.t2 22.7032
R94 X.n2 X.t1 22.7032
R95 X X.n5 12.9944
R96 X.n1 X 11.8308
R97 X X.n0 11.249
R98 X X.n3 8.72777
R99 X.n3 X 5.62474
R100 X X.n0 3.10353
R101 X.n1 X 2.52171
R102 X.n5 X 1.35808
R103 VPWR.n34 VPWR.n1 316.943
R104 VPWR.n11 VPWR.t1 266.226
R105 VPWR.n21 VPWR.t2 259.171
R106 VPWR.n10 VPWR.n9 119.267
R107 VPWR.n9 VPWR.t3 75.9978
R108 VPWR.n9 VPWR.t0 59.6916
R109 VPWR.n1 VPWR.t5 48.2655
R110 VPWR.n1 VPWR.t4 39.4005
R111 VPWR.n22 VPWR.n4 36.1417
R112 VPWR.n26 VPWR.n4 36.1417
R113 VPWR.n27 VPWR.n26 36.1417
R114 VPWR.n28 VPWR.n27 36.1417
R115 VPWR.n28 VPWR.n2 36.1417
R116 VPWR.n32 VPWR.n2 36.1417
R117 VPWR.n33 VPWR.n32 36.1417
R118 VPWR.n14 VPWR.n8 36.1417
R119 VPWR.n15 VPWR.n14 36.1417
R120 VPWR.n16 VPWR.n15 36.1417
R121 VPWR.n16 VPWR.n6 36.1417
R122 VPWR.n20 VPWR.n6 36.1417
R123 VPWR.n22 VPWR.n21 29.3652
R124 VPWR.n21 VPWR.n20 24.0946
R125 VPWR.n35 VPWR.n34 11.092
R126 VPWR.n12 VPWR.n8 9.3005
R127 VPWR.n14 VPWR.n13 9.3005
R128 VPWR.n15 VPWR.n7 9.3005
R129 VPWR.n17 VPWR.n16 9.3005
R130 VPWR.n18 VPWR.n6 9.3005
R131 VPWR.n20 VPWR.n19 9.3005
R132 VPWR.n21 VPWR.n5 9.3005
R133 VPWR.n23 VPWR.n22 9.3005
R134 VPWR.n24 VPWR.n4 9.3005
R135 VPWR.n26 VPWR.n25 9.3005
R136 VPWR.n27 VPWR.n3 9.3005
R137 VPWR.n29 VPWR.n28 9.3005
R138 VPWR.n30 VPWR.n2 9.3005
R139 VPWR.n32 VPWR.n31 9.3005
R140 VPWR.n33 VPWR.n0 9.3005
R141 VPWR.n34 VPWR.n33 7.90638
R142 VPWR.n11 VPWR.n10 6.8559
R143 VPWR.n10 VPWR.n8 4.14168
R144 VPWR.n12 VPWR.n11 0.565232
R145 VPWR VPWR.n35 0.163644
R146 VPWR.n35 VPWR.n0 0.144205
R147 VPWR.n13 VPWR.n12 0.122949
R148 VPWR.n13 VPWR.n7 0.122949
R149 VPWR.n17 VPWR.n7 0.122949
R150 VPWR.n18 VPWR.n17 0.122949
R151 VPWR.n19 VPWR.n18 0.122949
R152 VPWR.n19 VPWR.n5 0.122949
R153 VPWR.n23 VPWR.n5 0.122949
R154 VPWR.n24 VPWR.n23 0.122949
R155 VPWR.n25 VPWR.n24 0.122949
R156 VPWR.n25 VPWR.n3 0.122949
R157 VPWR.n29 VPWR.n3 0.122949
R158 VPWR.n30 VPWR.n29 0.122949
R159 VPWR.n31 VPWR.n30 0.122949
R160 VPWR.n31 VPWR.n0 0.122949
R161 VPB.t2 VPB.t5 1460.75
R162 VPB.t4 VPB.t2 824.866
R163 VPB.t5 VPB.t0 457.125
R164 VPB VPB.t7 334.543
R165 VPB.t7 VPB.t8 303.899
R166 VPB.t6 VPB.t4 273.253
R167 VPB.t8 VPB.t9 273.253
R168 VPB.t9 VPB.t3 257.93
R169 VPB.t0 VPB.t1 229.839
R170 VPB.t3 VPB.t6 229.839
R171 a_440_315.t0 a_440_315.n3 323.281
R172 a_440_315.n3 a_440_315.n2 272.488
R173 a_440_315.n0 a_440_315.t4 266.171
R174 a_440_315.n1 a_440_315.n0 236.214
R175 a_440_315.n3 a_440_315.t1 207.703
R176 a_440_315.n0 a_440_315.t2 186.374
R177 a_440_315.n2 a_440_315.t3 169.602
R178 a_440_315.n1 a_440_315.t5 159.06
R179 a_440_315.n2 a_440_315.n1 132.704
R180 a_416_113.n2 a_416_113.n1 588.88
R181 a_416_113.n1 a_416_113.t4 418.627
R182 a_416_113.n1 a_416_113.n0 278.825
R183 a_416_113.n2 a_416_113.t3 72.3364
R184 a_416_113.n3 a_416_113.n2 66.7802
R185 a_416_113.n0 a_416_113.t2 60.7549
R186 a_416_113.n2 a_416_113.t1 35.1315
R187 a_416_113.n0 a_416_113.t0 25.9831
R188 a_27_134.n2 a_27_134.n0 615.837
R189 a_27_134.t4 a_27_134.n3 412.753
R190 a_27_134.n2 a_27_134.n1 209.163
R191 a_27_134.n3 a_27_134.n2 194.421
R192 a_27_134.n3 a_27_134.t5 125.329
R193 a_27_134.n1 a_27_134.t2 58.1255
R194 a_27_134.n1 a_27_134.t0 46.7416
R195 a_27_134.n0 a_27_134.t3 46.1724
R196 a_27_134.n0 a_27_134.t1 46.1724
R197 a_1162_379.t1 a_1162_379.n2 655.798
R198 a_1162_379.n2 a_1162_379.n1 379.735
R199 a_1162_379.n2 a_1162_379.t0 337.269
R200 a_1162_379.n1 a_1162_379.n0 329.409
R201 a_1162_379.n1 a_1162_379.t2 181.596
R202 B.n2 B.n0 1028.15
R203 B.n2 B.n1 714.967
R204 B.n1 B.t0 578.4
R205 B.n0 B.t3 445.582
R206 B.n4 B.t5 279.293
R207 B.n0 B.t1 217.971
R208 B.n1 B.t4 202.44
R209 B.n3 B.t2 162.274
R210 B B.n4 158.788
R211 B.n3 B.n2 117.287
R212 B.n4 B.n3 9.6405
R213 C.n0 C.t2 303.661
R214 C.n2 C.n1 289.712
R215 C.n3 C.n0 215.293
R216 C.n0 C.t0 196.549
R217 C C.n3 167.873
R218 C.n2 C.t1 138.173
R219 C.n3 C.n2 20.449
C0 VPWR B 0.121293f
C1 A a_372_419# 2.85e-20
C2 X VGND 0.164715f
C3 A VPWR 0.015729f
C4 VPB a_372_419# 0.03022f
C5 a_372_419# a_1195_424# 0.121285f
C6 C a_372_419# 0.109813f
C7 VPWR VPB 0.236416f
C8 A B 0.007533f
C9 VPWR a_1195_424# 0.217866f
C10 VPWR C 0.012332f
C11 VPB B 0.482501f
C12 B a_1195_424# 3.75e-19
C13 C B 0.003379f
C14 VGND a_372_419# 0.50665f
C15 A VPB 0.051339f
C16 VPWR VGND 0.09074f
C17 X VPWR 0.189682f
C18 VPB a_1195_424# 0.101955f
C19 C VPB 0.13944f
C20 VGND B 0.082305f
C21 C a_1195_424# 0.115006f
C22 X B 1.51e-19
C23 A VGND 0.013826f
C24 VGND VPB 0.015295f
C25 VGND a_1195_424# 0.127979f
C26 VGND C 0.027103f
C27 VPWR a_372_419# 0.028535f
C28 X VPB 0.005552f
C29 X a_1195_424# 0.148414f
C30 X C 0.001518f
C31 B a_372_419# 0.097732f
C32 X VNB 0.03125f
C33 C VNB 0.345932f
C34 VGND VNB 1.13314f
C35 VPWR VNB 0.919777f
C36 A VNB 0.114753f
C37 B VNB 0.848326f
C38 VPB VNB 2.22754f
C39 a_1195_424# VNB 0.283368f
C40 a_372_419# VNB 0.087749f
.ends

* NGSPICE file created from sky130_fd_sc_hs__xor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor3_4 VNB VPB VPWR VGND X B C A
X0 VGND.t1 B.t0 a_397_320.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.42 pd=2.67 as=0.2072 ps=2.04 w=0.74 l=0.15
X1 a_416_118.t0 B.t1 a_74_294.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10375 pd=0.99 as=0.2208 ps=1.33 w=0.64 l=0.15
X2 VPWR.t4 a_74_294.t6 a_27_118.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X3 VGND.t2 a_1218_388.t4 X.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 X.t3 a_1218_388.t5 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2128 ps=1.5 w=1.12 l=0.15
X5 VGND.t3 a_1218_388.t6 X.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_27_118.t5 a_397_320.t2 a_416_118.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.09 as=0.10375 ps=0.99 w=0.42 l=0.15
X7 a_323_392.t0 B.t2 a_27_118.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.145875 pd=1.115 as=0.122 ps=1.09 w=0.64 l=0.15
X8 a_1218_388.t3 a_1155_284# a_416_118.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2226 pd=1.37 as=0.3822 ps=2.59 w=0.84 l=0.15
X9 a_323_392.t1 B.t3 a_74_294.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1527 pd=1.225 as=0.1853 ps=1.385 w=0.84 l=0.15
X10 VPWR.t2 a_1218_388.t7 X.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2128 pd=1.5 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t0 B.t4 a_397_320.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X12 X.t1 a_1218_388.t8 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4012 ps=1.875 w=1.12 l=0.15
X13 a_74_294.t3 A.t0 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.175 ps=1.35 w=1 l=0.15
X14 a_74_294.t4 a_397_320.t3 a_416_118.t5 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.546 pd=2.98 as=0.152625 ps=1.225 w=0.84 l=0.15
X15 a_323_392.t2 C.t0 a_1218_388.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2226 ps=1.37 w=0.84 l=0.15
X16 a_74_294.t0 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2208 pd=1.33 as=0.24225 ps=1.57 w=0.64 l=0.15
X17 a_27_118.t4 a_397_320.t4 a_323_392.t4 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.149875 pd=1.215 as=0.1527 ps=1.225 w=0.64 l=0.15
X18 a_74_294.t5 a_397_320.t5 a_323_392.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2848 pd=2.17 as=0.145875 ps=1.115 w=0.64 l=0.15
X19 a_416_118.t1 B.t5 a_27_118.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.152625 pd=1.225 as=0.149875 ps=1.215 w=0.64 l=0.15
X20 VGND C a_1155_284# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1471 pd=1.17 as=0.2121 ps=1.85 w=0.42 l=0.15
X21 VPWR.t6 a_1218_388.t9 X.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X22 VPWR C a_1155_284# VPB sky130_fd_pr__pfet_01v8 ad=0.4012 pd=1.875 as=0.1888 ps=1.87 w=0.64 l=0.15
X23 VGND.t4 a_74_294.t7 a_27_118.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.24225 pd=1.57 as=0.1824 ps=1.85 w=0.64 l=0.15
X24 a_1218_388.t2 a_1155_284# a_323_392.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.17 as=0.176 ps=1.83 w=0.64 l=0.15
X25 a_416_118.t2 C.t1 a_1218_388.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1696 ps=1.17 w=0.64 l=0.15
R0 B.n2 B.n1 1005.77
R1 B.n2 B.n0 772.808
R2 B.n0 B.t1 563.941
R3 B.n1 B.t3 537.966
R4 B.n3 B.t4 269.074
R5 B.n1 B.t5 219.31
R6 B.n0 B.t2 210.474
R7 B.n4 B.t0 170.638
R8 B B.n4 158.788
R9 B.n3 B.n2 125.32
R10 B.n4 B.n3 8.94483
R11 a_397_320.t1 a_397_320.n3 319.158
R12 a_397_320.n0 a_397_320.t4 292.413
R13 a_397_320.n3 a_397_320.n2 278.781
R14 a_397_320.n1 a_397_320.n0 215.732
R15 a_397_320.n3 a_397_320.t0 207.703
R16 a_397_320.n0 a_397_320.t2 186.374
R17 a_397_320.n2 a_397_320.t5 169.602
R18 a_397_320.n1 a_397_320.t3 159.06
R19 a_397_320.n2 a_397_320.n1 138.018
R20 VGND.n26 VGND.t1 271.027
R21 VGND.n1 VGND.n0 270.947
R22 VGND.n12 VGND.t3 181.082
R23 VGND.n11 VGND.t2 169.915
R24 VGND.n0 VGND.t0 48.7505
R25 VGND.n0 VGND.t4 48.7505
R26 VGND.n12 VGND.n11 36.1737
R27 VGND.n14 VGND.n13 36.1417
R28 VGND.n19 VGND.n18 36.1417
R29 VGND.n20 VGND.n19 36.1417
R30 VGND.n20 VGND.n7 36.1417
R31 VGND.n24 VGND.n7 36.1417
R32 VGND.n25 VGND.n24 36.1417
R33 VGND.n27 VGND.n5 36.1417
R34 VGND.n31 VGND.n5 36.1417
R35 VGND.n32 VGND.n31 36.1417
R36 VGND.n33 VGND.n32 36.1417
R37 VGND.n33 VGND.n3 36.1417
R38 VGND.n37 VGND.n3 36.1417
R39 VGND.n38 VGND.n37 36.1417
R40 VGND.n39 VGND.n38 36.1417
R41 VGND.n18 VGND.n9 30.8711
R42 VGND.n39 VGND.n1 17.725
R43 VGND.n14 VGND.n9 16.5652
R44 VGND.n27 VGND.n26 15.8123
R45 VGND.n41 VGND.n1 10.3987
R46 VGND.n40 VGND.n39 9.3005
R47 VGND.n38 VGND.n2 9.3005
R48 VGND.n37 VGND.n36 9.3005
R49 VGND.n35 VGND.n3 9.3005
R50 VGND.n34 VGND.n33 9.3005
R51 VGND.n32 VGND.n4 9.3005
R52 VGND.n31 VGND.n30 9.3005
R53 VGND.n29 VGND.n5 9.3005
R54 VGND.n28 VGND.n27 9.3005
R55 VGND.n25 VGND.n6 9.3005
R56 VGND.n24 VGND.n23 9.3005
R57 VGND.n22 VGND.n7 9.3005
R58 VGND.n21 VGND.n20 9.3005
R59 VGND.n19 VGND.n8 9.3005
R60 VGND.n18 VGND.n17 9.3005
R61 VGND.n16 VGND.n9 9.3005
R62 VGND.n13 VGND.n10 9.3005
R63 VGND.n15 VGND.n14 9.3005
R64 VGND.n13 VGND.n12 4.89462
R65 VGND.n11 VGND.n10 2.32491
R66 VGND.n26 VGND.n25 1.50638
R67 VGND VGND.n41 0.161675
R68 VGND.n41 VGND.n40 0.146149
R69 VGND.n15 VGND.n10 0.122949
R70 VGND.n16 VGND.n15 0.122949
R71 VGND.n17 VGND.n16 0.122949
R72 VGND.n17 VGND.n8 0.122949
R73 VGND.n21 VGND.n8 0.122949
R74 VGND.n22 VGND.n21 0.122949
R75 VGND.n23 VGND.n22 0.122949
R76 VGND.n23 VGND.n6 0.122949
R77 VGND.n28 VGND.n6 0.122949
R78 VGND.n29 VGND.n28 0.122949
R79 VGND.n30 VGND.n29 0.122949
R80 VGND.n30 VGND.n4 0.122949
R81 VGND.n34 VGND.n4 0.122949
R82 VGND.n35 VGND.n34 0.122949
R83 VGND.n36 VGND.n35 0.122949
R84 VGND.n36 VGND.n2 0.122949
R85 VGND.n40 VGND.n2 0.122949
R86 VNB.t4 VNB.t7 5635.7
R87 VNB.t3 VNB.t5 2817.85
R88 VNB.t9 VNB.t3 2713.91
R89 VNB.t7 VNB.t6 1986.35
R90 VNB.t0 VNB.t2 1940.16
R91 VNB.t5 VNB.t4 1570.6
R92 VNB.t8 VNB.t0 1547.51
R93 VNB.t10 VNB.t1 1385.83
R94 VNB.t1 VNB.t9 1362.73
R95 VNB.t2 VNB.t10 1154.86
R96 VNB VNB.t8 1143.31
R97 a_74_294.n7 a_74_294.n6 585
R98 a_74_294.n1 a_74_294.t4 397.92
R99 a_74_294.n1 a_74_294.t5 305.791
R100 a_74_294.n5 a_74_294.n0 289.146
R101 a_74_294.n4 a_74_294.n3 252.766
R102 a_74_294.n2 a_74_294.t6 231.629
R103 a_74_294.n2 a_74_294.t7 204.048
R104 a_74_294.n6 a_74_294.n1 202.726
R105 a_74_294.n4 a_74_294.n2 192.982
R106 a_74_294.n3 a_74_294.t1 73.1255
R107 a_74_294.n3 a_74_294.t0 56.2505
R108 a_74_294.n0 a_74_294.t2 55.1136
R109 a_74_294.n8 a_74_294.n7 43.4073
R110 a_74_294.n0 a_74_294.t3 29.5767
R111 a_74_294.n6 a_74_294.n5 20.6747
R112 a_74_294.n5 a_74_294.n4 13.6928
R113 a_74_294.n7 a_74_294.n0 11.1901
R114 a_416_118.n2 a_416_118.n1 585
R115 a_416_118.t3 a_416_118.n3 371.288
R116 a_416_118.n3 a_416_118.t2 313.591
R117 a_416_118.n2 a_416_118.n0 254.686
R118 a_416_118.n1 a_416_118.t1 72.3364
R119 a_416_118.n0 a_416_118.t4 60.7404
R120 a_416_118.n1 a_416_118.t5 32.3585
R121 a_416_118.n3 a_416_118.n2 29.4398
R122 a_416_118.n0 a_416_118.t0 25.9975
R123 a_27_118.n2 a_27_118.n1 621.096
R124 a_27_118.t2 a_27_118.n3 416.836
R125 a_27_118.n2 a_27_118.n0 222.632
R126 a_27_118.n3 a_27_118.n2 186.261
R127 a_27_118.n3 a_27_118.t3 126.305
R128 a_27_118.n1 a_27_118.t1 99.8903
R129 a_27_118.n0 a_27_118.t0 76.2951
R130 a_27_118.n1 a_27_118.t4 40.7889
R131 a_27_118.n0 a_27_118.t5 40.0005
R132 VPWR.n40 VPWR.n1 316.964
R133 VPWR.n12 VPWR.t6 264.714
R134 VPWR.n27 VPWR.t0 250.081
R135 VPWR.n11 VPWR.n10 243.916
R136 VPWR.n16 VPWR.t5 179.311
R137 VPWR.n10 VPWR.t2 40.4559
R138 VPWR.n12 VPWR.n11 40.1055
R139 VPWR.n1 VPWR.t3 39.4005
R140 VPWR.n28 VPWR.n4 36.1417
R141 VPWR.n32 VPWR.n4 36.1417
R142 VPWR.n33 VPWR.n32 36.1417
R143 VPWR.n34 VPWR.n33 36.1417
R144 VPWR.n34 VPWR.n2 36.1417
R145 VPWR.n38 VPWR.n2 36.1417
R146 VPWR.n39 VPWR.n38 36.1417
R147 VPWR.n20 VPWR.n8 36.1417
R148 VPWR.n21 VPWR.n20 36.1417
R149 VPWR.n22 VPWR.n21 36.1417
R150 VPWR.n22 VPWR.n6 36.1417
R151 VPWR.n26 VPWR.n6 36.1417
R152 VPWR.n15 VPWR.n14 36.1417
R153 VPWR.n1 VPWR.t4 29.5505
R154 VPWR.n16 VPWR.n15 28.6123
R155 VPWR.n10 VPWR.t1 26.3844
R156 VPWR.n28 VPWR.n27 25.977
R157 VPWR.n40 VPWR.n39 22.9652
R158 VPWR.n27 VPWR.n26 21.4593
R159 VPWR.n14 VPWR.n13 9.3005
R160 VPWR.n15 VPWR.n9 9.3005
R161 VPWR.n17 VPWR.n16 9.3005
R162 VPWR.n18 VPWR.n8 9.3005
R163 VPWR.n20 VPWR.n19 9.3005
R164 VPWR.n21 VPWR.n7 9.3005
R165 VPWR.n23 VPWR.n22 9.3005
R166 VPWR.n24 VPWR.n6 9.3005
R167 VPWR.n26 VPWR.n25 9.3005
R168 VPWR.n27 VPWR.n5 9.3005
R169 VPWR.n29 VPWR.n28 9.3005
R170 VPWR.n30 VPWR.n4 9.3005
R171 VPWR.n32 VPWR.n31 9.3005
R172 VPWR.n33 VPWR.n3 9.3005
R173 VPWR.n35 VPWR.n34 9.3005
R174 VPWR.n36 VPWR.n2 9.3005
R175 VPWR.n38 VPWR.n37 9.3005
R176 VPWR.n39 VPWR.n0 9.3005
R177 VPWR.n41 VPWR.n40 7.27223
R178 VPWR.n13 VPWR.n12 2.0514
R179 VPWR.n16 VPWR.n8 1.88285
R180 VPWR.n14 VPWR.n11 1.50638
R181 VPWR VPWR.n41 0.157962
R182 VPWR.n41 VPWR.n0 0.149814
R183 VPWR.n13 VPWR.n9 0.122949
R184 VPWR.n17 VPWR.n9 0.122949
R185 VPWR.n18 VPWR.n17 0.122949
R186 VPWR.n19 VPWR.n18 0.122949
R187 VPWR.n19 VPWR.n7 0.122949
R188 VPWR.n23 VPWR.n7 0.122949
R189 VPWR.n24 VPWR.n23 0.122949
R190 VPWR.n25 VPWR.n24 0.122949
R191 VPWR.n25 VPWR.n5 0.122949
R192 VPWR.n29 VPWR.n5 0.122949
R193 VPWR.n30 VPWR.n29 0.122949
R194 VPWR.n31 VPWR.n30 0.122949
R195 VPWR.n31 VPWR.n3 0.122949
R196 VPWR.n35 VPWR.n3 0.122949
R197 VPWR.n36 VPWR.n35 0.122949
R198 VPWR.n37 VPWR.n36 0.122949
R199 VPWR.n37 VPWR.n0 0.122949
R200 VPB.t3 VPB.t9 985.754
R201 VPB.t12 VPB.t1 837.635
R202 VPB.t1 VPB.t4 597.582
R203 VPB.t4 VPB.t3 347.312
R204 VPB.t11 VPB.t0 303.899
R205 VPB.t0 VPB.t12 273.253
R206 VPB.t2 VPB.t11 273.253
R207 VPB.t7 VPB.t2 273.253
R208 VPB.t6 VPB.t5 270.7
R209 VPB VPB.t8 257.93
R210 VPB.t8 VPB.t7 255.376
R211 VPB.t5 VPB.t10 229.839
R212 VPB.t9 VPB.t6 229.839
R213 a_1218_388.n11 a_1218_388.n10 298.973
R214 a_1218_388.n9 a_1218_388.t8 256.628
R215 a_1218_388.n3 a_1218_388.t9 252.248
R216 a_1218_388.n5 a_1218_388.t5 252.248
R217 a_1218_388.n7 a_1218_388.t7 252.248
R218 a_1218_388.n10 a_1218_388.n0 250.76
R219 a_1218_388.n3 a_1218_388.t4 167.679
R220 a_1218_388.n8 a_1218_388.n1 165.488
R221 a_1218_388.n6 a_1218_388.t6 165.488
R222 a_1218_388.n4 a_1218_388.n2 165.488
R223 a_1218_388.n10 a_1218_388.n9 115.29
R224 a_1218_388.n11 a_1218_388.t3 89.1195
R225 a_1218_388.n0 a_1218_388.t2 73.1255
R226 a_1218_388.n4 a_1218_388.n3 60.6157
R227 a_1218_388.n6 a_1218_388.n5 57.6944
R228 a_1218_388.n8 a_1218_388.n7 43.0884
R229 a_1218_388.t0 a_1218_388.n11 35.1791
R230 a_1218_388.n0 a_1218_388.t1 26.2505
R231 a_1218_388.n7 a_1218_388.n6 19.7187
R232 a_1218_388.n9 a_1218_388.n8 17.9155
R233 a_1218_388.n5 a_1218_388.n4 5.11262
R234 X.n5 X.n4 585
R235 X.n4 X.n0 290.923
R236 X.n2 X.n1 238.042
R237 X.n3 X.t5 167.357
R238 X.n2 X.t4 164.405
R239 X.n3 X.n2 38.024
R240 X.n4 X.t0 26.3844
R241 X.n4 X.t3 26.3844
R242 X.n1 X.t2 26.3844
R243 X.n1 X.t1 26.3844
R244 X X.n5 12.9944
R245 X X.n3 8.84414
R246 X X.n0 8.65194
R247 X.n0 X 5.59489
R248 X.n5 X 1.35808
R249 a_323_392.n2 a_323_392.t2 636.069
R250 a_323_392.n1 a_323_392.n0 17.1792
R251 a_323_392.n2 a_323_392.t3 257
R252 a_323_392.n4 a_323_392.n2 242.306
R253 a_323_392.n1 a_323_392.n4 520.63
R254 a_323_392.n4 a_323_392.n3 85.7805
R255 a_323_392.n0 a_323_392.t4 72.3364
R256 a_323_392.n0 a_323_392.t1 34.2334
R257 a_323_392.n3 a_323_392.t0 33.7864
R258 a_323_392.n5 a_323_392.n1 50.1414
R259 a_323_392.n3 a_323_392.t5 33.3106
R260 A.n0 A.t0 266.44
R261 A.n0 A.t1 162.274
R262 A A.n0 162.07
R263 C.n2 C.n1 526.987
R264 C.n2 C.n0 282.774
R265 C.n3 C.t0 192.776
R266 C.n3 C.t1 165.488
R267 C C.n4 154.522
R268 C.n4 C.n2 49.6611
R269 C.n4 C.n3 24.8308
C0 VPB C 0.149678f
C1 A VPWR 0.018662f
C2 VGND B 0.078185f
C3 VPWR C 0.012253f
C4 VGND a_1155_284# 0.096777f
C5 VGND X 0.34513f
C6 VPB VPWR 0.265346f
C7 B a_1155_284# 0.016518f
C8 B X 3.32e-19
C9 VGND A 0.009399f
C10 X a_1155_284# 0.003253f
C11 VGND C 0.030472f
C12 A B 0.01723f
C13 B C 0.004374f
C14 VGND VPB 0.015525f
C15 C a_1155_284# 0.090832f
C16 C X 0.002383f
C17 VGND VPWR 0.095889f
C18 VPB B 0.520497f
C19 VPB a_1155_284# 0.102314f
C20 VPB X 0.013943f
C21 B VPWR 0.130581f
C22 VPWR a_1155_284# 0.288952f
C23 VPWR X 0.444428f
C24 VPB A 0.041779f
C25 VGND VNB 1.24232f
C26 X VNB 0.040085f
C27 C VNB 0.361891f
C28 VPWR VNB 0.991161f
C29 B VNB 0.8543f
C30 A VNB 0.111957f
C31 VPB VNB 2.44181f
C32 a_1155_284# VNB 0.135432f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2111a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2111a_1 VNB VPB VPWR VGND A1 A2 B1 C1 D1 X
X0 VPWR.t3 a_82_48.t5 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.241575 pd=1.6 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t2 A2.t0 a_471_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1332 ps=1.1 w=0.74 l=0.15
X2 a_471_74.t1 A1.t0 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1443 ps=1.13 w=0.74 l=0.15
X3 VPWR.t4 A1.t1 a_600_381.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t0 C1.t0 a_82_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2541 pd=1.445 as=0.147 ps=1.19 w=0.84 l=0.15
X5 a_600_381.t1 A2.t1 a_82_48.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.1853 ps=1.385 w=1 l=0.15
X6 VGND.t0 a_82_48.t6 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.2035 ps=2.03 w=0.74 l=0.15
X7 a_471_74.t0 B1.t0 a_393_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X8 a_82_48.t1 D1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.241575 ps=1.6 w=0.84 l=0.15
X9 a_321_74.t1 D1.t1 a_82_48.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.259 ps=2.18 w=0.74 l=0.15
X10 a_393_74.t0 C1.t1 a_321_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.0777 ps=0.95 w=0.74 l=0.15
X11 a_82_48.t3 B1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2541 ps=1.445 w=0.84 l=0.15
R0 a_82_48.n4 a_82_48.n3 373.745
R1 a_82_48.n3 a_82_48.n2 300.755
R2 a_82_48.n0 a_82_48.t5 284.022
R3 a_82_48.n1 a_82_48.t4 178.989
R4 a_82_48.n0 a_82_48.t6 176.643
R5 a_82_48.n1 a_82_48.n0 152
R6 a_82_48.n3 a_82_48.n1 82.4583
R7 a_82_48.n4 a_82_48.t3 55.1136
R8 a_82_48.n5 a_82_48.n4 53.4242
R9 a_82_48.n2 a_82_48.t0 46.9053
R10 a_82_48.n2 a_82_48.t1 35.1791
R11 a_82_48.n4 a_82_48.t2 30.4598
R12 X.n1 X 589.572
R13 X.n1 X.n0 585
R14 X.n2 X.n1 585
R15 X X.t0 191.04
R16 X.n1 X.t1 26.3844
R17 X X.n2 12.2519
R18 X X.n0 10.6062
R19 X X.n0 2.92621
R20 X.n2 X 1.2805
R21 VPWR.n3 VPWR.n2 601.524
R22 VPWR.n8 VPWR.n1 314.961
R23 VPWR.n4 VPWR.t4 261.077
R24 VPWR.n2 VPWR.t0 71.5303
R25 VPWR.n2 VPWR.t2 70.3576
R26 VPWR.n1 VPWR.t1 65.6672
R27 VPWR.n1 VPWR.t3 38.3849
R28 VPWR.n7 VPWR.n6 36.1417
R29 VPWR.n8 VPWR.n7 19.2005
R30 VPWR.n6 VPWR.n5 9.3005
R31 VPWR.n7 VPWR.n0 9.3005
R32 VPWR.n9 VPWR.n8 7.43488
R33 VPWR.n4 VPWR.n3 7.19642
R34 VPWR.n6 VPWR.n3 4.51815
R35 VPWR.n5 VPWR.n4 0.2368
R36 VPWR VPWR.n9 0.160103
R37 VPWR.n9 VPWR.n0 0.1477
R38 VPWR.n5 VPWR.n0 0.122949
R39 VPB.t0 VPB.t3 385.618
R40 VPB.t4 VPB.t1 321.774
R41 VPB.t3 VPB.t2 273.253
R42 VPB VPB.t4 257.93
R43 VPB.t1 VPB.t0 255.376
R44 VPB.t2 VPB.t5 214.517
R45 A2.n0 A2.t0 241
R46 A2.n0 A2.t1 231.629
R47 A2 A2.n0 157.436
R48 a_471_74.n0 a_471_74.t1 297.421
R49 a_471_74.t0 a_471_74.n0 30.8113
R50 a_471_74.n0 a_471_74.t2 27.5681
R51 VGND.n1 VGND.n0 213.466
R52 VGND.n1 VGND.t0 144.395
R53 VGND.n0 VGND.t1 34.0546
R54 VGND.n0 VGND.t2 29.1897
R55 VGND VGND.n1 0.190488
R56 VNB.t2 VNB.t1 2413.65
R57 VNB.t5 VNB.t4 1247.24
R58 VNB.t3 VNB.t5 1177.95
R59 VNB VNB.t2 1120.21
R60 VNB.t0 VNB.t3 900.788
R61 VNB.t1 VNB.t0 831.496
R62 A1.n0 A1.t1 254.892
R63 A1.n0 A1.t0 196.516
R64 A1 A1.n0 156.462
R65 a_600_381.t0 a_600_381.t1 53.1905
R66 C1.n0 C1.t1 285.642
R67 C1.n0 C1.t0 202.096
R68 C1 C1.n0 158.012
R69 B1.n0 B1.t1 248.767
R70 B1.n0 B1.t0 241
R71 B1 B1.n0 161.293
R72 a_393_74.t0 a_393_74.t1 38.9194
R73 D1.n0 D1.t1 322.94
R74 D1.n0 D1.t0 212.617
R75 D1 D1.n0 157.237
R76 a_321_74.t0 a_321_74.t1 34.0546
C0 X VPWR 0.089318f
C1 VPWR B1 0.018227f
C2 B1 A2 0.083661f
C3 VPWR D1 0.013879f
C4 X VGND 0.088641f
C5 VPWR A1 0.05442f
C6 X VPB 0.013254f
C7 C1 B1 0.109312f
C8 A1 A2 0.096574f
C9 VGND B1 0.017416f
C10 B1 VPB 0.055638f
C11 D1 C1 0.117789f
C12 VGND D1 0.010929f
C13 A1 C1 0.002282f
C14 A1 VGND 0.016715f
C15 D1 VPB 0.062079f
C16 A1 VPB 0.046636f
C17 X D1 0.001501f
C18 A1 B1 1.96e-19
C19 VPWR A2 0.022433f
C20 VPWR C1 0.017347f
C21 VPWR VGND 0.062945f
C22 VPWR VPB 0.124052f
C23 C1 A2 9.19e-19
C24 VGND A2 0.017568f
C25 A2 VPB 0.03836f
C26 VGND C1 0.039266f
C27 C1 VPB 0.060196f
C28 VGND VPB 0.009677f
C29 VGND VNB 0.497373f
C30 A1 VNB 0.1727f
C31 A2 VNB 0.105217f
C32 B1 VNB 0.103821f
C33 C1 VNB 0.115785f
C34 D1 VNB 0.134845f
C35 VPWR VNB 0.423041f
C36 X VNB 0.112276f
C37 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o311ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311ai_4 VNB VPB VPWR VGND Y C1 B1 A3 A2 A1
X0 Y.t10 C1.t0 VPWR.t5 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.294 pd=1.645 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_841_368.t6 A2.t0 a_1350_368.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_459_74.t4 A3.t0 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19445 ps=2.05 w=0.74 l=0.15
X3 VGND.t1 A3.t1 a_459_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1773 pd=1.28 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 Y.t5 A3.t2 a_841_368.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2688 pd=1.6 as=0.2072 ps=1.49 w=1.12 l=0.15
X5 VPWR.t2 A1.t0 a_1350_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_459_74.t7 B1.t0 a_27_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_1350_368.t6 A1.t1 VPWR.t6 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8 VGND.t5 A1.t2 a_459_74.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10915 ps=1.035 w=0.74 l=0.15
X9 VGND.t3 A2.t1 a_459_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 Y.t6 C1.t1 a_27_74.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 a_459_74.t2 A3.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1773 ps=1.28 w=0.74 l=0.15
X12 a_27_74.t2 B1.t1 a_459_74.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.19515 pd=2.05 as=0.1073 ps=1.03 w=0.74 l=0.15
X13 a_1350_368.t4 A2.t2 a_841_368.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR.t0 B1.t2 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=1.8984 pd=5.63 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_841_368.t0 A3.t4 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2688 ps=1.6 w=1.12 l=0.15
X16 Y.t4 B1.t3 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X17 a_841_368.t4 A2.t3 a_1350_368.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_27_74.t1 B1.t4 a_459_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_1350_368.t2 A2.t4 a_841_368.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X20 VPWR.t7 A1.t3 a_1350_368.t7 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_27_74.t6 C1.t2 Y.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_459_74.t10 A1.t4 VGND.t6 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_27_74.t5 C1.t3 Y.t11 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.10545 ps=1.025 w=0.74 l=0.15
X24 VPWR.t4 C1.t4 Y.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.294 ps=1.645 w=1.12 l=0.15
X25 a_841_368.t1 A3.t5 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2072 pd=1.49 as=0.196 ps=1.47 w=1.12 l=0.15
X26 a_459_74.t1 B1.t5 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 VGND.t7 A1.t5 a_459_74.t11 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.31265 pd=1.585 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 a_1350_368.t5 A1.t6 VPWR.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 Y.t8 C1.t5 a_27_74.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 VGND.t4 A2.t5 a_459_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.13135 ps=1.095 w=0.74 l=0.15
X31 Y.t2 A3.t6 a_841_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 C1.n1 C1.t2 281.168
R1 C1.n2 C1.t4 240.197
R2 C1.n6 C1.t0 240.197
R3 C1.n8 C1.n7 162.832
R4 C1.n4 C1.n3 161.067
R5 C1.n5 C1.n4 152
R6 C1.n1 C1.t5 142.994
R7 C1.n7 C1.t1 142.994
R8 C1.n0 C1.t3 142.994
R9 C1.n2 C1.n1 38.6688
R10 C1.n6 C1.n5 24.9129
R11 C1.n5 C1.n0 21.1218
R12 C1.n3 C1.n0 15.7061
R13 C1.n3 C1.n2 11.3735
R14 C1.n8 C1 6.4005
R15 C1 C1.n8 6.4005
R16 C1.n4 C1 2.66717
R17 C1.n7 C1.n6 1.08365
R18 VPWR.n35 VPWR.n34 353.183
R19 VPWR.n12 VPWR.t6 342.69
R20 VPWR.n15 VPWR.n14 316.305
R21 VPWR.n2 VPWR.n1 315.928
R22 VPWR.n45 VPWR.n44 292.5
R23 VPWR.n43 VPWR.n42 292.5
R24 VPWR.n41 VPWR.n5 292.5
R25 VPWR.n34 VPWR.n6 292.5
R26 VPWR.n13 VPWR.t7 266.168
R27 VPWR.n52 VPWR.t5 248.744
R28 VPWR.n34 VPWR.n5 61.563
R29 VPWR.n43 VPWR.n5 60.6835
R30 VPWR.n44 VPWR.n43 60.6835
R31 VPWR.n51 VPWR.n50 36.1417
R32 VPWR.n47 VPWR.n46 36.1417
R33 VPWR.n21 VPWR.n20 36.1417
R34 VPWR.n22 VPWR.n21 36.1417
R35 VPWR.n22 VPWR.n10 36.1417
R36 VPWR.n26 VPWR.n10 36.1417
R37 VPWR.n27 VPWR.n26 36.1417
R38 VPWR.n28 VPWR.n27 36.1417
R39 VPWR.n28 VPWR.n8 36.1417
R40 VPWR.n32 VPWR.n8 36.1417
R41 VPWR.n33 VPWR.n32 36.1417
R42 VPWR.n1 VPWR.t1 35.1791
R43 VPWR.n20 VPWR.n12 29.7417
R44 VPWR.n44 VPWR.t0 26.3844
R45 VPWR.n1 VPWR.t4 26.3844
R46 VPWR.n14 VPWR.t3 26.3844
R47 VPWR.n14 VPWR.t2 26.3844
R48 VPWR.n16 VPWR.n15 25.224
R49 VPWR.n52 VPWR.n51 20.7064
R50 VPWR.n16 VPWR.n12 17.6946
R51 VPWR.n35 VPWR.n33 15.0543
R52 VPWR.n17 VPWR.n16 9.3005
R53 VPWR.n18 VPWR.n12 9.3005
R54 VPWR.n20 VPWR.n19 9.3005
R55 VPWR.n21 VPWR.n11 9.3005
R56 VPWR.n23 VPWR.n22 9.3005
R57 VPWR.n24 VPWR.n10 9.3005
R58 VPWR.n26 VPWR.n25 9.3005
R59 VPWR.n27 VPWR.n9 9.3005
R60 VPWR.n29 VPWR.n28 9.3005
R61 VPWR.n30 VPWR.n8 9.3005
R62 VPWR.n32 VPWR.n31 9.3005
R63 VPWR.n33 VPWR.n7 9.3005
R64 VPWR.n37 VPWR.n36 9.3005
R65 VPWR.n40 VPWR.n39 9.3005
R66 VPWR.n38 VPWR.n4 9.3005
R67 VPWR.n46 VPWR.n3 9.3005
R68 VPWR.n48 VPWR.n47 9.3005
R69 VPWR.n50 VPWR.n49 9.3005
R70 VPWR.n51 VPWR.n0 9.3005
R71 VPWR.n53 VPWR.n52 9.3005
R72 VPWR.n47 VPWR.n2 8.28285
R73 VPWR.n46 VPWR.n45 7.33247
R74 VPWR.n15 VPWR.n13 6.59649
R75 VPWR.n42 VPWR.n41 3.92583
R76 VPWR.n45 VPWR.n4 3.24317
R77 VPWR.n40 VPWR.n6 3.12939
R78 VPWR.n50 VPWR.n2 3.01226
R79 VPWR.n36 VPWR.n6 2.33294
R80 VPWR.n36 VPWR.n35 1.59339
R81 VPWR.n41 VPWR.n40 0.853833
R82 VPWR.n42 VPWR.n4 0.683167
R83 VPWR.n17 VPWR.n13 0.612104
R84 VPWR.n18 VPWR.n17 0.122949
R85 VPWR.n19 VPWR.n18 0.122949
R86 VPWR.n19 VPWR.n11 0.122949
R87 VPWR.n23 VPWR.n11 0.122949
R88 VPWR.n24 VPWR.n23 0.122949
R89 VPWR.n25 VPWR.n24 0.122949
R90 VPWR.n25 VPWR.n9 0.122949
R91 VPWR.n29 VPWR.n9 0.122949
R92 VPWR.n30 VPWR.n29 0.122949
R93 VPWR.n31 VPWR.n30 0.122949
R94 VPWR.n31 VPWR.n7 0.122949
R95 VPWR.n37 VPWR.n7 0.122949
R96 VPWR.n39 VPWR.n37 0.122949
R97 VPWR.n39 VPWR.n38 0.122949
R98 VPWR.n38 VPWR.n3 0.122949
R99 VPWR.n48 VPWR.n3 0.122949
R100 VPWR.n49 VPWR.n48 0.122949
R101 VPWR.n49 VPWR.n0 0.122949
R102 VPWR.n53 VPWR.n0 0.122949
R103 VPWR VPWR.n53 0.0617245
R104 Y Y.n9 354.493
R105 Y.n6 Y.n5 299.95
R106 Y.n2 Y.n0 255.935
R107 Y.n9 Y.n7 216.463
R108 Y.n2 Y.n1 203.127
R109 Y.n4 Y.n3 201.392
R110 Y.n4 Y.n2 196.894
R111 Y.n9 Y.n8 185
R112 Y.n0 Y.t10 57.1657
R113 Y.n5 Y.t0 52.7684
R114 Y Y.n6 51.6752
R115 Y.n6 Y.n4 50.4476
R116 Y.n0 Y.t9 35.1791
R117 Y.n3 Y.t2 35.1791
R118 Y.n5 Y.t5 31.6612
R119 Y.n1 Y.t3 26.3844
R120 Y.n1 Y.t4 26.3844
R121 Y.n3 Y.t1 26.3844
R122 Y.n7 Y.t11 23.514
R123 Y.n8 Y.t7 22.7032
R124 Y.n8 Y.t8 22.7032
R125 Y.n7 Y.t6 22.7032
R126 VPB.t4 VPB.t3 1248.79
R127 VPB.t7 VPB.t14 515.861
R128 VPB.t13 VPB.t12 344.759
R129 VPB.t11 VPB.t1 321.774
R130 VPB.t10 VPB.t0 280.914
R131 VPB.t2 VPB.t11 265.591
R132 VPB VPB.t13 257.93
R133 VPB.t8 VPB.t10 255.376
R134 VPB.t3 VPB.t2 255.376
R135 VPB.t12 VPB.t5 255.376
R136 VPB.t9 VPB.t15 229.839
R137 VPB.t6 VPB.t9 229.839
R138 VPB.t14 VPB.t6 229.839
R139 VPB.t0 VPB.t7 229.839
R140 VPB.t1 VPB.t8 229.839
R141 VPB.t5 VPB.t4 229.839
R142 A2.n7 A2.t2 250.909
R143 A2.n3 A2.t4 248.316
R144 A2.n0 A2.t3 237.519
R145 A2.n9 A2.t0 226.809
R146 A2.n2 A2.n1 218.507
R147 A2.n10 A2.t1 196.013
R148 A2.n7 A2.n6 196.013
R149 A2 A2.n4 159.591
R150 A2.n0 A2.t5 156.662
R151 A2.n11 A2.n10 152
R152 A2.n8 A2.n5 152
R153 A2.n10 A2.n4 49.6611
R154 A2.n2 A2.n0 39.4369
R155 A2.n9 A2.n8 35.7853
R156 A2.n3 A2.n2 31.6183
R157 A2.n10 A2.n9 13.8763
R158 A2.n8 A2.n7 13.146
R159 A2.n11 A2.n5 10.1214
R160 A2.n4 A2.n3 6.90744
R161 A2 A2.n11 2.53073
R162 A2.n5 A2 1.63771
R163 a_1350_368.n2 a_1350_368.n0 350.735
R164 a_1350_368.n2 a_1350_368.n1 298.154
R165 a_1350_368.n4 a_1350_368.n3 247.745
R166 a_1350_368.n5 a_1350_368.n4 206.941
R167 a_1350_368.n4 a_1350_368.n2 79.0705
R168 a_1350_368.n0 a_1350_368.t4 35.1791
R169 a_1350_368.n3 a_1350_368.t7 26.3844
R170 a_1350_368.n3 a_1350_368.t5 26.3844
R171 a_1350_368.n0 a_1350_368.t1 26.3844
R172 a_1350_368.n1 a_1350_368.t3 26.3844
R173 a_1350_368.n1 a_1350_368.t2 26.3844
R174 a_1350_368.t0 a_1350_368.n5 26.3844
R175 a_1350_368.n5 a_1350_368.t6 26.3844
R176 a_841_368.n1 a_841_368.t2 379.57
R177 a_841_368.n4 a_841_368.t4 376.183
R178 a_841_368.n1 a_841_368.n0 302.74
R179 a_841_368.n3 a_841_368.n2 302.74
R180 a_841_368.n5 a_841_368.n4 302.74
R181 a_841_368.n3 a_841_368.n1 57.977
R182 a_841_368.n4 a_841_368.n3 50.4476
R183 a_841_368.n0 a_841_368.t1 35.1791
R184 a_841_368.n5 a_841_368.t3 35.1791
R185 a_841_368.t6 a_841_368.n5 35.1791
R186 a_841_368.n0 a_841_368.t7 29.9023
R187 a_841_368.n2 a_841_368.t5 26.3844
R188 a_841_368.n2 a_841_368.t0 26.3844
R189 A3.n5 A3.t6 240.685
R190 A3.n1 A3.t4 226.809
R191 A3.n12 A3.t2 226.809
R192 A3.n6 A3.t5 226.809
R193 A3.n1 A3.n0 198.204
R194 A3.n7 A3.t0 196.013
R195 A3.n4 A3.t1 196.013
R196 A3.n3 A3.t3 196.013
R197 A3.n9 A3.n5 172.725
R198 A3 A3.n2 156.207
R199 A3.n9 A3.n8 152
R200 A3.n14 A3.n13 152
R201 A3.n11 A3.n10 152
R202 A3.n12 A3.n11 35.7853
R203 A3.n3 A3.n2 32.1338
R204 A3.n8 A3.n7 32.1338
R205 A3.n2 A3.n1 28.4823
R206 A3.n6 A3.n4 21.1793
R207 A3.n11 A3.n4 18.9884
R208 A3.n13 A3.n3 17.5278
R209 A3.n7 A3.n5 17.5278
R210 A3.n10 A3.n9 16.7015
R211 A3.n13 A3.n12 13.8763
R212 A3.n8 A3.n6 9.49444
R213 A3.n14 A3 9.32621
R214 A3 A3.n14 8.22907
R215 A3.n10 A3 3.10907
R216 VGND.n12 VGND.n11 276.623
R217 VGND.n20 VGND.t3 233.304
R218 VGND.n28 VGND.t2 231.137
R219 VGND.n26 VGND.n2 201.097
R220 VGND.n13 VGND.n12 185
R221 VGND.n7 VGND.t5 169.025
R222 VGND.n16 VGND.n15 124.29
R223 VGND.n2 VGND.t0 35.6762
R224 VGND.n2 VGND.t1 35.6762
R225 VGND.n11 VGND.n7 30.9646
R226 VGND.n16 VGND.n4 28.2358
R227 VGND.n22 VGND.n1 27.8593
R228 VGND.n21 VGND.n20 27.1064
R229 VGND.n16 VGND.n14 25.224
R230 VGND.n26 VGND.n1 24.0946
R231 VGND.n27 VGND.n26 23.3417
R232 VGND.n14 VGND.n13 23.1201
R233 VGND.n12 VGND.t7 22.7032
R234 VGND.n15 VGND.t6 22.7032
R235 VGND.n15 VGND.t4 22.7032
R236 VGND.n28 VGND.n27 22.5887
R237 VGND.n20 VGND.n4 20.3299
R238 VGND.n22 VGND.n21 18.824
R239 VGND.n27 VGND.n0 9.3005
R240 VGND.n26 VGND.n25 9.3005
R241 VGND.n24 VGND.n1 9.3005
R242 VGND.n23 VGND.n22 9.3005
R243 VGND.n21 VGND.n3 9.3005
R244 VGND.n20 VGND.n19 9.3005
R245 VGND.n18 VGND.n4 9.3005
R246 VGND.n17 VGND.n16 9.3005
R247 VGND.n10 VGND.n9 9.3005
R248 VGND.n8 VGND.n6 9.3005
R249 VGND.n14 VGND.n5 9.3005
R250 VGND.n29 VGND.n28 7.20603
R251 VGND.n10 VGND.n6 7.02221
R252 VGND.n9 VGND.n7 2.34593
R253 VGND VGND.n29 1.13555
R254 VGND.n11 VGND.n10 0.658786
R255 VGND.n13 VGND.n6 0.585643
R256 VGND.n29 VGND.n0 0.156478
R257 VGND.n9 VGND.n8 0.122949
R258 VGND.n8 VGND.n5 0.122949
R259 VGND.n17 VGND.n5 0.122949
R260 VGND.n18 VGND.n17 0.122949
R261 VGND.n19 VGND.n18 0.122949
R262 VGND.n19 VGND.n3 0.122949
R263 VGND.n23 VGND.n3 0.122949
R264 VGND.n24 VGND.n23 0.122949
R265 VGND.n25 VGND.n24 0.122949
R266 VGND.n25 VGND.n0 0.122949
R267 a_459_74.n1 a_459_74.t9 237.489
R268 a_459_74.n7 a_459_74.n5 229.288
R269 a_459_74.n4 a_459_74.t2 207.703
R270 a_459_74.n7 a_459_74.n6 185
R271 a_459_74.n9 a_459_74.n8 185
R272 a_459_74.n3 a_459_74.t6 143.052
R273 a_459_74.n2 a_459_74.t5 141.873
R274 a_459_74.n8 a_459_74.n7 116.085
R275 a_459_74.n1 a_459_74.n0 102.019
R276 a_459_74.n2 a_459_74.n1 78.7732
R277 a_459_74.n3 a_459_74.n2 76.8659
R278 a_459_74.n4 a_459_74.n3 59.7954
R279 a_459_74.n8 a_459_74.n4 59.364
R280 a_459_74.n6 a_459_74.t8 23.514
R281 a_459_74.n6 a_459_74.t7 23.514
R282 a_459_74.n5 a_459_74.t0 22.7032
R283 a_459_74.n5 a_459_74.t1 22.7032
R284 a_459_74.n0 a_459_74.t11 22.7032
R285 a_459_74.n0 a_459_74.t10 22.7032
R286 a_459_74.n9 a_459_74.t3 22.7032
R287 a_459_74.t4 a_459_74.n9 22.7032
R288 VNB.t2 VNB.t6 3372.18
R289 VNB.t15 VNB.t13 3325.98
R290 VNB.t8 VNB.t4 2933.33
R291 VNB.t6 VNB.t5 2251.97
R292 VNB.t3 VNB.t2 1362.73
R293 VNB VNB.t12 1143.31
R294 VNB.t7 VNB.t8 1016.27
R295 VNB.t12 VNB.t10 1004.72
R296 VNB.t14 VNB.t15 993.177
R297 VNB.t5 VNB.t14 993.177
R298 VNB.t4 VNB.t3 993.177
R299 VNB.t0 VNB.t7 993.177
R300 VNB.t1 VNB.t0 993.177
R301 VNB.t11 VNB.t1 993.177
R302 VNB.t9 VNB.t11 993.177
R303 VNB.t10 VNB.t9 993.177
R304 A1.n6 A1.t4 378.882
R305 A1.n5 A1.t0 226.809
R306 A1.n7 A1.t1 226.809
R307 A1.n4 A1.t6 225.838
R308 A1.n0 A1.t3 206.876
R309 A1.n6 A1.t5 196.013
R310 A1 A1.n1 155.423
R311 A1.n13 A1.n12 152
R312 A1.n11 A1.n10 152
R313 A1.n9 A1.n8 152
R314 A1.n0 A1.t2 149.317
R315 A1.n3 A1.n2 147.814
R316 A1.n12 A1.n11 49.6611
R317 A1.n8 A1.n5 44.549
R318 A1.n3 A1.n1 25.1047
R319 A1.n8 A1.n7 21.1793
R320 A1.n1 A1.n0 18.0781
R321 A1.n7 A1.n6 11.6853
R322 A1.n10 A1.n9 10.1214
R323 A1.n13 A1 7.5912
R324 A1.n12 A1.n4 7.19579
R325 A1 A1.n13 6.69817
R326 A1.n11 A1.n5 5.11262
R327 A1.n10 A1 2.53073
R328 A1.n9 A1 1.63771
R329 A1.n4 A1.n3 1.43996
R330 B1.n2 B1.t3 324.82
R331 B1.n2 B1.t2 218.602
R332 B1.n9 B1.t1 207.582
R333 B1.n3 B1.t5 196.013
R334 B1.n1 B1.t4 196.013
R335 B1.n7 B1.t0 196.013
R336 B1 B1.n4 157.304
R337 B1.n10 B1.n9 152
R338 B1.n8 B1.n0 152
R339 B1.n6 B1.n5 152
R340 B1.n9 B1.n8 43.7018
R341 B1.n7 B1.n6 42.4165
R342 B1.n4 B1.n1 30.8485
R343 B1.n4 B1.n3 24.4218
R344 B1.n6 B1.n1 12.8538
R345 B1.n10 B1.n0 12.4348
R346 B1.n5 B1 10.4234
R347 B1.n5 B1 7.13193
R348 B1.n3 B1.n2 6.09085
R349 B1 B1.n10 3.10907
R350 B1 B1.n0 2.01193
R351 B1.n8 B1.n7 1.28583
R352 a_27_74.n4 a_27_74.t2 276.978
R353 a_27_74.n1 a_27_74.t7 189.156
R354 a_27_74.n1 a_27_74.n0 185
R355 a_27_74.n3 a_27_74.n2 185
R356 a_27_74.n5 a_27_74.n4 185
R357 a_27_74.n4 a_27_74.n3 73.4123
R358 a_27_74.n3 a_27_74.n1 46.6678
R359 a_27_74.n2 a_27_74.t0 22.7032
R360 a_27_74.n2 a_27_74.t6 22.7032
R361 a_27_74.n0 a_27_74.t4 22.7032
R362 a_27_74.n0 a_27_74.t5 22.7032
R363 a_27_74.t3 a_27_74.n5 22.7032
R364 a_27_74.n5 a_27_74.t1 22.7032
C0 VGND A3 0.056577f
C1 VPB B1 0.149566f
C2 Y A2 0.052686f
C3 A1 Y 1.75e-19
C4 VPWR C1 0.078602f
C5 Y VPB 0.031383f
C6 B1 A3 0.034381f
C7 VGND B1 0.025792f
C8 VPWR A2 0.025901f
C9 Y A3 0.43758f
C10 Y VGND 0.045397f
C11 A1 VPWR 0.084207f
C12 VPWR VPB 0.289994f
C13 VPB C1 0.101554f
C14 A1 A2 0.050151f
C15 Y B1 0.426069f
C16 VPWR A3 0.026132f
C17 C1 A3 1.83e-19
C18 VPB A2 0.150944f
C19 VPWR VGND 0.191716f
C20 C1 VGND 0.025922f
C21 A1 VPB 0.167886f
C22 A3 A2 0.048681f
C23 VGND A2 0.072102f
C24 VPWR B1 0.051781f
C25 VPB A3 0.164605f
C26 C1 B1 0.074059f
C27 A1 VGND 0.082469f
C28 VPB VGND 0.015233f
C29 VPWR Y 0.585832f
C30 Y C1 0.182121f
C31 VGND VNB 1.26414f
C32 Y VNB 0.060312f
C33 VPWR VNB 1.05187f
C34 A1 VNB 0.500495f
C35 A2 VNB 0.414243f
C36 A3 VNB 0.44122f
C37 B1 VNB 0.40081f
C38 C1 VNB 0.40776f
C39 VPB VNB 2.54894f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o311ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311ai_2 VNB VPB VPWR VGND A2 A3 C1 B1 Y A1
X0 a_28_368.t2 A1.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.1736 ps=1.43 w=1.12 l=0.15
X1 a_27_74.t1 A3.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1147 ps=1.05 w=0.74 l=0.15
X2 VPWR.t2 A1.t1 a_28_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_670_74.t1 C1.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 VGND.t5 A1.t2 a_27_74.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 Y.t3 C1.t1 a_670_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VPWR.t4 C1.t2 Y.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_307_368.t3 A2.t0 a_28_368.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2072 pd=1.49 as=0.1904 ps=1.46 w=1.12 l=0.15
X8 Y.t4 B1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t1 C1.t3 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VPWR.t5 B1.t1 Y.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t5 A3.t1 a_307_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_307_368.t0 A3.t2 Y.t6 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X13 VGND.t2 A2.t1 a_27_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1258 ps=1.08 w=0.74 l=0.15
X14 VGND.t0 A3.t3 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X15 a_27_74.t5 B1.t2 a_670_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 a_27_74.t3 A2.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1073 ps=1.03 w=0.74 l=0.15
X17 a_27_74.t6 A1.t3 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1258 ps=1.08 w=0.74 l=0.15
X18 a_28_368.t0 A2.t3 a_307_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2072 ps=1.49 w=1.12 l=0.15
X19 a_670_74.t2 B1.t3 a_27_74.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A1.n0 A1.t0 226.809
R1 A1.n1 A1.t1 226.809
R2 A1.n1 A1.t2 198.204
R3 A1.n0 A1.t3 198.204
R4 A1.n3 A1.n2 152
R5 A1.n2 A1.n0 56.2338
R6 A1.n3 A1 12.8005
R7 A1.n2 A1.n1 10.955
R8 A1 A1.n3 1.48887
R9 VPWR.n7 VPWR.n6 329.116
R10 VPWR.n17 VPWR.n1 323.406
R11 VPWR.n5 VPWR.n4 315.928
R12 VPWR.n10 VPWR.n9 36.1417
R13 VPWR.n11 VPWR.n10 36.1417
R14 VPWR.n11 VPWR.n2 36.1417
R15 VPWR.n15 VPWR.n2 36.1417
R16 VPWR.n16 VPWR.n15 36.1417
R17 VPWR.n1 VPWR.t3 28.1434
R18 VPWR.n1 VPWR.t2 26.3844
R19 VPWR.n4 VPWR.t1 26.3844
R20 VPWR.n4 VPWR.t5 26.3844
R21 VPWR.n6 VPWR.t0 26.3844
R22 VPWR.n6 VPWR.t4 26.3844
R23 VPWR.n9 VPWR.n5 26.3534
R24 VPWR.n17 VPWR.n16 22.5887
R25 VPWR.n9 VPWR.n8 9.3005
R26 VPWR.n10 VPWR.n3 9.3005
R27 VPWR.n12 VPWR.n11 9.3005
R28 VPWR.n13 VPWR.n2 9.3005
R29 VPWR.n15 VPWR.n14 9.3005
R30 VPWR.n16 VPWR.n0 9.3005
R31 VPWR.n18 VPWR.n17 7.53404
R32 VPWR.n7 VPWR.n5 6.51247
R33 VPWR.n8 VPWR.n7 0.610428
R34 VPWR VPWR.n18 0.161409
R35 VPWR.n18 VPWR.n0 0.146411
R36 VPWR.n8 VPWR.n3 0.122949
R37 VPWR.n12 VPWR.n3 0.122949
R38 VPWR.n13 VPWR.n12 0.122949
R39 VPWR.n14 VPWR.n13 0.122949
R40 VPWR.n14 VPWR.n0 0.122949
R41 a_28_368.n0 a_28_368.t0 432.118
R42 a_28_368.n0 a_28_368.t1 278.553
R43 a_28_368.n1 a_28_368.n0 205.486
R44 a_28_368.t2 a_28_368.n1 33.4201
R45 a_28_368.n1 a_28_368.t3 26.3844
R46 VPB.t3 VPB.t0 515.861
R47 VPB.t8 VPB.t3 265.591
R48 VPB VPB.t5 260.485
R49 VPB.t6 VPB.t8 250.269
R50 VPB.t5 VPB.t6 234.946
R51 VPB.t7 VPB.t1 229.839
R52 VPB.t2 VPB.t7 229.839
R53 VPB.t9 VPB.t2 229.839
R54 VPB.t4 VPB.t9 229.839
R55 VPB.t0 VPB.t4 229.839
R56 A3.n0 A3.t1 344.932
R57 A3.n2 A3.t3 235.216
R58 A3.n0 A3.t2 203.612
R59 A3.n1 A3.t0 196.013
R60 A3.n3 A3.n2 152
R61 A3.n1 A3.n0 26.1078
R62 A3.n2 A3.n1 19.9232
R63 A3 A3.n3 10.2703
R64 A3.n3 A3 4.0191
R65 VGND.n2 VGND.n1 213.653
R66 VGND.n4 VGND.n3 208.079
R67 VGND.n7 VGND.n6 208.079
R68 VGND.n6 VGND.t4 32.4329
R69 VGND.n1 VGND.t0 27.5681
R70 VGND.n5 VGND.n4 25.224
R71 VGND.n7 VGND.n5 24.4711
R72 VGND.n3 VGND.t2 24.3248
R73 VGND.n1 VGND.t1 22.7032
R74 VGND.n3 VGND.t3 22.7032
R75 VGND.n6 VGND.t5 22.7032
R76 VGND.n5 VGND.n0 9.3005
R77 VGND.n8 VGND.n7 7.19894
R78 VGND.n4 VGND.n2 6.62585
R79 VGND.n2 VGND.n0 0.566682
R80 VGND VGND.n8 0.156997
R81 VGND.n8 VGND.n0 0.150766
R82 a_27_74.n4 a_27_74.t5 267.265
R83 a_27_74.n1 a_27_74.t7 208.529
R84 a_27_74.n1 a_27_74.n0 104.579
R85 a_27_74.n3 a_27_74.n2 104.579
R86 a_27_74.n5 a_27_74.n4 104.579
R87 a_27_74.n3 a_27_74.n1 51.2005
R88 a_27_74.n4 a_27_74.n3 51.2005
R89 a_27_74.n0 a_27_74.t2 32.4329
R90 a_27_74.n2 a_27_74.t0 29.1897
R91 a_27_74.n0 a_27_74.t6 22.7032
R92 a_27_74.n2 a_27_74.t3 22.7032
R93 a_27_74.n5 a_27_74.t4 22.7032
R94 a_27_74.t1 a_27_74.n5 22.7032
R95 VNB.t7 VNB.t0 2286.61
R96 VNB.t6 VNB.t7 1316.54
R97 VNB VNB.t9 1143.31
R98 VNB.t8 VNB.t3 1131.76
R99 VNB.t9 VNB.t8 1131.76
R100 VNB.t4 VNB.t1 1085.56
R101 VNB.t1 VNB.t2 1062.47
R102 VNB.t3 VNB.t4 1016.27
R103 VNB.t0 VNB.t5 993.177
R104 VNB.t2 VNB.t6 993.177
R105 C1.n3 C1.t2 246.769
R106 C1.n2 C1.t3 240.197
R107 C1.n3 C1.t0 179.947
R108 C1.n1 C1.t1 179.947
R109 C1.n1 C1.n0 176.101
R110 C1.n5 C1.n4 152
R111 C1.n4 C1.n3 37.246
R112 C1.n4 C1.n2 21.9096
R113 C1.n5 C1.n0 9.06717
R114 C1.n2 C1.n1 3.65202
R115 C1 C1.n5 3.6005
R116 C1.n0 C1 0.133833
R117 Y.n1 Y.t6 418.31
R118 Y.n2 Y.t1 274.788
R119 Y.n5 Y.t0 210.159
R120 Y.n1 Y.n0 208.776
R121 Y.n4 Y.n3 208.274
R122 Y.n6 Y.t3 199.569
R123 Y.n2 Y.n1 48.9417
R124 Y.n0 Y.t7 26.3844
R125 Y.n0 Y.t5 26.3844
R126 Y.n3 Y.t2 26.3844
R127 Y.n3 Y.t4 26.3844
R128 Y Y.n4 16.9549
R129 Y Y.n6 6.4005
R130 Y.n5 Y 4.65505
R131 Y.n6 Y.n5 3.29747
R132 Y.n5 Y 2.63064
R133 Y.n4 Y.n2 0.691466
R134 a_670_74.n1 a_670_74.n0 476.154
R135 a_670_74.n0 a_670_74.t3 34.0546
R136 a_670_74.n0 a_670_74.t2 34.0546
R137 a_670_74.n1 a_670_74.t0 22.7032
R138 a_670_74.t1 a_670_74.n1 22.7032
R139 A2.n0 A2.t3 236.303
R140 A2.n1 A2.t0 228.877
R141 A2.n1 A2.t1 196.013
R142 A2.n0 A2.t2 196.013
R143 A2.n5 A2.n4 152
R144 A2.n3 A2.n2 152
R145 A2.n4 A2.n3 49.6611
R146 A2.n2 A2 13.3958
R147 A2.n3 A2.n1 13.146
R148 A2.n5 A2 9.22841
R149 A2 A2.n5 5.06097
R150 A2.n4 A2.n0 1.46111
R151 A2.n2 A2 0.893523
R152 a_307_368.n1 a_307_368.n0 706.144
R153 a_307_368.n0 a_307_368.t3 38.6969
R154 a_307_368.n0 a_307_368.t2 26.3844
R155 a_307_368.t1 a_307_368.n1 26.3844
R156 a_307_368.n1 a_307_368.t0 26.3844
R157 B1.n1 B1.t3 302.053
R158 B1.n0 B1.t0 295.091
R159 B1.n0 B1.t1 237.762
R160 B1.n1 B1.t2 153.948
R161 B1.n3 B1.n2 152
R162 B1.n2 B1.n1 37.246
R163 B1.n2 B1.n0 13.146
R164 B1.n3 B1 12.5028
R165 B1 B1.n3 1.78655
C0 A2 Y 2.43e-19
C1 A3 VPWR 0.018669f
C2 B1 C1 0.037933f
C3 Y VGND 0.050235f
C4 Y A1 1.32e-19
C5 A2 VPB 0.072144f
C6 A3 B1 0.10549f
C7 VGND VPB 0.0087f
C8 VPB A1 0.066845f
C9 A2 VPWR 0.017954f
C10 VPWR VGND 0.090547f
C11 Y VPB 0.025613f
C12 VPWR A1 0.036714f
C13 VPWR Y 0.402606f
C14 B1 VGND 0.019242f
C15 C1 VGND 0.017192f
C16 VPWR VPB 0.143624f
C17 B1 Y 0.138f
C18 C1 Y 0.239956f
C19 A2 A3 0.083363f
C20 A3 VGND 0.037882f
C21 B1 VPB 0.068174f
C22 C1 VPB 0.077024f
C23 B1 VPWR 0.042248f
C24 A3 Y 0.094136f
C25 C1 VPWR 0.037168f
C26 A2 VGND 0.038099f
C27 A3 VPB 0.096177f
C28 A2 A1 0.083765f
C29 VGND A1 0.037138f
C30 VGND VNB 0.668183f
C31 Y VNB 0.110368f
C32 VPWR VNB 0.542914f
C33 C1 VNB 0.274293f
C34 B1 VNB 0.25019f
C35 A3 VNB 0.22619f
C36 A2 VNB 0.201606f
C37 A1 VNB 0.244366f
C38 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o311ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311ai_1 VNB VPB VPWR VGND A2 A1 C1 B1 Y A3
X0 Y.t1 C1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X1 a_128_74.t3 A3.t0 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.222 ps=1.34 w=0.74 l=0.15
X2 a_128_74.t2 A1.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.2627 ps=2.19 w=0.74 l=0.15
X3 a_222_368.t1 A2.t0 a_138_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X4 VGND.t0 A2.t1 a_128_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=1.34 as=0.11285 ps=1.045 w=0.74 l=0.15
X5 a_138_368.t0 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 Y.t2 A3.t1 a_222_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X7 a_469_74.t1 B1.t0 a_128_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 VPWR.t2 B1.t1 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X9 Y.t0 C1.t1 a_469_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1147 ps=1.05 w=0.74 l=0.15
R0 C1.n0 C1.t0 261.62
R1 C1 C1.n0 209.179
R2 C1.n0 C1.t1 156.431
R3 VPWR.n1 VPWR.t1 255.061
R4 VPWR.n1 VPWR.n0 228.386
R5 VPWR.n0 VPWR.t0 38.6969
R6 VPWR.n0 VPWR.t2 35.1791
R7 VPWR VPWR.n1 0.114608
R8 Y.n4 Y.n3 585
R9 Y.n3 Y.n0 291.286
R10 Y.n2 Y.n1 252.492
R11 Y.n2 Y.t0 193.363
R12 Y.n1 Y.t2 47.4916
R13 Y.n3 Y.t1 26.3844
R14 Y.n1 Y.t3 26.3844
R15 Y Y.n2 14.4815
R16 Y Y.n4 9.97259
R17 Y Y.n0 6.65358
R18 Y.n0 Y 4.29935
R19 Y.n4 Y 1.04236
R20 VPB VPB.t2 314.113
R21 VPB.t4 VPB.t0 291.13
R22 VPB.t1 VPB.t4 291.13
R23 VPB.t3 VPB.t1 291.13
R24 VPB.t2 VPB.t3 214.517
R25 A3.n0 A3.t1 285.719
R26 A3.n0 A3.t0 178.34
R27 A3 A3.n0 158.788
R28 VGND.n1 VGND.n0 190.899
R29 VGND.n1 VGND.t1 161.46
R30 VGND.n0 VGND.t0 50.2708
R31 VGND.n0 VGND.t2 47.0275
R32 VGND VGND.n1 0.328559
R33 a_128_74.n1 a_128_74.n0 264.375
R34 a_128_74.n1 a_128_74.t3 34.0546
R35 a_128_74.n0 a_128_74.t1 26.7573
R36 a_128_74.n0 a_128_74.t2 22.7032
R37 a_128_74.t0 a_128_74.n1 22.7032
R38 VNB.t2 VNB.t4 1732.28
R39 VNB VNB.t3 1304.99
R40 VNB.t4 VNB.t0 1154.86
R41 VNB.t0 VNB.t1 1062.47
R42 VNB.t3 VNB.t2 1050.92
R43 A1.n0 A1.t1 250.909
R44 A1.n0 A1.t0 220.113
R45 A1 A1.n0 163.46
R46 A2.n0 A2.t0 250.909
R47 A2.n0 A2.t1 220.113
R48 A2 A2.n0 154.25
R49 a_138_368.t0 a_138_368.t1 47.4916
R50 a_222_368.t0 a_222_368.t1 73.8755
R51 B1.n0 B1.t1 285.719
R52 B1.n0 B1.t0 178.34
R53 B1 B1.n0 158.054
R54 a_469_74.t0 a_469_74.t1 50.2708
C0 VGND VPWR 0.055981f
C1 B1 VPWR 0.017068f
C2 A2 VPWR 0.08544f
C3 VPWR VPB 0.104796f
C4 VGND B1 0.014466f
C5 VGND A2 0.017834f
C6 B1 A2 5.28e-19
C7 VGND VPB 0.007281f
C8 B1 VPB 0.032224f
C9 A2 VPB 0.037432f
C10 C1 VPWR 0.018547f
C11 Y VPWR 0.281111f
C12 VGND C1 0.009746f
C13 B1 C1 0.051084f
C14 A3 VPWR 0.013642f
C15 A1 VPWR 0.056467f
C16 C1 VPB 0.046338f
C17 Y VGND 0.06319f
C18 VGND A3 0.015438f
C19 Y B1 0.092293f
C20 VGND A1 0.04753f
C21 Y A2 0.055261f
C22 A3 B1 0.077833f
C23 A3 A2 0.071594f
C24 A1 A2 0.095021f
C25 Y VPB 0.026332f
C26 A3 VPB 0.032733f
C27 A1 VPB 0.03984f
C28 Y C1 0.131946f
C29 Y A3 0.020386f
C30 Y A1 1.61e-19
C31 A3 A1 3.79e-19
C32 VGND VNB 0.466617f
C33 Y VNB 0.099359f
C34 VPWR VNB 0.391062f
C35 C1 VNB 0.180891f
C36 B1 VNB 0.107206f
C37 A3 VNB 0.114802f
C38 A2 VNB 0.111858f
C39 A1 VNB 0.15394f
C40 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o311a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311a_4 VNB VPB VPWR VGND C1 B1 A3 A2 A1 X
X0 VPWR.t6 a_83_244.t7 X.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.2716 ps=1.605 w=1.12 l=0.15
X1 X.t5 a_83_244.t8 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_564_78.t4 A3.t0 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0912 pd=0.925 as=0.1232 ps=1.025 w=0.64 l=0.15
X3 VPWR.t7 C1.t0 a_83_244.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3575 pd=1.715 as=0.21 ps=1.42 w=1 l=0.15
X4 a_1034_392.t1 A2.t0 a_1338_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.325 pd=2.65 as=0.16 ps=1.32 w=1 l=0.15
X5 VPWR.t1 B1.t0 a_83_244.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X6 X.t7 a_83_244.t9 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.20165 ps=1.285 w=0.74 l=0.15
X7 a_83_244.t2 C1.t1 a_651_78.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.171975 pd=1.295 as=0.2544 ps=1.435 w=0.64 l=0.15
X8 a_564_78.t5 A1.t0 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1216 pd=1.02 as=0.12 ps=1.015 w=0.64 l=0.15
X9 X.t4 a_83_244.t10 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2716 pd=1.605 as=0.196 ps=1.47 w=1.12 l=0.15
X10 a_1338_392.t1 A2.t1 a_1034_392.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.1525 ps=1.305 w=1 l=0.15
X11 X.t6 a_83_244.t11 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X12 a_1338_392.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.15 ps=1.3 w=1 l=0.15
X13 VPWR.t9 A1.t2 a_1338_392.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.21 ps=1.42 w=1 l=0.15
X14 a_83_244.t3 C1.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.3575 ps=1.715 w=1 l=0.15
X15 a_564_78.t6 B1.t1 a_651_78.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1216 pd=1.02 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 a_83_244.t1 A3.t1 a_1034_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.445 ps=2.89 w=1 l=0.15
X17 VGND.t6 A3.t2 a_564_78.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1232 pd=1.025 as=0.1216 ps=1.02 w=0.64 l=0.15
X18 VPWR.t3 a_83_244.t12 X.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VGND.t4 A2.t2 a_564_78.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12 pd=1.015 as=0.0912 ps=0.925 w=0.64 l=0.15
X20 VGND.t1 a_83_244.t13 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.20165 pd=1.285 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 a_651_78.t2 C1.t3 a_83_244.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.171975 ps=1.295 w=0.64 l=0.15
X22 a_651_78.t0 B1.t2 a_564_78.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2544 pd=1.435 as=0.178025 ps=1.85 w=0.64 l=0.15
X23 a_83_244.t6 B1.t3 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.1934 ps=1.475 w=1 l=0.15
X24 VGND.t0 a_83_244.t14 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X25 a_564_78.t2 A2.t3 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0944 ps=0.935 w=0.64 l=0.15
R0 a_83_244.n2 a_83_244.t1 815.446
R1 a_83_244.n2 a_83_244.n1 346.247
R2 a_83_244.n5 a_83_244.t8 270.384
R3 a_83_244.n0 a_83_244.t7 261.62
R4 a_83_244.n9 a_83_244.t10 261.62
R5 a_83_244.n6 a_83_244.t12 261.62
R6 a_83_244.n13 a_83_244.n3 205.202
R7 a_83_244.n15 a_83_244.n14 204.425
R8 a_83_244.n0 a_83_244.t14 167.386
R9 a_83_244.n8 a_83_244.n4 165.189
R10 a_83_244.n5 a_83_244.t11 154.24
R11 a_83_244.n7 a_83_244.t13 154.24
R12 a_83_244.n10 a_83_244.t9 154.24
R13 a_83_244.n11 a_83_244.n4 152
R14 a_83_244.n12 a_83_244.n0 152
R15 a_83_244.n14 a_83_244.n2 89.3033
R16 a_83_244.n14 a_83_244.n13 83.9763
R17 a_83_244.n8 a_83_244.n7 62.0763
R18 a_83_244.n13 a_83_244.n12 60.5895
R19 a_83_244.n6 a_83_244.n5 56.9641
R20 a_83_244.n3 a_83_244.t5 53.1905
R21 a_83_244.n0 a_83_244.n11 49.6611
R22 a_83_244.n1 a_83_244.t4 41.2505
R23 a_83_244.n1 a_83_244.t2 41.2505
R24 a_83_244.t0 a_83_244.n15 39.4005
R25 a_83_244.n10 a_83_244.n9 34.3247
R26 a_83_244.n3 a_83_244.t6 29.5505
R27 a_83_244.n15 a_83_244.t3 29.5505
R28 a_83_244.n12 a_83_244.n4 13.1884
R29 a_83_244.n11 a_83_244.n10 10.2247
R30 a_83_244.n7 a_83_244.n6 5.84292
R31 a_83_244.n9 a_83_244.n8 5.11262
R32 X.n5 X.n3 261.149
R33 X.n5 X.n4 210.702
R34 X.n2 X.n0 158.917
R35 X.n2 X.n1 96.6686
R36 X.n3 X.t0 50.13
R37 X.n6 X.n5 44.0431
R38 X.n3 X.t4 35.1791
R39 X.n0 X.t1 34.0546
R40 X.n6 X.n2 29.6618
R41 X.n4 X.t3 26.3844
R42 X.n4 X.t5 26.3844
R43 X.n1 X.t2 22.7032
R44 X.n1 X.t6 22.7032
R45 X.n0 X.t7 22.7032
R46 X X.n6 0.835283
R47 VPWR.n7 VPWR.n6 748.833
R48 VPWR.n7 VPWR.t1 318.791
R49 VPWR.n19 VPWR.t5 259.171
R50 VPWR.n17 VPWR.n2 221.766
R51 VPWR.n4 VPWR.n3 221.766
R52 VPWR.n10 VPWR.n9 139.442
R53 VPWR.n9 VPWR.t7 65.4173
R54 VPWR.n9 VPWR.t2 65.417
R55 VPWR.n3 VPWR.t8 40.3855
R56 VPWR.n12 VPWR.n11 36.1417
R57 VPWR.n16 VPWR.n4 35.3887
R58 VPWR.n2 VPWR.t3 35.1791
R59 VPWR.n8 VPWR.n7 32.5777
R60 VPWR.n6 VPWR.t0 29.5505
R61 VPWR.n6 VPWR.t9 29.5505
R62 VPWR.n3 VPWR.t6 27.6909
R63 VPWR.n19 VPWR.n18 26.7299
R64 VPWR.n2 VPWR.t4 26.3844
R65 VPWR.n18 VPWR.n17 25.977
R66 VPWR.n17 VPWR.n16 21.4593
R67 VPWR.n12 VPWR.n4 12.0476
R68 VPWR.n11 VPWR.n5 9.3005
R69 VPWR.n13 VPWR.n12 9.3005
R70 VPWR.n14 VPWR.n4 9.3005
R71 VPWR.n16 VPWR.n15 9.3005
R72 VPWR.n17 VPWR.n1 9.3005
R73 VPWR.n18 VPWR.n0 9.3005
R74 VPWR.n20 VPWR.n19 9.3005
R75 VPWR.n11 VPWR.n10 7.90638
R76 VPWR.n10 VPWR.n8 5.96639
R77 VPWR.n8 VPWR.n5 0.486035
R78 VPWR.n13 VPWR.n5 0.122949
R79 VPWR.n14 VPWR.n13 0.122949
R80 VPWR.n15 VPWR.n14 0.122949
R81 VPWR.n15 VPWR.n1 0.122949
R82 VPWR.n1 VPWR.n0 0.122949
R83 VPWR.n20 VPWR.n0 0.122949
R84 VPWR VPWR.n20 0.0617245
R85 VPB.t1 VPB.t2 592.473
R86 VPB.t2 VPB.t10 472.447
R87 VPB.t9 VPB.t3 441.801
R88 VPB.t6 VPB.t8 324.329
R89 VPB.t10 VPB.t12 291.13
R90 VPB.t11 VPB.t9 291.13
R91 VPB.t8 VPB.t11 257.93
R92 VPB VPB.t7 257.93
R93 VPB.t3 VPB.t1 255.376
R94 VPB.t5 VPB.t6 255.376
R95 VPB.t0 VPB.t4 240.054
R96 VPB.t12 VPB.t0 229.839
R97 VPB.t7 VPB.t5 229.839
R98 A3.n1 A3.t0 237.151
R99 A3.n2 A3.t2 230.339
R100 A3.n1 A3.n0 220.917
R101 A3.n2 A3.t1 220.917
R102 A3 A3.n3 156.268
R103 A3.n3 A3.n2 50.3914
R104 A3.n3 A3.n1 18.2581
R105 VGND.n8 VGND.t5 282.632
R106 VGND.n10 VGND.n9 205.752
R107 VGND.n13 VGND.n12 205.752
R108 VGND.n30 VGND.n2 199.488
R109 VGND.n25 VGND.t0 154.839
R110 VGND.n32 VGND.t2 140.934
R111 VGND.n2 VGND.t3 44.5951
R112 VGND.n2 VGND.t1 43.7843
R113 VGND.n9 VGND.t4 39.3755
R114 VGND.n12 VGND.t7 38.438
R115 VGND.n17 VGND.n6 36.1417
R116 VGND.n18 VGND.n17 36.1417
R117 VGND.n19 VGND.n18 36.1417
R118 VGND.n19 VGND.n4 36.1417
R119 VGND.n23 VGND.n4 36.1417
R120 VGND.n24 VGND.n23 36.1417
R121 VGND.n26 VGND.n1 36.1417
R122 VGND.n12 VGND.t6 33.7505
R123 VGND.n9 VGND.t8 30.938
R124 VGND.n31 VGND.n30 29.7417
R125 VGND.n13 VGND.n11 28.9887
R126 VGND.n11 VGND.n10 21.4593
R127 VGND.n32 VGND.n31 20.7064
R128 VGND.n13 VGND.n6 18.4476
R129 VGND.n33 VGND.n32 9.3005
R130 VGND.n31 VGND.n0 9.3005
R131 VGND.n30 VGND.n29 9.3005
R132 VGND.n28 VGND.n1 9.3005
R133 VGND.n27 VGND.n26 9.3005
R134 VGND.n11 VGND.n7 9.3005
R135 VGND.n14 VGND.n13 9.3005
R136 VGND.n15 VGND.n6 9.3005
R137 VGND.n17 VGND.n16 9.3005
R138 VGND.n18 VGND.n5 9.3005
R139 VGND.n20 VGND.n19 9.3005
R140 VGND.n21 VGND.n4 9.3005
R141 VGND.n23 VGND.n22 9.3005
R142 VGND.n24 VGND.n3 9.3005
R143 VGND.n30 VGND.n1 8.28285
R144 VGND.n10 VGND.n8 6.88087
R145 VGND.n26 VGND.n25 6.02403
R146 VGND.n25 VGND.n24 5.27109
R147 VGND.n8 VGND.n7 0.513127
R148 VGND.n14 VGND.n7 0.122949
R149 VGND.n15 VGND.n14 0.122949
R150 VGND.n16 VGND.n15 0.122949
R151 VGND.n16 VGND.n5 0.122949
R152 VGND.n20 VGND.n5 0.122949
R153 VGND.n21 VGND.n20 0.122949
R154 VGND.n22 VGND.n21 0.122949
R155 VGND.n22 VGND.n3 0.122949
R156 VGND.n27 VGND.n3 0.122949
R157 VGND.n28 VGND.n27 0.122949
R158 VGND.n29 VGND.n28 0.122949
R159 VGND.n29 VGND.n0 0.122949
R160 VGND.n33 VGND.n0 0.122949
R161 VGND VGND.n33 0.0617245
R162 a_564_78.n1 a_564_78.t0 398.193
R163 a_564_78.n2 a_564_78.t2 185.756
R164 a_564_78.n2 a_564_78.t5 130.553
R165 a_564_78.n4 a_564_78.n3 95.7887
R166 a_564_78.n1 a_564_78.n0 89.3175
R167 a_564_78.n3 a_564_78.n1 56.8151
R168 a_564_78.n3 a_564_78.n2 50.4476
R169 a_564_78.n0 a_564_78.t6 39.3755
R170 a_564_78.n0 a_564_78.t3 31.8755
R171 a_564_78.t4 a_564_78.n4 27.188
R172 a_564_78.n4 a_564_78.t1 26.2505
R173 VNB.t3 VNB.t0 2286.61
R174 VNB.t11 VNB.t8 2251.97
R175 VNB.t0 VNB.t1 2182.68
R176 VNB.t4 VNB.t6 1605.25
R177 VNB.t1 VNB.t2 1362.73
R178 VNB VNB.t5 1304.99
R179 VNB.t9 VNB.t10 1235.7
R180 VNB.t12 VNB.t9 1224.15
R181 VNB.t7 VNB.t11 1212.6
R182 VNB.t6 VNB.t3 1154.86
R183 VNB.t10 VNB.t7 1004.72
R184 VNB.t2 VNB.t12 993.177
R185 VNB.t5 VNB.t4 993.177
R186 C1.n0 C1.t3 369.625
R187 C1.n2 C1.t0 331.976
R188 C1.n1 C1.t2 216.9
R189 C1.n0 C1.t1 196.013
R190 C1 C1.n2 157.381
R191 C1.n2 C1.n1 40.0769
R192 C1.n1 C1.n0 10.2904
R193 A2.n2 A2.t0 312.125
R194 A2.n0 A2.t1 298.572
R195 A2.n1 A2.n0 255.714
R196 A2.n0 A2.t2 187.981
R197 A2.n2 A2.t3 154.405
R198 A2.n3 A2.n2 152
R199 A2 A2.n3 10.6672
R200 A2.n3 A2.n1 3.49141
R201 A2.n1 A2 0.194439
R202 a_1338_392.n1 a_1338_392.n0 951.438
R203 a_1338_392.n0 a_1338_392.t1 45.3105
R204 a_1338_392.n0 a_1338_392.t3 37.4305
R205 a_1338_392.n1 a_1338_392.t2 33.4905
R206 a_1338_392.t0 a_1338_392.n1 29.5505
R207 a_1034_392.n0 a_1034_392.t0 807.837
R208 a_1034_392.n0 a_1034_392.t2 781.587
R209 a_1034_392.t1 a_1034_392.n0 374.07
R210 B1.n0 B1.t0 365.2
R211 B1 B1.n1 338.467
R212 B1.n1 B1.t3 298.572
R213 B1.n1 B1.t2 287.885
R214 B1.n0 B1.t1 268.313
R215 B1 B1.n0 161.31
R216 a_651_78.n1 a_651_78.n0 328.635
R217 a_651_78.n0 a_651_78.t0 75.2294
R218 a_651_78.n0 a_651_78.t3 59.0447
R219 a_651_78.t1 a_651_78.n1 26.2505
R220 a_651_78.n1 a_651_78.t2 26.2505
R221 A1.n1 A1.n0 253.708
R222 A1.n2 A1.t0 246.405
R223 A1.n1 A1.t1 207.529
R224 A1.n2 A1.t2 207.529
R225 A1.n3 A1 155.298
R226 A1.n5 A1.n4 152
R227 A1.n4 A1.n3 49.6611
R228 A1.n3 A1.n2 12.4157
R229 A1.n5 A1 9.89141
R230 A1 A1.n5 8.72777
R231 A1.n4 A1.n1 3.65202
C0 C1 VGND 0.014109f
C1 VGND A1 0.027515f
C2 B1 X 0.003085f
C3 A3 A2 0.081676f
C4 A2 VPWR 0.054012f
C5 VPWR X 0.453021f
C6 B1 A3 0.053656f
C7 VPB A2 0.090182f
C8 VPB X 0.014436f
C9 B1 VPWR 0.041606f
C10 VPB B1 0.139765f
C11 A2 VGND 0.034841f
C12 VGND X 0.34081f
C13 B1 VGND 0.032405f
C14 A2 A1 0.265411f
C15 C1 X 1.14e-20
C16 A3 VPWR 0.036365f
C17 B1 C1 0.233235f
C18 VPB A3 0.080136f
C19 VPB VPWR 0.23422f
C20 A3 VGND 0.027311f
C21 VGND VPWR 0.142805f
C22 VPB VGND 0.013973f
C23 C1 VPWR 0.03984f
C24 A3 A1 0.00592f
C25 A1 VPWR 0.06706f
C26 VPB C1 0.124517f
C27 VPB A1 0.080317f
C28 VGND VNB 1.02863f
C29 X VNB 0.052121f
C30 VPWR VNB 0.821352f
C31 A1 VNB 0.210822f
C32 A2 VNB 0.320472f
C33 A3 VNB 0.209545f
C34 C1 VNB 0.299689f
C35 B1 VNB 0.330266f
C36 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o311a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311a_2 VNB VPB VPWR VGND X A1 A2 A3 B1 C1
X0 VPWR.t0 A1.t0 a_444_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=1.555 as=0.2184 ps=1.51 w=1.12 l=0.15
X1 a_135_74.t0 C1.t0 a_32_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0999 pd=1.01 as=0.2701 ps=2.21 w=0.74 l=0.15
X2 a_219_74.t2 A2.t0 VGND.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2487 ps=1.49 w=0.74 l=0.15
X3 VGND.t2 a_32_74.t4 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2775 pd=2.23 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_219_74.t3 B1.t0 a_135_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0999 ps=1.01 w=0.74 l=0.15
X5 VGND.t0 A3.t0 a_219_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2487 pd=1.49 as=0.1443 ps=1.13 w=0.74 l=0.15
X6 VGND.t1 A1.t1 a_219_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.16465 pd=1.185 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t1 a_32_74.t5 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t0 a_32_74.t6 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2436 ps=1.555 w=1.12 l=0.15
X9 X.t2 a_32_74.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.16465 ps=1.185 w=0.74 l=0.15
X10 VPWR.t3 C1.t1 a_32_74.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.295 ps=2.59 w=1 l=0.15
X11 a_32_74.t3 B1.t1 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2127 pd=1.51 as=0.21 ps=1.42 w=1 l=0.15
X12 a_444_368.t1 A2.t1 a_360_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1512 ps=1.39 w=1.12 l=0.15
X13 a_360_368.t0 A3.t1 a_32_74.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.2127 ps=1.51 w=1.12 l=0.15
R0 A1.n0 A1.t0 250.909
R1 A1.n0 A1.t1 220.113
R2 A1 A1.n0 158.102
R3 a_444_368.t0 a_444_368.t1 68.5987
R4 VPWR.n12 VPWR.n1 319.615
R5 VPWR.n3 VPWR.t1 263.45
R6 VPWR.n5 VPWR.n4 222.361
R7 VPWR.n4 VPWR.t2 50.13
R8 VPWR.n1 VPWR.t3 49.2505
R9 VPWR.n6 VPWR.n2 36.1417
R10 VPWR.n10 VPWR.n2 36.1417
R11 VPWR.n11 VPWR.n10 36.1417
R12 VPWR.n1 VPWR.t4 33.4905
R13 VPWR.n4 VPWR.t0 26.3844
R14 VPWR.n13 VPWR.n12 11.845
R15 VPWR.n5 VPWR.n3 10.5879
R16 VPWR.n7 VPWR.n6 9.3005
R17 VPWR.n8 VPWR.n2 9.3005
R18 VPWR.n10 VPWR.n9 9.3005
R19 VPWR.n11 VPWR.n0 9.3005
R20 VPWR.n6 VPWR.n5 7.90638
R21 VPWR.n12 VPWR.n11 7.15344
R22 VPWR.n7 VPWR.n3 0.576242
R23 VPWR VPWR.n13 0.163644
R24 VPWR.n13 VPWR.n0 0.144205
R25 VPWR.n8 VPWR.n7 0.122949
R26 VPWR.n9 VPWR.n8 0.122949
R27 VPWR.n9 VPWR.n0 0.122949
R28 VPB VPB.t4 314.113
R29 VPB.t0 VPB.t3 298.791
R30 VPB.t4 VPB.t6 291.13
R31 VPB.t2 VPB.t0 275.807
R32 VPB.t6 VPB.t5 275.807
R33 VPB.t3 VPB.t1 229.839
R34 VPB.t5 VPB.t2 214.517
R35 C1.n0 C1.t1 244.53
R36 C1 C1.n0 206.988
R37 C1.n0 C1.t0 154.24
R38 a_32_74.n3 a_32_74.n2 348.894
R39 a_32_74.n1 a_32_74.t6 266.731
R40 a_32_74.n0 a_32_74.t5 261.62
R41 a_32_74.n5 a_32_74.n4 252.547
R42 a_32_74.n4 a_32_74.t0 231.577
R43 a_32_74.n0 a_32_74.t4 156.431
R44 a_32_74.n1 a_32_74.t7 154.24
R45 a_32_74.n3 a_32_74.t1 127.956
R46 a_32_74.n4 a_32_74.n3 59.4829
R47 a_32_74.n2 a_32_74.n0 54.7732
R48 a_32_74.n5 a_32_74.t3 47.2805
R49 a_32_74.t2 a_32_74.n5 26.8503
R50 a_32_74.n2 a_32_74.n1 5.84292
R51 a_135_74.t0 a_135_74.t1 43.7843
R52 VNB.t0 VNB.t2 1662.99
R53 VNB VNB.t5 1385.83
R54 VNB.t1 VNB.t3 1374.28
R55 VNB.t6 VNB.t0 1247.24
R56 VNB.t3 VNB.t4 993.177
R57 VNB.t2 VNB.t1 993.177
R58 VNB.t5 VNB.t6 970.08
R59 A2.n0 A2.t1 250.909
R60 A2.n0 A2.t0 220.113
R61 A2 A2.n0 154.522
R62 VGND.n3 VGND.t2 282.464
R63 VGND.n5 VGND.n4 208.079
R64 VGND.n1 VGND.n0 195
R65 VGND.n0 VGND.t4 46.2167
R66 VGND.n0 VGND.t0 46.2167
R67 VGND.n4 VGND.t3 38.1086
R68 VGND.n7 VGND.n6 36.1417
R69 VGND.n4 VGND.t1 34.0546
R70 VGND.n6 VGND.n5 14.3064
R71 VGND.n9 VGND.n1 13.4361
R72 VGND.n8 VGND.n7 9.3005
R73 VGND.n6 VGND.n2 9.3005
R74 VGND.n5 VGND.n3 7.0997
R75 VGND.n7 VGND.n1 5.78592
R76 VGND.n3 VGND.n2 0.580021
R77 VGND VGND.n9 0.404642
R78 VGND.n9 VGND.n8 0.149306
R79 VGND.n8 VGND.n2 0.122949
R80 a_219_74.n1 a_219_74.n0 440.363
R81 a_219_74.n1 a_219_74.t3 40.541
R82 a_219_74.n0 a_219_74.t1 22.7032
R83 a_219_74.n0 a_219_74.t2 22.7032
R84 a_219_74.t0 a_219_74.n1 22.7032
R85 X X.n0 246.19
R86 X X.n1 115.844
R87 X.n0 X.t1 26.3844
R88 X.n0 X.t0 26.3844
R89 X.n1 X.t3 22.7032
R90 X.n1 X.t2 22.7032
R91 B1.n0 B1.t1 231.629
R92 B1.n0 B1.t0 220.113
R93 B1 B1.n0 154.25
R94 A3.n0 A3.t1 250.909
R95 A3.n0 A3.t0 220.113
R96 A3 A3.n0 154.522
R97 a_360_368.t0 a_360_368.t1 47.4916
C0 VPWR VGND 0.072555f
C1 A3 VGND 0.011424f
C2 A1 VPWR 0.0407f
C3 A2 X 0.003953f
C4 VPB VGND 0.008987f
C5 B1 VPWR 0.015074f
C6 A1 VPB 0.035919f
C7 A3 B1 0.083755f
C8 VPB B1 0.038258f
C9 VPWR X 0.222653f
C10 A3 X 2.77e-20
C11 A2 VPWR 0.080736f
C12 VPB X 0.011311f
C13 C1 VPWR 0.012266f
C14 A3 A2 0.092078f
C15 A2 VPB 0.035365f
C16 VPB C1 0.049224f
C17 A3 VPWR 0.011294f
C18 VPB VPWR 0.134995f
C19 A3 VPB 0.035071f
C20 A1 VGND 0.01504f
C21 B1 VGND 0.010985f
C22 X VGND 0.128687f
C23 A1 X 0.007254f
C24 A2 VGND 0.012401f
C25 C1 VGND 0.008639f
C26 B1 X 8.13e-20
C27 A2 A1 0.098829f
C28 A2 B1 5.78e-19
C29 C1 B1 0.056523f
C30 VGND VNB 0.541911f
C31 X VNB 0.072834f
C32 VPWR VNB 0.471085f
C33 A1 VNB 0.105746f
C34 A2 VNB 0.105112f
C35 A3 VNB 0.107626f
C36 B1 VNB 0.102541f
C37 C1 VNB 0.177507f
C38 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o311a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311a_1 VNB VPB VPWR VGND C1 B1 A3 A2 A1 X
X0 a_31_387.t2 B1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X1 a_209_74.t1 A3.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2976 pd=1.57 as=0.1824 ps=1.21 w=0.64 l=0.15
X2 X.t1 a_31_387.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2519 ps=1.59 w=1.12 l=0.15
X3 a_536_387.t0 A2.t0 a_320_387.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.465 ps=1.93 w=1 l=0.15
X4 X.t0 a_31_387.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1277 ps=1.1 w=0.74 l=0.15
X5 VPWR.t3 A1.t0 a_536_387.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2519 pd=1.59 as=0.21 ps=1.42 w=1 l=0.15
X6 a_209_74.t2 B1.t1 a_131_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
X7 VGND.t3 A2.t1 a_209_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.21 as=0.1248 ps=1.03 w=0.64 l=0.15
X8 a_131_74.t1 C1.t0 a_31_387.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X9 VGND.t1 A1.t1 a_209_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1277 pd=1.1 as=0.2976 ps=1.57 w=0.64 l=0.15
X10 VPWR.t1 C1.t1 a_31_387.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.295 ps=2.59 w=1 l=0.15
X11 a_320_387.t1 A3.t1 a_31_387.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.465 pd=1.93 as=0.15 ps=1.3 w=1 l=0.15
R0 B1.n0 B1.t0 313.3
R1 B1.n0 B1.t1 168.701
R2 B1 B1.n0 155.332
R3 VPWR.n2 VPWR.n1 228.875
R4 VPWR.n2 VPWR.n0 228.714
R5 VPWR.n0 VPWR.t3 53.1905
R6 VPWR.n1 VPWR.t2 39.4005
R7 VPWR.n1 VPWR.t1 39.4005
R8 VPWR.n0 VPWR.t0 34.3618
R9 VPWR VPWR.n2 0.200869
R10 a_31_387.n2 a_31_387.n1 411.959
R11 a_31_387.t0 a_31_387.n3 260.865
R12 a_31_387.n1 a_31_387.t4 250.909
R13 a_31_387.n1 a_31_387.t5 220.113
R14 a_31_387.n3 a_31_387.t3 193.22
R15 a_31_387.n2 a_31_387.n0 189.034
R16 a_31_387.n3 a_31_387.n2 62.6126
R17 a_31_387.n0 a_31_387.t1 29.5505
R18 a_31_387.n0 a_31_387.t2 29.5505
R19 VPB.t3 VPB.t1 551.614
R20 VPB.t5 VPB.t0 316.668
R21 VPB.t1 VPB.t5 291.13
R22 VPB.t2 VPB.t4 280.914
R23 VPB VPB.t2 268.146
R24 VPB.t4 VPB.t3 229.839
R25 A3.n0 A3.t1 461.113
R26 A3.n0 A3.t0 156.139
R27 A3.n1 A3.n0 152
R28 A3.n1 A3 11.4429
R29 A3 A3.n1 2.90959
R30 VGND.n2 VGND.n0 303.736
R31 VGND.n2 VGND.n1 89.2272
R32 VGND.n0 VGND.t2 53.438
R33 VGND.n0 VGND.t3 53.438
R34 VGND.n1 VGND.t0 37.6611
R35 VGND VGND.n2 33.1958
R36 VGND.n1 VGND.t1 26.2505
R37 a_209_74.n1 a_209_74.n0 218.924
R38 a_209_74.t0 a_209_74.n1 85.6107
R39 a_209_74.n1 a_209_74.t1 65.8753
R40 a_209_74.n0 a_209_74.t3 39.3755
R41 a_209_74.n0 a_209_74.t2 33.7505
R42 VNB.t2 VNB.t1 2494.49
R43 VNB.t4 VNB.t2 1662.99
R44 VNB VNB.t5 1339.63
R45 VNB.t3 VNB.t4 1247.24
R46 VNB.t1 VNB.t0 1177.95
R47 VNB.t5 VNB.t3 900.788
R48 X.n0 X.t1 301.562
R49 X.t0 X.n0 279.738
R50 X.n1 X.t0 279.738
R51 X.n1 X 11.3978
R52 X.n0 X 4.38406
R53 X X.n1 1.57858
R54 A2.n0 A2.t0 544.357
R55 A2.n0 A2.t1 320.7
R56 A2 A2.n0 3.47479
R57 a_320_387.t0 a_320_387.t1 183.21
R58 a_536_387.t0 a_536_387.t1 82.7405
R59 A1.n0 A1.t0 318.656
R60 A1.n0 A1.t1 162.274
R61 A1 A1.n0 159.177
R62 a_131_74.t0 a_131_74.t1 45.0005
R63 C1.n0 C1.t1 303.661
R64 C1.n0 C1.t0 159.06
R65 C1 C1.n0 156.462
C0 X VGND 0.090721f
C1 VGND A2 0.05233f
C2 X A1 0.008869f
C3 A2 A1 0.035684f
C4 C1 VGND 0.01201f
C5 B1 X 4.54e-20
C6 B1 A2 0.065361f
C7 C1 B1 0.064398f
C8 VPWR VGND 0.069854f
C9 VPWR A1 0.011799f
C10 X A2 7.64e-20
C11 VGND A3 0.042399f
C12 A3 A1 0.020948f
C13 VPB VGND 0.008478f
C14 B1 VPWR 0.020198f
C15 VPB A1 0.039345f
C16 B1 A3 0.024604f
C17 VPB B1 0.036014f
C18 VPWR X 0.128322f
C19 X A3 1.82e-19
C20 VPWR A2 0.014548f
C21 A3 A2 0.261243f
C22 VPB X 0.015365f
C23 C1 VPWR 0.021048f
C24 VPB A2 0.050179f
C25 VPB C1 0.048652f
C26 VPWR A3 0.009948f
C27 VPB VPWR 0.119785f
C28 VPB A3 0.07681f
C29 VGND A1 0.053744f
C30 B1 VGND 0.014905f
C31 VGND VNB 0.538077f
C32 X VNB 0.115052f
C33 VPWR VNB 0.427323f
C34 A1 VNB 0.132855f
C35 A2 VNB 0.151801f
C36 A3 VNB 0.153561f
C37 B1 VNB 0.114962f
C38 C1 VNB 0.186117f
C39 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o221ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221ai_4 VNB VPB VPWR VGND B1 A2 C1 B2 Y A1
X0 VPWR.t4 A1.t0 a_1288_368# VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t12 C1.t0 a_27_84.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 Y.t8 C1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 VPWR.t8 B1.t0 a_508_368.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_1288_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_27_84.t2 B1.t1 a_483_74.t13 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_508_368.t5 B1.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7 Y.t4 A2.t0 a_1288_368# VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_1288_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_508_368.t0 B2.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X10 Y.t3 A2.t1 a_1288_368# VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1988 ps=1.475 w=1.12 l=0.15
X11 a_27_84.t9 B1.t3 a_483_74.t12 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 VGND.t7 A1.t1 a_483_74.t9 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 a_483_74.t4 B2.t1 a_27_84.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_483_74.t8 A1.t2 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1073 ps=1.03 w=0.74 l=0.15
X15 a_1288_368# A1.t3 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.475 as=0.224 ps=1.52 w=1.12 l=0.15
X16 a_27_84.t3 C1.t2 Y.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 Y.t1 B2.t2 a_508_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_483_74.t11 B1.t4 a_27_84.t10 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 VPWR.t5 C1.t3 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.182 ps=1.445 w=1.12 l=0.15
X20 a_508_368.t2 B2.t3 Y.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_27_84.t6 C1.t4 Y.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 Y.t13 B2.t4 a_508_368.t7 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_483_74.t10 B1.t5 a_27_84.t11 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_483_74.t3 A2.t2 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X25 a_508_368.t4 B1.t6 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X26 Y.t6 C1.t5 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.182 pd=1.445 as=0.2156 ps=1.505 w=1.12 l=0.15
X27 Y.t9 C1.t6 a_27_84.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VGND.t2 A2.t3 a_483_74.t2 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 VPWR.t7 C1.t7 Y.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2156 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X30 VPWR.t2 A1.t4 a_1288_368# VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X31 a_483_74.t5 B2.t5 a_27_84.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 VGND.t1 A2.t4 a_483_74.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 a_483_74.t7 A1.t5 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X34 a_27_84.t7 B2.t6 a_483_74.t14 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X35 VPWR.t10 B1.t7 a_508_368.t3 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.196 ps=1.47 w=1.12 l=0.15
X36 a_1288_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X37 a_27_84.t8 B2.t7 a_483_74.t15 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X38 a_483_74.t0 A2.t5 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X39 VGND.t4 A1.t6 a_483_74.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
R0 A1.n12 A1.n0 299.339
R1 A1.n0 A1.t3 275.009
R2 A1.n3 A1.t4 250.909
R3 A1.n2 A1.n1 250.909
R4 A1.n9 A1.t0 250.909
R5 A1.n0 A1.t1 191.194
R6 A1.n9 A1.t2 169.285
R7 A1.n3 A1.t5 169.285
R8 A1.n4 A1.t6 167.094
R9 A1.n11 A1.n10 152
R10 A1.n8 A1.n7 152
R11 A1.n6 A1.n5 152
R12 A1.n10 A1.n8 49.6611
R13 A1.n5 A1.n4 39.4369
R14 A1.n5 A1.n3 21.1793
R15 A1.n10 A1.n9 10.955
R16 A1.n12 A1.n11 9.23127
R17 A1.n6 A1 8.12358
R18 A1.n7 A1 7.13896
R19 A1.n4 A1.n2 5.11262
R20 A1.n8 A1.n2 5.11262
R21 A1.n7 A1 4.67742
R22 A1 A1.n6 3.69281
R23 A1 A1.n12 1.35435
R24 A1.n11 A1 1.23127
R25 VPWR.n32 VPWR.n6 604.976
R26 VPWR.n14 VPWR.t4 349.789
R27 VPWR.n38 VPWR.n2 315.928
R28 VPWR.n4 VPWR.n3 315.738
R29 VPWR.n10 VPWR.n9 315.738
R30 VPWR.n13 VPWR.t2 264.493
R31 VPWR.n40 VPWR.t1 257.433
R32 VPWR.n26 VPWR.n25 36.1417
R33 VPWR.n27 VPWR.n26 36.1417
R34 VPWR.n27 VPWR.n7 36.1417
R35 VPWR.n31 VPWR.n7 36.1417
R36 VPWR.n15 VPWR.n12 36.1417
R37 VPWR.n19 VPWR.n12 36.1417
R38 VPWR.n20 VPWR.n19 36.1417
R39 VPWR.n21 VPWR.n20 36.1417
R40 VPWR.n2 VPWR.t7 35.1791
R41 VPWR.n3 VPWR.t0 35.1791
R42 VPWR.n6 VPWR.t9 35.1791
R43 VPWR.n6 VPWR.t8 35.1791
R44 VPWR.n9 VPWR.t3 35.1791
R45 VPWR.n9 VPWR.t10 35.1791
R46 VPWR.n2 VPWR.t6 32.5407
R47 VPWR.n25 VPWR.n10 30.4946
R48 VPWR.n33 VPWR.n32 28.9887
R49 VPWR.n40 VPWR.n39 26.7299
R50 VPWR.n3 VPWR.t5 26.3844
R51 VPWR.n39 VPWR.n38 25.977
R52 VPWR.n37 VPWR.n4 25.977
R53 VPWR.n15 VPWR.n14 24.8476
R54 VPWR.n38 VPWR.n37 21.4593
R55 VPWR.n33 VPWR.n4 21.4593
R56 VPWR.n32 VPWR.n31 18.4476
R57 VPWR.n21 VPWR.n10 16.9417
R58 VPWR.n16 VPWR.n15 9.3005
R59 VPWR.n17 VPWR.n12 9.3005
R60 VPWR.n19 VPWR.n18 9.3005
R61 VPWR.n20 VPWR.n11 9.3005
R62 VPWR.n22 VPWR.n21 9.3005
R63 VPWR.n23 VPWR.n10 9.3005
R64 VPWR.n25 VPWR.n24 9.3005
R65 VPWR.n26 VPWR.n8 9.3005
R66 VPWR.n28 VPWR.n27 9.3005
R67 VPWR.n29 VPWR.n7 9.3005
R68 VPWR.n31 VPWR.n30 9.3005
R69 VPWR.n32 VPWR.n5 9.3005
R70 VPWR.n34 VPWR.n33 9.3005
R71 VPWR.n35 VPWR.n4 9.3005
R72 VPWR.n37 VPWR.n36 9.3005
R73 VPWR.n38 VPWR.n1 9.3005
R74 VPWR.n39 VPWR.n0 9.3005
R75 VPWR.n41 VPWR.n40 9.3005
R76 VPWR.n14 VPWR.n13 6.97336
R77 VPWR.n16 VPWR.n13 0.546712
R78 VPWR.n17 VPWR.n16 0.122949
R79 VPWR.n18 VPWR.n17 0.122949
R80 VPWR.n18 VPWR.n11 0.122949
R81 VPWR.n22 VPWR.n11 0.122949
R82 VPWR.n23 VPWR.n22 0.122949
R83 VPWR.n24 VPWR.n23 0.122949
R84 VPWR.n24 VPWR.n8 0.122949
R85 VPWR.n28 VPWR.n8 0.122949
R86 VPWR.n29 VPWR.n28 0.122949
R87 VPWR.n30 VPWR.n29 0.122949
R88 VPWR.n30 VPWR.n5 0.122949
R89 VPWR.n34 VPWR.n5 0.122949
R90 VPWR.n35 VPWR.n34 0.122949
R91 VPWR.n36 VPWR.n35 0.122949
R92 VPWR.n36 VPWR.n1 0.122949
R93 VPWR.n1 VPWR.n0 0.122949
R94 VPWR.n41 VPWR.n0 0.122949
R95 VPWR VPWR.n41 0.0617245
R96 VPB.t6 VPB.t4 459.678
R97 VPB.t12 VPB.t6 459.678
R98 VPB.t11 VPB.t12 459.678
R99 VPB.t15 VPB.t5 280.914
R100 VPB.t13 VPB.t14 280.914
R101 VPB.t9 VPB.t8 273.253
R102 VPB.t5 VPB.t11 257.93
R103 VPB VPB.t2 257.93
R104 VPB.t0 VPB.t15 255.376
R105 VPB.t3 VPB.t0 255.376
R106 VPB.t7 VPB.t1 255.376
R107 VPB.t8 VPB.t7 242.608
R108 VPB.t10 VPB.t3 229.839
R109 VPB.t16 VPB.t10 229.839
R110 VPB.t14 VPB.t16 229.839
R111 VPB.t1 VPB.t13 229.839
R112 VPB.t2 VPB.t9 229.839
R113 C1.n0 C1.t3 262.666
R114 C1.n1 C1.t5 226.809
R115 C1.n4 C1.t7 226.809
R116 C1.n6 C1.t1 226.809
R117 C1.n6 C1.t0 181.407
R118 C1.n5 C1.t4 179.947
R119 C1.n2 C1.t6 179.947
R120 C1.n0 C1.t2 179.947
R121 C1 C1.n3 155.721
R122 C1.n10 C1.n9 152
R123 C1.n8 C1.n7 152
R124 C1.n9 C1.n8 49.6611
R125 C1.n1 C1.n0 43.0884
R126 C1.n4 C1.n3 41.6278
R127 C1.n2 C1.n1 19.7187
R128 C1.n3 C1.n2 16.7975
R129 C1.n7 C1 12.0563
R130 C1.n8 C1.n6 8.03383
R131 C1.n10 C1 7.88887
R132 C1 C1.n10 6.4005
R133 C1.n5 C1.n4 4.38232
R134 C1.n9 C1.n5 3.65202
R135 C1.n7 C1 2.23306
R136 a_27_84.n2 a_27_84.n0 229.611
R137 a_27_84.n4 a_27_84.t4 206.721
R138 a_27_84.n4 a_27_84.n3 206.559
R139 a_27_84.n7 a_27_84.n6 185
R140 a_27_84.n2 a_27_84.n1 185
R141 a_27_84.n9 a_27_84.n8 185
R142 a_27_84.n5 a_27_84.t3 137.606
R143 a_27_84.n5 a_27_84.n4 67.8611
R144 a_27_84.n8 a_27_84.n7 50.2088
R145 a_27_84.n8 a_27_84.n2 42.2184
R146 a_27_84.n7 a_27_84.n5 34.8226
R147 a_27_84.n6 a_27_84.t10 22.7032
R148 a_27_84.n6 a_27_84.t9 22.7032
R149 a_27_84.n3 a_27_84.t5 22.7032
R150 a_27_84.n3 a_27_84.t6 22.7032
R151 a_27_84.n1 a_27_84.t1 22.7032
R152 a_27_84.n1 a_27_84.t8 22.7032
R153 a_27_84.n0 a_27_84.t11 22.7032
R154 a_27_84.n0 a_27_84.t7 22.7032
R155 a_27_84.t0 a_27_84.n9 22.7032
R156 a_27_84.n9 a_27_84.t2 22.7032
R157 Y.n12 Y.t3 772.15
R158 Y Y.t3 704.741
R159 Y.n6 Y.n1 585
R160 Y.n12 Y.t4 419.534
R161 Y.n8 Y.n1 311.286
R162 Y.n9 Y.n0 298.943
R163 Y.n11 Y.n10 296.659
R164 Y.n7 Y.n2 256.688
R165 Y.n9 Y.n8 174.306
R166 Y.n5 Y.n3 138.5
R167 Y.n13 Y.n11 119.719
R168 Y.n5 Y.n4 98.418
R169 Y.n6 Y.n5 59.8367
R170 Y.n11 Y.n9 59.1064
R171 Y.n10 Y.t1 35.1791
R172 Y.n1 Y.t6 30.7817
R173 Y.n0 Y.t2 26.3844
R174 Y.n0 Y.t13 26.3844
R175 Y.n1 Y.t7 26.3844
R176 Y.n2 Y.t5 26.3844
R177 Y.n2 Y.t8 26.3844
R178 Y.n10 Y.t0 26.3844
R179 Y.n4 Y.t11 22.7032
R180 Y.n4 Y.t9 22.7032
R181 Y.n3 Y.t10 22.7032
R182 Y.n3 Y.t12 22.7032
R183 Y Y.n13 5.70652
R184 Y.n8 Y.n7 5.1205
R185 Y.n7 Y.n6 2.5605
R186 Y.n13 Y.n12 0.617367
R187 VNB.t11 VNB.t17 2286.61
R188 VNB.t7 VNB.t3 1316.54
R189 VNB.t6 VNB.t4 1154.86
R190 VNB.t16 VNB.t1 1154.86
R191 VNB.t19 VNB.t7 1154.86
R192 VNB VNB.t12 1143.31
R193 VNB.t15 VNB.t6 1016.27
R194 VNB.t4 VNB.t5 993.177
R195 VNB.t1 VNB.t15 993.177
R196 VNB.t3 VNB.t16 993.177
R197 VNB.t13 VNB.t19 993.177
R198 VNB.t2 VNB.t13 993.177
R199 VNB.t14 VNB.t2 993.177
R200 VNB.t0 VNB.t14 993.177
R201 VNB.t8 VNB.t0 993.177
R202 VNB.t18 VNB.t8 993.177
R203 VNB.t17 VNB.t18 993.177
R204 VNB.t9 VNB.t11 993.177
R205 VNB.t10 VNB.t9 993.177
R206 VNB.t12 VNB.t10 993.177
R207 B1.n2 B1.t2 262.594
R208 B1.n0 B1.t7 250.909
R209 B1.n7 B1.t6 245.522
R210 B1.n4 B1.t0 226.809
R211 B1.n0 B1.t5 220.113
R212 B1.n3 B1.t3 196.013
R213 B1.n6 B1.t1 168.701
R214 B1 B1.n0 161.661
R215 B1.n2 B1.n1 160.212
R216 B1.n8 B1.n7 152
R217 B1.n5 B1.n1 152
R218 B1.n6 B1.t4 151.5
R219 B1 B1.n8 144.005
R220 B1.n7 B1.n6 28.9205
R221 B1.n4 B1.n3 20.449
R222 B1.n5 B1.n4 19.7187
R223 B1.n7 B1.n5 11.6853
R224 B1.n3 B1.n2 9.49444
R225 B1.n8 B1.n1 8.21182
R226 a_508_368.n2 a_508_368.n0 352.997
R227 a_508_368.n5 a_508_368.n4 352.729
R228 a_508_368.n2 a_508_368.n1 302.55
R229 a_508_368.n4 a_508_368.n3 289.24
R230 a_508_368.n4 a_508_368.n2 56.227
R231 a_508_368.n0 a_508_368.t0 35.1791
R232 a_508_368.n3 a_508_368.t7 26.3844
R233 a_508_368.n3 a_508_368.t4 26.3844
R234 a_508_368.n0 a_508_368.t3 26.3844
R235 a_508_368.n1 a_508_368.t1 26.3844
R236 a_508_368.n1 a_508_368.t2 26.3844
R237 a_508_368.t6 a_508_368.n5 26.3844
R238 a_508_368.n5 a_508_368.t5 26.3844
R239 A2.n3 A2.t0 226.809
R240 A2.n5 A2.n4 226.809
R241 A2.n7 A2.t1 226.809
R242 A2.n1 A2.n0 204.678
R243 A2.n7 A2.t5 198.204
R244 A2.n1 A2.t3 196.714
R245 A2.n6 A2.t4 196.013
R246 A2.n2 A2.t2 196.013
R247 A2.n13 A2.n12 152
R248 A2.n11 A2.n10 152
R249 A2.n9 A2.n8 152
R250 A2.n2 A2.n1 62.106
R251 A2.n12 A2.n11 49.6611
R252 A2.n8 A2.n6 40.1672
R253 A2.n8 A2.n7 20.449
R254 A2.n10 A2.n9 12.4348
R255 A2.n13 A2 12.2519
R256 A2.n12 A2.n3 11.6853
R257 A2 A2.n13 5.30336
R258 A2.n6 A2.n5 5.11262
R259 A2.n9 A2 4.93764
R260 A2.n11 A2.n5 4.38232
R261 A2.n3 A2.n2 2.19141
R262 A2.n10 A2 0.183357
R263 a_483_74.n12 a_483_74.t12 323.769
R264 a_483_74.n1 a_483_74.t7 202.599
R265 a_483_74.n3 a_483_74.n2 185
R266 a_483_74.n5 a_483_74.n4 185
R267 a_483_74.n9 a_483_74.n8 185
R268 a_483_74.n11 a_483_74.n10 185
R269 a_483_74.n13 a_483_74.n12 185
R270 a_483_74.n1 a_483_74.n0 95.2869
R271 a_483_74.n7 a_483_74.n6 90.3626
R272 a_483_74.n7 a_483_74.n5 60.2159
R273 a_483_74.n5 a_483_74.n3 56.8145
R274 a_483_74.n3 a_483_74.n1 56.2361
R275 a_483_74.n9 a_483_74.n7 46.6708
R276 a_483_74.n11 a_483_74.n9 44.0325
R277 a_483_74.n12 a_483_74.n11 44.0325
R278 a_483_74.n6 a_483_74.t10 34.0546
R279 a_483_74.n0 a_483_74.t8 34.0546
R280 a_483_74.n10 a_483_74.t15 22.7032
R281 a_483_74.n10 a_483_74.t4 22.7032
R282 a_483_74.n8 a_483_74.t14 22.7032
R283 a_483_74.n8 a_483_74.t5 22.7032
R284 a_483_74.n6 a_483_74.t9 22.7032
R285 a_483_74.n4 a_483_74.t1 22.7032
R286 a_483_74.n4 a_483_74.t0 22.7032
R287 a_483_74.n2 a_483_74.t2 22.7032
R288 a_483_74.n2 a_483_74.t3 22.7032
R289 a_483_74.n0 a_483_74.t6 22.7032
R290 a_483_74.t13 a_483_74.n13 22.7032
R291 a_483_74.n13 a_483_74.t11 22.7032
R292 B2.n2 B2.t0 261.62
R293 B2.n5 B2.t2 261.62
R294 B2.n1 B2.t4 227.762
R295 B2.n1 B2.t3 219.766
R296 B2.n2 B2.t6 160.083
R297 B2 B2.n10 156.445
R298 B2.n3 B2 154.667
R299 B2.n9 B2.t1 154.24
R300 B2.n4 B2.t5 154.24
R301 B2.n6 B2.n0 152
R302 B2.n8 B2.t7 136.567
R303 B2.n9 B2.n8 75.7434
R304 B2.n3 B2.n2 41.6278
R305 B2.n10 B2.n1 29.6318
R306 B2.n7 B2.n6 26.2914
R307 B2.n8 B2.n7 23.0527
R308 B2.n6 B2.n5 18.2581
R309 B2.n10 B2.n9 17.1037
R310 B2.n5 B2.n4 16.0672
R311 B2.n4 B2.n3 15.3369
R312 B2 B2.n0 9.42272
R313 B2.n10 B2.n7 8.03383
R314 B2 B2.n0 7.64494
R315 VGND.n6 VGND.n5 211.964
R316 VGND.n9 VGND.n2 204.201
R317 VGND.n12 VGND.n11 204.201
R318 VGND.n4 VGND.n3 203.636
R319 VGND.n2 VGND.t3 34.0546
R320 VGND.n11 VGND.t0 34.0546
R321 VGND.n11 VGND.t7 34.0546
R322 VGND.n10 VGND.n9 28.2358
R323 VGND.n4 VGND.n1 25.977
R324 VGND.n3 VGND.t6 23.514
R325 VGND.n3 VGND.t2 23.514
R326 VGND.n5 VGND.t5 22.7032
R327 VGND.n5 VGND.t4 22.7032
R328 VGND.n2 VGND.t1 22.7032
R329 VGND.n9 VGND.n1 19.2005
R330 VGND.n12 VGND.n10 16.9417
R331 VGND.n10 VGND.n0 9.3005
R332 VGND.n9 VGND.n8 9.3005
R333 VGND.n7 VGND.n1 9.3005
R334 VGND.n13 VGND.n12 7.45461
R335 VGND.n6 VGND.n4 6.5391
R336 VGND VGND.n13 1.63166
R337 VGND.n7 VGND.n6 0.568197
R338 VGND.n13 VGND.n0 0.152559
R339 VGND.n8 VGND.n7 0.122949
R340 VGND.n8 VGND.n0 0.122949
C0 VGND B1 0.030661f
C1 VPWR B2 0.022419f
C2 VGND A2 0.054118f
C3 A1 a_1288_368# 0.155274f
C4 Y a_1288_368# 0.268486f
C5 C1 B1 0.034405f
C6 A1 B1 0.073479f
C7 Y B1 0.344704f
C8 A1 A2 0.303498f
C9 VGND C1 0.025386f
C10 VGND A1 0.077465f
C11 Y A2 0.162529f
C12 VPB a_1288_368# 0.017029f
C13 Y VGND 0.029627f
C14 VPWR a_1288_368# 0.54686f
C15 VPB B1 0.155511f
C16 A2 VPB 0.133355f
C17 B2 B1 0.274685f
C18 VGND VPB 0.008462f
C19 VPWR B1 0.070449f
C20 Y C1 0.327999f
C21 VGND B2 0.025324f
C22 Y A1 0.041468f
C23 VPWR A2 0.024399f
C24 VPWR VGND 0.160517f
C25 VPB C1 0.14764f
C26 B2 C1 5.75e-20
C27 A1 VPB 0.134643f
C28 VPWR C1 0.103457f
C29 Y VPB 0.015121f
C30 B2 A1 0.004536f
C31 Y B2 0.056173f
C32 VPWR A1 0.099723f
C33 VPWR Y 0.509156f
C34 B1 a_1288_368# 4.69e-19
C35 A2 a_1288_368# 0.049173f
C36 VGND a_1288_368# 0.007365f
C37 B2 VPB 0.129106f
C38 A2 B1 0.005656f
C39 VPWR VPB 0.253535f
C40 VGND VNB 1.11939f
C41 Y VNB 0.037629f
C42 VPWR VNB 0.971153f
C43 A2 VNB 0.392043f
C44 A1 VNB 0.483219f
C45 B2 VNB 0.400762f
C46 B1 VNB 0.437774f
C47 C1 VNB 0.444284f
C48 VPB VNB 2.33467f
C49 a_1288_368# VNB 0.011145f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o221ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221ai_2 VNB VPB VPWR VGND Y B1 A1 C1 B2 A2
X0 VPWR.t2 C1.t0 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3696 pd=1.78 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_311_85.t7 B1.t0 a_27_74.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.14985 ps=1.145 w=0.74 l=0.15
X2 VPWR.t3 B1.t1 a_376_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.196 ps=1.47 w=1.12 l=0.15
X3 a_27_74.t3 B2.t0 a_311_85.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.14985 pd=1.145 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_776_368.t2 A2.t0 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VGND.t1 A1.t0 a_311_85.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1406 pd=1.12 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 Y.t1 C1.t1 a_27_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 Y.t5 A2.t1 a_776_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8 VPWR.t4 A1.t1 a_776_368.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_311_85.t1 A2.t2 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1406 ps=1.12 w=0.74 l=0.15
X10 a_311_85.t4 A1.t2 VGND.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1258 ps=1.08 w=0.74 l=0.15
X11 Y.t2 C1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X12 a_376_368.t1 B2.t1 Y.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1764 ps=1.435 w=1.12 l=0.15
X13 a_311_85.t0 B2.t2 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_776_368.t0 A1.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.224 ps=1.52 w=1.12 l=0.15
X15 VGND.t2 A2.t3 a_311_85.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1221 ps=1.07 w=0.74 l=0.15
X16 a_27_74.t1 C1.t3 Y.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_376_368.t2 B1.t2 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.3696 ps=1.78 w=1.12 l=0.15
X18 a_27_74.t4 B1.t3 a_311_85.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X19 Y.t6 B2.t3 a_376_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
R0 C1.n0 C1.t0 262.543
R1 C1.n1 C1.t2 240.197
R2 C1 C1.n2 187.93
R3 C1.n0 C1.t3 179.947
R4 C1.n2 C1.t1 179.947
R5 C1.n1 C1.n0 61.346
R6 C1.n2 C1.n1 7.30353
R7 Y.n2 Y.n0 720.234
R8 Y.n8 Y 591.4
R9 Y.n2 Y.n1 585
R10 Y.n8 Y.n6 585
R11 Y.n9 Y.n8 585
R12 Y.n5 Y.n4 185
R13 Y.n3 Y.n2 116.934
R14 Y.n1 Y.t6 29.0228
R15 Y.n1 Y.t7 26.3844
R16 Y.n0 Y.t4 26.3844
R17 Y.n0 Y.t5 26.3844
R18 Y.n8 Y.t3 26.3844
R19 Y.n8 Y.t2 26.3844
R20 Y.n4 Y.t0 22.7032
R21 Y.n4 Y.t1 22.7032
R22 Y Y.n5 16.5931
R23 Y Y.n9 15.882
R24 Y Y.n7 11.7765
R25 Y.n7 Y 7.1685
R26 Y.n7 Y.n6 2.84494
R27 Y Y.n3 2.60791
R28 Y.n9 Y 1.65976
R29 Y.n6 Y.n3 1.18569
R30 Y.n5 Y 0.948648
R31 VPWR.n5 VPWR.n4 605.365
R32 VPWR.n11 VPWR.n1 585
R33 VPWR.n13 VPWR.n12 585
R34 VPWR.n6 VPWR.t4 358.493
R35 VPWR.n19 VPWR.t1 257.433
R36 VPWR.n12 VPWR.n11 63.3219
R37 VPWR.n9 VPWR.n3 36.1417
R38 VPWR.n10 VPWR.n9 36.1417
R39 VPWR.n14 VPWR.n10 35.2569
R40 VPWR.n4 VPWR.t0 35.1791
R41 VPWR.n4 VPWR.t3 35.1791
R42 VPWR.n18 VPWR.n17 27.5884
R43 VPWR.n12 VPWR.t5 26.3844
R44 VPWR.n11 VPWR.t2 26.3844
R45 VPWR.n19 VPWR.n18 23.7181
R46 VPWR.n5 VPWR.n3 18.4476
R47 VPWR.n7 VPWR.n3 9.3005
R48 VPWR.n9 VPWR.n8 9.3005
R49 VPWR.n10 VPWR.n2 9.3005
R50 VPWR.n15 VPWR.n14 9.3005
R51 VPWR.n17 VPWR.n16 9.3005
R52 VPWR.n18 VPWR.n0 9.3005
R53 VPWR.n20 VPWR.n19 9.3005
R54 VPWR.n6 VPWR.n5 7.38057
R55 VPWR.n13 VPWR.n1 5.87056
R56 VPWR.n14 VPWR.n13 1.63107
R57 VPWR.n17 VPWR.n1 0.326615
R58 VPWR.n7 VPWR.n6 0.167197
R59 VPWR.n8 VPWR.n7 0.122949
R60 VPWR.n8 VPWR.n2 0.122949
R61 VPWR.n15 VPWR.n2 0.122949
R62 VPWR.n16 VPWR.n15 0.122949
R63 VPWR.n16 VPWR.n0 0.122949
R64 VPWR.n20 VPWR.n0 0.122949
R65 VPWR VPWR.n20 0.0617245
R66 VPB.t2 VPB.t9 413.711
R67 VPB.t5 VPB.t0 280.914
R68 VPB VPB.t1 278.361
R69 VPB.t0 VPB.t4 255.376
R70 VPB.t8 VPB.t5 255.376
R71 VPB.t9 VPB.t6 247.715
R72 VPB.t6 VPB.t8 237.5
R73 VPB.t3 VPB.t7 229.839
R74 VPB.t4 VPB.t3 229.839
R75 VPB.t1 VPB.t2 229.839
R76 B1.n1 B1.t2 250.909
R77 B1.n0 B1.t1 250.909
R78 B1 B1.n0 235.731
R79 B1.n0 B1.t0 202.44
R80 B1.n1 B1.t3 191.903
R81 B1.n2 B1.n1 152
R82 B1 B1.n2 4.65505
R83 B1.n2 B1 3.32518
R84 a_27_74.t2 a_27_74.n3 226.339
R85 a_27_74.n2 a_27_74.n0 194.412
R86 a_27_74.n2 a_27_74.n1 155.135
R87 a_27_74.n3 a_27_74.t1 134.338
R88 a_27_74.n3 a_27_74.n2 79.839
R89 a_27_74.n1 a_27_74.t3 38.5257
R90 a_27_74.n1 a_27_74.t5 27.1503
R91 a_27_74.n0 a_27_74.t0 22.7032
R92 a_27_74.n0 a_27_74.t4 22.7032
R93 a_311_85.t6 a_311_85.n5 263.565
R94 a_311_85.n1 a_311_85.t4 199.077
R95 a_311_85.n5 a_311_85.n4 185
R96 a_311_85.n1 a_311_85.n0 99.7274
R97 a_311_85.n3 a_311_85.n2 87.1354
R98 a_311_85.n5 a_311_85.n3 81.5874
R99 a_311_85.n3 a_311_85.n1 65.2752
R100 a_311_85.n0 a_311_85.t1 29.1897
R101 a_311_85.n0 a_311_85.t5 24.3248
R102 a_311_85.n4 a_311_85.t2 22.7032
R103 a_311_85.n4 a_311_85.t0 22.7032
R104 a_311_85.n2 a_311_85.t3 22.7032
R105 a_311_85.n2 a_311_85.t7 22.7032
R106 VNB.t2 VNB.t8 2286.61
R107 VNB.t4 VNB.t9 1281.89
R108 VNB.t5 VNB.t1 1224.15
R109 VNB VNB.t3 1143.31
R110 VNB.t7 VNB.t6 1131.76
R111 VNB.t1 VNB.t7 1108.66
R112 VNB.t9 VNB.t5 993.177
R113 VNB.t0 VNB.t4 993.177
R114 VNB.t8 VNB.t0 993.177
R115 VNB.t3 VNB.t2 993.177
R116 a_376_368.n1 a_376_368.n0 1234.8
R117 a_376_368.n0 a_376_368.t1 35.1791
R118 a_376_368.n1 a_376_368.t0 32.5407
R119 a_376_368.n0 a_376_368.t3 26.3844
R120 a_376_368.t2 a_376_368.n1 26.3844
R121 B2.n1 B2.t3 235.637
R122 B2.n0 B2.t1 226.809
R123 B2.n0 B2.t0 181.262
R124 B2.n1 B2.t2 178.34
R125 B2 B2.n2 155.87
R126 B2.n2 B2.n1 49.6611
R127 B2.n2 B2.n0 10.2247
R128 A2.n0 A2.t0 226.809
R129 A2.n1 A2.t1 226.809
R130 A2.n1 A2.t2 180.531
R131 A2.n0 A2.t3 180.531
R132 A2 A2.n2 154.522
R133 A2.n2 A2.n0 35.7853
R134 A2.n2 A2.n1 29.9429
R135 a_776_368.n1 a_776_368.n0 941.597
R136 a_776_368.n0 a_776_368.t1 35.1791
R137 a_776_368.n0 a_776_368.t0 26.3844
R138 a_776_368.n1 a_776_368.t3 26.3844
R139 a_776_368.t2 a_776_368.n1 26.3844
R140 A1 A1.n0 251.903
R141 A1.n1 A1.t1 250.909
R142 A1.n0 A1.t3 250.909
R143 A1.n1 A1.t2 202.44
R144 A1.n0 A1.t0 202.44
R145 A1 A1.n1 153.173
R146 VGND.n2 VGND.n0 216.202
R147 VGND.n2 VGND.n1 215.886
R148 VGND.n1 VGND.t1 34.0546
R149 VGND.n0 VGND.t2 32.4329
R150 VGND.n1 VGND.t3 27.5681
R151 VGND.n0 VGND.t0 22.7032
R152 VGND VGND.n2 1.32628
C0 VPWR VPB 0.154731f
C1 VGND B1 0.01783f
C2 A1 VPWR 0.080188f
C3 B2 Y 0.02251f
C4 VPWR Y 0.297989f
C5 VPB B1 0.079191f
C6 A1 B1 0.104032f
C7 Y B1 0.274669f
C8 VGND C1 0.014675f
C9 B2 VPWR 0.010491f
C10 A2 VGND 0.030957f
C11 VPB C1 0.084205f
C12 A2 VPB 0.060328f
C13 B2 B1 0.21727f
C14 Y C1 0.118244f
C15 VPWR B1 0.054048f
C16 VGND VPB 0.006339f
C17 A1 A2 0.21082f
C18 A1 VGND 0.033712f
C19 A2 Y 0.01426f
C20 Y VGND 0.013567f
C21 A1 VPB 0.078175f
C22 VPWR C1 0.06142f
C23 Y VPB 0.007522f
C24 A1 Y 0.0973f
C25 B2 VGND 0.010429f
C26 A2 VPWR 0.011521f
C27 VPWR VGND 0.09251f
C28 C1 B1 0.036857f
C29 B2 VPB 0.060963f
C30 VGND VNB 0.674517f
C31 Y VNB 0.02347f
C32 VPWR VNB 0.599622f
C33 A2 VNB 0.185264f
C34 A1 VNB 0.265481f
C35 B2 VNB 0.181196f
C36 B1 VNB 0.225894f
C37 C1 VNB 0.285994f
C38 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o221ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221ai_1 VNB VPB VPWR VGND Y B1 A1 C1 B2 A2
X0 VGND.t1 A2.t0 a_239_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2368 pd=1.38 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 a_114_74.t2 C1.t0 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 a_239_74.t0 B2.t0 a_114_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 Y.t0 B2.t1 a_324_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X4 VPWR.t2 C1.t1 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.4256 pd=1.88 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 a_324_368.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.4256 ps=1.88 w=1.12 l=0.15
X6 a_522_368.t1 A2.t1 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X7 a_114_74.t1 B1.t1 a_239_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VPWR.t1 A1.t0 a_522_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X9 a_239_74.t2 A1.t1 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2368 ps=1.38 w=0.74 l=0.15
R0 A2.n0 A2.t1 250.909
R1 A2.n0 A2.t0 220.113
R2 A2 A2.n0 154.522
R3 A2.n1 A2 13.8245
R4 A2 A2.n1 5.1205
R5 A2.n1 A2 3.87929
R6 a_239_74.n0 a_239_74.t1 337.682
R7 a_239_74.n0 a_239_74.t2 214.216
R8 a_239_74.n1 a_239_74.n0 99.7716
R9 a_239_74.t0 a_239_74.n1 34.0546
R10 a_239_74.n1 a_239_74.t3 22.7032
R11 VGND VGND.n0 99.4656
R12 VGND.n0 VGND.t0 47.9151
R13 VGND.n0 VGND.t1 47.9151
R14 VNB.t1 VNB.t2 2448.29
R15 VNB.t4 VNB.t3 1824.67
R16 VNB.t0 VNB.t4 1154.86
R17 VNB.t2 VNB.t0 1154.86
R18 VNB VNB.t1 1143.31
R19 C1.n0 C1.t1 265.363
R20 C1.n0 C1.t0 197.05
R21 C1 C1.n0 155.067
R22 Y.n1 Y.n0 306.005
R23 Y.t3 Y.n2 279.738
R24 Y.n3 Y.t3 279.738
R25 Y.n1 Y.t2 243.82
R26 Y.n2 Y.n1 83.2918
R27 Y.n0 Y.t1 47.4916
R28 Y.n0 Y.t0 26.3844
R29 Y.n3 Y 12.6066
R30 Y.n2 Y 4.84898
R31 Y Y.n3 1.74595
R32 a_114_74.n0 a_114_74.t2 462.394
R33 a_114_74.n0 a_114_74.t1 34.0546
R34 a_114_74.t0 a_114_74.n0 22.7032
R35 B2.n0 B2.t1 250.909
R36 B2.n0 B2.t0 220.113
R37 B2 B2.n0 154.081
R38 a_324_368.t0 a_324_368.t1 47.4916
R39 VPB.t4 VPB.t0 464.786
R40 VPB VPB.t4 324.329
R41 VPB.t3 VPB.t1 291.13
R42 VPB.t2 VPB.t3 291.13
R43 VPB.t0 VPB.t2 214.517
R44 VPWR.n1 VPWR.n0 586.256
R45 VPWR.n2 VPWR.n0 585
R46 VPWR.n4 VPWR.n3 273.582
R47 VPWR.n5 VPWR.t1 255.972
R48 VPWR.n3 VPWR.n2 37.8396
R49 VPWR.n3 VPWR.n1 37.8396
R50 VPWR.n1 VPWR.t0 26.3844
R51 VPWR.n2 VPWR.t2 26.3844
R52 VPWR.n5 VPWR.n4 11.7037
R53 VPWR.n4 VPWR.n0 5.65449
R54 VPWR VPWR.n5 0.290733
R55 B1.n0 B1.t0 226.809
R56 B1.n0 B1.t1 197.475
R57 B1 B1.n0 101.273
R58 a_522_368.t0 a_522_368.t1 73.8755
R59 A1.n1 A1.t0 251.151
R60 A1.n0 A1.t1 179.947
R61 A1.n0 A1 177.695
R62 A1.n2 A1.n1 152
R63 A1.n1 A1.n0 24.1005
R64 A1.n2 A1 8.93383
R65 A1 A1.n2 3.86717
C0 Y VGND 0.045907f
C1 VGND VPB 0.009529f
C2 B2 A2 0.086191f
C3 VGND B1 0.008442f
C4 VPWR C1 0.02075f
C5 Y A2 0.08892f
C6 VPWR B2 0.014822f
C7 VPB A2 0.039109f
C8 A1 VGND 0.019094f
C9 B1 A2 3.61e-19
C10 Y VPWR 0.263563f
C11 VPWR VPB 0.121685f
C12 Y C1 0.133516f
C13 VPB C1 0.057907f
C14 A1 A2 0.080857f
C15 Y B2 0.053607f
C16 VPWR B1 0.024707f
C17 C1 B1 0.032111f
C18 VPB B2 0.033095f
C19 B1 B2 0.085595f
C20 A1 VPWR 0.058637f
C21 Y VPB 0.016842f
C22 VGND A2 0.014711f
C23 Y B1 0.102296f
C24 A1 B2 1.11e-19
C25 VPB B1 0.053899f
C26 VPWR VGND 0.062913f
C27 VGND C1 0.01095f
C28 A1 Y 8.4e-19
C29 A1 VPB 0.060574f
C30 VGND B2 0.00899f
C31 A1 B1 5.52e-20
C32 VPWR A2 0.0786f
C33 VGND VNB 0.47734f
C34 VPWR VNB 0.424563f
C35 Y VNB 0.10014f
C36 A1 VNB 0.193422f
C37 A2 VNB 0.111178f
C38 B2 VNB 0.105078f
C39 B1 VNB 0.147508f
C40 C1 VNB 0.186016f
C41 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2111a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2111a_2 VNB VPB VPWR VGND A1 A2 B1 C1 D1 X
X0 a_236_368.t0 A2.t0 a_152_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X1 a_152_368.t1 A1.t0 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X2 VPWR.t2 a_236_368.t5 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_369_74.t0 B1.t0 a_54_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 a_461_74.t1 C1.t0 a_369_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1147 ps=1.05 w=0.74 l=0.15
X5 VPWR.t4 B1.t1 a_236_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.245 pd=1.49 as=0.21 ps=1.42 w=1 l=0.15
X6 X.t0 a_236_368.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4309 ps=1.95 w=1.12 l=0.15
X7 VGND.t3 a_236_368.t7 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=2.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_54_74.t0 A2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 VPWR.t5 D1.t0 a_236_368.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.4309 pd=1.95 as=0.175 ps=1.35 w=1 l=0.15
X10 X.t2 a_236_368.t8 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X11 VGND.t1 A1.t1 a_54_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2627 ps=2.19 w=0.74 l=0.15
X12 a_236_368.t1 C1.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.245 ps=1.49 w=1 l=0.15
X13 a_236_368.t2 D1.t1 a_461_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
R0 A2.n0 A2.t0 266.44
R1 A2.n0 A2.t1 178.34
R2 A2 A2.n0 158.788
R3 a_152_368.t0 a_152_368.t1 53.1905
R4 a_236_368.n6 a_236_368.n5 259.11
R5 a_236_368.n0 a_236_368.t5 240.197
R6 a_236_368.n2 a_236_368.t6 240.197
R7 a_236_368.n5 a_236_368.n4 202.178
R8 a_236_368.n3 a_236_368.t2 196.202
R9 a_236_368.n0 a_236_368.t7 187.412
R10 a_236_368.n1 a_236_368.t8 179.947
R11 a_236_368.n3 a_236_368.n2 168.798
R12 a_236_368.n5 a_236_368.n3 97.8829
R13 a_236_368.n1 a_236_368.n0 56.2338
R14 a_236_368.t0 a_236_368.n6 53.1905
R15 a_236_368.n4 a_236_368.t4 39.4005
R16 a_236_368.n4 a_236_368.t1 29.5505
R17 a_236_368.n6 a_236_368.t3 29.5505
R18 a_236_368.n2 a_236_368.n1 9.49444
R19 VPB.t6 VPB.t1 500.538
R20 VPB VPB.t5 349.866
R21 VPB.t4 VPB.t3 326.882
R22 VPB.t0 VPB.t4 291.13
R23 VPB.t3 VPB.t6 255.376
R24 VPB.t1 VPB.t2 229.839
R25 VPB.t5 VPB.t0 214.517
R26 A1.n0 A1.t0 242.339
R27 A1.n0 A1.t1 156.431
R28 A1.n1 A1.n0 94.8376
R29 A1 A1.n1 10.4704
R30 A1.n1 A1 5.75841
R31 VPWR.n8 VPWR.n7 319.616
R32 VPWR.n3 VPWR.t2 265.825
R33 VPWR.n15 VPWR.t0 256.668
R34 VPWR.n5 VPWR.n4 136.951
R35 VPWR.n4 VPWR.t1 78.103
R36 VPWR.n4 VPWR.t5 70.2531
R37 VPWR.n7 VPWR.t3 57.1305
R38 VPWR.n7 VPWR.t4 39.4005
R39 VPWR.n13 VPWR.n1 36.1417
R40 VPWR.n14 VPWR.n13 36.1417
R41 VPWR.n9 VPWR.n6 36.1417
R42 VPWR.n6 VPWR.n5 17.6946
R43 VPWR.n16 VPWR.n15 13.4417
R44 VPWR.n6 VPWR.n2 9.3005
R45 VPWR.n10 VPWR.n9 9.3005
R46 VPWR.n11 VPWR.n1 9.3005
R47 VPWR.n13 VPWR.n12 9.3005
R48 VPWR.n14 VPWR.n0 9.3005
R49 VPWR.n8 VPWR.n1 7.90638
R50 VPWR.n15 VPWR.n14 7.15344
R51 VPWR.n5 VPWR.n3 3.84167
R52 VPWR.n9 VPWR.n8 3.38874
R53 VPWR.n3 VPWR.n2 0.45173
R54 VPWR.n10 VPWR.n2 0.122949
R55 VPWR.n11 VPWR.n10 0.122949
R56 VPWR.n12 VPWR.n11 0.122949
R57 VPWR.n12 VPWR.n0 0.122949
R58 VPWR.n16 VPWR.n0 0.122949
R59 VPWR VPWR.n16 0.0617245
R60 X.n1 X.n0 268.474
R61 X.n2 X.n1 185
R62 X.n3 X.n2 185
R63 X.n0 X.t1 26.3844
R64 X.n0 X.t0 26.3844
R65 X.n2 X.t3 22.7032
R66 X.n2 X.t2 22.7032
R67 X.n3 X 12.6066
R68 X.n1 X 4.84898
R69 X X.n3 1.74595
R70 B1.n0 B1.t1 266.44
R71 B1.n0 B1.t0 178.34
R72 B1 B1.n0 158.4
R73 a_54_74.n0 a_54_74.t2 288.014
R74 a_54_74.t0 a_54_74.n0 34.0546
R75 a_54_74.n0 a_54_74.t1 22.7032
R76 a_369_74.t0 a_369_74.t1 50.2708
R77 VNB.t5 VNB.t3 2448.29
R78 VNB VNB.t2 1616.8
R79 VNB.t6 VNB.t5 1316.54
R80 VNB.t2 VNB.t0 1316.54
R81 VNB.t0 VNB.t1 1154.86
R82 VNB.t1 VNB.t6 1062.47
R83 VNB.t3 VNB.t4 993.177
R84 C1.n0 C1.t1 231.629
R85 C1.n0 C1.t0 220.113
R86 C1 C1.n0 158.995
R87 a_461_74.t0 a_461_74.t1 68.1086
R88 VGND.n3 VGND.t2 232.139
R89 VGND.n11 VGND.n10 199.844
R90 VGND.n2 VGND.t3 174.583
R91 VGND.n4 VGND.n1 36.1417
R92 VGND.n8 VGND.n1 36.1417
R93 VGND.n9 VGND.n8 36.1417
R94 VGND.n11 VGND.n9 34.6358
R95 VGND.n10 VGND.t0 34.0546
R96 VGND.n10 VGND.t1 34.0546
R97 VGND.n4 VGND.n3 21.8358
R98 VGND.n9 VGND.n0 9.3005
R99 VGND.n8 VGND.n7 9.3005
R100 VGND.n6 VGND.n1 9.3005
R101 VGND.n5 VGND.n4 9.3005
R102 VGND.n3 VGND.n2 6.79888
R103 VGND.n12 VGND.n11 4.77522
R104 VGND.n5 VGND.n2 0.584371
R105 VGND VGND.n12 0.237916
R106 VGND.n12 VGND.n0 0.192318
R107 VGND.n6 VGND.n5 0.122949
R108 VGND.n7 VGND.n6 0.122949
R109 VGND.n7 VGND.n0 0.122949
R110 D1.n0 D1.t0 222.534
R111 D1.n0 D1.t1 211.019
R112 D1 D1.n0 154.522
C0 X VGND 0.142586f
C1 D1 VPWR 0.022022f
C2 D1 B1 4.21e-19
C3 VPWR A2 0.018588f
C4 VPB VPWR 0.172816f
C5 A2 B1 0.076099f
C6 VPB B1 0.034058f
C7 C1 VPWR 0.016249f
C8 VGND VPWR 0.093034f
C9 C1 B1 0.06557f
C10 VPWR A1 0.050584f
C11 VGND B1 0.014068f
C12 VPB D1 0.049658f
C13 VPB A2 0.031631f
C14 VGND D1 0.012999f
C15 C1 D1 0.094945f
C16 X VPWR 0.195277f
C17 C1 A2 5.21e-19
C18 VGND A2 0.015525f
C19 VPB C1 0.038466f
C20 VGND VPB 0.011667f
C21 A1 A2 0.087828f
C22 VPB A1 0.052803f
C23 VGND C1 0.021666f
C24 X D1 5.48e-19
C25 C1 A1 2.95e-19
C26 VGND A1 0.018764f
C27 X VPB 0.005949f
C28 VPWR B1 0.013664f
C29 VGND VNB 0.64239f
C30 X VNB 0.029702f
C31 VPWR VNB 0.55281f
C32 D1 VNB 0.130758f
C33 C1 VNB 0.113758f
C34 B1 VNB 0.109089f
C35 A2 VNB 0.10597f
C36 A1 VNB 0.190715f
C37 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2111a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2111a_4 VNB VPB VPWR VGND D1 C1 B1 A2 A1 X
X0 VPWR.t10 D1.t0 a_27_392.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VPWR.t5 C1.t0 a_27_392.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.126 ps=1.14 w=0.84 l=0.15
X2 a_27_392.t7 D1.t1 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X3 X.t3 a_27_392.t10 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4 a_477_198.t1 A1.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_27_392.t9 D1.t2 a_27_74.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6 a_27_392.t2 A2.t0 a_747_392.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X7 VPWR.t3 a_27_392.t11 X.t7 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_477_198.t3 A2.t1 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2183 pd=2.07 as=0.1258 ps=1.08 w=0.74 l=0.15
X9 X.t6 a_27_392.t12 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t0 a_27_392.t13 X.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t1 a_27_392.t14 X.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X12 a_287_74.t1 B1.t0 a_477_198.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.21835 ps=2.21 w=0.74 l=0.15
X13 a_27_74.t1 C1.t1 a_287_74.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.24285 pd=2.49 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_747_392.t2 A2.t2 a_27_392.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.2103 ps=1.435 w=1 l=0.15
X15 X.t1 a_27_392.t15 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 X.t4 a_27_392.t16 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2084 ps=1.505 w=1.12 l=0.15
X17 a_27_74.t2 D1.t3 a_27_392.t8 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_477_198.t5 B1.t1 a_287_74.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_27_392.t4 C1.t2 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1974 pd=1.31 as=0.147 ps=1.19 w=0.84 l=0.15
X20 VPWR.t7 A1.t1 a_747_392.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2084 pd=1.505 as=0.15 ps=1.3 w=1 l=0.15
X21 a_287_74.t2 C1.t3 a_27_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_747_392.t0 A1.t2 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.345 ps=2.69 w=1 l=0.15
X23 VGND.t2 a_27_392.t17 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_27_392.t5 B1.t2 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2103 pd=1.435 as=0.126 ps=1.14 w=0.84 l=0.15
X25 VGND.t7 A1.t3 a_477_198.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 VPWR.t4 B1.t3 a_27_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1974 ps=1.31 w=0.84 l=0.15
X27 VGND.t4 A2.t3 a_477_198.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 D1.n0 D1.t3 285.988
R1 D1.n2 D1.t2 249.356
R2 D1.n0 D1.t1 227.344
R3 D1.n1 D1.t0 196.817
R4 D1 D1.n2 160.922
R5 D1.n1 D1.n0 107.647
R6 D1.n2 D1.n1 11.5685
R7 a_27_392.t2 a_27_392.n21 879.801
R8 a_27_392.n21 a_27_392.n20 593.566
R9 a_27_392.n1 a_27_392.t6 417.976
R10 a_27_392.n3 a_27_392.n2 300.748
R11 a_27_392.n5 a_27_392.n4 300.454
R12 a_27_392.n19 a_27_392.n18 289.051
R13 a_27_392.n7 a_27_392.t11 287.861
R14 a_27_392.n1 a_27_392.n0 253.518
R15 a_27_392.n8 a_27_392.t12 226.809
R16 a_27_392.n11 a_27_392.t14 226.809
R17 a_27_392.n14 a_27_392.t16 226.809
R18 a_27_392.n17 a_27_392.n16 217.851
R19 a_27_392.n14 a_27_392.t15 209.359
R20 a_27_392.n7 a_27_392.t13 196.013
R21 a_27_392.n13 a_27_392.t17 196.013
R22 a_27_392.n9 a_27_392.t10 196.013
R23 a_27_392.n10 a_27_392.n6 165.189
R24 a_27_392.n16 a_27_392.n15 152
R25 a_27_392.n12 a_27_392.n6 152
R26 a_27_392.n8 a_27_392.n7 115.972
R27 a_27_392.n17 a_27_392.n5 55.7181
R28 a_27_392.n19 a_27_392.t5 55.1136
R29 a_27_392.n4 a_27_392.t0 55.1136
R30 a_27_392.n4 a_27_392.t4 55.1136
R31 a_27_392.n5 a_27_392.n3 53.0829
R32 a_27_392.n15 a_27_392.n13 41.6278
R33 a_27_392.n11 a_27_392.n10 37.246
R34 a_27_392.n2 a_27_392.t1 35.1791
R35 a_27_392.n2 a_27_392.t7 35.1791
R36 a_27_392.n20 a_27_392.t3 33.8801
R37 a_27_392.n10 a_27_392.n9 25.5611
R38 a_27_392.n3 a_27_392.n1 23.3417
R39 a_27_392.n0 a_27_392.t8 22.7032
R40 a_27_392.n0 a_27_392.t9 22.7032
R41 a_27_392.n21 a_27_392.n18 20.0884
R42 a_27_392.n16 a_27_392.n6 13.1884
R43 a_27_392.n12 a_27_392.n11 12.4157
R44 a_27_392.n15 a_27_392.n14 10.955
R45 a_27_392.n18 a_27_392.n17 10.0035
R46 a_27_392.n13 a_27_392.n12 8.03383
R47 a_27_392.n20 a_27_392.n19 5.8636
R48 a_27_392.n9 a_27_392.n8 2.92171
R49 VPWR.n17 VPWR.t11 802.365
R50 VPWR.n32 VPWR.n1 617.971
R51 VPWR.n30 VPWR.n3 617.971
R52 VPWR.n24 VPWR.n23 617.971
R53 VPWR.n11 VPWR.n10 316.116
R54 VPWR.n15 VPWR.n9 315.928
R55 VPWR.n12 VPWR.t3 265.527
R56 VPWR.n1 VPWR.t9 46.9053
R57 VPWR.n1 VPWR.t10 46.9053
R58 VPWR.n3 VPWR.t5 46.9053
R59 VPWR.n9 VPWR.t7 46.2955
R60 VPWR.n29 VPWR.n4 36.1417
R61 VPWR.n21 VPWR.n6 36.1417
R62 VPWR.n22 VPWR.n21 36.1417
R63 VPWR.n25 VPWR.n22 36.1417
R64 VPWR.n3 VPWR.t6 35.1791
R65 VPWR.n23 VPWR.t8 35.1791
R66 VPWR.n23 VPWR.t4 35.1791
R67 VPWR.n31 VPWR.n30 31.2476
R68 VPWR.n17 VPWR.n16 30.8711
R69 VPWR.n9 VPWR.t0 27.5507
R70 VPWR.n10 VPWR.t2 26.3844
R71 VPWR.n10 VPWR.t1 26.3844
R72 VPWR.n15 VPWR.n14 25.224
R73 VPWR.n16 VPWR.n15 22.2123
R74 VPWR.n14 VPWR.n11 21.4593
R75 VPWR.n32 VPWR.n31 19.2005
R76 VPWR.n17 VPWR.n6 16.5652
R77 VPWR.n30 VPWR.n29 16.1887
R78 VPWR.n14 VPWR.n13 9.3005
R79 VPWR.n15 VPWR.n8 9.3005
R80 VPWR.n16 VPWR.n7 9.3005
R81 VPWR.n18 VPWR.n17 9.3005
R82 VPWR.n19 VPWR.n6 9.3005
R83 VPWR.n21 VPWR.n20 9.3005
R84 VPWR.n22 VPWR.n5 9.3005
R85 VPWR.n26 VPWR.n25 9.3005
R86 VPWR.n27 VPWR.n4 9.3005
R87 VPWR.n29 VPWR.n28 9.3005
R88 VPWR.n30 VPWR.n2 9.3005
R89 VPWR.n31 VPWR.n0 9.3005
R90 VPWR.n25 VPWR.n24 7.90638
R91 VPWR.n33 VPWR.n32 7.43488
R92 VPWR.n12 VPWR.n11 6.75308
R93 VPWR.n24 VPWR.n4 3.38874
R94 VPWR.n13 VPWR.n12 0.636608
R95 VPWR VPWR.n33 0.160103
R96 VPWR.n33 VPWR.n0 0.1477
R97 VPWR.n13 VPWR.n8 0.122949
R98 VPWR.n8 VPWR.n7 0.122949
R99 VPWR.n18 VPWR.n7 0.122949
R100 VPWR.n19 VPWR.n18 0.122949
R101 VPWR.n20 VPWR.n19 0.122949
R102 VPWR.n20 VPWR.n5 0.122949
R103 VPWR.n26 VPWR.n5 0.122949
R104 VPWR.n27 VPWR.n26 0.122949
R105 VPWR.n28 VPWR.n27 0.122949
R106 VPWR.n28 VPWR.n2 0.122949
R107 VPWR.n2 VPWR.n0 0.122949
R108 VPB.t6 VPB.t13 541.399
R109 VPB.t8 VPB.t4 316.668
R110 VPB.t10 VPB.t7 298.791
R111 VPB.t12 VPB.t11 280.914
R112 VPB.t9 VPB.t0 273.253
R113 VPB VPB.t12 257.93
R114 VPB.t0 VPB.t1 255.376
R115 VPB.t7 VPB.t6 255.376
R116 VPB.t5 VPB.t8 255.376
R117 VPB.t2 VPB.t3 229.839
R118 VPB.t1 VPB.t2 229.839
R119 VPB.t13 VPB.t9 229.839
R120 VPB.t4 VPB.t10 229.839
R121 VPB.t11 VPB.t5 229.839
R122 C1.n1 C1.t2 221.756
R123 C1.n1 C1.t0 204.851
R124 C1.n0 C1.t3 158.089
R125 C1.n2 C1.n1 152
R126 C1.n0 C1.t1 148.26
R127 C1.n1 C1.n0 40.3544
R128 C1.n2 C1 18.0369
R129 C1 C1.n2 0.582318
R130 VGND.n5 VGND.t0 250.821
R131 VGND.n1 VGND.n0 213.315
R132 VGND.n7 VGND.n6 210.213
R133 VGND.n14 VGND.t6 138.363
R134 VGND.n10 VGND.n9 116.644
R135 VGND.n16 VGND.n15 36.1417
R136 VGND.n10 VGND.n8 35.0123
R137 VGND.n6 VGND.t1 34.0546
R138 VGND.n6 VGND.t2 34.0546
R139 VGND.n9 VGND.t3 34.0546
R140 VGND.n0 VGND.t5 32.4329
R141 VGND.n14 VGND.n3 27.4829
R142 VGND.n9 VGND.t7 22.7032
R143 VGND.n0 VGND.t4 22.7032
R144 VGND.n15 VGND.n14 19.9534
R145 VGND.n18 VGND.n1 17.8152
R146 VGND.n8 VGND.n7 15.4358
R147 VGND.n10 VGND.n3 12.424
R148 VGND.n17 VGND.n16 9.3005
R149 VGND.n15 VGND.n2 9.3005
R150 VGND.n14 VGND.n13 9.3005
R151 VGND.n12 VGND.n3 9.3005
R152 VGND.n8 VGND.n4 9.3005
R153 VGND.n11 VGND.n10 9.3005
R154 VGND.n7 VGND.n5 7.03723
R155 VGND.n16 VGND.n1 1.12991
R156 VGND VGND.n18 0.896606
R157 VGND.n5 VGND.n4 0.600107
R158 VGND.n18 VGND.n17 0.149471
R159 VGND.n11 VGND.n4 0.122949
R160 VGND.n12 VGND.n11 0.122949
R161 VGND.n13 VGND.n12 0.122949
R162 VGND.n13 VGND.n2 0.122949
R163 VGND.n17 VGND.n2 0.122949
R164 X.n2 X.n0 237.975
R165 X.n2 X.n1 201.84
R166 X.n5 X.n3 152.159
R167 X.n5 X.n4 101.71
R168 X X.n2 54.4613
R169 X.n0 X.t4 35.1791
R170 X X.n5 28.2358
R171 X.n1 X.t7 26.3844
R172 X.n1 X.t6 26.3844
R173 X.n0 X.t5 26.3844
R174 X.n3 X.t0 22.7032
R175 X.n3 X.t1 22.7032
R176 X.n4 X.t2 22.7032
R177 X.n4 X.t3 22.7032
R178 VNB.t8 VNB.t9 2390.55
R179 VNB.t5 VNB.t6 2379
R180 VNB.t0 VNB.t3 1316.54
R181 VNB.t12 VNB.t1 1154.86
R182 VNB VNB.t11 1154.86
R183 VNB.t4 VNB.t5 1131.76
R184 VNB.t3 VNB.t2 993.177
R185 VNB.t1 VNB.t0 993.177
R186 VNB.t6 VNB.t12 993.177
R187 VNB.t13 VNB.t4 993.177
R188 VNB.t9 VNB.t13 993.177
R189 VNB.t7 VNB.t8 993.177
R190 VNB.t10 VNB.t7 993.177
R191 VNB.t11 VNB.t10 993.177
R192 A1.n1 A1.t0 230.339
R193 A1.n0 A1.t3 228.148
R194 A1.n0 A1.t1 218.362
R195 A1.n1 A1.t2 212.883
R196 A1 A1.n2 154.133
R197 A1.n2 A1.n1 39.4369
R198 A1.n2 A1.n0 21.1793
R199 a_477_198.n1 a_477_198.t4 268.022
R200 a_477_198.n3 a_477_198.n2 175.555
R201 a_477_198.n2 a_477_198.t3 143.228
R202 a_477_198.n1 a_477_198.n0 100.257
R203 a_477_198.n2 a_477_198.n1 52.7365
R204 a_477_198.n0 a_477_198.t2 22.7032
R205 a_477_198.n0 a_477_198.t5 22.7032
R206 a_477_198.n3 a_477_198.t0 22.7032
R207 a_477_198.t1 a_477_198.n3 22.7032
R208 a_27_74.n0 a_27_74.t1 338.115
R209 a_27_74.n0 a_27_74.t3 174.082
R210 a_27_74.n1 a_27_74.n0 98.896
R211 a_27_74.n1 a_27_74.t0 22.7032
R212 a_27_74.t2 a_27_74.n1 22.7032
R213 A2.n3 A2.t2 216.536
R214 A2.n1 A2.t0 212.883
R215 A2.n1 A2.t1 175.712
R216 A2.n3 A2.t3 173.52
R217 A2.n2 A2.n0 152
R218 A2.n5 A2.n4 152
R219 A2.n4 A2.n2 49.6611
R220 A2.n0 A2 15.5157
R221 A2.n2 A2.n1 12.4157
R222 A2 A2.n5 10.0853
R223 A2.n5 A2 8.53383
R224 A2.n4 A2.n3 7.30353
R225 A2 A2.n0 3.10353
R226 a_747_392.n1 a_747_392.n0 981.412
R227 a_747_392.n0 a_747_392.t3 39.4005
R228 a_747_392.n0 a_747_392.t2 29.5505
R229 a_747_392.t1 a_747_392.n1 29.5505
R230 a_747_392.n1 a_747_392.t0 29.5505
R231 B1.n0 B1.t3 229.462
R232 B1.n2 B1.t1 188.857
R233 B1.n1 B1.t2 187.178
R234 B1.n0 B1.t0 173.52
R235 B1 B1.n2 156.462
R236 B1.n1 B1.n0 36.5157
R237 B1.n2 B1.n1 10.955
R238 a_287_74.n1 a_287_74.n0 465.274
R239 a_287_74.n0 a_287_74.t3 22.7032
R240 a_287_74.n0 a_287_74.t2 22.7032
R241 a_287_74.n1 a_287_74.t0 22.7032
R242 a_287_74.t1 a_287_74.n1 22.7032
C0 D1 VPWR 0.031677f
C1 VPWR VGND 0.132594f
C2 B1 VPWR 0.028568f
C3 D1 VGND 0.011262f
C4 A1 VPWR 0.032374f
C5 B1 VGND 0.014398f
C6 VPWR X 0.399269f
C7 VPWR VPB 0.249774f
C8 C1 VPWR 0.034147f
C9 D1 X 2.13e-21
C10 A1 VGND 0.042044f
C11 X VGND 0.340904f
C12 D1 VPB 0.098882f
C13 VGND VPB 0.015949f
C14 A2 VPWR 0.014513f
C15 D1 C1 0.065098f
C16 B1 X 5.79e-20
C17 C1 VGND 0.014144f
C18 B1 VPB 0.091519f
C19 C1 B1 0.032862f
C20 A1 X 0.002109f
C21 A2 VGND 0.030645f
C22 A1 VPB 0.083615f
C23 X VPB 0.012854f
C24 A1 C1 0.00147f
C25 A2 B1 0.074218f
C26 C1 X 1.22e-20
C27 C1 VPB 0.086646f
C28 A2 A1 0.051784f
C29 A2 X 2.91e-19
C30 A2 VPB 0.096588f
C31 VGND VNB 0.983282f
C32 X VNB 0.063877f
C33 VPWR VNB 0.786805f
C34 B1 VNB 0.18987f
C35 C1 VNB 0.219298f
C36 D1 VNB 0.261256f
C37 A1 VNB 0.205947f
C38 A2 VNB 0.197956f
C39 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2111ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2111ai_1 VNB VPB VPWR VGND Y D1 C1 B1 A2 A1
X0 VPWR.t1 A1.t0 a_490_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1708 ps=1.425 w=1.12 l=0.15
X1 a_368_74.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1628 ps=1.18 w=0.74 l=0.15
X2 Y.t3 B1.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.182 pd=1.445 as=0.2688 ps=1.6 w=1.12 l=0.15
X3 a_368_74.t2 B1.t1 a_260_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.1443 ps=1.13 w=0.74 l=0.15
X4 a_182_74.t0 D1.t0 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.4625 ps=2.73 w=0.74 l=0.15
X5 VGND.t1 A2.t0 a_368_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.1332 ps=1.1 w=0.74 l=0.15
X6 a_260_74.t0 C1.t0 a_182_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0888 ps=0.98 w=0.74 l=0.15
X7 VPWR.t2 C1.t1 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2688 pd=1.6 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_490_368.t1 A2.t1 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.182 ps=1.445 w=1.12 l=0.15
X9 Y.t0 D1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
R0 A1.n0 A1.t0 277.062
R1 A1.n0 A1.t1 169.684
R2 A1 A1.n0 158.788
R3 a_490_368.t0 a_490_368.t1 53.6478
R4 VPWR.n3 VPWR.t1 257.144
R5 VPWR.n7 VPWR.t0 256.943
R6 VPWR.n2 VPWR.n1 221.766
R7 VPWR.n1 VPWR.t2 53.6478
R8 VPWR.n6 VPWR.n5 36.1417
R9 VPWR.n1 VPWR.t3 30.7817
R10 VPWR.n5 VPWR.n2 21.4593
R11 VPWR.n8 VPWR.n7 19.8417
R12 VPWR.n5 VPWR.n4 9.3005
R13 VPWR.n6 VPWR.n0 9.3005
R14 VPWR.n3 VPWR.n2 7.17169
R15 VPWR.n7 VPWR.n6 0.753441
R16 VPWR.n4 VPWR.n3 0.243906
R17 VPWR.n4 VPWR.n0 0.122949
R18 VPWR.n8 VPWR.n0 0.122949
R19 VPWR VPWR.n8 0.0617245
R20 VPB VPB.t0 418.817
R21 VPB.t2 VPB.t4 321.774
R22 VPB.t4 VPB.t3 242.608
R23 VPB.t3 VPB.t1 232.393
R24 VPB.t0 VPB.t2 229.839
R25 VGND VGND.n0 206.742
R26 VGND.n0 VGND.t0 41.3519
R27 VGND.n0 VGND.t1 30.0005
R28 a_368_74.t0 a_368_74.n0 292.69
R29 a_368_74.n0 a_368_74.t1 34.0546
R30 a_368_74.n0 a_368_74.t2 24.3248
R31 VNB VNB.t4 1928.61
R32 VNB.t1 VNB.t0 1362.73
R33 VNB.t3 VNB.t2 1247.24
R34 VNB.t2 VNB.t1 1177.95
R35 VNB.t4 VNB.t3 900.788
R36 B1.n0 B1.t0 285.719
R37 B1.n0 B1.t1 178.34
R38 B1 B1.n0 159.958
R39 Y.n3 Y 588.678
R40 Y.n3 Y.n0 585
R41 Y.n4 Y.n3 585
R42 Y.n2 Y.n1 261.149
R43 Y.n2 Y.t2 173.951
R44 Y.n1 Y.t3 30.7817
R45 Y.n3 Y.t1 26.3844
R46 Y.n3 Y.t0 26.3844
R47 Y.n1 Y.t4 26.3844
R48 Y Y.n4 9.85797
R49 Y Y.n0 8.53383
R50 Y Y.n2 4.26717
R51 Y Y.n0 2.35452
R52 Y.n4 Y 1.03039
R53 a_260_74.t0 a_260_74.t1 63.2437
R54 D1.n0 D1.t1 285.719
R55 D1.n0 D1.t0 178.34
R56 D1 D1.n0 158.788
R57 a_182_74.t0 a_182_74.t1 38.9194
R58 A2.n0 A2.t1 285.719
R59 A2.n0 A2.t0 178.34
R60 A2 A2.n0 158.573
R61 C1.n0 C1.t1 285.719
R62 C1.n0 C1.t0 178.34
R63 C1 C1.n0 158.589
C0 B1 VPWR 0.023131f
C1 VPB VPWR 0.120197f
C2 B1 VPB 0.031612f
C3 A1 VGND 0.015194f
C4 C1 VGND 0.034067f
C5 A1 C1 1.9e-19
C6 Y VGND 0.08015f
C7 A1 Y 0.005706f
C8 A2 VGND 0.016729f
C9 A2 A1 0.09433f
C10 D1 VGND 0.012664f
C11 C1 Y 0.092859f
C12 A2 C1 4.47e-19
C13 D1 C1 0.100245f
C14 VPWR VGND 0.056469f
C15 A1 VPWR 0.049371f
C16 B1 VGND 0.014702f
C17 A2 Y 0.024925f
C18 D1 Y 0.1028f
C19 VPB VGND 0.008153f
C20 C1 VPWR 0.009366f
C21 A1 VPB 0.041533f
C22 B1 C1 0.085898f
C23 VPB C1 0.031139f
C24 VPWR Y 0.446027f
C25 B1 Y 0.056897f
C26 A2 VPWR 0.023843f
C27 B1 A2 0.08466f
C28 D1 VPWR 0.019498f
C29 VPB Y 0.026559f
C30 A2 VPB 0.030865f
C31 VPB D1 0.034597f
C32 VGND VNB 0.431477f
C33 Y VNB 0.096522f
C34 VPWR VNB 0.417862f
C35 A1 VNB 0.170352f
C36 A2 VNB 0.107762f
C37 B1 VNB 0.107256f
C38 C1 VNB 0.110628f
C39 D1 VNB 0.133908f
C40 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2111ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2111ai_2 VNB VPB VPWR VGND D1 C1 B1 A2 A1 Y
X0 VPWR.t3 D1.t0 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_510_74.t2 B1.t0 a_299_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2 a_697_368.t3 A1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X3 a_510_74.t4 A1.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 VPWR.t0 A1.t2 a_697_368.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_299_74.t0 B1.t1 a_510_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_510_74.t0 A2.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.111 ps=1.04 w=0.74 l=0.15
X7 a_697_368.t1 A2.t1 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Y.t0 A2.t2 a_697_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X9 Y.t3 D1.t1 a_40_74.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 Y.t4 D1.t2 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X11 VGND.t2 A1.t3 a_510_74.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VPWR.t6 B1.t2 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X13 Y.t9 B1.t3 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR.t4 C1.t0 Y.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Y.t7 C1.t1 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X16 a_40_74.t3 C1.t2 a_299_74.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 VGND.t1 A2.t3 a_510_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_40_74.t1 D1.t3 Y.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_299_74.t2 C1.t3 a_40_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 D1.n0 D1.t0 262.349
R1 D1.n2 D1.t2 261.62
R2 D1 D1.n2 198.956
R3 D1.n1 D1.t1 154.24
R4 D1.n0 D1.t3 154.24
R5 D1.n1 D1.n0 62.8066
R6 D1.n2 D1.n1 2.19141
R7 Y.n8 Y 589.85
R8 Y.n8 Y.n0 585
R9 Y.n9 Y.n8 585
R10 Y.n3 Y.n1 385.033
R11 Y.n3 Y.n2 205.487
R12 Y Y.n6 202.601
R13 Y.n5 Y.n4 202.457
R14 Y.n7 Y.n5 51.8262
R15 Y.n5 Y.n3 43.5898
R16 Y.n8 Y.t5 26.3844
R17 Y.n8 Y.t4 26.3844
R18 Y.n4 Y.t6 26.3844
R19 Y.n4 Y.t7 26.3844
R20 Y.n1 Y.t1 26.3844
R21 Y.n1 Y.t0 26.3844
R22 Y.n2 Y.t8 26.3844
R23 Y.n2 Y.t9 26.3844
R24 Y.n6 Y.t2 22.7032
R25 Y.n6 Y.t3 22.7032
R26 Y Y.n9 12.9944
R27 Y.n7 Y 11.8308
R28 Y Y.n0 11.249
R29 Y Y.n0 3.10353
R30 Y Y.n7 2.52171
R31 Y.n9 Y 1.35808
R32 VPWR.n6 VPWR.t6 349.789
R33 VPWR.n8 VPWR.n7 331.5
R34 VPWR.n14 VPWR.n2 325.255
R35 VPWR.n5 VPWR.n4 322.154
R36 VPWR.n16 VPWR.t2 259.171
R37 VPWR.n13 VPWR.n3 36.1417
R38 VPWR.n9 VPWR.n8 35.3887
R39 VPWR.n2 VPWR.t3 35.1791
R40 VPWR.n4 VPWR.t1 35.1791
R41 VPWR.n15 VPWR.n14 28.9887
R42 VPWR.n2 VPWR.t5 26.3844
R43 VPWR.n7 VPWR.t7 26.3844
R44 VPWR.n7 VPWR.t4 26.3844
R45 VPWR.n4 VPWR.t0 26.3844
R46 VPWR.n9 VPWR.n6 25.977
R47 VPWR.n14 VPWR.n13 24.4711
R48 VPWR.n16 VPWR.n15 23.7181
R49 VPWR.n10 VPWR.n9 9.3005
R50 VPWR.n11 VPWR.n3 9.3005
R51 VPWR.n13 VPWR.n12 9.3005
R52 VPWR.n14 VPWR.n1 9.3005
R53 VPWR.n15 VPWR.n0 9.3005
R54 VPWR.n17 VPWR.n16 9.3005
R55 VPWR.n6 VPWR.n5 7.31736
R56 VPWR.n8 VPWR.n3 0.753441
R57 VPWR.n10 VPWR.n5 0.167001
R58 VPWR.n11 VPWR.n10 0.122949
R59 VPWR.n12 VPWR.n11 0.122949
R60 VPWR.n12 VPWR.n1 0.122949
R61 VPWR.n1 VPWR.n0 0.122949
R62 VPWR.n17 VPWR.n0 0.122949
R63 VPWR VPWR.n17 0.0617245
R64 VPB.t8 VPB.t2 515.861
R65 VPB VPB.t4 278.361
R66 VPB.t0 VPB.t1 255.376
R67 VPB.t5 VPB.t7 255.376
R68 VPB.t3 VPB.t0 229.839
R69 VPB.t2 VPB.t3 229.839
R70 VPB.t9 VPB.t8 229.839
R71 VPB.t6 VPB.t9 229.839
R72 VPB.t7 VPB.t6 229.839
R73 VPB.t4 VPB.t5 229.839
R74 B1.n0 B1.t3 343.356
R75 B1.n0 B1.t2 227.712
R76 B1.n4 B1.t0 213.542
R77 B1.n1 B1.t1 196.013
R78 B1.n5 B1.n4 152
R79 B1.n3 B1.n2 152
R80 B1.n4 B1.n3 49.6611
R81 B1.n2 B1 11.7586
R82 B1.n1 B1.n0 7.9791
R83 B1.n5 B1 7.5912
R84 B1 B1.n5 6.69817
R85 B1.n3 B1.n1 5.84292
R86 B1.n2 B1 2.53073
R87 a_299_74.n1 a_299_74.n0 482.2
R88 a_299_74.n0 a_299_74.t3 34.0546
R89 a_299_74.t0 a_299_74.n1 34.0546
R90 a_299_74.n0 a_299_74.t2 22.7032
R91 a_299_74.n1 a_299_74.t1 22.7032
R92 a_510_74.n2 a_510_74.t1 274.418
R93 a_510_74.n1 a_510_74.t4 203.258
R94 a_510_74.n1 a_510_74.n0 104.579
R95 a_510_74.n3 a_510_74.n2 103.65
R96 a_510_74.n2 a_510_74.n1 59.8593
R97 a_510_74.n0 a_510_74.t5 22.7032
R98 a_510_74.n0 a_510_74.t0 22.7032
R99 a_510_74.n3 a_510_74.t3 22.7032
R100 a_510_74.t2 a_510_74.n3 22.7032
R101 VNB.t9 VNB.t1 2286.61
R102 VNB VNB.t7 1293.44
R103 VNB.t8 VNB.t4 1154.86
R104 VNB.t1 VNB.t2 1154.86
R105 VNB.t5 VNB.t9 1154.86
R106 VNB.t3 VNB.t0 1039.37
R107 VNB.t0 VNB.t8 993.177
R108 VNB.t2 VNB.t3 993.177
R109 VNB.t6 VNB.t5 993.177
R110 VNB.t7 VNB.t6 993.177
R111 A1.n2 A1.t0 250.909
R112 A1.n0 A1.t2 230.825
R113 A1.n1 A1.t1 218.654
R114 A1.n0 A1.t3 201.998
R115 A1.n3 A1.n2 152
R116 A1.n1 A1.n0 50.4957
R117 A1.n3 A1 8.7819
R118 A1 A1.n3 5.50748
R119 A1.n2 A1.n1 1.46111
R120 a_697_368.n0 a_697_368.t0 425.627
R121 a_697_368.n0 a_697_368.t3 315.962
R122 a_697_368.n1 a_697_368.n0 183.911
R123 a_697_368.t2 a_697_368.n1 26.3844
R124 a_697_368.n1 a_697_368.t1 26.3844
R125 VGND.n2 VGND.n0 213.803
R126 VGND.n2 VGND.n1 213.524
R127 VGND.n0 VGND.t2 34.0546
R128 VGND.n1 VGND.t0 25.9464
R129 VGND.n0 VGND.t3 22.7032
R130 VGND.n1 VGND.t1 22.7032
R131 VGND VGND.n2 1.36436
R132 A2.n0 A2.t1 229
R133 A2.n1 A2.t2 226.809
R134 A2.n1 A2.t3 198.204
R135 A2.n0 A2.t0 196.013
R136 A2.n3 A2.n2 152
R137 A2.n2 A2.n1 40.1672
R138 A2.n2 A2.n0 23.3702
R139 A2 A2.n3 10.2703
R140 A2.n3 A2 4.0191
R141 a_40_74.n1 a_40_74.t3 280.728
R142 a_40_74.t2 a_40_74.n1 217.006
R143 a_40_74.n1 a_40_74.n0 86.7629
R144 a_40_74.n0 a_40_74.t0 22.7032
R145 a_40_74.n0 a_40_74.t1 22.7032
R146 C1.n1 C1.t0 243.849
R147 C1.n3 C1.t1 240.197
R148 C1.n3 C1.t3 190.901
R149 C1.n1 C1.t2 179.947
R150 C1.n2 C1.n0 158.595
R151 C1 C1.n4 155.298
R152 C1.n4 C1.n2 49.6611
R153 C1.n2 C1.n1 10.2247
R154 C1.n0 C1 5.0092
R155 C1 C1.n0 3.29747
R156 C1.n4 C1.n3 2.19141
C0 VPWR Y 0.614205f
C1 VGND Y 0.015498f
C2 Y B1 0.145684f
C3 VPWR A2 0.013359f
C4 VPWR D1 0.059219f
C5 Y VPB 0.028192f
C6 VGND A2 0.037027f
C7 B1 A2 0.081869f
C8 VGND D1 0.015447f
C9 D1 B1 1.52e-19
C10 VPB A2 0.065901f
C11 VPB D1 0.076402f
C12 A1 Y 8.65e-20
C13 VGND VPWR 0.093095f
C14 A1 A2 0.095541f
C15 Y C1 0.119731f
C16 VPWR B1 0.035072f
C17 VPWR VPB 0.171176f
C18 VGND B1 0.019263f
C19 C1 A2 1.8e-19
C20 VGND VPB 0.009401f
C21 VPB B1 0.096861f
C22 D1 C1 0.057779f
C23 A1 VPWR 0.04048f
C24 VGND A1 0.036553f
C25 VPWR C1 0.031404f
C26 A1 VPB 0.073443f
C27 VGND C1 0.015543f
C28 C1 B1 0.050045f
C29 VPB C1 0.061534f
C30 A1 C1 9.18e-20
C31 Y A2 0.053769f
C32 Y D1 0.114909f
C33 VGND VNB 0.667695f
C34 Y VNB 0.030642f
C35 VPWR VNB 0.585444f
C36 A1 VNB 0.254373f
C37 A2 VNB 0.19043f
C38 B1 VNB 0.251609f
C39 C1 VNB 0.215426f
C40 D1 VNB 0.273993f
C41 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2_1 VNB VPB VPWR VGND B A X
X0 VGND.t2 A.t0 a_63_368.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.130625 ps=1.025 w=0.55 l=0.15
X1 VPWR.t1 A.t1 a_152_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3346 pd=1.76 as=0.1134 ps=1.11 w=0.84 l=0.15
X2 a_152_368.t0 B.t0 a_63_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.2478 ps=2.27 w=0.84 l=0.15
X3 X.t0 a_63_368.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X4 X.t1 a_63_368.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3346 ps=1.76 w=1.12 l=0.15
X5 a_63_368.t1 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.130625 pd=1.025 as=0.2695 ps=2.08 w=0.55 l=0.15
R0 A.n0 A.t1 204.041
R1 A.n0 A.t0 187.889
R2 A A.n0 154.828
R3 a_63_368.t0 a_63_368.n2 500.592
R4 a_63_368.n1 a_63_368.t4 263.25
R5 a_63_368.n2 a_63_368.n0 246.553
R6 a_63_368.n1 a_63_368.t3 203
R7 a_63_368.n2 a_63_368.n1 152
R8 a_63_368.n0 a_63_368.t1 65.455
R9 a_63_368.n0 a_63_368.t2 38.1823
R10 VGND.n1 VGND.t1 251.845
R11 VGND.n1 VGND.n0 217.077
R12 VGND.n0 VGND.t2 48.0005
R13 VGND.n0 VGND.t0 35.7351
R14 VGND VGND.n1 0.311433
R15 VNB VNB.t1 1616.8
R16 VNB.t1 VNB.t2 1443.57
R17 VNB.t2 VNB.t0 1339.63
R18 a_152_368.t0 a_152_368.t1 63.3219
R19 VPWR.n4 VPWR.n3 641.586
R20 VPWR.n1 VPWR.n0 589.067
R21 VPWR.n2 VPWR.n0 586.653
R22 VPWR.n3 VPWR.n2 59.8041
R23 VPWR.n2 VPWR.t1 35.1791
R24 VPWR.n1 VPWR.t0 23.9385
R25 VPWR VPWR.n4 14.7079
R26 VPWR.n3 VPWR.n1 13.5656
R27 VPWR.n4 VPWR.n0 7.43276
R28 VPB.t2 VPB.t0 403.495
R29 VPB VPB.t1 349.866
R30 VPB.t1 VPB.t2 214.517
R31 B.n0 B.t0 216.632
R32 B.n0 B.t1 125.904
R33 B B.n0 105.308
R34 X.n1 X 589.508
R35 X.n1 X.n0 585
R36 X.n2 X.n1 585
R37 X X.t0 206.401
R38 X.n1 X.t1 26.3844
R39 X X.n2 12.0794
R40 X X.n0 10.4568
R41 X X.n0 2.88501
R42 X.n2 X 1.26247
C0 VPWR B 0.011359f
C1 VGND VPWR 0.041037f
C2 X B 2.15e-19
C3 X VGND 0.082342f
C4 X VPWR 0.100256f
C5 VPB A 0.042005f
C6 VPB B 0.052677f
C7 VPB VGND 0.008221f
C8 B A 0.065928f
C9 VGND A 0.012653f
C10 VPB VPWR 0.083418f
C11 VPB X 0.013593f
C12 VPWR A 0.01531f
C13 X A 0.001932f
C14 VGND B 0.057552f
C15 VGND VNB 0.374027f
C16 X VNB 0.111556f
C17 A VNB 0.122737f
C18 B VNB 0.192791f
C19 VPWR VNB 0.273255f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2_2 VNB VPB VPWR VGND X B A
X0 VPWR.t2 A.t0 a_114_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2127 pd=1.51 as=0.12 ps=1.24 w=1 l=0.15
X1 X.t1 a_27_368.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.2127 ps=1.51 w=1.12 l=0.15
X2 X.t3 a_27_368.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1276 ps=1.095 w=0.74 l=0.15
X3 VGND.t3 A.t1 a_27_368.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1276 pd=1.095 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 VGND.t0 a_27_368.t5 X.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2479 pd=2.15 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_114_368.t1 B.t0 a_27_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.285 ps=2.57 w=1 l=0.15
X6 a_27_368.t0 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1792 ps=1.84 w=0.64 l=0.15
X7 VPWR.t1 a_27_368.t6 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1792 ps=1.44 w=1.12 l=0.15
R0 A.n0 A.t0 231.629
R1 A.n0 A.t1 204.048
R2 A A.n0 153.892
R3 a_114_368.t0 a_114_368.t1 47.2805
R4 VPWR.n1 VPWR.t1 866.831
R5 VPWR.n1 VPWR.n0 611.698
R6 VPWR.n0 VPWR.t2 47.2805
R7 VPWR.n0 VPWR.t0 26.8503
R8 VPWR VPWR.n1 0.721008
R9 VPB.t2 VPB.t0 275.807
R10 VPB VPB.t3 252.823
R11 VPB.t0 VPB.t1 240.054
R12 VPB.t3 VPB.t2 199.195
R13 a_27_368.n4 a_27_368.n3 313.195
R14 a_27_368.t2 a_27_368.n4 293.562
R15 a_27_368.n3 a_27_368.t6 240.197
R16 a_27_368.n1 a_27_368.t3 240.197
R17 a_27_368.n4 a_27_368.n0 221.643
R18 a_27_368.n1 a_27_368.t4 179.947
R19 a_27_368.n2 a_27_368.t5 179.947
R20 a_27_368.n2 a_27_368.n1 62.8066
R21 a_27_368.n0 a_27_368.t1 26.2505
R22 a_27_368.n0 a_27_368.t0 26.2505
R23 a_27_368.n3 a_27_368.n2 5.84292
R24 X X.n0 586.601
R25 X.n2 X.n1 185
R26 X.n3 X.n2 185
R27 X.n0 X.t0 28.1434
R28 X.n0 X.t1 28.1434
R29 X.n2 X.t2 22.7032
R30 X.n2 X.t3 22.7032
R31 X.n3 X 17.3338
R32 X.n1 X 13.0672
R33 X.n1 X 6.66717
R34 X X.n3 2.4005
R35 VGND.n5 VGND.t2 243.638
R36 VGND.n3 VGND.n2 210.213
R37 VGND.n1 VGND.t0 163.69
R38 VGND.n2 VGND.t3 40.313
R39 VGND.n4 VGND.n3 24.4711
R40 VGND.n2 VGND.t1 21.3967
R41 VGND.n5 VGND.n4 21.0829
R42 VGND.n6 VGND.n5 9.3005
R43 VGND.n4 VGND.n0 9.3005
R44 VGND.n3 VGND.n1 6.57757
R45 VGND.n1 VGND.n0 0.660337
R46 VGND.n6 VGND.n0 0.122949
R47 VGND VGND.n6 0.0617245
R48 VNB.t3 VNB.t1 1166.4
R49 VNB VNB.t2 1131.76
R50 VNB.t1 VNB.t0 993.177
R51 VNB.t2 VNB.t3 993.177
R52 B.n0 B.t0 258.909
R53 B B.n0 158.788
R54 B.n0 B.t1 154.743
C0 A VPWR 0.017402f
C1 VGND VPWR 0.041304f
C2 VPB A 0.037211f
C3 VPB VGND 0.005702f
C4 VGND A 0.015903f
C5 VPWR X 0.014924f
C6 VPB X 0.002356f
C7 B VPWR 0.00965f
C8 VPB B 0.038664f
C9 A X 4.57e-19
C10 VGND X 0.133512f
C11 B A 0.094233f
C12 VPB VPWR 0.075246f
C13 B VGND 0.050201f
C14 VGND VNB 0.397173f
C15 X VNB 0.01237f
C16 VPWR VNB 0.278991f
C17 A VNB 0.114764f
C18 B VNB 0.165724f
C19 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2_4 VNB VPB VPWR VGND X B A
X0 X.t3 a_83_260.t4 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t5 B.t0 a_83_260.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.9287 pd=3.99 as=0.12395 ps=1.075 w=0.74 l=0.15
X2 X.t7 a_83_260.t5 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_83_260.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12395 pd=1.075 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 VPWR.t5 A.t1 a_493_388.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.64 as=0.175 ps=1.35 w=1 l=0.15
X5 VPWR.t1 a_83_260.t6 X.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t3 a_83_260.t7 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.13505 ps=1.105 w=0.74 l=0.15
X7 X.t1 a_83_260.t8 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t3 a_83_260.t9 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VGND.t2 a_83_260.t10 X.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_493_388.t3 B.t1 a_83_260.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X11 a_83_260.t3 B.t2 a_493_388.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X12 a_493_388.t0 A.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2102 ps=1.505 w=1 l=0.15
X13 X.t4 a_83_260.t11 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.13505 pd=1.105 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_83_260.n15 a_83_260.n14 848.005
R1 a_83_260.n1 a_83_260.t6 240.197
R2 a_83_260.n9 a_83_260.t8 240.197
R3 a_83_260.n2 a_83_260.t9 240.197
R4 a_83_260.n4 a_83_260.t4 240.197
R5 a_83_260.n1 a_83_260.t7 182.138
R6 a_83_260.n4 a_83_260.t5 181.407
R7 a_83_260.n3 a_83_260.t10 179.947
R8 a_83_260.n8 a_83_260.t11 179.947
R9 a_83_260.n6 a_83_260.n5 165.189
R10 a_83_260.n7 a_83_260.n6 152
R11 a_83_260.n10 a_83_260.n0 152
R12 a_83_260.n12 a_83_260.n11 152
R13 a_83_260.n14 a_83_260.n13 101.71
R14 a_83_260.n14 a_83_260.n12 50.8354
R15 a_83_260.n11 a_83_260.n10 49.6611
R16 a_83_260.n8 a_83_260.n7 37.246
R17 a_83_260.n5 a_83_260.n4 37.246
R18 a_83_260.n13 a_83_260.t1 31.6221
R19 a_83_260.t2 a_83_260.n15 29.5505
R20 a_83_260.n15 a_83_260.t3 29.5505
R21 a_83_260.n5 a_83_260.n3 24.1005
R22 a_83_260.n13 a_83_260.t0 22.7032
R23 a_83_260.n7 a_83_260.n2 21.1793
R24 a_83_260.n12 a_83_260.n0 13.1884
R25 a_83_260.n6 a_83_260.n0 13.1884
R26 a_83_260.n11 a_83_260.n1 10.955
R27 a_83_260.n9 a_83_260.n8 7.30353
R28 a_83_260.n10 a_83_260.n9 5.11262
R29 a_83_260.n3 a_83_260.n2 4.38232
R30 VPWR.n5 VPWR.t5 836.072
R31 VPWR.n11 VPWR.t2 351.637
R32 VPWR.n9 VPWR.n1 334.173
R33 VPWR.n4 VPWR.n3 325.5
R34 VPWR.n3 VPWR.t4 46.2955
R35 VPWR.n8 VPWR.n2 36.1417
R36 VPWR.n10 VPWR.n9 34.6358
R37 VPWR.n11 VPWR.n10 26.7299
R38 VPWR.n1 VPWR.t0 26.3844
R39 VPWR.n1 VPWR.t3 26.3844
R40 VPWR.n3 VPWR.t1 25.3542
R41 VPWR.n4 VPWR.n2 23.7181
R42 VPWR.n6 VPWR.n2 9.3005
R43 VPWR.n8 VPWR.n7 9.3005
R44 VPWR.n10 VPWR.n0 9.3005
R45 VPWR.n12 VPWR.n11 9.3005
R46 VPWR.n5 VPWR.n4 7.41279
R47 VPWR.n9 VPWR.n8 1.50638
R48 VPWR.n6 VPWR.n5 0.165146
R49 VPWR.n7 VPWR.n6 0.122949
R50 VPWR.n7 VPWR.n0 0.122949
R51 VPWR.n12 VPWR.n0 0.122949
R52 VPWR VPWR.n12 0.0617245
R53 X.n2 X.n0 250.518
R54 X.n2 X.n1 207.6
R55 X.n5 X.n3 146.538
R56 X.n5 X.n4 102.019
R57 X.n3 X.t6 33.2437
R58 X X.n2 32.7862
R59 X.n0 X.t2 26.3844
R60 X.n0 X.t1 26.3844
R61 X.n1 X.t0 26.3844
R62 X.n1 X.t3 26.3844
R63 X.n3 X.t4 25.9464
R64 X X.n5 23.489
R65 X.n4 X.t5 22.7032
R66 X.n4 X.t7 22.7032
R67 VPB.t2 VPB.t6 273.253
R68 VPB VPB.t3 257.93
R69 VPB.t4 VPB.t7 255.376
R70 VPB.t5 VPB.t4 229.839
R71 VPB.t6 VPB.t5 229.839
R72 VPB.t1 VPB.t2 229.839
R73 VPB.t0 VPB.t1 229.839
R74 VPB.t3 VPB.t0 229.839
R75 B.n1 B.t1 236.966
R76 B.n0 B.t0 228.148
R77 B.n0 B.t2 209.107
R78 B B.n1 154.133
R79 B.n1 B.n0 34.3247
R80 VGND.n10 VGND.t4 285.764
R81 VGND.n8 VGND.n2 214.185
R82 VGND.n4 VGND.n3 211.183
R83 VGND.n5 VGND.t5 118.507
R84 VGND.n8 VGND.n1 34.2593
R85 VGND.n3 VGND.t0 34.0546
R86 VGND.n10 VGND.n9 26.7299
R87 VGND.n3 VGND.t3 22.7032
R88 VGND.n2 VGND.t1 22.7032
R89 VGND.n2 VGND.t2 22.7032
R90 VGND.n9 VGND.n8 19.2005
R91 VGND.n4 VGND.n1 18.0711
R92 VGND.n11 VGND.n10 9.3005
R93 VGND.n6 VGND.n1 9.3005
R94 VGND.n8 VGND.n7 9.3005
R95 VGND.n9 VGND.n0 9.3005
R96 VGND.n5 VGND.n4 7.17842
R97 VGND.n6 VGND.n5 0.35955
R98 VGND.n7 VGND.n6 0.122949
R99 VGND.n7 VGND.n0 0.122949
R100 VGND.n11 VGND.n0 0.122949
R101 VGND VGND.n11 0.0617245
R102 VNB.t1 VNB.t3 1189.5
R103 VNB.t3 VNB.t0 1154.86
R104 VNB VNB.t4 1143.31
R105 VNB.t0 VNB.t5 1120.21
R106 VNB.t2 VNB.t1 993.177
R107 VNB.t4 VNB.t2 993.177
R108 A A.t1 481.851
R109 A.n0 A.t2 258.406
R110 A.n0 A.t0 220.113
R111 A A.n0 153.528
R112 a_493_388.n1 a_493_388.n0 942.571
R113 a_493_388.n1 a_493_388.t3 39.4005
R114 a_493_388.n0 a_493_388.t2 29.5505
R115 a_493_388.n0 a_493_388.t0 29.5505
R116 a_493_388.t1 a_493_388.n1 29.5505
C0 VPB A 0.096576f
C1 X VGND 0.279912f
C2 VPWR X 0.399379f
C3 VPWR VGND 0.074948f
C4 B VGND 0.022379f
C5 VPB X 0.015635f
C6 VPB VGND 0.0068f
C7 X A 0.016299f
C8 VPWR B 0.010778f
C9 A VGND 0.022355f
C10 VPB VPWR 0.125028f
C11 VPB B 0.069537f
C12 VPWR A 0.048587f
C13 A B 0.201503f
C14 VGND VNB 0.569986f
C15 B VNB 0.161217f
C16 A VNB 0.188338f
C17 X VNB 0.06869f
C18 VPWR VNB 0.471543f
C19 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2b_1 VNB VPB VPWR VGND X B_N A
X0 a_264_368.t1 a_27_112.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.174625 ps=1.185 w=0.55 l=0.15
X1 VGND.t3 B_N.t0 a_27_112.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.174625 pd=1.185 as=0.3685 ps=2.44 w=0.55 l=0.15
X2 X.t0 a_264_368.t3 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2382 ps=1.555 w=1.12 l=0.15
X3 X.t1 a_264_368.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.193225 ps=1.32 w=0.74 l=0.15
X4 VGND.t2 A.t0 a_264_368.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.193225 pd=1.32 as=0.077 ps=0.83 w=0.55 l=0.15
X5 VPWR.t1 B_N.t1 a_27_112.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2898 pd=2.37 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 VPWR.t2 A.t1 a_353_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.135 ps=1.27 w=1 l=0.15
X7 a_353_368.t0 a_27_112.t3 a_264_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
R0 a_27_112.t0 a_27_112.n1 438.252
R1 a_27_112.n0 a_27_112.t3 224.276
R2 a_27_112.n1 a_27_112.n0 220.404
R3 a_27_112.n1 a_27_112.t1 167.5
R4 a_27_112.n0 a_27_112.t2 149.421
R5 VGND.n2 VGND.n0 211.375
R6 VGND.n2 VGND.n1 102.374
R7 VGND.n1 VGND.t0 64.7156
R8 VGND.n0 VGND.t2 64.3641
R9 VGND.n1 VGND.t3 61.4429
R10 VGND.n0 VGND.t1 52.0988
R11 VGND VGND.n2 0.459094
R12 a_264_368.t0 a_264_368.n2 297.731
R13 a_264_368.n0 a_264_368.t3 264.298
R14 a_264_368.n2 a_264_368.n0 209.609
R15 a_264_368.n0 a_264_368.t4 204.048
R16 a_264_368.n2 a_264_368.n1 194.51
R17 a_264_368.n1 a_264_368.t2 30.546
R18 a_264_368.n1 a_264_368.t1 30.546
R19 VNB VNB.t3 2032.55
R20 VNB.t3 VNB.t0 1813.12
R21 VNB.t2 VNB.t1 1686.09
R22 VNB.t0 VNB.t2 993.177
R23 B_N.n0 B_N.t1 294.824
R24 B_N.n0 B_N.t0 235.888
R25 B_N B_N.n0 188
R26 VPWR.n1 VPWR.t1 402.017
R27 VPWR.n1 VPWR.n0 229.296
R28 VPWR.n0 VPWR.t2 46.2955
R29 VPWR.n0 VPWR.t0 35.2408
R30 VPWR VPWR.n1 0.224282
R31 X.n1 X 588.077
R32 X.n1 X.n0 585
R33 X.n2 X.n1 585
R34 X X.t1 203.812
R35 X.n1 X.t0 26.3844
R36 X X.n2 8.24665
R37 X X.n0 7.13896
R38 X X.n0 1.96973
R39 X.n2 X 0.862038
R40 VPB.t2 VPB.t0 605.242
R41 VPB.t3 VPB.t1 298.791
R42 VPB VPB.t2 257.93
R43 VPB.t0 VPB.t3 214.517
R44 A.n0 A.t1 230.581
R45 A.n0 A.t0 188.54
R46 A A.n0 155.721
R47 a_353_368.t0 a_353_368.t1 53.1905
C0 A VPB 0.037679f
C1 VGND VPWR 0.056031f
C2 X VGND 0.085557f
C3 VGND B_N 0.018013f
C4 X VPWR 0.14477f
C5 B_N VPWR 0.02274f
C6 A VGND 0.01161f
C7 VGND VPB 0.010357f
C8 A VPWR 0.033223f
C9 X B_N 2.03e-19
C10 VPB VPWR 0.118707f
C11 X VPB 0.023313f
C12 A X 0.006331f
C13 VPB B_N 0.084012f
C14 VGND VNB 0.462841f
C15 X VNB 0.114093f
C16 A VNB 0.111086f
C17 VPWR VNB 0.353682f
C18 B_N VNB 0.217773f
C19 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2b_2 VNB VPB VPWR VGND X B_N A
X0 VPWR.t0 B_N.t0 a_27_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VGND.t0 B_N.t1 a_27_368.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 VGND.t1 a_27_368.t2 a_187_48.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2336 pd=2.01 as=0.1104 ps=0.985 w=0.64 l=0.15
X3 VPWR.t2 a_187_48.t3 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.54 as=0.2884 ps=1.635 w=1.12 l=0.15
X4 VGND.t2 a_187_48.t4 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2349 pd=1.435 as=0.10545 ps=1.025 w=0.74 l=0.15
X5 a_187_48.t2 A.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1104 pd=0.985 as=0.2349 ps=1.435 w=0.64 l=0.15
X6 a_187_48.t1 a_27_368.t3 a_470_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.415 pd=2.83 as=0.135 ps=1.27 w=1 l=0.15
X7 a_470_368.t1 A.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2277 ps=1.54 w=1 l=0.15
X8 X.t2 a_187_48.t5 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2884 pd=1.635 as=0.203 ps=1.505 w=1.12 l=0.15
X9 X.t0 a_187_48.t6 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.126075 ps=1.1 w=0.74 l=0.15
R0 B_N.n0 B_N.t0 203.03
R1 B_N.n0 B_N.t1 186.696
R2 B_N B_N.n0 158.847
R3 a_27_368.t0 a_27_368.n1 343.495
R4 a_27_368.n1 a_27_368.n0 334.329
R5 a_27_368.n1 a_27_368.t1 310.337
R6 a_27_368.n0 a_27_368.t3 239.661
R7 a_27_368.n0 a_27_368.t2 226.541
R8 VPWR.n2 VPWR.n1 678.652
R9 VPWR.n2 VPWR.n0 613.028
R10 VPWR.n1 VPWR.t0 55.1136
R11 VPWR.n0 VPWR.t1 53.1905
R12 VPWR.n1 VPWR.t3 29.6087
R13 VPWR.n0 VPWR.t2 27.0196
R14 VPWR VPWR.n2 0.377872
R15 VPB.t4 VPB.t3 339.651
R16 VPB.t3 VPB.t2 291.13
R17 VPB.t0 VPB.t4 273.253
R18 VPB VPB.t0 257.93
R19 VPB.t2 VPB.t1 214.517
R20 VGND.n3 VGND.t1 242.995
R21 VGND.n10 VGND.n9 219.871
R22 VGND.n7 VGND.n6 185
R23 VGND.n5 VGND.n4 185
R24 VGND.n6 VGND.n5 76.8755
R25 VGND.n9 VGND.t0 47.6797
R26 VGND.n8 VGND.n7 28.5366
R27 VGND.n5 VGND.t3 27.188
R28 VGND.n10 VGND.n8 24.0946
R29 VGND.n6 VGND.t2 22.6611
R30 VGND.n9 VGND.t4 21.551
R31 VGND.n2 VGND.n1 9.3005
R32 VGND.n8 VGND.n0 9.3005
R33 VGND.n4 VGND.n3 8.33638
R34 VGND.n11 VGND.n10 7.47871
R35 VGND.n4 VGND.n1 5.57815
R36 VGND.n3 VGND.n2 0.576964
R37 VGND.n7 VGND.n1 0.286534
R38 VGND VGND.n11 0.16068
R39 VGND.n11 VGND.n0 0.14713
R40 VGND.n2 VGND.n0 0.122949
R41 VNB.t2 VNB.t3 1951.71
R42 VNB.t0 VNB.t4 1177.95
R43 VNB VNB.t0 1154.86
R44 VNB.t3 VNB.t1 1143.31
R45 VNB.t4 VNB.t2 1004.72
R46 a_187_48.t1 a_187_48.n4 344.377
R47 a_187_48.n2 a_187_48.t3 251.151
R48 a_187_48.n0 a_187_48.t5 240.197
R49 a_187_48.n4 a_187_48.n2 222.024
R50 a_187_48.n0 a_187_48.t6 185.041
R51 a_187_48.n1 a_187_48.t4 179.947
R52 a_187_48.n4 a_187_48.n3 103.532
R53 a_187_48.n1 a_187_48.n0 59.155
R54 a_187_48.n3 a_187_48.t2 38.438
R55 a_187_48.n2 a_187_48.n1 27.0217
R56 a_187_48.n3 a_187_48.t0 26.2505
R57 X.n1 X.n0 654.874
R58 X.n2 X.n1 185
R59 X.n3 X.n2 185
R60 X.n0 X.t3 45.7326
R61 X.n0 X.t2 44.8532
R62 X.n2 X.t1 23.514
R63 X.n2 X.t0 22.7032
R64 X.n3 X 12.6066
R65 X.n1 X 4.84898
R66 X X.n3 1.74595
R67 A.n0 A.t0 236.18
R68 A.n0 A.t1 231.629
R69 A A.n0 155.721
R70 a_470_368.t0 a_470_368.t1 53.1905
C0 X A 0.005732f
C1 VPWR X 0.026287f
C2 VPB A 0.036825f
C3 VPB VPWR 0.105045f
C4 VPB X 0.004962f
C5 B_N VGND 0.012215f
C6 A VGND 0.018405f
C7 VPWR VGND 0.056718f
C8 VPWR B_N 0.009234f
C9 X VGND 0.122384f
C10 VPWR A 0.014052f
C11 VPB VGND 0.007942f
C12 B_N X 0.001169f
C13 VPB B_N 0.04437f
C14 VGND VNB 0.462616f
C15 A VNB 0.117533f
C16 X VNB 0.006483f
C17 B_N VNB 0.162031f
C18 VPWR VNB 0.357943f
C19 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2b_4 VNB VPB VPWR VGND A B_N X
X0 a_81_296.t3 a_676_48.t2 a_489_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.29 ps=2.58 w=1 l=0.15
X1 VGND.t7 a_81_296.t6 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.11285 ps=1.045 w=0.74 l=0.15
X2 VPWR.t4 a_81_296.t7 X.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2046 pd=1.495 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X.t3 a_81_296.t8 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_81_296.t5 a_676_48.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
X5 VPWR.t2 a_81_296.t9 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 X.t6 a_81_296.t10 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 a_81_296.t1 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.144 pd=1.09 as=0.1165 ps=1.065 w=0.64 l=0.15
X8 a_676_48.t0 B_N.t0 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.29 ps=2.58 w=1 l=0.15
X9 X.t5 a_81_296.t11 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 VGND.t0 A.t1 a_81_296.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.144 ps=1.09 w=0.64 l=0.15
X11 X.t1 a_81_296.t12 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X12 a_676_48.t1 B_N.t1 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.6272 pd=3.24 as=0.112 ps=0.99 w=0.64 l=0.15
X13 VGND.t4 a_81_296.t13 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t6 A.t2 a_489_392.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.15 ps=1.3 w=1 l=0.15
X15 a_489_392.t0 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2046 ps=1.495 w=1 l=0.15
X16 VGND.t2 a_676_48.t4 a_81_296.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X17 a_489_392.t1 a_676_48.t5 a_81_296.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.15 ps=1.3 w=1 l=0.15
R0 a_676_48.n2 a_676_48.t3 358.288
R1 a_676_48.t0 a_676_48.n8 298.514
R2 a_676_48.n2 a_676_48.t2 255.728
R3 a_676_48.n3 a_676_48.t4 242.607
R4 a_676_48.n5 a_676_48.n4 221.724
R5 a_676_48.n4 a_676_48.t5 207.529
R6 a_676_48.n5 a_676_48.n1 185
R7 a_676_48.n8 a_676_48.n7 185
R8 a_676_48.n4 a_676_48.n3 106.332
R9 a_676_48.n7 a_676_48.n6 90.6969
R10 a_676_48.n1 a_676_48.n0 90.6713
R11 a_676_48.n3 a_676_48.n2 22.4938
R12 a_676_48.n7 a_676_48.t1 21.4291
R13 a_676_48.n1 a_676_48.t1 20.2046
R14 a_676_48.n6 a_676_48.n0 7.26921
R15 a_676_48.n8 a_676_48.n0 3.66048
R16 a_676_48.n6 a_676_48.n5 3.60923
R17 a_489_392.n0 a_489_392.t1 316.296
R18 a_489_392.n1 a_489_392.n0 275.491
R19 a_489_392.n0 a_489_392.t2 216.737
R20 a_489_392.n1 a_489_392.t3 29.5505
R21 a_489_392.t0 a_489_392.n1 29.5505
R22 a_81_296.n15 a_81_296.n14 352.99
R23 a_81_296.n2 a_81_296.t12 260.281
R24 a_81_296.n2 a_81_296.t10 257.87
R25 a_81_296.n1 a_81_296.t7 240.197
R26 a_81_296.n6 a_81_296.t8 240.197
R27 a_81_296.n4 a_81_296.t9 240.197
R28 a_81_296.n1 a_81_296.t6 185.06
R29 a_81_296.n3 a_81_296.t13 179.947
R30 a_81_296.n7 a_81_296.t11 179.947
R31 a_81_296.n5 a_81_296.n0 165.189
R32 a_81_296.n8 a_81_296.n0 152
R33 a_81_296.n10 a_81_296.n9 152
R34 a_81_296.n14 a_81_296.n13 113.671
R35 a_81_296.n12 a_81_296.n11 108.576
R36 a_81_296.n3 a_81_296.n2 96.1084
R37 a_81_296.n14 a_81_296.n12 52.7064
R38 a_81_296.n9 a_81_296.n8 49.6611
R39 a_81_296.n11 a_81_296.t0 45.0005
R40 a_81_296.n12 a_81_296.n10 43.2262
R41 a_81_296.n6 a_81_296.n5 41.6278
R42 a_81_296.n11 a_81_296.t1 39.3755
R43 a_81_296.n15 a_81_296.t2 29.5505
R44 a_81_296.t3 a_81_296.n15 29.5505
R45 a_81_296.n13 a_81_296.t4 26.2505
R46 a_81_296.n13 a_81_296.t5 26.2505
R47 a_81_296.n5 a_81_296.n4 24.1005
R48 a_81_296.n10 a_81_296.n0 13.1884
R49 a_81_296.n9 a_81_296.n1 8.03383
R50 a_81_296.n7 a_81_296.n6 4.38232
R51 a_81_296.n8 a_81_296.n7 3.65202
R52 a_81_296.n4 a_81_296.n3 2.92171
R53 VPB.t1 VPB.t7 510.753
R54 VPB.t8 VPB.t2 508.2
R55 VPB.t6 VPB.t0 268.146
R56 VPB VPB.t3 252.823
R57 VPB.t2 VPB.t1 229.839
R58 VPB.t0 VPB.t8 229.839
R59 VPB.t5 VPB.t6 229.839
R60 VPB.t4 VPB.t5 229.839
R61 VPB.t3 VPB.t4 229.839
R62 X.n5 X.n3 256.541
R63 X.n5 X.n4 215.559
R64 X.n2 X.n0 150.971
R65 X.n2 X.n1 102.019
R66 X.n6 X.n5 36.4748
R67 X X.n6 28.1048
R68 X.n0 X.t7 26.7573
R69 X.n4 X.t2 26.3844
R70 X.n4 X.t1 26.3844
R71 X.n3 X.t0 26.3844
R72 X.n3 X.t3 26.3844
R73 X.n1 X.t4 22.7032
R74 X.n1 X.t6 22.7032
R75 X.n0 X.t5 22.7032
R76 X.n6 X.n2 7.13511
R77 VGND.n14 VGND.n2 208.274
R78 VGND.n16 VGND.t6 145.216
R79 VGND.n5 VGND.n4 121.325
R80 VGND.n7 VGND.n6 115.659
R81 VGND.n10 VGND.n9 115.659
R82 VGND.n4 VGND.t8 39.3755
R83 VGND.n6 VGND.t3 39.3755
R84 VGND.n2 VGND.t5 34.0546
R85 VGND.n9 VGND.t7 31.0986
R86 VGND.n14 VGND.n1 28.2358
R87 VGND.n8 VGND.n7 27.4829
R88 VGND.n16 VGND.n15 26.7299
R89 VGND.n4 VGND.t2 26.2505
R90 VGND.n6 VGND.t0 26.2505
R91 VGND.n9 VGND.t1 26.2505
R92 VGND.n10 VGND.n8 25.224
R93 VGND.n2 VGND.t4 22.7032
R94 VGND.n10 VGND.n1 22.2123
R95 VGND.n15 VGND.n14 19.2005
R96 VGND.n17 VGND.n16 9.3005
R97 VGND.n8 VGND.n3 9.3005
R98 VGND.n11 VGND.n10 9.3005
R99 VGND.n12 VGND.n1 9.3005
R100 VGND.n14 VGND.n13 9.3005
R101 VGND.n15 VGND.n0 9.3005
R102 VGND.n7 VGND.n5 6.49816
R103 VGND.n5 VGND.n3 0.56347
R104 VGND.n11 VGND.n3 0.122949
R105 VGND.n12 VGND.n11 0.122949
R106 VGND.n13 VGND.n12 0.122949
R107 VGND.n13 VGND.n0 0.122949
R108 VGND.n17 VGND.n0 0.122949
R109 VGND VGND.n17 0.0617245
R110 VNB.t1 VNB.t0 1385.83
R111 VNB.t2 VNB.t8 1154.86
R112 VNB.t0 VNB.t3 1154.86
R113 VNB.t4 VNB.t5 1154.86
R114 VNB VNB.t6 1143.31
R115 VNB.t7 VNB.t1 1097.11
R116 VNB.t5 VNB.t7 1050.92
R117 VNB.t3 VNB.t2 993.177
R118 VNB.t6 VNB.t4 993.177
R119 VPWR.n6 VPWR.t6 352.957
R120 VPWR.n12 VPWR.n2 325.255
R121 VPWR.n5 VPWR.t5 258.104
R122 VPWR.n14 VPWR.t1 250.081
R123 VPWR.n4 VPWR.n3 231.184
R124 VPWR.n3 VPWR.t0 44.3255
R125 VPWR.n12 VPWR.n11 32.0005
R126 VPWR.n7 VPWR.n4 30.4946
R127 VPWR.n3 VPWR.t4 27.2574
R128 VPWR.n2 VPWR.t3 26.3844
R129 VPWR.n2 VPWR.t2 26.3844
R130 VPWR.n7 VPWR.n6 24.0946
R131 VPWR.n11 VPWR.n4 22.9652
R132 VPWR.n13 VPWR.n12 21.4593
R133 VPWR.n14 VPWR.n13 21.4593
R134 VPWR.n8 VPWR.n7 9.3005
R135 VPWR.n9 VPWR.n4 9.3005
R136 VPWR.n11 VPWR.n10 9.3005
R137 VPWR.n12 VPWR.n1 9.3005
R138 VPWR.n13 VPWR.n0 9.3005
R139 VPWR.n15 VPWR.n14 9.3005
R140 VPWR.n6 VPWR.n5 7.39937
R141 VPWR.n8 VPWR.n5 0.163603
R142 VPWR.n9 VPWR.n8 0.122949
R143 VPWR.n10 VPWR.n9 0.122949
R144 VPWR.n10 VPWR.n1 0.122949
R145 VPWR.n1 VPWR.n0 0.122949
R146 VPWR.n15 VPWR.n0 0.122949
R147 VPWR VPWR.n15 0.0617245
R148 A.n0 A.t3 283.844
R149 A.n0 A.t0 261.084
R150 A.n1 A.t1 251.956
R151 A.n2 A.t2 236.983
R152 A.n3 A.n2 152
R153 A.n1 A.n0 77.1205
R154 A.n2 A.n1 14.6066
R155 A.n3 A 12.0247
R156 A A.n3 6.59444
R157 B_N.n1 B_N.t1 308.365
R158 B_N.n0 B_N.t0 231.454
R159 B_N B_N.n0 153.745
R160 B_N.n2 B_N.n1 152
R161 B_N.n1 B_N.n0 39.0195
R162 B_N B_N.n2 11.4429
R163 B_N.n2 B_N 2.90959
C0 VGND B_N 0.022108f
C1 VPWR VPB 0.184859f
C2 VGND X 0.310919f
C3 VPWR B_N 0.05462f
C4 VPB A 0.095844f
C5 B_N A 3.49e-19
C6 VGND VPWR 0.095701f
C7 VPWR X 0.423334f
C8 VGND A 0.037614f
C9 X A 0.005808f
C10 B_N VPB 0.064217f
C11 VGND VPB 0.012539f
C12 VPWR A 0.038462f
C13 X VPB 0.01479f
C14 VGND VNB 0.717158f
C15 B_N VNB 0.226033f
C16 X VNB 0.051768f
C17 VPWR VNB 0.585585f
C18 A VNB 0.232525f
C19 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2111ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2111ai_4 VNB VPB VPWR VGND Y B1 A1 A2 C1 D1
X0 a_954_368.t2 A1.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_472_74.t5 B1.t0 a_841_74.t11 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t2 A1.t1 a_954_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_954_368.t6 A2.t0 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X4 a_954_368.t0 A1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1764 ps=1.435 w=1.12 l=0.15
X5 Y.t4 B1.t1 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6 a_472_74.t0 C1.t0 a_27_74.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VGND.t3 A1.t3 a_841_74.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 Y.t10 D1.t0 a_27_74.t7 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_472_74.t4 B1.t2 a_841_74.t10 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_841_74.t0 A2.t1 VGND.t7 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 Y.t7 A2.t2 a_954_368.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X12 a_472_74.t1 C1.t1 a_27_74.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 Y.t6 A2.t3 a_954_368.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.1764 ps=1.435 w=1.12 l=0.15
X14 Y.t1 D1.t1 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_841_74.t9 B1.t3 a_472_74.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VPWR.t8 D1.t2 Y.t13 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=1.176 ps=4.34 w=1.12 l=0.15
X17 a_27_74.t3 C1.t2 a_472_74.t6 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VGND.t6 A2.t4 a_841_74.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_27_74.t0 D1.t3 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_954_368.t3 A2.t5 Y.t5 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1876 ps=1.455 w=1.12 l=0.15
X21 VGND.t2 A1.t4 a_841_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_841_74.t6 A2.t6 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 VPWR.t0 B1.t4 Y.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_841_74.t8 B1.t5 a_472_74.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 a_27_74.t6 D1.t4 Y.t9 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X26 Y.t11 C1.t3 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4032 ps=1.84 w=1.12 l=0.15
X27 a_841_74.t2 A1.t5 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VPWR.t7 C1.t4 Y.t12 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.4032 pd=1.84 as=0.168 ps=1.42 w=1.12 l=0.15
X29 a_27_74.t2 C1.t5 a_472_74.t7 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 Y.t2 D1.t5 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X31 a_841_74.t1 A1.t6 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X32 VGND.t4 A2.t7 a_841_74.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1332 ps=1.1 w=0.74 l=0.15
R0 A1.n6 A1.n5 239.528
R1 A1.n0 A1.t0 226.809
R2 A1.n3 A1.t1 226.809
R3 A1.n4 A1.t2 226.809
R4 A1.n0 A1.t5 202.655
R5 A1.n6 A1.t3 186.374
R6 A1.n11 A1.t6 186.374
R7 A1.n2 A1.t4 186.374
R8 A1 A1.n1 155.423
R9 A1.n13 A1.n12 152
R10 A1.n10 A1.n9 152
R11 A1.n8 A1.n7 152
R12 A1.n12 A1.n11 36.8199
R13 A1.n7 A1.n4 36.8199
R14 A1.n2 A1.n1 24.7699
R15 A1.n1 A1.n0 20.7533
R16 A1.n3 A1.n2 14.7283
R17 A1.n7 A1.n6 12.7199
R18 A1.n9 A1.n8 10.1214
R19 A1.n11 A1.n10 8.70328
R20 A1.n10 A1.n4 8.70328
R21 A1.n13 A1 7.5912
R22 A1 A1.n13 6.69817
R23 A1.n12 A1.n3 6.0255
R24 A1.n9 A1 2.53073
R25 A1.n8 A1 1.63771
R26 VPWR.n9 VPWR.t1 865.167
R27 VPWR.n8 VPWR.n7 626.366
R28 VPWR.n17 VPWR.n16 315.928
R29 VPWR.n25 VPWR.n1 315.926
R30 VPWR.n23 VPWR.n3 142.464
R31 VPWR.n3 VPWR.t7 59.182
R32 VPWR.n3 VPWR.t6 59.1816
R33 VPWR.n22 VPWR.n4 36.1417
R34 VPWR.n10 VPWR.n6 36.1417
R35 VPWR.n14 VPWR.n6 36.1417
R36 VPWR.n15 VPWR.n14 36.1417
R37 VPWR.n18 VPWR.n15 36.1417
R38 VPWR.n1 VPWR.t4 35.1791
R39 VPWR.n1 VPWR.t8 35.1791
R40 VPWR.n16 VPWR.t5 35.1791
R41 VPWR.n16 VPWR.t0 35.1791
R42 VPWR.n25 VPWR.n24 34.6358
R43 VPWR.n7 VPWR.t3 26.3844
R44 VPWR.n7 VPWR.t2 26.3844
R45 VPWR.n10 VPWR.n9 25.224
R46 VPWR.n24 VPWR.n23 15.8123
R47 VPWR.n11 VPWR.n10 9.3005
R48 VPWR.n12 VPWR.n6 9.3005
R49 VPWR.n14 VPWR.n13 9.3005
R50 VPWR.n15 VPWR.n5 9.3005
R51 VPWR.n19 VPWR.n18 9.3005
R52 VPWR.n20 VPWR.n4 9.3005
R53 VPWR.n22 VPWR.n21 9.3005
R54 VPWR.n23 VPWR.n2 9.3005
R55 VPWR.n24 VPWR.n0 9.3005
R56 VPWR.n23 VPWR.n22 7.52991
R57 VPWR.n9 VPWR.n8 6.98058
R58 VPWR.n17 VPWR.n4 6.77697
R59 VPWR.n26 VPWR.n25 6.36235
R60 VPWR.n18 VPWR.n17 4.51815
R61 VPWR.n11 VPWR.n8 0.536037
R62 VPWR VPWR.n26 0.384136
R63 VPWR.n26 VPWR.n0 0.169491
R64 VPWR.n12 VPWR.n11 0.122949
R65 VPWR.n13 VPWR.n12 0.122949
R66 VPWR.n13 VPWR.n5 0.122949
R67 VPWR.n19 VPWR.n5 0.122949
R68 VPWR.n20 VPWR.n19 0.122949
R69 VPWR.n21 VPWR.n20 0.122949
R70 VPWR.n21 VPWR.n2 0.122949
R71 VPWR.n2 VPWR.n0 0.122949
R72 a_954_368.n3 a_954_368.n0 351.974
R73 a_954_368.n2 a_954_368.n1 302.74
R74 a_954_368.n2 a_954_368.t6 294.469
R75 a_954_368.n4 a_954_368.n3 289.051
R76 a_954_368.n3 a_954_368.n2 64.1354
R77 a_954_368.n1 a_954_368.t3 35.1791
R78 a_954_368.n4 a_954_368.t5 29.0228
R79 a_954_368.n0 a_954_368.t1 26.3844
R80 a_954_368.n0 a_954_368.t0 26.3844
R81 a_954_368.n1 a_954_368.t4 26.3844
R82 a_954_368.t2 a_954_368.n4 26.3844
R83 VPB.t9 VPB.t1 1325.4
R84 VPB VPB.t12 643.548
R85 VPB.t11 VPB.t10 444.356
R86 VPB.t0 VPB.t9 280.914
R87 VPB.t12 VPB.t5 280.914
R88 VPB.t6 VPB.t8 255.376
R89 VPB.t4 VPB.t6 255.376
R90 VPB.t7 VPB.t4 247.715
R91 VPB.t3 VPB.t7 237.5
R92 VPB.t2 VPB.t3 229.839
R93 VPB.t1 VPB.t2 229.839
R94 VPB.t10 VPB.t0 229.839
R95 VPB.t5 VPB.t11 229.839
R96 B1.n1 B1.t4 376.567
R97 B1.n9 B1.t3 219.149
R98 B1.n1 B1.t1 204.048
R99 B1.n0 B1.t5 196.013
R100 B1.n2 B1.t0 196.013
R101 B1.n8 B1.t2 196.013
R102 B1.n10 B1.n9 152
R103 B1.n7 B1.n6 152
R104 B1.n5 B1.n0 152
R105 B1.n4 B1.n3 152
R106 B1.n2 B1.n1 119.233
R107 B1.n7 B1.n0 43.7018
R108 B1.n3 B1.n0 43.7018
R109 B1.n9 B1.n8 32.1338
R110 B1.n8 B1.n7 11.5685
R111 B1.n3 B1.n2 11.5685
R112 B1.n6 B1.n5 10.1214
R113 B1 B1.n4 8.93073
R114 B1 B1.n10 7.14469
R115 B1.n10 B1 7.14469
R116 B1.n4 B1 5.35864
R117 B1.n6 B1 2.97724
R118 B1.n5 B1 1.1912
R119 a_841_74.n3 a_841_74.t11 310.755
R120 a_841_74.n8 a_841_74.t6 204.012
R121 a_841_74.n3 a_841_74.n2 185
R122 a_841_74.n7 a_841_74.n6 104.579
R123 a_841_74.n9 a_841_74.n8 104.579
R124 a_841_74.n5 a_841_74.n0 103.65
R125 a_841_74.n4 a_841_74.n1 95.6388
R126 a_841_74.n5 a_841_74.n4 64.0005
R127 a_841_74.n7 a_841_74.n5 58.3534
R128 a_841_74.n8 a_841_74.n7 51.2005
R129 a_841_74.n4 a_841_74.n3 36.0732
R130 a_841_74.n9 a_841_74.t7 35.6762
R131 a_841_74.n1 a_841_74.t9 34.0546
R132 a_841_74.n2 a_841_74.t10 22.7032
R133 a_841_74.n2 a_841_74.t8 22.7032
R134 a_841_74.n1 a_841_74.t4 22.7032
R135 a_841_74.n0 a_841_74.t3 22.7032
R136 a_841_74.n0 a_841_74.t1 22.7032
R137 a_841_74.n6 a_841_74.t5 22.7032
R138 a_841_74.n6 a_841_74.t2 22.7032
R139 a_841_74.t0 a_841_74.n9 22.7032
R140 a_472_74.n3 a_472_74.n1 222.315
R141 a_472_74.n4 a_472_74.n0 221.556
R142 a_472_74.n3 a_472_74.n2 185
R143 a_472_74.n5 a_472_74.n4 185
R144 a_472_74.n4 a_472_74.n3 61.6141
R145 a_472_74.n1 a_472_74.t6 22.7032
R146 a_472_74.n1 a_472_74.t1 22.7032
R147 a_472_74.n2 a_472_74.t7 22.7032
R148 a_472_74.n2 a_472_74.t0 22.7032
R149 a_472_74.n0 a_472_74.t3 22.7032
R150 a_472_74.n0 a_472_74.t4 22.7032
R151 a_472_74.n5 a_472_74.t2 22.7032
R152 a_472_74.t5 a_472_74.n5 22.7032
R153 VNB.t19 VNB.t15 2286.61
R154 VNB.t0 VNB.t9 1177.95
R155 VNB.t7 VNB.t0 1154.86
R156 VNB.t6 VNB.t3 1154.86
R157 VNB.t13 VNB.t6 1154.86
R158 VNB.t18 VNB.t17 1154.86
R159 VNB VNB.t18 1143.31
R160 VNB.t9 VNB.t8 993.177
R161 VNB.t4 VNB.t7 993.177
R162 VNB.t5 VNB.t4 993.177
R163 VNB.t3 VNB.t5 993.177
R164 VNB.t14 VNB.t13 993.177
R165 VNB.t12 VNB.t14 993.177
R166 VNB.t15 VNB.t12 993.177
R167 VNB.t10 VNB.t19 993.177
R168 VNB.t16 VNB.t10 993.177
R169 VNB.t11 VNB.t16 993.177
R170 VNB.t1 VNB.t11 993.177
R171 VNB.t2 VNB.t1 993.177
R172 VNB.t17 VNB.t2 993.177
R173 A2.n6 A2.t3 232.635
R174 A2.n5 A2.t5 226.809
R175 A2.n0 A2.t0 204.048
R176 A2.n3 A2.t2 204.048
R177 A2.n0 A2.t6 156.739
R178 A2 A2.n1 155.87
R179 A2.n6 A2.t4 155.847
R180 A2.n4 A2.t1 155.847
R181 A2.n2 A2.t7 155.847
R182 A2.n12 A2.n11 152
R183 A2.n10 A2.n9 152
R184 A2.n8 A2.n7 152
R185 A2.n11 A2.n10 34.6841
R186 A2.n7 A2.n6 25.4247
R187 A2.n2 A2.n1 22.3153
R188 A2.n7 A2.n5 20.128
R189 A2.n1 A2.n0 15.1746
R190 A2.n9 A2.n8 10.1214
R191 A2.n10 A2.n4 8.47523
R192 A2.n12 A2 8.03771
R193 A2.n5 A2.n4 7.41588
R194 A2.n3 A2.n2 7.14124
R195 A2 A2.n12 6.25166
R196 A2.n9 A2 2.08422
R197 A2.n8 A2 2.08422
R198 A2.n11 A2.n3 0.893093
R199 Y.n2 Y.n0 350.397
R200 Y.n2 Y.n1 299.95
R201 Y.n3 Y.n2 275.954
R202 Y.n3 Y.t4 231.87
R203 Y.n11 Y.n9 215.578
R204 Y.n5 Y.n4 202.457
R205 Y.n7 Y.n6 202.457
R206 Y.n11 Y.n10 185
R207 Y.n7 Y.t13 174.227
R208 Y.n8 Y.n5 79.685
R209 Y.n5 Y.n3 51.1192
R210 Y.n0 Y.t7 35.1791
R211 Y.n9 Y.t10 34.0546
R212 Y.n1 Y.t6 32.5407
R213 Y.n6 Y.t12 26.3844
R214 Y.n6 Y.t2 26.3844
R215 Y.n4 Y.t3 26.3844
R216 Y.n4 Y.t11 26.3844
R217 Y.n0 Y.t8 26.3844
R218 Y.n1 Y.t5 26.3844
R219 Y Y.n11 25.6005
R220 Y.n9 Y.t9 22.7032
R221 Y.n10 Y.t0 22.7032
R222 Y.n10 Y.t1 22.7032
R223 Y Y.n8 17.6845
R224 Y.n8 Y.n7 5.14381
R225 C1.n2 C1.t5 263.762
R226 C1.n0 C1.t4 216.012
R227 C1.n3 C1.t3 214.758
R228 C1.n6 C1.n5 152
R229 C1.n4 C1.t2 142.994
R230 C1.n0 C1.t1 142.994
R231 C1.n2 C1.t0 142.994
R232 C1.n6 C1.n1 85.4362
R233 C1 C1.n6 36.4611
R234 C1.n5 C1.n4 30.3486
R235 C1.n1 C1.n0 22.4592
R236 C1.n4 C1.n1 13.2742
R237 C1.n5 C1.n3 6.69494
R238 C1.n3 C1.n2 1.33939
R239 a_27_74.n4 a_27_74.t2 308.368
R240 a_27_74.n1 a_27_74.n0 185
R241 a_27_74.n5 a_27_74.n4 185
R242 a_27_74.n1 a_27_74.t7 184.821
R243 a_27_74.n3 a_27_74.n2 88.6236
R244 a_27_74.n3 a_27_74.n1 51.7878
R245 a_27_74.n4 a_27_74.n3 42.7019
R246 a_27_74.n0 a_27_74.t1 22.7032
R247 a_27_74.n0 a_27_74.t6 22.7032
R248 a_27_74.n2 a_27_74.t4 22.7032
R249 a_27_74.n2 a_27_74.t0 22.7032
R250 a_27_74.t5 a_27_74.n5 22.7032
R251 a_27_74.n5 a_27_74.t3 22.7032
R252 VGND.n6 VGND.n3 216.046
R253 VGND.n5 VGND.n4 210.406
R254 VGND.n9 VGND.n2 210.406
R255 VGND.n12 VGND.n11 210.406
R256 VGND.n4 VGND.t6 34.0546
R257 VGND.n11 VGND.t3 34.0546
R258 VGND.n10 VGND.n9 28.2358
R259 VGND.n5 VGND.n1 25.977
R260 VGND.n3 VGND.t5 22.7032
R261 VGND.n3 VGND.t4 22.7032
R262 VGND.n4 VGND.t7 22.7032
R263 VGND.n2 VGND.t1 22.7032
R264 VGND.n2 VGND.t2 22.7032
R265 VGND.n11 VGND.t0 22.7032
R266 VGND.n9 VGND.n1 19.2005
R267 VGND.n12 VGND.n10 11.6711
R268 VGND.n7 VGND.n1 9.3005
R269 VGND.n9 VGND.n8 9.3005
R270 VGND.n10 VGND.n0 9.3005
R271 VGND.n13 VGND.n12 7.6387
R272 VGND.n6 VGND.n5 6.59375
R273 VGND VGND.n13 1.63461
R274 VGND.n7 VGND.n6 0.559358
R275 VGND.n13 VGND.n0 0.149657
R276 VGND.n8 VGND.n7 0.122949
R277 VGND.n8 VGND.n0 0.122949
R278 D1.n0 D1.t5 233.502
R279 D1.n2 D1.t2 226.809
R280 D1 D1.n3 154.084
R281 D1.n8 D1.n7 152
R282 D1.n6 D1.n5 152
R283 D1.n0 D1.t3 148.037
R284 D1.n6 D1.t0 143.968
R285 D1.n1 D1.t1 142.994
R286 D1.n4 D1.t4 142.994
R287 D1.n1 D1.n0 39.4835
R288 D1.n7 D1.n6 33.1076
R289 D1.n4 D1.n3 18.5015
R290 D1.n2 D1.n1 16.4556
R291 D1.n7 D1.n4 14.6066
R292 D1.n5 D1 10.4191
R293 D1 D1.n8 8.03771
R294 D1.n3 D1.n2 7.30353
R295 D1.n8 D1 6.25166
R296 D1.n5 D1 3.87027
C0 VGND VPWR 0.158121f
C1 VGND B1 0.027532f
C2 A2 Y 0.201441f
C3 A2 C1 6.9e-20
C4 VPB Y 0.051068f
C5 VPB C1 0.098244f
C6 VPWR A1 0.056137f
C7 B1 A1 0.085768f
C8 VPB D1 0.120141f
C9 VGND Y 0.032816f
C10 VGND C1 0.026806f
C11 D1 VGND 0.027079f
C12 VPB A2 0.147768f
C13 Y A1 0.142866f
C14 VPWR B1 0.038231f
C15 C1 A1 1.42e-19
C16 VGND A2 0.075321f
C17 VPB VGND 0.012228f
C18 Y VPWR 0.81774f
C19 VPWR C1 0.047297f
C20 Y B1 0.191731f
C21 A2 A1 0.09985f
C22 C1 B1 0.097635f
C23 D1 VPWR 0.039897f
C24 VPB A1 0.142523f
C25 VGND A1 0.069209f
C26 A2 VPWR 0.026913f
C27 Y C1 0.230299f
C28 D1 Y 0.319349f
C29 VPB VPWR 0.246046f
C30 D1 C1 0.055932f
C31 VPB B1 0.16897f
C32 VGND VNB 1.11927f
C33 VPWR VNB 0.894287f
C34 Y VNB 0.05895f
C35 A2 VNB 0.451805f
C36 A1 VNB 0.397513f
C37 B1 VNB 0.424111f
C38 C1 VNB 0.35869f
C39 D1 VNB 0.400701f
C40 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3b_1 VNB VPB VPWR VGND A B C_N X
X0 a_452_391.t1 B.t0 a_368_391.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_368_391.t0 a_124_424.t2 a_239_74.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X2 VGND.t0 A.t0 a_239_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.190125 pd=1.345 as=0.086625 ps=0.865 w=0.55 l=0.15
X3 a_124_424.t1 C_N.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1595 pd=1.68 as=0.1925 ps=1.8 w=0.55 l=0.15
X4 VGND.t4 a_124_424.t3 a_239_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.15675 ps=1.67 w=0.55 l=0.15
X5 X.t1 a_239_74.t4 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2382 ps=1.555 w=1.12 l=0.15
X6 a_239_74.t1 B.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.086625 pd=0.865 as=0.1155 ps=0.97 w=0.55 l=0.15
X7 VPWR.t0 A.t1 a_452_391.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.135 ps=1.27 w=1 l=0.15
X8 X.t0 a_239_74.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.190125 ps=1.345 w=0.74 l=0.15
X9 a_124_424.t0 C_N.t1 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2562 pd=2.29 as=0.2814 ps=2.35 w=0.84 l=0.15
R0 B.n0 B.t0 305.267
R1 B.n0 B.t1 199.227
R2 B B.n0 160
R3 a_368_391.t0 a_368_391.t1 53.1905
R4 a_452_391.t0 a_452_391.t1 53.1905
R5 VPB.t1 VPB.t3 623.119
R6 VPB.t2 VPB.t0 298.791
R7 VPB VPB.t1 278.361
R8 VPB.t4 VPB.t2 214.517
R9 VPB.t3 VPB.t4 214.517
R10 a_124_424.t0 a_124_424.n3 414.45
R11 a_124_424.n2 a_124_424.t2 377.86
R12 a_124_424.n1 a_124_424.t3 307.166
R13 a_124_424.n0 a_124_424.t1 253.321
R14 a_124_424.n3 a_124_424.n2 152
R15 a_124_424.n1 a_124_424.n0 152
R16 a_124_424.n2 a_124_424.n1 49.6611
R17 a_124_424.n3 a_124_424.n0 10.1214
R18 a_239_74.t3 a_239_74.n3 273.928
R19 a_239_74.n0 a_239_74.t4 263.938
R20 a_239_74.n3 a_239_74.t2 238.556
R21 a_239_74.n2 a_239_74.n0 229.913
R22 a_239_74.n0 a_239_74.t5 203.688
R23 a_239_74.n2 a_239_74.n1 185
R24 a_239_74.n3 a_239_74.n2 50.9645
R25 a_239_74.n1 a_239_74.t0 38.1823
R26 a_239_74.n1 a_239_74.t1 30.546
R27 A.n0 A.t1 275.812
R28 A.n0 A.t0 234.573
R29 A A.n0 155.333
R30 VGND.n8 VGND.t2 254.745
R31 VGND.n2 VGND.n1 204.976
R32 VGND.n4 VGND.n3 191.118
R33 VGND.n3 VGND.t1 63.2753
R34 VGND.n3 VGND.t0 62.1823
R35 VGND.n1 VGND.t3 45.8187
R36 VGND.n1 VGND.t4 45.8187
R37 VGND.n7 VGND.n6 36.1417
R38 VGND.n6 VGND.n2 35.7652
R39 VGND.n8 VGND.n7 20.7064
R40 VGND.n9 VGND.n8 9.3005
R41 VGND.n6 VGND.n5 9.3005
R42 VGND.n7 VGND.n0 9.3005
R43 VGND.n4 VGND.n2 6.0321
R44 VGND.n5 VGND.n4 0.380851
R45 VGND.n5 VGND.n0 0.122949
R46 VGND.n9 VGND.n0 0.122949
R47 VGND VGND.n9 0.0617245
R48 VNB.t2 VNB.t4 2298.16
R49 VNB.t0 VNB.t1 1743.83
R50 VNB.t4 VNB.t3 1316.54
R51 VNB VNB.t2 1293.44
R52 VNB.t3 VNB.t0 1074.02
R53 C_N.n0 C_N.t1 252.113
R54 C_N.n1 C_N.t0 171.512
R55 C_N C_N.n0 152.934
R56 C_N.n2 C_N.n1 152
R57 C_N.n1 C_N.n0 45.5227
R58 C_N C_N.n2 8.13383
R59 C_N.n2 C_N 1.73383
R60 VPWR.n1 VPWR.t2 405.568
R61 VPWR.n1 VPWR.n0 229.379
R62 VPWR.n0 VPWR.t0 46.2955
R63 VPWR.n0 VPWR.t1 32.6283
R64 VPWR VPWR.n1 0.0997027
R65 X.n0 X.t1 289.135
R66 X.t0 X.n0 279.738
R67 X.n1 X.t0 279.738
R68 X.n1 X 11.5561
R69 X.n0 X 4.44494
R70 X X.n1 1.6005
C0 A VGND 0.014637f
C1 VPB VGND 0.010523f
C2 B A 0.116865f
C3 VPB B 0.041982f
C4 VPWR X 0.14283f
C5 C_N VPWR 0.045245f
C6 B VGND 0.013733f
C7 C_N X 8.35e-20
C8 VPWR A 0.033109f
C9 VPB VPWR 0.124734f
C10 VPWR VGND 0.062738f
C11 A X 0.006566f
C12 VPB X 0.023102f
C13 VPWR B 0.078334f
C14 VPB C_N 0.069638f
C15 X VGND 0.070951f
C16 C_N VGND 0.052499f
C17 B X 0.003677f
C18 VPB A 0.043097f
C19 C_N B 2.1e-19
C20 VGND VNB 0.520012f
C21 X VNB 0.11236f
C22 A VNB 0.127334f
C23 B VNB 0.129335f
C24 VPWR VNB 0.429874f
C25 C_N VNB 0.203943f
C26 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4_2 VNB VPB VPWR VGND X D A B C
X0 a_258_392.t0 C.t0 a_174_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t3 a_85_392.t5 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2382 ps=1.555 w=1.12 l=0.15
X2 a_174_392.t1 D.t0 a_85_392.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X3 VGND.t5 A.t0 a_85_392.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1805 pd=1.265 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 X.t1 a_85_392.t6 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1805 ps=1.265 w=0.74 l=0.15
X5 VPWR.t2 A.t1 a_342_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.215 ps=1.43 w=1 l=0.15
X6 a_85_392.t2 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1943 ps=1.255 w=0.64 l=0.15
X7 a_85_392.t4 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.284075 ps=2.19 w=0.64 l=0.15
X8 VGND.t1 C.t1 a_85_392.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1943 pd=1.255 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 a_342_392.t1 B.t1 a_258_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t3 a_85_392.t7 X.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t1 a_85_392.t8 X.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
R0 C.n0 C.t0 312.591
R1 C.n0 C.t1 176.025
R2 C C.n0 161.697
R3 a_174_392.t0 a_174_392.t1 53.1905
R4 a_258_392.t0 a_258_392.t1 53.1905
R5 VPB VPB.t5 406.048
R6 VPB.t3 VPB.t2 298.791
R7 VPB.t4 VPB.t3 296.238
R8 VPB.t2 VPB.t1 229.839
R9 VPB.t0 VPB.t4 214.517
R10 VPB.t5 VPB.t0 214.517
R11 a_85_392.t3 a_85_392.n6 363.14
R12 a_85_392.n2 a_85_392.t5 251.151
R13 a_85_392.n0 a_85_392.t8 240.197
R14 a_85_392.n4 a_85_392.n2 213.764
R15 a_85_392.n0 a_85_392.t7 198.127
R16 a_85_392.n1 a_85_392.t6 179.947
R17 a_85_392.n6 a_85_392.n5 97.8183
R18 a_85_392.n4 a_85_392.n3 97.5208
R19 a_85_392.n6 a_85_392.n4 63.2476
R20 a_85_392.n1 a_85_392.n0 48.9308
R21 a_85_392.n3 a_85_392.t0 26.2505
R22 a_85_392.n3 a_85_392.t2 26.2505
R23 a_85_392.n5 a_85_392.t1 26.2505
R24 a_85_392.n5 a_85_392.t4 26.2505
R25 a_85_392.n2 a_85_392.n1 5.84292
R26 VPWR.n1 VPWR.t1 359.94
R27 VPWR.n1 VPWR.n0 227.627
R28 VPWR.n0 VPWR.t2 46.2955
R29 VPWR.n0 VPWR.t0 35.2408
R30 VPWR VPWR.n1 0.996835
R31 X X.n0 246.786
R32 X X.n1 131.531
R33 X.n0 X.t2 26.3844
R34 X.n0 X.t3 26.3844
R35 X.n1 X.t0 22.7032
R36 X.n1 X.t1 22.7032
R37 D.n0 D.t1 265.101
R38 D.n0 D.t0 228.186
R39 D D.n0 164.333
R40 A.n0 A.t1 263.762
R41 A.n0 A.t0 236.18
R42 A A.n0 158.4
R43 VGND.n10 VGND.t0 248.691
R44 VGND.n4 VGND.t3 237.993
R45 VGND.n3 VGND.n2 203.98
R46 VGND.n8 VGND.n7 198.067
R47 VGND.n7 VGND.t2 55.313
R48 VGND.n7 VGND.t1 55.313
R49 VGND.n2 VGND.t5 50.6255
R50 VGND.n2 VGND.t4 44.2236
R51 VGND.n8 VGND.n1 36.1417
R52 VGND.n9 VGND.n8 36.1417
R53 VGND.n10 VGND.n9 15.8123
R54 VGND.n3 VGND.n1 15.0593
R55 VGND.n11 VGND.n10 9.3005
R56 VGND.n9 VGND.n0 9.3005
R57 VGND.n5 VGND.n1 9.3005
R58 VGND.n4 VGND.n3 6.6595
R59 VGND.n8 VGND.n6 4.62059
R60 VGND.n5 VGND.n4 0.655456
R61 VGND.n6 VGND.n5 0.184273
R62 VGND.n6 VGND.n0 0.184273
R63 VGND.n11 VGND.n0 0.122949
R64 VGND VGND.n11 0.0617245
R65 VNB.t1 VNB.t2 1709.19
R66 VNB.t5 VNB.t4 1559.06
R67 VNB VNB.t0 1478.22
R68 VNB.t4 VNB.t3 993.177
R69 VNB.t2 VNB.t5 993.177
R70 VNB.t0 VNB.t1 993.177
R71 a_342_392.t0 a_342_392.t1 84.7105
R72 B.n0 B.t1 263.053
R73 B.n0 B.t0 235.471
R74 B B.n0 154.522
C0 A VGND 0.015482f
C1 VGND C 0.015588f
C2 VPB VGND 0.00925f
C3 A X 0.005728f
C4 VPWR B 0.074855f
C5 VPB X 0.0123f
C6 VGND D 0.014574f
C7 A VPWR 0.035358f
C8 A B 0.109525f
C9 VPWR C 0.033557f
C10 VPB VPWR 0.115033f
C11 C B 0.177884f
C12 VPB B 0.044964f
C13 X VGND 0.143959f
C14 A C 4.07e-19
C15 VPWR D 0.011538f
C16 VPB A 0.048149f
C17 VPB C 0.039806f
C18 VPWR VGND 0.064311f
C19 VGND B 0.014809f
C20 D C 0.129525f
C21 VPB D 0.056407f
C22 VPWR X 0.232757f
C23 X B 0.003691f
C24 VGND VNB 0.516053f
C25 X VNB 0.063636f
C26 VPWR VNB 0.420299f
C27 A VNB 0.116436f
C28 B VNB 0.11257f
C29 C VNB 0.120271f
C30 D VNB 0.156052f
C31 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4_1 VNB VPB VPWR VGND D C A X B
X0 VPWR.t1 A.t0 a_331_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2859 pd=1.66 as=0.21 ps=1.42 w=1 l=0.15
X1 VGND.t3 C.t0 a_44_392.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1674 pd=1.165 as=0.077 ps=0.83 w=0.55 l=0.15
X2 VGND.t4 A.t1 a_44_392.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.121 ps=0.99 w=0.55 l=0.15
X3 X.t0 a_44_392.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.126075 ps=1.1 w=0.74 l=0.15
X4 a_44_392.t1 D.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.19525 ps=1.81 w=0.55 l=0.15
X5 a_44_392.t0 B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.121 pd=0.99 as=0.1674 ps=1.165 w=0.55 l=0.15
X6 X.t1 a_44_392.t6 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2859 ps=1.66 w=1.12 l=0.15
X7 a_217_392.t1 C.t1 a_133_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X8 a_133_392.t1 D.t1 a_44_392.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X9 a_331_392.t0 B.t1 a_217_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
R0 A.n0 A.t0 263.401
R1 A.n0 A.t1 189.227
R2 A A.n0 156.465
R3 a_331_392.t0 a_331_392.t1 82.7405
R4 VPWR VPWR.n0 316.538
R5 VPWR.n0 VPWR.t0 74.8307
R6 VPWR.n0 VPWR.t1 29.5505
R7 VPB.t4 VPB.t2 352.42
R8 VPB VPB.t3 301.344
R9 VPB.t1 VPB.t4 291.13
R10 VPB.t0 VPB.t1 291.13
R11 VPB.t3 VPB.t0 214.517
R12 C.n0 C.t1 245.018
R13 C.n0 C.t0 212.081
R14 C C.n0 153.067
R15 a_44_392.t2 a_44_392.n4 424.01
R16 a_44_392.n2 a_44_392.n0 267.279
R17 a_44_392.n3 a_44_392.t6 264.298
R18 a_44_392.n3 a_44_392.t5 204.048
R19 a_44_392.n2 a_44_392.n1 185
R20 a_44_392.n4 a_44_392.n3 152
R21 a_44_392.n4 a_44_392.n2 52.2266
R22 a_44_392.n1 a_44_392.t4 48.0005
R23 a_44_392.n1 a_44_392.t0 48.0005
R24 a_44_392.n0 a_44_392.t3 30.546
R25 a_44_392.n0 a_44_392.t1 30.546
R26 VGND.n6 VGND.t2 247.934
R27 VGND.n2 VGND.n1 217.5
R28 VGND.n4 VGND.n3 203.19
R29 VGND.n3 VGND.t0 64.3641
R30 VGND.n3 VGND.t3 63.2732
R31 VGND.n1 VGND.t4 47.6797
R32 VGND.n5 VGND.n4 30.4946
R33 VGND.n1 VGND.t1 21.551
R34 VGND.n6 VGND.n5 20.7064
R35 VGND.n7 VGND.n6 9.3005
R36 VGND.n5 VGND.n0 9.3005
R37 VGND.n4 VGND.n2 5.37113
R38 VGND.n2 VGND.n0 0.309716
R39 VGND.n7 VGND.n0 0.122949
R40 VGND VGND.n7 0.0617245
R41 VNB.t3 VNB.t0 1697.64
R42 VNB.t0 VNB.t4 1362.73
R43 VNB VNB.t2 1304.99
R44 VNB.t4 VNB.t1 1177.95
R45 VNB.t2 VNB.t3 993.177
R46 X.n1 X 589.268
R47 X.n1 X.n0 585
R48 X.n2 X.n1 585
R49 X X.t0 207.392
R50 X.n1 X.t1 26.3844
R51 X X.n2 11.4352
R52 X X.n0 9.89917
R53 X X.n0 2.73117
R54 X.n2 X 1.19517
R55 D.n0 D.t1 248.304
R56 D.n0 D.t0 212.081
R57 D D.n0 163.733
R58 B.n0 B.t1 245.018
R59 B.n0 B.t0 212.081
R60 B B.n0 154.133
R61 a_133_392.t0 a_133_392.t1 53.1905
R62 a_217_392.t0 a_217_392.t1 82.7405
C0 A VPWR 0.017693f
C1 X A 0.001508f
C2 VGND B 0.012157f
C3 C A 1.33e-19
C4 D VPWR 0.011748f
C5 VGND VPB 0.008588f
C6 X D 7.21e-20
C7 D C 0.08773f
C8 B VPWR 0.012462f
C9 X B 2.21e-19
C10 VPB VPWR 0.089281f
C11 C B 0.075304f
C12 D A 7.46e-20
C13 X VPB 0.014573f
C14 VPB C 0.04105f
C15 B A 0.079089f
C16 VPB A 0.046703f
C17 VGND VPWR 0.055333f
C18 VPB D 0.048809f
C19 X VGND 0.077359f
C20 VGND C 0.013273f
C21 VPB B 0.042882f
C22 X VPWR 0.085688f
C23 VGND A 0.012935f
C24 C VPWR 0.01204f
C25 VGND D 0.039887f
C26 X C 1.16e-19
C27 VGND VNB 0.49439f
C28 X VNB 0.115371f
C29 VPWR VNB 0.352831f
C30 A VNB 0.113427f
C31 B VNB 0.108384f
C32 C VNB 0.106904f
C33 D VNB 0.153141f
C34 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3b_4 VNB VPB VPWR VGND A B C_N X
X0 VGND.t7 A.t0 a_409_392.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 X.t3 a_409_392.t5 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2 VGND.t3 a_409_392.t6 X.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 X.t7 a_409_392.t7 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t0 C_N.t0 a_27_392.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.66075 pd=3.58 as=0.1824 ps=1.85 w=0.64 l=0.15
X5 VGND.t6 a_409_392.t8 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.11285 ps=1.045 w=0.74 l=0.15
X6 a_217_392.t1 B.t0 a_307_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X7 a_307_392.t3 a_27_392.t2 a_409_392.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1625 ps=1.325 w=1 l=0.15
X8 VPWR.t3 a_409_392.t9 X.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VPWR.t2 a_409_392.t10 X.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VPWR.t6 A.t1 a_217_392.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1959 pd=1.48 as=0.18 ps=1.36 w=1 l=0.15
X11 X.t4 a_409_392.t11 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1959 ps=1.48 w=1.12 l=0.15
X12 a_409_392.t3 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 a_307_392.t0 B.t2 a_217_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X14 a_217_392.t2 A.t2 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.18 ps=1.36 w=1 l=0.15
X15 a_409_392.t1 a_27_392.t3 a_307_392.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.18 ps=1.36 w=1 l=0.15
X16 VGND.t1 a_27_392.t4 a_409_392.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2072 ps=2.04 w=0.74 l=0.15
X17 X.t0 a_409_392.t12 VGND.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1332 ps=1.1 w=0.74 l=0.15
X18 VPWR.t0 C_N.t1 a_27_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.29 ps=2.58 w=1 l=0.15
R0 A A.t2 551.149
R1 A.n0 A.t1 298.572
R2 A.n0 A.t0 178.34
R3 A A.n0 171.194
R4 a_409_392.n15 a_409_392.n14 727.615
R5 a_409_392.n5 a_409_392.t10 240.197
R6 a_409_392.n4 a_409_392.t7 240.197
R7 a_409_392.n0 a_409_392.t9 240.197
R8 a_409_392.n11 a_409_392.t11 240.197
R9 a_409_392.n2 a_409_392.t2 187.185
R10 a_409_392.n11 a_409_392.t12 182.138
R11 a_409_392.n5 a_409_392.t6 179.947
R12 a_409_392.n0 a_409_392.t8 179.947
R13 a_409_392.n6 a_409_392.t5 179.947
R14 a_409_392.n8 a_409_392.n7 165.189
R15 a_409_392.n13 a_409_392.n12 152
R16 a_409_392.n10 a_409_392.n3 152
R17 a_409_392.n9 a_409_392.n8 152
R18 a_409_392.n2 a_409_392.n1 97.1225
R19 a_409_392.n14 a_409_392.n2 58.7299
R20 a_409_392.n12 a_409_392.n10 49.6611
R21 a_409_392.n0 a_409_392.n9 44.549
R22 a_409_392.n7 a_409_392.n5 37.246
R23 a_409_392.t0 a_409_392.n15 32.5055
R24 a_409_392.n15 a_409_392.t1 31.5205
R25 a_409_392.n7 a_409_392.n6 25.5611
R26 a_409_392.n1 a_409_392.t4 22.7032
R27 a_409_392.n1 a_409_392.t3 22.7032
R28 a_409_392.n9 a_409_392.n4 21.1793
R29 a_409_392.n8 a_409_392.n3 13.1884
R30 a_409_392.n13 a_409_392.n3 13.1884
R31 a_409_392.n12 a_409_392.n11 10.955
R32 a_409_392.n14 a_409_392.n13 7.3702
R33 a_409_392.n10 a_409_392.n0 5.11262
R34 a_409_392.n6 a_409_392.n4 2.92171
R35 VGND.n17 VGND.t0 365.646
R36 VGND.n6 VGND.t3 238.641
R37 VGND.n5 VGND.n4 215.464
R38 VGND.n2 VGND.n1 205.752
R39 VGND.n10 VGND.n9 204.388
R40 VGND.n16 VGND.n15 36.1417
R41 VGND.n9 VGND.t7 34.8654
R42 VGND.n1 VGND.t1 34.0546
R43 VGND.n15 VGND.n2 31.624
R44 VGND.n4 VGND.t4 30.8113
R45 VGND.n11 VGND.n10 29.3652
R46 VGND.n8 VGND.n5 24.4711
R47 VGND.n9 VGND.t5 23.514
R48 VGND.n4 VGND.t6 22.7032
R49 VGND.n1 VGND.t2 22.7032
R50 VGND.n17 VGND.n16 20.3299
R51 VGND.n10 VGND.n8 17.3181
R52 VGND.n11 VGND.n2 15.8123
R53 VGND.n16 VGND.n0 9.3005
R54 VGND.n15 VGND.n14 9.3005
R55 VGND.n13 VGND.n2 9.3005
R56 VGND.n12 VGND.n11 9.3005
R57 VGND.n10 VGND.n3 9.3005
R58 VGND.n8 VGND.n7 9.3005
R59 VGND.n6 VGND.n5 6.92167
R60 VGND.n18 VGND.n17 6.72455
R61 VGND.n7 VGND.n6 0.602654
R62 VGND VGND.n18 0.268037
R63 VGND.n18 VGND.n0 0.162655
R64 VGND.n7 VGND.n3 0.122949
R65 VGND.n12 VGND.n3 0.122949
R66 VGND.n13 VGND.n12 0.122949
R67 VGND.n14 VGND.n13 0.122949
R68 VGND.n14 VGND.n0 0.122949
R69 VNB.t0 VNB.t1 4492.39
R70 VNB VNB.t0 1189.5
R71 VNB.t7 VNB.t3 1177.95
R72 VNB.t1 VNB.t2 1154.86
R73 VNB.t4 VNB.t6 1108.66
R74 VNB.t3 VNB.t4 1050.92
R75 VNB.t6 VNB.t5 993.177
R76 VNB.t2 VNB.t7 993.177
R77 X.n2 X.n0 268.01
R78 X.n2 X.n1 207.6
R79 X.n5 X.n3 156.275
R80 X.n5 X.n4 102.019
R81 X X.n2 32.0332
R82 X X.n5 29.5125
R83 X.n3 X.t0 26.7573
R84 X.n0 X.t6 26.3844
R85 X.n0 X.t4 26.3844
R86 X.n1 X.t5 26.3844
R87 X.n1 X.t7 26.3844
R88 X.n3 X.t1 22.7032
R89 X.n4 X.t2 22.7032
R90 X.n4 X.t3 22.7032
R91 VPWR.n8 VPWR.t2 358.748
R92 VPWR.n7 VPWR.n6 325.255
R93 VPWR.n11 VPWR.n5 315.738
R94 VPWR.n19 VPWR.n1 222.463
R95 VPWR.n1 VPWR.t5 41.3705
R96 VPWR.n5 VPWR.t6 37.4305
R97 VPWR.n13 VPWR.n12 36.1417
R98 VPWR.n13 VPWR.n2 36.1417
R99 VPWR.n17 VPWR.n2 36.1417
R100 VPWR.n18 VPWR.n17 36.1417
R101 VPWR.n5 VPWR.t1 31.4907
R102 VPWR.n1 VPWR.t0 29.5505
R103 VPWR.n12 VPWR.n11 28.9887
R104 VPWR.n6 VPWR.t4 26.3844
R105 VPWR.n6 VPWR.t3 26.3844
R106 VPWR.n10 VPWR.n7 25.977
R107 VPWR.n19 VPWR.n18 23.3417
R108 VPWR.n11 VPWR.n10 18.4476
R109 VPWR.n10 VPWR.n9 9.3005
R110 VPWR.n11 VPWR.n4 9.3005
R111 VPWR.n12 VPWR.n3 9.3005
R112 VPWR.n14 VPWR.n13 9.3005
R113 VPWR.n15 VPWR.n2 9.3005
R114 VPWR.n17 VPWR.n16 9.3005
R115 VPWR.n18 VPWR.n0 9.3005
R116 VPWR.n20 VPWR.n19 7.25439
R117 VPWR.n8 VPWR.n7 6.92649
R118 VPWR.n9 VPWR.n8 0.547078
R119 VPWR VPWR.n20 0.157727
R120 VPWR.n20 VPWR.n0 0.150046
R121 VPWR.n9 VPWR.n4 0.122949
R122 VPWR.n4 VPWR.n3 0.122949
R123 VPWR.n14 VPWR.n3 0.122949
R124 VPWR.n15 VPWR.n14 0.122949
R125 VPWR.n16 VPWR.n15 0.122949
R126 VPWR.n16 VPWR.n0 0.122949
R127 VPB.t10 VPB.t5 260.485
R128 VPB.t4 VPB.t10 260.485
R129 VPB.t1 VPB.t3 260.485
R130 VPB.t0 VPB.t9 260.485
R131 VPB VPB.t0 255.376
R132 VPB.t3 VPB.t2 242.608
R133 VPB.t8 VPB.t6 229.839
R134 VPB.t7 VPB.t8 229.839
R135 VPB.t5 VPB.t7 229.839
R136 VPB.t2 VPB.t4 229.839
R137 VPB.t9 VPB.t1 229.839
R138 C_N.t0 C_N.t1 442.904
R139 C_N C_N.t0 233.162
R140 a_27_392.n0 a_27_392.t2 352.128
R141 a_27_392.n1 a_27_392.t3 352.128
R142 a_27_392.n2 a_27_392.n1 283.839
R143 a_27_392.t0 a_27_392.n2 283.089
R144 a_27_392.n2 a_27_392.t1 211.25
R145 a_27_392.n0 a_27_392.t4 163.077
R146 a_27_392.n1 a_27_392.n0 94.7938
R147 B B.t2 387.344
R148 B.n0 B.t1 258.673
R149 B.n0 B.t0 231.629
R150 B B.n0 170.177
R151 B.n1 B 20.7365
R152 B B.n1 3.8405
R153 B.n1 B 3.09727
R154 a_307_392.n1 a_307_392.n0 1212.29
R155 a_307_392.n1 a_307_392.t0 41.3705
R156 a_307_392.n0 a_307_392.t1 29.5505
R157 a_307_392.n0 a_307_392.t3 29.5505
R158 a_307_392.t2 a_307_392.n1 29.5505
R159 a_217_392.n1 a_217_392.n0 616.073
R160 a_217_392.t1 a_217_392.n1 39.4005
R161 a_217_392.n1 a_217_392.t3 31.5205
R162 a_217_392.n0 a_217_392.t0 29.5505
R163 a_217_392.n0 a_217_392.t2 29.5505
C0 B X 3.16e-19
C1 VPWR VGND 0.096562f
C2 VPWR A 0.054106f
C3 A VGND 0.039385f
C4 B VPWR 0.020325f
C5 B A 0.269547f
C6 VPWR C_N 0.025654f
C7 B VGND 0.018963f
C8 X VPB 0.014054f
C9 C_N A 0.04571f
C10 C_N VGND 0.123125f
C11 VPWR VPB 0.159428f
C12 B C_N 1.28e-19
C13 VPB VGND 0.009791f
C14 VPB A 0.082676f
C15 VPWR X 0.37059f
C16 B VPB 0.085763f
C17 X VGND 0.256217f
C18 X A 0.002265f
C19 VPB C_N 0.039839f
C20 VGND VNB 0.707296f
C21 X VNB 0.074764f
C22 VPWR VNB 0.574796f
C23 B VNB 0.158651f
C24 A VNB 0.18833f
C25 C_N VNB 0.230448f
C26 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3b_2 VNB VPB VPWR VGND X A B C_N
X0 VPWR.t3 C_N.t0 a_27_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 a_190_260.t0 a_27_368.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1344 ps=1.06 w=0.64 l=0.15
X2 X.t3 a_190_260.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.126075 ps=1.1 w=0.74 l=0.15
X3 a_542_368.t1 B.t0 a_458_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X4 a_190_260.t1 a_27_368.t3 a_542_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.195 ps=1.39 w=1 l=0.15
X5 VGND.t4 C_N.t1 a_27_368.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X6 VGND.t3 B.t1 a_190_260.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.112 ps=0.99 w=0.64 l=0.15
X7 a_458_368.t0 A.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.318575 ps=1.705 w=1 l=0.15
X8 VGND.t2 a_190_260.t5 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1965 pd=1.315 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t0 a_190_260.t6 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.318575 pd=1.705 as=0.168 ps=1.42 w=1.12 l=0.15
X10 X.t0 a_190_260.t7 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.203 ps=1.505 w=1.12 l=0.15
X11 a_190_260.t3 A.t1 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1965 ps=1.315 w=0.64 l=0.15
R0 C_N.n0 C_N.t0 217.538
R1 C_N.n0 C_N.t1 170.583
R2 C_N C_N.n0 155.067
R3 a_27_368.n1 a_27_368.n0 363.966
R4 a_27_368.t0 a_27_368.n1 327.127
R5 a_27_368.n1 a_27_368.t1 295.211
R6 a_27_368.n0 a_27_368.t3 226.15
R7 a_27_368.n0 a_27_368.t2 204.048
R8 VPWR.n2 VPWR.n1 678.558
R9 VPWR.n2 VPWR.n0 604.751
R10 VPWR.n0 VPWR.t2 57.1305
R11 VPWR.n1 VPWR.t3 55.1136
R12 VPWR.n0 VPWR.t0 46.2544
R13 VPWR.n1 VPWR.t1 29.6087
R14 VPWR VPWR.n2 0.464004
R15 VPB.t1 VPB.t4 370.296
R16 VPB.t3 VPB.t0 275.807
R17 VPB.t5 VPB.t2 273.253
R18 VPB VPB.t5 257.93
R19 VPB.t2 VPB.t1 229.839
R20 VPB.t4 VPB.t3 214.517
R21 VGND.n1 VGND.n0 221.828
R22 VGND.n3 VGND.n2 215.784
R23 VGND.n5 VGND.n4 201.315
R24 VGND.n4 VGND.t2 56.4111
R25 VGND.n4 VGND.t5 47.813
R26 VGND.n0 VGND.t4 47.6797
R27 VGND.n2 VGND.t0 39.3755
R28 VGND.n2 VGND.t3 39.3755
R29 VGND.n6 VGND.n5 32.0005
R30 VGND.n6 VGND.n1 25.6005
R31 VGND.n0 VGND.t1 21.551
R32 VGND.n8 VGND.n1 18.245
R33 VGND.n7 VGND.n6 9.3005
R34 VGND.n5 VGND.n3 4.47495
R35 VGND.n7 VGND.n3 0.385337
R36 VGND VGND.n8 0.163644
R37 VGND.n8 VGND.n7 0.144205
R38 a_190_260.t1 a_190_260.n5 412.485
R39 a_190_260.n0 a_190_260.t7 299.644
R40 a_190_260.n2 a_190_260.t6 263.938
R41 a_190_260.n4 a_190_260.n2 214.639
R42 a_190_260.n1 a_190_260.t5 190.738
R43 a_190_260.n0 a_190_260.t4 179.947
R44 a_190_260.n5 a_190_260.t0 136.16
R45 a_190_260.n1 a_190_260.n0 104.433
R46 a_190_260.n4 a_190_260.n3 100.817
R47 a_190_260.n5 a_190_260.n4 50.4476
R48 a_190_260.n3 a_190_260.t3 39.3755
R49 a_190_260.n3 a_190_260.t2 26.2505
R50 a_190_260.n2 a_190_260.n1 12.9498
R51 VNB.t1 VNB.t5 1674.54
R52 VNB.t3 VNB.t0 1316.54
R53 VNB VNB.t4 1304.99
R54 VNB.t4 VNB.t2 1177.95
R55 VNB.t5 VNB.t3 1154.86
R56 VNB.t2 VNB.t1 993.177
R57 X.n3 X.n2 585
R58 X.n1 X.n0 154.03
R59 X.n2 X.t1 26.3844
R60 X.n2 X.t0 26.3844
R61 X.n0 X.t2 22.7032
R62 X.n0 X.t3 22.7032
R63 X X.n3 12.8005
R64 X.n3 X.n1 4.46111
R65 X.n1 X 1.35808
R66 B.n0 B.t0 231.629
R67 B.n0 B.t1 204.048
R68 B B.n0 155.721
R69 a_458_368.t0 a_458_368.t1 53.1905
R70 a_542_368.t0 a_542_368.t1 76.8305
R71 A.n0 A.t0 231.629
R72 A.n0 A.t1 204.048
R73 A A.n0 154.522
C0 VPB VPWR 0.116041f
C1 VPWR C_N 0.008618f
C2 VPWR A 0.016889f
C3 X VGND 0.117216f
C4 B VGND 0.01262f
C5 VPB VGND 0.0087f
C6 C_N VGND 0.009547f
C7 A VGND 0.014355f
C8 VPB X 0.004914f
C9 VPB B 0.033021f
C10 C_N X 7.22e-19
C11 VPWR VGND 0.064479f
C12 X A 0.032847f
C13 A B 0.092454f
C14 VPB C_N 0.050327f
C15 VPB A 0.039223f
C16 VPWR X 0.022558f
C17 C_N A 2.11e-19
C18 VPWR B 0.006581f
C19 VGND VNB 0.511682f
C20 B VNB 0.104229f
C21 A VNB 0.109332f
C22 X VNB 0.009566f
C23 C_N VNB 0.180283f
C24 VPWR VNB 0.397188f
C25 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4b_1 VNB VPB VPWR VGND D_N A B C X
X0 a_440_368.t1 C.t0 a_356_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t1 A.t0 a_524_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2907 pd=1.66 as=0.195 ps=1.39 w=1 l=0.15
X2 VGND.t5 A.t1 a_228_74.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.159875 pd=1.235 as=0.077 ps=0.83 w=0.55 l=0.15
X3 VGND.t1 D_N.t0 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.15675 ps=1.67 w=0.55 l=0.15
X4 a_356_368.t0 a_27_74.t2 a_228_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5 X.t0 a_228_74.t5 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2907 ps=1.66 w=1.12 l=0.15
X6 a_228_74.t2 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.1155 ps=0.97 w=0.55 l=0.15
X7 X.t1 a_228_74.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.159875 ps=1.235 w=0.74 l=0.15
X8 VPWR.t0 D_N.t1 a_27_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2898 pd=2.37 as=0.2478 ps=2.27 w=0.84 l=0.15
X9 a_228_74.t1 a_27_74.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.254375 pd=1.475 as=0.1155 ps=0.97 w=0.55 l=0.15
X10 VGND.t4 C.t1 a_228_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.254375 ps=1.475 w=0.55 l=0.15
X11 a_524_368.t0 B.t1 a_440_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
R0 C.n0 C.t0 313.3
R1 C.n0 C.t1 152.633
R2 C C.n0 152
R3 a_356_368.t0 a_356_368.t1 53.1905
R4 a_440_368.t0 a_440_368.t1 53.1905
R5 VPB.t2 VPB.t0 610.35
R6 VPB.t5 VPB.t4 352.42
R7 VPB.t1 VPB.t5 275.807
R8 VPB VPB.t2 260.485
R9 VPB.t3 VPB.t1 214.517
R10 VPB.t0 VPB.t3 214.517
R11 A.n0 A.t1 250.641
R12 A.n0 A.t0 231.629
R13 A A.n0 155.721
R14 a_524_368.t0 a_524_368.t1 76.8305
R15 VPWR.n1 VPWR.t0 368.615
R16 VPWR.n1 VPWR.n0 322.332
R17 VPWR.n0 VPWR.t1 66.9805
R18 VPWR.n0 VPWR.t2 35.2408
R19 VPWR VPWR.n1 0.198961
R20 a_228_74.n1 a_228_74.t5 264.298
R21 a_228_74.n2 a_228_74.n0 255.59
R22 a_228_74.t0 a_228_74.n4 230.768
R23 a_228_74.n1 a_228_74.t6 204.048
R24 a_228_74.n4 a_228_74.n2 175.737
R25 a_228_74.n2 a_228_74.n1 152
R26 a_228_74.n4 a_228_74.n3 117.097
R27 a_228_74.n3 a_228_74.t3 83.6754
R28 a_228_74.n3 a_228_74.t1 81.1792
R29 a_228_74.n0 a_228_74.t4 30.546
R30 a_228_74.n0 a_228_74.t2 30.546
R31 VGND.n5 VGND.n2 213.417
R32 VGND.n11 VGND.n10 210.018
R33 VGND.n4 VGND.n3 208.661
R34 VGND.n2 VGND.t5 53.455
R35 VGND.n2 VGND.t3 48.0026
R36 VGND.n3 VGND.t2 45.8187
R37 VGND.n3 VGND.t4 45.8187
R38 VGND.n10 VGND.t0 45.8187
R39 VGND.n10 VGND.t1 45.8187
R40 VGND.n8 VGND.n1 36.1417
R41 VGND.n9 VGND.n8 36.1417
R42 VGND.n11 VGND.n9 19.2005
R43 VGND.n5 VGND.n4 10.9526
R44 VGND.n6 VGND.n1 9.3005
R45 VGND.n8 VGND.n7 9.3005
R46 VGND.n9 VGND.n0 9.3005
R47 VGND.n4 VGND.n1 7.52991
R48 VGND.n12 VGND.n11 7.43488
R49 VGND.n6 VGND.n5 0.57347
R50 VGND VGND.n12 0.160103
R51 VGND.n12 VGND.n0 0.1477
R52 VGND.n7 VGND.n6 0.122949
R53 VGND.n7 VGND.n0 0.122949
R54 VNB.t0 VNB.t4 2482.94
R55 VNB.t5 VNB.t3 1489.76
R56 VNB.t4 VNB.t2 1316.54
R57 VNB.t1 VNB.t0 1316.54
R58 VNB VNB.t1 1143.31
R59 VNB.t2 VNB.t5 993.177
R60 D_N.n0 D_N.t0 282.774
R61 D_N.n0 D_N.t1 252.296
R62 D_N D_N.n0 161.697
R63 a_27_74.t0 a_27_74.n1 441.423
R64 a_27_74.n0 a_27_74.t2 377.276
R65 a_27_74.n0 a_27_74.t3 300.447
R66 a_27_74.n1 a_27_74.t1 299.75
R67 a_27_74.n1 a_27_74.n0 165.145
R68 X.n1 X 589
R69 X.n1 X.n0 585
R70 X.n2 X.n1 585
R71 X X.t1 204.773
R72 X.n1 X.t0 26.3844
R73 X X.n2 10.7205
R74 X X.n0 9.2805
R75 X X.n0 2.5605
R76 X.n2 X 1.1205
R77 B.n0 B.t1 277.151
R78 B.n0 B.t0 196.013
R79 B.n1 B.n0 152
R80 B B.n1 9.11565
R81 B.n1 B 5.23686
C0 VPB A 0.038226f
C1 VPWR C 0.008103f
C2 X B 2.3e-19
C3 VGND C 0.021348f
C4 B A 0.097314f
C5 VGND VPWR 0.069727f
C6 VPB B 0.031323f
C7 D_N VPWR 0.018158f
C8 X C 1.4e-19
C9 X VPWR 0.104887f
C10 VGND D_N 0.016608f
C11 VPB C 0.028316f
C12 VPWR A 0.012973f
C13 VPB VPWR 0.140433f
C14 X VGND 0.082836f
C15 VGND A 0.011245f
C16 C B 0.11568f
C17 X D_N 5.91e-20
C18 VGND VPB 0.011152f
C19 VPWR B 0.009962f
C20 VPB D_N 0.068197f
C21 VGND B 0.028116f
C22 X A 0.001995f
C23 X VPB 0.015925f
C24 VGND VNB 0.549511f
C25 X VNB 0.114232f
C26 A VNB 0.123203f
C27 B VNB 0.119886f
C28 C VNB 0.139474f
C29 VPWR VNB 0.436155f
C30 D_N VNB 0.177692f
C31 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4_4 VNB VPB VPWR VGND X D C B A
X0 X.t7 a_83_264.t6 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_83_264.t4 B.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1835 ps=1.27 w=0.74 l=0.15
X2 VGND.t3 a_83_264.t7 X.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1835 pd=1.27 as=0.22385 ps=1.345 w=0.74 l=0.15
X3 VGND.t6 D.t0 a_83_264.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.3445 pd=3.08 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 a_588_392.t3 A.t0 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.15 ps=1.3 w=1 l=0.15
X5 a_499_392.t3 C.t0 a_962_392.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.15 ps=1.3 w=1 l=0.15
X6 VPWR.t4 A.t1 a_588_392.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X7 a_962_392.t1 D.t1 a_83_264.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X8 X.t2 a_83_264.t8 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X9 a_588_392.t1 B.t1 a_499_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X10 a_83_264.t3 D.t2 a_962_392.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X11 a_83_264.t5 C.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.5035 ps=2.07 w=0.74 l=0.15
X12 X.t1 a_83_264.t9 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.22385 pd=1.345 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 VPWR.t3 a_83_264.t10 X.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X14 X.t5 a_83_264.t11 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_962_392.t3 C.t2 a_499_392.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X16 VPWR.t1 a_83_264.t12 X.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 VGND.t5 A.t2 a_83_264.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.5035 pd=2.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VGND.t0 a_83_264.t13 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_499_392.t0 B.t2 a_588_392.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
R0 a_83_264.n15 a_83_264.n14 836.763
R1 a_83_264.n2 a_83_264.t6 267.832
R2 a_83_264.n3 a_83_264.t12 256.264
R3 a_83_264.n9 a_83_264.t10 234.841
R4 a_83_264.n5 a_83_264.t11 234.841
R5 a_83_264.n10 a_83_264.t7 199.519
R6 a_83_264.n2 a_83_264.t8 186.374
R7 a_83_264.n4 a_83_264.t13 186.374
R8 a_83_264.n7 a_83_264.t9 186.374
R9 a_83_264.n6 a_83_264.n1 165.189
R10 a_83_264.n8 a_83_264.n1 152
R11 a_83_264.n11 a_83_264.n10 152
R12 a_83_264.n14 a_83_264.n13 116.24
R13 a_83_264.n13 a_83_264.n12 95.8655
R14 a_83_264.n14 a_83_264.n0 95.0012
R15 a_83_264.n13 a_83_264.n11 81.4094
R16 a_83_264.n3 a_83_264.n2 75.1925
R17 a_83_264.n5 a_83_264.n4 74.842
R18 a_83_264.n8 a_83_264.n7 47.4702
R19 a_83_264.n10 a_83_264.n9 44.549
R20 a_83_264.n0 a_83_264.t1 34.0546
R21 a_83_264.t2 a_83_264.n15 29.5505
R22 a_83_264.n15 a_83_264.t3 29.5505
R23 a_83_264.n0 a_83_264.t5 22.7032
R24 a_83_264.n12 a_83_264.t0 22.7032
R25 a_83_264.n12 a_83_264.t4 22.7032
R26 a_83_264.n11 a_83_264.n1 13.1884
R27 a_83_264.n6 a_83_264.n5 10.955
R28 a_83_264.n4 a_83_264.n3 7.7125
R29 a_83_264.n9 a_83_264.n8 5.11262
R30 a_83_264.n7 a_83_264.n6 2.19141
R31 VPWR.n5 VPWR.n4 610.986
R32 VPWR.n3 VPWR.t3 342.784
R33 VPWR.n10 VPWR.t0 342.783
R34 VPWR.n8 VPWR.n2 316.399
R35 VPWR.n4 VPWR.t5 29.5505
R36 VPWR.n4 VPWR.t4 29.5505
R37 VPWR.n2 VPWR.t2 26.3844
R38 VPWR.n2 VPWR.t1 26.3844
R39 VPWR.n8 VPWR.n7 25.224
R40 VPWR.n9 VPWR.n8 22.2123
R41 VPWR.n10 VPWR.n9 20.7064
R42 VPWR.n7 VPWR.n3 17.6946
R43 VPWR.n7 VPWR.n6 9.3005
R44 VPWR.n8 VPWR.n1 9.3005
R45 VPWR.n9 VPWR.n0 9.3005
R46 VPWR.n11 VPWR.n10 9.3005
R47 VPWR.n5 VPWR.n3 7.35647
R48 VPWR.n6 VPWR.n5 0.220535
R49 VPWR.n6 VPWR.n1 0.122949
R50 VPWR.n1 VPWR.n0 0.122949
R51 VPWR.n11 VPWR.n0 0.122949
R52 VPWR VPWR.n11 0.0617245
R53 X.n6 X.n2 204.335
R54 X.n1 X.n0 203.242
R55 X.n5 X.n3 150.994
R56 X.n5 X.n4 100.547
R57 X.n3 X.t3 64.0546
R58 X.n3 X.t1 34.0546
R59 X.n0 X.t6 26.3844
R60 X.n0 X.t5 26.3844
R61 X.n2 X.t4 26.3844
R62 X.n2 X.t7 26.3844
R63 X.n4 X.t0 22.7032
R64 X.n4 X.t2 22.7032
R65 X X.n5 19.262
R66 X.n1 X 17.2611
R67 X X.n6 6.59444
R68 X X.n1 1.35808
R69 X.n6 X 0.546841
R70 VPB.t2 VPB.t6 515.861
R71 VPB VPB.t3 257.93
R72 VPB.t9 VPB.t5 255.376
R73 VPB.t7 VPB.t9 255.376
R74 VPB.t10 VPB.t7 240.054
R75 VPB.t4 VPB.t11 229.839
R76 VPB.t5 VPB.t4 229.839
R77 VPB.t8 VPB.t10 229.839
R78 VPB.t6 VPB.t8 229.839
R79 VPB.t1 VPB.t2 229.839
R80 VPB.t0 VPB.t1 229.839
R81 VPB.t3 VPB.t0 229.839
R82 B B.t2 525.755
R83 B.n0 B.t1 298.572
R84 B.n0 B.t0 178.34
R85 B.n1 B.n0 152
R86 B.n1 B 7.77193
R87 B.n2 B.n1 5.02907
R88 B.n2 B 2.74336
R89 B B.n2 1.82907
R90 VGND.n23 VGND.n2 207.498
R91 VGND.n18 VGND.n17 201.179
R92 VGND.n10 VGND.n4 185
R93 VGND.n12 VGND.n11 185
R94 VGND.n9 VGND.n8 185
R95 VGND.n7 VGND.t6 156.976
R96 VGND.n25 VGND.t2 154.727
R97 VGND.n11 VGND.n9 62.2505
R98 VGND.n11 VGND.n10 62.2505
R99 VGND.n17 VGND.t4 38.1086
R100 VGND.n17 VGND.t3 38.1086
R101 VGND.n19 VGND.n1 36.1417
R102 VGND.n2 VGND.t0 34.0546
R103 VGND.n10 VGND.t5 33.9127
R104 VGND.n9 VGND.t7 33.9127
R105 VGND.n24 VGND.n23 29.7417
R106 VGND.n18 VGND.n16 28.6123
R107 VGND.n16 VGND.n4 26.3374
R108 VGND.n2 VGND.t1 22.7032
R109 VGND.n25 VGND.n24 20.7064
R110 VGND.n23 VGND.n1 17.6946
R111 VGND.n19 VGND.n18 16.5652
R112 VGND.n8 VGND.n7 9.74573
R113 VGND.n26 VGND.n25 9.3005
R114 VGND.n6 VGND.n5 9.3005
R115 VGND.n14 VGND.n13 9.3005
R116 VGND.n16 VGND.n15 9.3005
R117 VGND.n18 VGND.n3 9.3005
R118 VGND.n20 VGND.n19 9.3005
R119 VGND.n21 VGND.n1 9.3005
R120 VGND.n23 VGND.n22 9.3005
R121 VGND.n24 VGND.n0 9.3005
R122 VGND.n13 VGND.n12 7.44447
R123 VGND.n8 VGND.n6 6.26433
R124 VGND.n12 VGND.n6 1.27142
R125 VGND.n7 VGND.n5 0.427083
R126 VGND.n14 VGND.n5 0.122949
R127 VGND.n15 VGND.n14 0.122949
R128 VGND.n15 VGND.n3 0.122949
R129 VGND.n20 VGND.n3 0.122949
R130 VGND.n21 VGND.n20 0.122949
R131 VGND.n22 VGND.n21 0.122949
R132 VGND.n22 VGND.n0 0.122949
R133 VGND.n26 VGND.n0 0.122949
R134 VGND.n13 VGND.n4 0.0912801
R135 VGND VGND.n26 0.0617245
R136 VNB.t5 VNB.t7 3279.79
R137 VNB.t1 VNB.t3 1743.83
R138 VNB.t3 VNB.t4 1432.02
R139 VNB VNB.t2 1304.99
R140 VNB.t7 VNB.t6 1154.86
R141 VNB.t0 VNB.t1 1154.86
R142 VNB.t4 VNB.t5 993.177
R143 VNB.t2 VNB.t0 993.177
R144 D D.n1 377.685
R145 D.n1 D.t1 291.878
R146 D.n0 D.t2 291.878
R147 D.n0 D.t0 145.404
R148 D.n1 D.n0 72.3005
R149 A.n0 A.t2 236.764
R150 A.n1 A.t0 236.011
R151 A.n0 A.t1 207.529
R152 A A.n1 154.133
R153 A.n1 A.n0 37.246
R154 a_588_392.n1 a_588_392.n0 637.018
R155 a_588_392.n0 a_588_392.t0 31.5205
R156 a_588_392.n0 a_588_392.t3 31.5205
R157 a_588_392.t2 a_588_392.n1 29.5505
R158 a_588_392.n1 a_588_392.t1 29.5505
R159 C C.t0 408.647
R160 C.n0 C.t1 249.034
R161 C.n0 C.t2 239.661
R162 C C.n0 157.825
R163 a_962_392.n1 a_962_392.n0 1211.14
R164 a_962_392.n0 a_962_392.t3 39.4005
R165 a_962_392.n0 a_962_392.t0 29.5505
R166 a_962_392.n1 a_962_392.t2 29.5505
R167 a_962_392.t1 a_962_392.n1 29.5505
R168 a_499_392.n1 a_499_392.t3 458.32
R169 a_499_392.t1 a_499_392.n1 366.974
R170 a_499_392.n1 a_499_392.n0 193.863
R171 a_499_392.n0 a_499_392.t0 39.4005
R172 a_499_392.n0 a_499_392.t2 29.5505
C0 B VGND 0.029538f
C1 C VPWR 0.020293f
C2 A X 0.001967f
C3 VPB X 0.024687f
C4 B C 0.067998f
C5 A VPB 0.075152f
C6 D VGND 0.120488f
C7 VPWR X 0.407698f
C8 B X 0.00237f
C9 C D 0.16437f
C10 A VPWR 0.026589f
C11 VPB VPWR 0.184606f
C12 B A 0.167509f
C13 B VPB 0.086029f
C14 D X 3.08e-19
C15 B VPWR 0.023027f
C16 C VGND 0.020597f
C17 A D 4.05e-20
C18 VPB D 0.074893f
C19 D VPWR 0.01176f
C20 X VGND 0.318226f
C21 B D 0.001396f
C22 A VGND 0.017322f
C23 C X 8.49e-20
C24 VPB VGND 0.013301f
C25 A C 0.009362f
C26 C VPB 0.091035f
C27 VPWR VGND 0.109687f
C28 VGND VNB 0.815311f
C29 X VNB 0.064279f
C30 VPWR VNB 0.642426f
C31 D VNB 0.412512f
C32 C VNB 0.188007f
C33 A VNB 0.155584f
C34 B VNB 0.207616f
C35 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3_4 VNB VPB VPWR VGND B A C X
X0 a_206_388.t2 B.t0 a_116_388.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X1 a_302_388.t1 C.t0 a_206_388.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR.t3 a_302_388.t5 X.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X.t5 a_302_388.t6 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2087 ps=1.505 w=1.12 l=0.15
X4 VGND.t4 a_302_388.t7 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VGND.t0 C.t1 a_302_388.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 X.t1 a_302_388.t8 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1258 ps=1.08 w=0.74 l=0.15
X7 a_116_388.t0 A.t0 VPWR.t4 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X8 X.t0 a_302_388.t9 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 VPWR.t5 A.t1 a_116_388.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2087 pd=1.505 as=0.175 ps=1.35 w=1 l=0.15
X10 VGND.t1 a_302_388.t10 X.t7 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.10545 ps=1.025 w=0.74 l=0.15
X11 VGND.t6 A.t2 a_302_388.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1258 ps=1.08 w=0.74 l=0.15
X12 a_116_388.t2 B.t1 a_206_388.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.1775 ps=1.355 w=1 l=0.15
X13 a_302_388.t3 B.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1332 ps=1.1 w=0.74 l=0.15
X14 VPWR.t1 a_302_388.t11 X.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_206_388.t3 C.t2 a_302_388.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1775 pd=1.355 as=0.15 ps=1.3 w=1 l=0.15
X16 X.t3 a_302_388.t12 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B.n1 B.t0 383.628
R1 B.n0 B.t2 252.248
R2 B.n0 B.t1 231.629
R3 B B.n0 163.831
R4 B.n1 B 12.9944
R5 B B.n1 5.62474
R6 a_116_388.n1 a_116_388.n0 621.463
R7 a_116_388.n0 a_116_388.t2 39.4005
R8 a_116_388.n0 a_116_388.t3 29.5505
R9 a_116_388.n1 a_116_388.t1 29.5505
R10 a_116_388.t0 a_116_388.n1 29.5505
R11 a_206_388.n1 a_206_388.n0 1218.13
R12 a_206_388.n0 a_206_388.t1 35.4605
R13 a_206_388.n0 a_206_388.t3 34.4755
R14 a_206_388.n1 a_206_388.t0 32.5055
R15 a_206_388.t2 a_206_388.n1 32.5055
R16 VPB.t9 VPB.t3 273.253
R17 VPB.t8 VPB.t4 257.93
R18 VPB VPB.t1 257.93
R19 VPB.t4 VPB.t9 255.376
R20 VPB.t5 VPB.t0 245.161
R21 VPB.t7 VPB.t6 229.839
R22 VPB.t2 VPB.t7 229.839
R23 VPB.t3 VPB.t2 229.839
R24 VPB.t0 VPB.t8 229.839
R25 VPB.t1 VPB.t5 229.839
R26 C C.n1 474.204
R27 C.n1 C.t0 322.091
R28 C.n0 C.t2 296.925
R29 C.n0 C.t1 227.76
R30 C.n1 C.n0 21.3433
R31 a_302_388.n16 a_302_388.n15 729.355
R32 a_302_388.n12 a_302_388.t6 240.928
R33 a_302_388.n4 a_302_388.t11 240.197
R34 a_302_388.n3 a_302_388.t12 240.197
R35 a_302_388.n9 a_302_388.t5 240.197
R36 a_302_388.n4 a_302_388.t7 181.407
R37 a_302_388.n12 a_302_388.t9 179.947
R38 a_302_388.n10 a_302_388.t10 179.947
R39 a_302_388.n5 a_302_388.t8 179.947
R40 a_302_388.n1 a_302_388.t2 168.834
R41 a_302_388.n7 a_302_388.n6 165.189
R42 a_302_388.n14 a_302_388.n13 152
R43 a_302_388.n11 a_302_388.n2 152
R44 a_302_388.n8 a_302_388.n7 152
R45 a_302_388.n1 a_302_388.n0 95.685
R46 a_302_388.n15 a_302_388.n1 59.4829
R47 a_302_388.n13 a_302_388.n11 49.6611
R48 a_302_388.n9 a_302_388.n8 44.549
R49 a_302_388.n6 a_302_388.n4 37.246
R50 a_302_388.n0 a_302_388.t3 32.4329
R51 a_302_388.n16 a_302_388.t0 29.5505
R52 a_302_388.t1 a_302_388.n16 29.5505
R53 a_302_388.n6 a_302_388.n5 24.1005
R54 a_302_388.n0 a_302_388.t4 22.7032
R55 a_302_388.n8 a_302_388.n3 21.1793
R56 a_302_388.n7 a_302_388.n2 13.1884
R57 a_302_388.n14 a_302_388.n2 13.1884
R58 a_302_388.n13 a_302_388.n12 10.2247
R59 a_302_388.n15 a_302_388.n14 7.3702
R60 a_302_388.n5 a_302_388.n3 4.38232
R61 a_302_388.n11 a_302_388.n10 3.65202
R62 a_302_388.n10 a_302_388.n9 1.46111
R63 X.n2 X.n0 268.01
R64 X.n2 X.n1 207.6
R65 X.n5 X.n3 157.029
R66 X.n5 X.n4 102.019
R67 X X.n2 32.7862
R68 X X.n5 29.5125
R69 X.n0 X.t6 26.3844
R70 X.n0 X.t5 26.3844
R71 X.n1 X.t4 26.3844
R72 X.n1 X.t3 26.3844
R73 X.n3 X.t0 23.514
R74 X.n3 X.t7 22.7032
R75 X.n4 X.t2 22.7032
R76 X.n4 X.t1 22.7032
R77 VPWR.n7 VPWR.t1 358.716
R78 VPWR.n6 VPWR.n5 325.255
R79 VPWR.n10 VPWR.n4 315.928
R80 VPWR.n18 VPWR.t4 261.757
R81 VPWR.n4 VPWR.t5 46.2955
R82 VPWR.n12 VPWR.n11 36.1417
R83 VPWR.n12 VPWR.n1 36.1417
R84 VPWR.n16 VPWR.n1 36.1417
R85 VPWR.n17 VPWR.n16 36.1417
R86 VPWR.n11 VPWR.n10 29.7417
R87 VPWR.n18 VPWR.n17 26.7299
R88 VPWR.n5 VPWR.t0 26.3844
R89 VPWR.n5 VPWR.t3 26.3844
R90 VPWR.n4 VPWR.t2 25.6649
R91 VPWR.n9 VPWR.n6 25.224
R92 VPWR.n10 VPWR.n9 17.6946
R93 VPWR.n9 VPWR.n8 9.3005
R94 VPWR.n10 VPWR.n3 9.3005
R95 VPWR.n11 VPWR.n2 9.3005
R96 VPWR.n13 VPWR.n12 9.3005
R97 VPWR.n14 VPWR.n1 9.3005
R98 VPWR.n16 VPWR.n15 9.3005
R99 VPWR.n17 VPWR.n0 9.3005
R100 VPWR.n19 VPWR.n18 9.3005
R101 VPWR.n7 VPWR.n6 6.95806
R102 VPWR.n8 VPWR.n7 0.546775
R103 VPWR.n8 VPWR.n3 0.122949
R104 VPWR.n3 VPWR.n2 0.122949
R105 VPWR.n13 VPWR.n2 0.122949
R106 VPWR.n14 VPWR.n13 0.122949
R107 VPWR.n15 VPWR.n14 0.122949
R108 VPWR.n15 VPWR.n0 0.122949
R109 VPWR.n19 VPWR.n0 0.122949
R110 VPWR VPWR.n19 0.0617245
R111 VGND.n5 VGND.t4 238.069
R112 VGND.n4 VGND.n3 214.185
R113 VGND.n8 VGND.n2 204.976
R114 VGND.n11 VGND.n10 204.976
R115 VGND.n2 VGND.t6 34.0546
R116 VGND.n10 VGND.t0 34.0546
R117 VGND.n3 VGND.t3 32.4329
R118 VGND.n9 VGND.n8 30.8711
R119 VGND.n10 VGND.t5 24.3248
R120 VGND.n4 VGND.n1 23.7181
R121 VGND.n3 VGND.t1 22.7032
R122 VGND.n2 VGND.t2 22.7032
R123 VGND.n11 VGND.n9 19.577
R124 VGND.n8 VGND.n1 16.5652
R125 VGND.n9 VGND.n0 9.3005
R126 VGND.n8 VGND.n7 9.3005
R127 VGND.n6 VGND.n1 9.3005
R128 VGND.n12 VGND.n11 7.34641
R129 VGND.n5 VGND.n4 6.96039
R130 VGND.n6 VGND.n5 0.594857
R131 VGND VGND.n12 0.522673
R132 VGND.n12 VGND.n0 0.154231
R133 VGND.n7 VGND.n6 0.122949
R134 VGND.n7 VGND.n0 0.122949
R135 VNB VNB.t0 4457.74
R136 VNB.t0 VNB.t5 1177.95
R137 VNB.t6 VNB.t2 1154.86
R138 VNB.t1 VNB.t3 1131.76
R139 VNB.t5 VNB.t6 1131.76
R140 VNB.t2 VNB.t1 1004.72
R141 VNB.t3 VNB.t4 993.177
R142 A.n1 A.n0 335.022
R143 A.n1 A.t0 328.216
R144 A.n0 A.t1 293.217
R145 A.n0 A.t2 178.34
R146 A A.n1 0.350511
C0 C VGND 0.067124f
C1 VGND A 0.095654f
C2 C VPB 0.07239f
C3 VPB A 0.090268f
C4 VPWR X 0.37611f
C5 X B 3.03e-19
C6 VGND VPB 0.009677f
C7 C X 7.5e-19
C8 X A 0.002008f
C9 VPWR B 0.020692f
C10 X VGND 0.256385f
C11 C VPWR 0.012155f
C12 VPWR A 0.059751f
C13 X VPB 0.014129f
C14 C B 0.138941f
C15 A B 0.303862f
C16 VPWR VGND 0.086266f
C17 VGND B 0.019796f
C18 C A 0.128201f
C19 VPWR VPB 0.158262f
C20 VPB B 0.085261f
C21 VGND VNB 0.656607f
C22 X VNB 0.074841f
C23 VPWR VNB 0.574654f
C24 C VNB 0.317912f
C25 B VNB 0.166073f
C26 A VNB 0.44126f
C27 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3_2 VNB VPB VPWR VGND X C A B
X0 VGND.t2 a_27_74.t4 X.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_27_74.t1 B.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1616 ps=1.145 w=0.64 l=0.15
X2 VGND.t0 C.t0 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1616 pd=1.145 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 X.t2 a_27_74.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1933 ps=1.305 w=0.74 l=0.15
X4 VPWR.t1 a_27_74.t6 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5 X.t1 a_27_74.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2459 ps=1.58 w=1.12 l=0.15
X6 a_234_392.t1 B.t1 a_150_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X7 a_150_392.t0 C.t1 a_27_74.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X8 VPWR.t2 A.t0 a_234_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2459 pd=1.58 as=0.21 ps=1.42 w=1 l=0.15
X9 VGND.t4 A.t1 a_27_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1933 pd=1.305 as=0.112 ps=0.99 w=0.64 l=0.15
R0 a_27_74.t2 a_27_74.n7 321.995
R1 a_27_74.n3 a_27_74.t7 245.31
R2 a_27_74.n0 a_27_74.t6 240.197
R3 a_27_74.n7 a_27_74.t0 219.113
R4 a_27_74.n0 a_27_74.t4 192.102
R5 a_27_74.n6 a_27_74.n5 185
R6 a_27_74.n2 a_27_74.t5 179.947
R7 a_27_74.n4 a_27_74.n1 165.189
R8 a_27_74.n4 a_27_74.n3 152
R9 a_27_74.n6 a_27_74.n4 82.3163
R10 a_27_74.n7 a_27_74.n6 60.3099
R11 a_27_74.n2 a_27_74.n1 41.6278
R12 a_27_74.n5 a_27_74.t3 39.3755
R13 a_27_74.n5 a_27_74.t1 26.2505
R14 a_27_74.n1 a_27_74.n0 10.955
R15 a_27_74.n3 a_27_74.n2 8.03383
R16 X X.n0 250.173
R17 X X.n1 128.53
R18 X.n0 X.t0 26.3844
R19 X.n0 X.t1 26.3844
R20 X.n1 X.t3 22.7032
R21 X.n1 X.t2 22.7032
R22 VGND.n3 VGND.t2 247.887
R23 VGND.n8 VGND.n7 200.885
R24 VGND.n2 VGND.n1 185
R25 VGND.n1 VGND.t1 56.4111
R26 VGND.n7 VGND.t3 47.813
R27 VGND.n7 VGND.t0 46.8755
R28 VGND.n1 VGND.t4 45.938
R29 VGND.n6 VGND.n5 36.1417
R30 VGND.n8 VGND.n6 12.8005
R31 VGND.n3 VGND.n2 10.5884
R32 VGND.n6 VGND.n0 9.3005
R33 VGND.n5 VGND.n4 9.3005
R34 VGND.n9 VGND.n8 7.43488
R35 VGND.n5 VGND.n2 6.55164
R36 VGND.n4 VGND.n3 0.579212
R37 VGND VGND.n9 0.160103
R38 VGND.n9 VGND.n0 0.1477
R39 VGND.n4 VGND.n0 0.122949
R40 VNB.t4 VNB.t1 1651.44
R41 VNB.t0 VNB.t3 1512.86
R42 VNB.t3 VNB.t4 1154.86
R43 VNB VNB.t0 1143.31
R44 VNB.t1 VNB.t2 993.177
R45 B.n0 B.t1 252.206
R46 B.n0 B.t0 187.85
R47 B B.n0 80.6631
R48 C.n0 C.t1 233.258
R49 C.n1 C.t0 161.226
R50 C C.n0 153.44
R51 C.n2 C.n1 152
R52 C.n1 C.n0 47.5019
R53 C C.n2 9.4405
R54 C.n2 C 2.4005
R55 VPWR.n1 VPWR.t1 359.882
R56 VPWR.n1 VPWR.n0 228.681
R57 VPWR.n0 VPWR.t0 59.0707
R58 VPWR.n0 VPWR.t2 29.5505
R59 VPWR VPWR.n1 0.668459
R60 VPB VPB.t2 344.759
R61 VPB.t3 VPB.t0 311.56
R62 VPB.t4 VPB.t3 291.13
R63 VPB.t0 VPB.t1 229.839
R64 VPB.t2 VPB.t4 214.517
R65 a_150_392.t0 a_150_392.t1 53.1905
R66 a_234_392.t0 a_234_392.t1 82.7405
R67 A.n0 A.t0 298.572
R68 A.n0 A.t1 194.407
R69 A A.n0 158.589
C0 C VPWR 0.011915f
C1 X VGND 0.138001f
C2 C B 0.133191f
C3 A VGND 0.014099f
C4 VPB X 0.014225f
C5 A VPB 0.043222f
C6 VPWR VGND 0.056915f
C7 A X 0.002664f
C8 B VGND 0.013267f
C9 VPB VPWR 0.105152f
C10 B VPB 0.047111f
C11 VPWR X 0.215124f
C12 A VPWR 0.032356f
C13 B X 0.005527f
C14 C VGND 0.015843f
C15 B A 0.102782f
C16 C VPB 0.047551f
C17 B VPWR 0.081147f
C18 C A 2.79e-20
C19 VPB VGND 0.008991f
C20 VGND VNB 0.453271f
C21 X VNB 0.063308f
C22 VPWR VNB 0.384094f
C23 A VNB 0.118983f
C24 B VNB 0.115871f
C25 C VNB 0.155202f
C26 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3_1 VNB VPB VPWR VGND A B C X
X0 a_116_368.t0 C.t0 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X1 VGND.t0 C.t1 a_27_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 VGND.t1 A.t0 a_27_74.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.13925 pd=1.16 as=0.182875 ps=1.215 w=0.55 l=0.15
X3 a_200_368.t1 B.t0 a_116_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t0 A.t1 a_200_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3809 pd=1.85 as=0.21 ps=1.42 w=1 l=0.15
X5 a_27_74.t3 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.182875 pd=1.215 as=0.09625 ps=0.9 w=0.55 l=0.15
X6 X.t0 a_27_74.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.13925 ps=1.16 w=0.74 l=0.15
X7 X.t1 a_27_74.t5 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3809 ps=1.85 w=1.12 l=0.15
R0 C.n0 C.t1 250.641
R1 C.n0 C.t0 233.697
R2 C C.n0 159.442
R3 a_27_74.t0 a_27_74.n5 556.308
R4 a_27_74.n0 a_27_74.t1 292.7
R5 a_27_74.n4 a_27_74.t5 263.589
R6 a_27_74.n4 a_27_74.t4 203.339
R7 a_27_74.n1 a_27_74.n0 185
R8 a_27_74.n3 a_27_74.n2 185
R9 a_27_74.n5 a_27_74.n4 152
R10 a_27_74.n2 a_27_74.n1 84.0005
R11 a_27_74.n5 a_27_74.n3 48.9823
R12 a_27_74.n2 a_27_74.t2 30.546
R13 a_27_74.n1 a_27_74.t3 30.546
R14 a_27_74.n3 a_27_74.n0 6.79774
R15 a_116_368.t0 a_116_368.t1 53.1905
R16 VPB.t1 VPB.t3 449.462
R17 VPB.t2 VPB.t1 291.13
R18 VPB VPB.t0 257.93
R19 VPB.t0 VPB.t2 214.517
R20 VGND.n2 VGND.n0 216.088
R21 VGND.n2 VGND.n1 215.81
R22 VGND.n0 VGND.t1 45.8187
R23 VGND.n1 VGND.t2 45.8187
R24 VGND.n0 VGND.t3 39.2753
R25 VGND.n1 VGND.t0 30.546
R26 VGND VGND.n2 0.252924
R27 VNB.t2 VNB.t1 1882.41
R28 VNB.t1 VNB.t3 1316.54
R29 VNB.t0 VNB.t2 1154.86
R30 VNB VNB.t0 1143.31
R31 A.n0 A.t0 243.109
R32 A.n0 A.t1 224.097
R33 A A.n0 154.522
R34 B.n0 B.t1 250.641
R35 B.n0 B.t0 231.629
R36 B B.n0 155.423
R37 a_200_368.t0 a_200_368.t1 82.7405
R38 VPWR.n2 VPWR.n0 585
R39 VPWR.n1 VPWR.n0 585
R40 VPWR.n4 VPWR.n3 272.753
R41 VPWR.n3 VPWR.n2 39.4965
R42 VPWR.n3 VPWR.n1 39.4965
R43 VPWR.n2 VPWR.t0 29.5505
R44 VPWR.n1 VPWR.t1 27.5507
R45 VPWR VPWR.n4 14.4445
R46 VPWR.n4 VPWR.n0 5.72682
R47 X.n0 X.t1 296.899
R48 X.t0 X.n0 279.738
R49 X.n1 X.t0 279.738
R50 X.n1 X 11.3978
R51 X.n0 X 4.38406
R52 X X.n1 1.57858
C0 A VGND 0.016397f
C1 B VGND 0.016608f
C2 C VPWR 0.010149f
C3 B A 0.086245f
C4 VPB X 0.013291f
C5 C VGND 0.01702f
C6 VPB VPWR 0.084971f
C7 VPWR X 0.090752f
C8 C B 0.090136f
C9 VPB VGND 0.006464f
C10 X VGND 0.080913f
C11 VPB A 0.047125f
C12 A X 0.001954f
C13 VPB B 0.034148f
C14 B X 1.59e-19
C15 VPWR VGND 0.047553f
C16 A VPWR 0.020659f
C17 VPB C 0.037151f
C18 B VPWR 0.012144f
C19 C X 9.38e-20
C20 VGND VNB 0.384969f
C21 X VNB 0.1141f
C22 VPWR VNB 0.307461f
C23 A VNB 0.14374f
C24 B VNB 0.123513f
C25 C VNB 0.171265f
C26 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4b_2 VNB VPB VPWR VGND A B C D_N X
X0 VPWR.t3 D_N.t0 a_27_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 X.t1 a_190_48.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.127925 ps=1.105 w=0.74 l=0.15
X2 a_536_392.t1 B.t0 a_452_392.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t1 a_190_48.t6 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1533 pd=1.18 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_190_48.t4 C.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.1584 ps=1.135 w=0.64 l=0.15
X5 a_638_392.t0 C.t1 a_536_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.18 ps=1.36 w=1 l=0.15
X6 a_452_392.t0 A.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2884 ps=1.665 w=1 l=0.15
X7 a_190_48.t1 a_27_368.t2 a_638_392.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.445 pd=2.89 as=0.195 ps=1.39 w=1 l=0.15
X8 VGND.t4 D_N.t1 a_27_368.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.127925 pd=1.105 as=0.15675 ps=1.67 w=0.55 l=0.15
X9 VPWR.t0 a_190_48.t7 X.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2884 pd=1.665 as=0.168 ps=1.42 w=1.12 l=0.15
X10 X.t2 a_190_48.t8 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.203 ps=1.505 w=1.12 l=0.15
X11 VGND.t3 a_27_368.t3 a_190_48.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.104 ps=0.965 w=0.64 l=0.15
X12 a_190_48.t3 A.t1 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1408 pd=1.08 as=0.1533 ps=1.18 w=0.64 l=0.15
X13 VGND.t0 B.t1 a_190_48.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1584 pd=1.135 as=0.1408 ps=1.08 w=0.64 l=0.15
R0 D_N.n0 D_N.t0 204.95
R1 D_N.n0 D_N.t1 187.276
R2 D_N D_N.n0 158.847
R3 a_27_368.n1 a_27_368.n0 448.853
R4 a_27_368.t0 a_27_368.n1 340.56
R5 a_27_368.n1 a_27_368.t1 309.584
R6 a_27_368.n0 a_27_368.t2 239.661
R7 a_27_368.n0 a_27_368.t3 232.968
R8 VPWR.n2 VPWR.n1 678.548
R9 VPWR.n2 VPWR.n0 591.159
R10 VPWR.n1 VPWR.t3 55.1136
R11 VPWR.n0 VPWR.t2 54.1755
R12 VPWR.n0 VPWR.t0 51.3309
R13 VPWR.n1 VPWR.t1 29.6087
R14 VPWR VPWR.n2 0.465093
R15 VPB.t1 VPB.t4 354.974
R16 VPB.t3 VPB.t5 275.807
R17 VPB.t6 VPB.t2 273.253
R18 VPB.t0 VPB.t3 260.485
R19 VPB VPB.t6 257.93
R20 VPB.t2 VPB.t1 229.839
R21 VPB.t4 VPB.t0 214.517
R22 a_190_48.t1 a_190_48.n6 355.885
R23 a_190_48.n0 a_190_48.t8 308.481
R24 a_190_48.n2 a_190_48.t7 262.921
R25 a_190_48.n4 a_190_48.n2 209.698
R26 a_190_48.n0 a_190_48.t5 200.03
R27 a_190_48.n1 a_190_48.t6 190.275
R28 a_190_48.n4 a_190_48.n3 98.8784
R29 a_190_48.n6 a_190_48.n5 98.8784
R30 a_190_48.n1 a_190_48.n0 80.3338
R31 a_190_48.n6 a_190_48.n4 65.5064
R32 a_190_48.n3 a_190_48.t0 41.2505
R33 a_190_48.n3 a_190_48.t3 41.2505
R34 a_190_48.n5 a_190_48.t4 34.688
R35 a_190_48.n5 a_190_48.t2 26.2505
R36 a_190_48.n2 a_190_48.n1 12.3948
R37 VGND.n3 VGND.t3 257.844
R38 VGND.n13 VGND.n12 215.464
R39 VGND.n10 VGND.n2 203.744
R40 VGND.n5 VGND.n4 200.138
R41 VGND.n4 VGND.t6 48.7505
R42 VGND.n12 VGND.t4 48.0005
R43 VGND.n2 VGND.t1 44.2236
R44 VGND.n4 VGND.t0 44.063
R45 VGND.n6 VGND.n1 36.1417
R46 VGND.n2 VGND.t5 34.688
R47 VGND.n11 VGND.n10 28.2358
R48 VGND.n13 VGND.n11 23.3417
R49 VGND.n12 VGND.t2 22.2054
R50 VGND.n10 VGND.n1 12.424
R51 VGND.n7 VGND.n6 9.3005
R52 VGND.n8 VGND.n1 9.3005
R53 VGND.n10 VGND.n9 9.3005
R54 VGND.n11 VGND.n0 9.3005
R55 VGND.n14 VGND.n13 7.5068
R56 VGND.n5 VGND.n3 6.96039
R57 VGND.n6 VGND.n5 3.38874
R58 VGND.n7 VGND.n3 0.594857
R59 VGND VGND.n14 0.16105
R60 VGND.n14 VGND.n0 0.146765
R61 VGND.n8 VGND.n7 0.122949
R62 VGND.n9 VGND.n8 0.122949
R63 VGND.n9 VGND.n0 0.122949
R64 X X.n0 586.212
R65 X X.n1 159.067
R66 X.n0 X.t3 26.3844
R67 X.n0 X.t2 26.3844
R68 X.n1 X.t0 22.7032
R69 X.n1 X.t1 22.7032
R70 VNB.t0 VNB.t6 1489.76
R71 VNB.t5 VNB.t0 1362.73
R72 VNB.t1 VNB.t5 1362.73
R73 VNB.t4 VNB.t2 1189.5
R74 VNB VNB.t4 1177.95
R75 VNB.t6 VNB.t3 1097.11
R76 VNB.t2 VNB.t1 993.177
R77 B.n0 B.t1 242.607
R78 B.n0 B.t0 231.629
R79 B.n1 B.n0 152
R80 B.n1 B 12.2187
R81 B B.n1 2.13383
R82 a_452_392.t0 a_452_392.t1 53.1905
R83 a_536_392.t0 a_536_392.t1 70.9205
R84 C.n0 C.t0 242.607
R85 C.n0 C.t1 231.629
R86 C.n1 C.n0 152
R87 C.n1 C 11.5205
R88 C C.n1 2.01193
R89 a_638_392.t0 a_638_392.t1 76.8305
R90 A.n0 A.t0 263.762
R91 A.n0 A.t1 204.048
R92 A A.n0 154.522
C0 B VPWR 0.008301f
C1 VGND C 0.01603f
C2 X VPWR 0.015659f
C3 VPB C 0.042791f
C4 A B 0.113635f
C5 VGND VPB 0.008676f
C6 X A 0.019941f
C7 B C 0.10971f
C8 VGND B 0.013075f
C9 D_N VPWR 0.00817f
C10 X C 3.39e-19
C11 X VGND 0.119756f
C12 VPB B 0.041018f
C13 D_N A 2.31e-19
C14 X VPB 0.003928f
C15 D_N VGND 0.012106f
C16 D_N VPB 0.044041f
C17 A VPWR 0.018619f
C18 D_N X 0.001208f
C19 C VPWR 0.010577f
C20 VGND VPWR 0.071376f
C21 VPB VPWR 0.118985f
C22 A C 7.15e-19
C23 VGND A 0.014378f
C24 VPB A 0.047008f
C25 VGND VNB 0.585509f
C26 X VNB 0.007748f
C27 D_N VNB 0.160869f
C28 VPWR VNB 0.433447f
C29 C VNB 0.10446f
C30 B VNB 0.106195f
C31 A VNB 0.111909f
C32 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4b_4 VNB VPB VPWR C VGND B A X D_N
X0 a_496_392.t3 C.t0 a_27_392.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X1 VGND.t8 D_N.t0 a_563_48.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.135 pd=1.115 as=0.32135 ps=2.98 w=0.64 l=0.15
X2 a_116_392.t2 B.t0 a_27_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X3 VGND.t4 C.t1 a_27_74.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.40885 ps=1.845 w=0.74 l=0.15
X4 X.t3 a_27_74.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.14985 pd=1.145 as=0.135 ps=1.115 w=0.74 l=0.15
X5 X.t5 a_27_74.t7 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t3 B.t1 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 X.t2 a_27_74.t8 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 a_27_392.t1 B.t2 a_116_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 VPWR.t2 D_N.t1 a_563_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.295 ps=2.59 w=1 l=0.15
X10 X.t4 a_27_74.t9 VPWR.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X11 a_27_74.t0 a_563_48.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X12 VGND.t6 a_27_74.t10 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VGND.t7 a_27_74.t11 X.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.14985 ps=1.145 w=0.74 l=0.15
X14 a_116_392.t0 A.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X15 VPWR.t1 A.t1 a_116_392.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X16 a_27_392.t2 C.t2 a_496_392.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X17 a_496_392.t0 a_563_48.t3 a_27_74.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X18 a_27_74.t1 a_563_48.t4 a_496_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X19 a_27_74.t4 A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.40885 pd=1.845 as=0.1554 ps=1.16 w=0.74 l=0.15
R0 C.n1 C.t2 482.471
R1 C.n0 C.t0 298.572
R2 C.n0 C.t1 178.34
R3 C.n1 C.n0 166.208
R4 C C.n1 0.0466957
R5 a_27_392.n1 a_27_392.t2 522.061
R6 a_27_392.t0 a_27_392.n1 364.44
R7 a_27_392.n1 a_27_392.n0 194.012
R8 a_27_392.n0 a_27_392.t1 39.4005
R9 a_27_392.n0 a_27_392.t3 29.5505
R10 a_496_392.n1 a_496_392.n0 1211.14
R11 a_496_392.n0 a_496_392.t3 39.4005
R12 a_496_392.n0 a_496_392.t1 29.5505
R13 a_496_392.t2 a_496_392.n1 29.5505
R14 a_496_392.n1 a_496_392.t0 29.5505
R15 VPB.t8 VPB.t0 515.861
R16 VPB.t10 VPB.t3 459.678
R17 VPB.t0 VPB.t10 273.253
R18 VPB VPB.t1 257.93
R19 VPB.t9 VPB.t6 255.376
R20 VPB.t4 VPB.t9 255.376
R21 VPB.t2 VPB.t4 255.376
R22 VPB.t5 VPB.t8 229.839
R23 VPB.t6 VPB.t5 229.839
R24 VPB.t7 VPB.t2 229.839
R25 VPB.t1 VPB.t7 229.839
R26 D_N.n0 D_N.t1 261.276
R27 D_N D_N.n0 158.054
R28 D_N.n0 D_N.t0 157.109
R29 a_563_48.n0 a_563_48.t1 783.351
R30 a_563_48.t0 a_563_48.n2 460.531
R31 a_563_48.n1 a_563_48.t2 236.764
R32 a_563_48.n0 a_563_48.t3 207.529
R33 a_563_48.n1 a_563_48.t4 207.529
R34 a_563_48.n2 a_563_48.n1 63.5369
R35 a_563_48.n2 a_563_48.n0 2.19141
R36 VGND.n6 VGND.n5 207.498
R37 VGND.n11 VGND.n10 206.333
R38 VGND.n26 VGND.n25 204.976
R39 VGND.n19 VGND.n18 203.57
R40 VGND.n7 VGND.t6 170.706
R41 VGND.n18 VGND.t0 43.7843
R42 VGND.n10 VGND.t8 41.2505
R43 VGND.n12 VGND.n3 36.1417
R44 VGND.n16 VGND.n3 36.1417
R45 VGND.n17 VGND.n16 36.1417
R46 VGND.n23 VGND.n1 36.1417
R47 VGND.n24 VGND.n23 36.1417
R48 VGND.n5 VGND.t5 34.0546
R49 VGND.n25 VGND.t2 34.0546
R50 VGND.n25 VGND.t3 34.0546
R51 VGND.n19 VGND.n17 29.7417
R52 VGND.n11 VGND.n9 27.4829
R53 VGND.n18 VGND.t4 24.3248
R54 VGND.n10 VGND.t1 23.252
R55 VGND.n9 VGND.n6 22.9652
R56 VGND.n5 VGND.t7 22.7032
R57 VGND.n12 VGND.n11 19.9534
R58 VGND.n26 VGND.n24 19.2005
R59 VGND.n19 VGND.n1 15.8123
R60 VGND.n24 VGND.n0 9.3005
R61 VGND.n23 VGND.n22 9.3005
R62 VGND.n21 VGND.n1 9.3005
R63 VGND.n20 VGND.n19 9.3005
R64 VGND.n17 VGND.n2 9.3005
R65 VGND.n16 VGND.n15 9.3005
R66 VGND.n14 VGND.n3 9.3005
R67 VGND.n13 VGND.n12 9.3005
R68 VGND.n11 VGND.n4 9.3005
R69 VGND.n9 VGND.n8 9.3005
R70 VGND.n27 VGND.n26 7.43488
R71 VGND.n7 VGND.n6 6.6595
R72 VGND.n8 VGND.n7 0.655456
R73 VGND VGND.n27 0.160103
R74 VGND.n27 VGND.n0 0.1477
R75 VGND.n8 VGND.n4 0.122949
R76 VGND.n13 VGND.n4 0.122949
R77 VGND.n14 VGND.n13 0.122949
R78 VGND.n15 VGND.n14 0.122949
R79 VGND.n15 VGND.n2 0.122949
R80 VGND.n20 VGND.n2 0.122949
R81 VGND.n21 VGND.n20 0.122949
R82 VGND.n22 VGND.n21 0.122949
R83 VGND.n22 VGND.n0 0.122949
R84 VNB.t0 VNB.t8 4169.03
R85 VNB.t2 VNB.t4 2898.69
R86 VNB.t4 VNB.t0 1316.54
R87 VNB.t3 VNB.t2 1316.54
R88 VNB.t1 VNB.t7 1281.89
R89 VNB.t8 VNB.t1 1212.6
R90 VNB.t7 VNB.t5 1154.86
R91 VNB VNB.t3 1143.31
R92 VNB.t5 VNB.t6 993.177
R93 B B.t2 529.266
R94 B.n0 B.t0 298.572
R95 B.n0 B.t1 178.34
R96 B.n1 B.n0 152
R97 B B.n1 8.0005
R98 B.n1 B 5.96414
R99 a_116_392.n1 a_116_392.n0 657.193
R100 a_116_392.n0 a_116_392.t0 39.4005
R101 a_116_392.n0 a_116_392.t1 29.5505
R102 a_116_392.n1 a_116_392.t3 29.5505
R103 a_116_392.t2 a_116_392.n1 29.5505
R104 a_27_74.n22 a_27_74.n21 668.938
R105 a_27_74.t0 a_27_74.n20 291.342
R106 a_27_74.n21 a_27_74.t0 279.738
R107 a_27_74.n3 a_27_74.n2 240.418
R108 a_27_74.n5 a_27_74.t7 234.841
R109 a_27_74.n7 a_27_74.n1 234.841
R110 a_27_74.n10 a_27_74.t9 234.841
R111 a_27_74.n11 a_27_74.t6 199.519
R112 a_27_74.n3 a_27_74.t10 187.864
R113 a_27_74.n8 a_27_74.t11 186.374
R114 a_27_74.n4 a_27_74.t8 185.704
R115 a_27_74.n15 a_27_74.t3 172.415
R116 a_27_74.n13 a_27_74.n12 168.18
R117 a_27_74.n6 a_27_74.n0 165.189
R118 a_27_74.n12 a_27_74.n11 152
R119 a_27_74.n9 a_27_74.n0 152
R120 a_27_74.n16 a_27_74.n15 92.5005
R121 a_27_74.n17 a_27_74.n14 92.5005
R122 a_27_74.n19 a_27_74.n18 92.5005
R123 a_27_74.n4 a_27_74.n3 63.6474
R124 a_27_74.n18 a_27_74.n17 61.6221
R125 a_27_74.n17 a_27_74.n16 60.8113
R126 a_27_74.n20 a_27_74.n19 55.9096
R127 a_27_74.n10 a_27_74.n9 43.8187
R128 a_27_74.n6 a_27_74.n5 37.9763
R129 a_27_74.n18 a_27_74.t5 34.0546
R130 a_27_74.t2 a_27_74.n22 29.5505
R131 a_27_74.n22 a_27_74.t1 29.5505
R132 a_27_74.n7 a_27_74.n6 27.752
R133 a_27_74.n16 a_27_74.t4 22.7032
R134 a_27_74.n9 a_27_74.n8 18.2581
R135 a_27_74.n12 a_27_74.n0 13.1884
R136 a_27_74.n19 a_27_74.n14 8.24457
R137 a_27_74.n15 a_27_74.n14 8.13609
R138 a_27_74.n11 a_27_74.n10 5.84292
R139 a_27_74.n8 a_27_74.n7 3.65202
R140 a_27_74.n5 a_27_74.n4 3.64028
R141 a_27_74.n20 a_27_74.n13 2.38983
R142 a_27_74.n21 a_27_74.n13 1.36583
R143 X X.t4 260.63
R144 X.n4 X.t5 229.895
R145 X.n2 X.n0 150.994
R146 X.n2 X.n1 103.043
R147 X.n3 X.n2 34.0747
R148 X.n0 X.t0 34.0546
R149 X.n0 X.t3 31.6221
R150 X.n1 X.t1 22.7032
R151 X.n1 X.t2 22.7032
R152 X.n3 X 14.1581
R153 X X.n4 3.10353
R154 X.n4 X.n3 1.35808
R155 VPWR.n1 VPWR.n0 605.365
R156 VPWR.n7 VPWR.t4 348.385
R157 VPWR.n6 VPWR.n5 232.787
R158 VPWR.n5 VPWR.t2 46.2955
R159 VPWR.n10 VPWR.n9 36.1417
R160 VPWR.n11 VPWR.n10 36.1417
R161 VPWR.n11 VPWR.n3 36.1417
R162 VPWR.n15 VPWR.n3 36.1417
R163 VPWR.n16 VPWR.n15 36.1417
R164 VPWR.n17 VPWR.n16 36.1417
R165 VPWR.n9 VPWR.n6 30.1181
R166 VPWR.n0 VPWR.t0 29.5505
R167 VPWR.n0 VPWR.t1 29.5505
R168 VPWR.n5 VPWR.t3 26.8503
R169 VPWR.n17 VPWR.n1 25.224
R170 VPWR.n9 VPWR.n8 9.3005
R171 VPWR.n10 VPWR.n4 9.3005
R172 VPWR.n12 VPWR.n11 9.3005
R173 VPWR.n13 VPWR.n3 9.3005
R174 VPWR.n15 VPWR.n14 9.3005
R175 VPWR.n16 VPWR.n2 9.3005
R176 VPWR.n18 VPWR.n17 9.3005
R177 VPWR.n19 VPWR.n1 7.06957
R178 VPWR.n7 VPWR.n6 6.74224
R179 VPWR.n8 VPWR.n7 0.520427
R180 VPWR VPWR.n19 0.273369
R181 VPWR.n19 VPWR.n18 0.157405
R182 VPWR.n8 VPWR.n4 0.122949
R183 VPWR.n12 VPWR.n4 0.122949
R184 VPWR.n13 VPWR.n12 0.122949
R185 VPWR.n14 VPWR.n13 0.122949
R186 VPWR.n14 VPWR.n2 0.122949
R187 VPWR.n18 VPWR.n2 0.122949
R188 A.n1 A.t0 247.208
R189 A.n0 A.t1 228.951
R190 A.n0 A.t2 228.148
R191 A A.n1 154.133
R192 A.n1 A.n0 15.3369
C0 VPB B 0.082895f
C1 X VPWR 0.401832f
C2 VGND C 0.084305f
C3 A VPWR 0.029308f
C4 VPB D_N 0.044588f
C5 B VPWR 0.022344f
C6 X VGND 0.297729f
C7 D_N VPWR 0.021279f
C8 X C 5.7e-19
C9 VGND A 0.014869f
C10 A C 0.009925f
C11 B VGND 0.023909f
C12 VPB VPWR 0.197864f
C13 B C 0.086059f
C14 D_N VGND 0.01395f
C15 D_N C 0.051294f
C16 VPB VGND 0.012619f
C17 B A 0.161243f
C18 VPB C 0.094872f
C19 D_N X 0.00175f
C20 VGND VPWR 0.089168f
C21 C VPWR 0.057569f
C22 VPB X 0.016387f
C23 VPB A 0.074675f
C24 VGND VNB 0.886012f
C25 X VNB 0.058761f
C26 D_N VNB 0.126449f
C27 VPWR VNB 0.686541f
C28 C VNB 0.232924f
C29 A VNB 0.162925f
C30 B VNB 0.255096f
C31 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4bb_1 VNB VPB VPWR VGND D_N C_N B A X
X0 a_216_424.t0 D_N.t0 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.1155 ps=0.97 w=0.55 l=0.15
X1 VGND.t6 C_N.t0 a_27_424.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 VGND.t5 A.t0 a_357_378.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.148875 pd=1.195 as=0.09625 ps=0.9 w=0.55 l=0.15
X3 X.t0 a_357_378.t5 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.148875 ps=1.195 w=0.74 l=0.15
X4 a_357_378.t2 B.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.114125 ps=0.965 w=0.55 l=0.15
X5 VPWR.t2 C_N.t1 a_27_424.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 a_626_378.t0 B.t1 a_530_378.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X7 VGND.t4 a_27_424.t2 a_357_378.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.114125 pd=0.965 as=0.092125 ps=0.885 w=0.55 l=0.15
X8 a_357_378.t1 a_216_424.t2 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.092125 pd=0.885 as=0.165 ps=1.7 w=0.55 l=0.15
X9 a_530_378.t1 a_27_424.t3 a_446_378.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10 X.t1 a_357_378.t6 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2362 ps=1.555 w=1.12 l=0.15
X11 a_216_424.t1 D_N.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.43785 pd=2.97 as=0.147 ps=1.19 w=0.84 l=0.15
X12 a_446_378.t0 a_216_424.t3 a_357_378.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X13 VPWR.t3 A.t1 a_626_378.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2362 pd=1.555 as=0.195 ps=1.39 w=1 l=0.15
R0 D_N.n0 D_N.t1 286.74
R1 D_N.n0 D_N.t0 169.302
R2 D_N D_N.n0 69.6965
R3 VGND.n1 VGND.t0 245.186
R4 VGND.n4 VGND.n3 213.571
R5 VGND.n14 VGND.n13 207.109
R6 VGND.n6 VGND.n5 201.69
R7 VGND.n5 VGND.t4 52.3641
R8 VGND.n3 VGND.t1 46.9117
R9 VGND.n3 VGND.t5 45.8187
R10 VGND.n13 VGND.t2 45.8187
R11 VGND.n13 VGND.t6 45.8187
R12 VGND.n5 VGND.t3 38.1823
R13 VGND.n8 VGND.n7 36.1417
R14 VGND.n12 VGND.n11 36.1417
R15 VGND.n14 VGND.n12 17.3181
R16 VGND.n11 VGND.n1 10.9181
R17 VGND.n7 VGND.n2 9.3005
R18 VGND.n9 VGND.n8 9.3005
R19 VGND.n11 VGND.n10 9.3005
R20 VGND.n12 VGND.n0 9.3005
R21 VGND.n7 VGND.n6 7.90638
R22 VGND.n15 VGND.n14 7.5068
R23 VGND.n6 VGND.n4 7.17299
R24 VGND.n8 VGND.n1 6.4005
R25 VGND.n4 VGND.n2 0.54632
R26 VGND VGND.n15 0.16105
R27 VGND.n15 VGND.n0 0.146765
R28 VGND.n9 VGND.n2 0.122949
R29 VGND.n10 VGND.n9 0.122949
R30 VGND.n10 VGND.n0 0.122949
R31 a_216_424.t1 a_216_424.n3 843.433
R32 a_216_424.n0 a_216_424.t0 238.268
R33 a_216_424.n2 a_216_424.t3 228.567
R34 a_216_424.n3 a_216_424.n2 152
R35 a_216_424.n1 a_216_424.n0 152
R36 a_216_424.n1 a_216_424.t2 136.141
R37 a_216_424.n2 a_216_424.n1 25.6068
R38 a_216_424.n3 a_216_424.n0 10.3624
R39 VNB.t1 VNB.t2 2425.2
R40 VNB.t5 VNB.t0 1397.38
R41 VNB.t6 VNB.t1 1316.54
R42 VNB.t4 VNB.t3 1304.99
R43 VNB VNB.t6 1201.05
R44 VNB.t3 VNB.t5 1154.86
R45 VNB.t2 VNB.t4 1120.21
R46 C_N.n0 C_N.t1 287.11
R47 C_N.n0 C_N.t0 227.395
R48 C_N C_N.n0 155.601
R49 a_27_424.t0 a_27_424.n1 402.029
R50 a_27_424.n1 a_27_424.n0 373.012
R51 a_27_424.n1 a_27_424.t1 322.168
R52 a_27_424.n0 a_27_424.t3 287.861
R53 a_27_424.n0 a_27_424.t2 199.227
R54 A.n0 A.t0 250.641
R55 A.n0 A.t1 245.018
R56 A A.n0 156.614
R57 a_357_378.t0 a_357_378.n4 463.322
R58 a_357_378.n0 a_357_378.t6 264.298
R59 a_357_378.n2 a_357_378.n0 206.833
R60 a_357_378.n0 a_357_378.t5 204.048
R61 a_357_378.n2 a_357_378.n1 196.249
R62 a_357_378.n4 a_357_378.n3 185
R63 a_357_378.n4 a_357_378.n2 58.4939
R64 a_357_378.n1 a_357_378.t2 45.8187
R65 a_357_378.n3 a_357_378.t1 42.546
R66 a_357_378.n3 a_357_378.t3 30.546
R67 a_357_378.n1 a_357_378.t4 30.546
R68 X.n0 X.t1 289.598
R69 X.t0 X.n0 279.738
R70 X.n1 X.t0 279.738
R71 X.n1 X 11.2437
R72 X.n0 X 4.32482
R73 X X.n1 1.55726
R74 B.n0 B.t0 250.641
R75 B.n0 B.t1 245.018
R76 B B.n0 154.522
R77 VPWR.n2 VPWR.n1 610.769
R78 VPWR.n2 VPWR.n0 228.911
R79 VPWR.n1 VPWR.t2 46.9053
R80 VPWR.n0 VPWR.t3 46.2955
R81 VPWR.n1 VPWR.t1 35.1791
R82 VPWR.n0 VPWR.t0 34.2292
R83 VPWR VPWR.n2 0.197993
R84 VPB.t2 VPB.t3 587.366
R85 VPB.t6 VPB.t1 298.791
R86 VPB.t0 VPB.t6 275.807
R87 VPB VPB.t4 257.93
R88 VPB.t4 VPB.t2 255.376
R89 VPB.t5 VPB.t0 245.161
R90 VPB.t3 VPB.t5 214.517
R91 a_530_378.t0 a_530_378.t1 65.0105
R92 a_626_378.t0 a_626_378.t1 76.8305
R93 a_446_378.t0 a_446_378.t1 53.1905
C0 VGND VPWR 0.076912f
C1 X B 0.003789f
C2 VPB VPWR 0.128686f
C3 VGND C_N 0.016226f
C4 X D_N 7.93e-20
C5 VPB C_N 0.06422f
C6 B A 0.107243f
C7 X VPWR 0.139646f
C8 VGND VPB 0.011578f
C9 VPWR A 0.031692f
C10 D_N B 1.46e-19
C11 X VGND 0.080445f
C12 X VPB 0.02126f
C13 VPWR B 0.07699f
C14 VGND A 0.014945f
C15 D_N VPWR 0.015744f
C16 VPB A 0.042037f
C17 C_N D_N 0.069026f
C18 X A 0.006876f
C19 VGND B 0.015166f
C20 VPB B 0.040641f
C21 C_N VPWR 0.014424f
C22 VGND D_N 0.024065f
C23 VPB D_N 0.066207f
C24 VGND VNB 0.598285f
C25 X VNB 0.113162f
C26 A VNB 0.123312f
C27 B VNB 0.116547f
C28 VPWR VNB 0.471774f
C29 D_N VNB 0.135821f
C30 C_N VNB 0.193971f
C31 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4bb_2 VNB VPB VPWR VGND X D_N C_N B A
X0 VPWR.t3 A.t0 a_689_392.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1874 pd=1.39 as=0.12 ps=1.24 w=1 l=0.15
X1 VPWR.t1 a_182_270.t5 X.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_587_392.t0 a_548_110.t2 a_503_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X3 a_548_110.t0 C_N.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=2.26 as=0.1874 ps=1.39 w=0.84 l=0.15
X4 X.t2 a_182_270.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1862 ps=1.475 w=1.12 l=0.15
X5 a_689_392.t1 B.t0 a_587_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.18 ps=1.36 w=1 l=0.15
X6 VGND.t4 A.t1 a_182_270.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.129925 pd=1.225 as=0.0928 ps=0.93 w=0.64 l=0.15
X7 VPWR.t4 D_N.t0 a_27_424.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2394 ps=2.25 w=0.84 l=0.15
X8 a_503_392.t0 a_27_424.t2 a_182_270.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X9 a_182_270.t1 a_27_424.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1668 pd=1.205 as=0.1997 ps=1.325 w=0.64 l=0.15
X10 VGND.t7 D_N.t1 a_27_424.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.127925 pd=1.105 as=0.15675 ps=1.67 w=0.55 l=0.15
X11 VGND.t3 a_548_110.t3 a_182_270.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.1668 ps=1.205 w=0.64 l=0.15
X12 a_548_110.t1 C_N.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.129925 ps=1.225 w=0.55 l=0.15
X13 X.t1 a_182_270.t7 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.127925 ps=1.105 w=0.74 l=0.15
X14 a_182_270.t4 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.1248 ps=1.03 w=0.64 l=0.15
X15 VGND.t5 a_182_270.t8 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1997 pd=1.325 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t0 231.629
R1 A.n0 A.t1 175.127
R2 A A.n0 164.412
R3 a_689_392.t0 a_689_392.t1 47.2805
R4 VPWR.n4 VPWR.t1 878.788
R5 VPWR.n6 VPWR.n1 605.753
R6 VPWR.n3 VPWR.n2 323.356
R7 VPWR.n2 VPWR.t0 56.2862
R8 VPWR.n1 VPWR.t4 46.9053
R9 VPWR.n1 VPWR.t2 32.1717
R10 VPWR.n2 VPWR.t3 30.7494
R11 VPWR.n5 VPWR.n4 23.3417
R12 VPWR.n6 VPWR.n5 19.9534
R13 VPWR.n5 VPWR.n0 9.3005
R14 VPWR.n7 VPWR.n6 7.40447
R15 VPWR.n4 VPWR.n3 7.16516
R16 VPWR VPWR.n7 0.159703
R17 VPWR.n3 VPWR.n0 0.159664
R18 VPWR.n7 VPWR.n0 0.148095
R19 VPB.t1 VPB.t4 505.646
R20 VPB.t5 VPB.t0 275.807
R21 VPB.t3 VPB.t6 260.485
R22 VPB.t7 VPB.t2 257.93
R23 VPB VPB.t7 252.823
R24 VPB.t2 VPB.t1 229.839
R25 VPB.t4 VPB.t3 214.517
R26 VPB.t6 VPB.t5 199.195
R27 a_182_270.t2 a_182_270.n5 934.744
R28 a_182_270.n0 a_182_270.t6 255.323
R29 a_182_270.n2 a_182_270.t5 248.303
R30 a_182_270.n5 a_182_270.n3 247.191
R31 a_182_270.n5 a_182_270.n2 212.236
R32 a_182_270.n1 a_182_270.t8 169.221
R33 a_182_270.n0 a_182_270.t7 154.24
R34 a_182_270.n5 a_182_270.n4 100.43
R35 a_182_270.n1 a_182_270.n0 70.7622
R36 a_182_270.n4 a_182_270.t0 39.8844
R37 a_182_270.n4 a_182_270.t1 34.479
R38 a_182_270.n3 a_182_270.t3 28.1255
R39 a_182_270.n3 a_182_270.t4 26.2505
R40 a_182_270.n2 a_182_270.n1 6.51401
R41 X.n1 X.n0 650.13
R42 X.n2 X.n1 185
R43 X.n3 X.n2 185
R44 X.n0 X.t3 26.3844
R45 X.n0 X.t2 26.3844
R46 X.n2 X.t0 22.7032
R47 X.n2 X.t1 22.7032
R48 X X.n3 9.78874
R49 X X.n1 8.78481
R50 X.n3 X 8.78481
R51 a_548_110.t0 a_548_110.n1 404.163
R52 a_548_110.n1 a_548_110.t1 312.615
R53 a_548_110.n1 a_548_110.n0 253.126
R54 a_548_110.n0 a_548_110.t2 231.629
R55 a_548_110.n0 a_548_110.t3 175.127
R56 a_503_392.t0 a_503_392.t1 53.1905
R57 a_587_392.t0 a_587_392.t1 70.9205
R58 C_N.n0 C_N.t0 243.742
R59 C_N.n0 C_N.t1 199.559
R60 C_N C_N.n0 157.662
R61 B.t1 B.t0 442.904
R62 B B.t1 322.401
R63 VGND.n6 VGND.n5 242.173
R64 VGND.n14 VGND.n13 231.207
R65 VGND.n4 VGND.n3 215.966
R66 VGND.n11 VGND.n2 206.983
R67 VGND.n3 VGND.t4 57.7602
R68 VGND.n2 VGND.t0 53.438
R69 VGND.n2 VGND.t5 52.6611
R70 VGND.n13 VGND.t7 48.0005
R71 VGND.n5 VGND.t1 46.8755
R72 VGND.n7 VGND.n1 36.1417
R73 VGND.n3 VGND.t2 30.5465
R74 VGND.n12 VGND.n11 28.2358
R75 VGND.n5 VGND.t3 26.2505
R76 VGND.n6 VGND.n4 24.2883
R77 VGND.n14 VGND.n12 24.0946
R78 VGND.n13 VGND.t6 22.2054
R79 VGND.n7 VGND.n6 19.2005
R80 VGND.n11 VGND.n1 9.41227
R81 VGND.n12 VGND.n0 9.3005
R82 VGND.n11 VGND.n10 9.3005
R83 VGND.n9 VGND.n1 9.3005
R84 VGND.n8 VGND.n7 9.3005
R85 VGND.n15 VGND.n14 7.47871
R86 VGND.n8 VGND.n4 0.438054
R87 VGND VGND.n15 0.16068
R88 VGND.n15 VGND.n0 0.14713
R89 VGND.n9 VGND.n8 0.122949
R90 VGND.n10 VGND.n9 0.122949
R91 VGND.n10 VGND.n0 0.122949
R92 VNB.t5 VNB.t0 1697.64
R93 VNB.t0 VNB.t3 1466.67
R94 VNB.t3 VNB.t1 1247.24
R95 VNB.t7 VNB.t6 1189.5
R96 VNB.t4 VNB.t2 1177.95
R97 VNB VNB.t7 1154.86
R98 VNB.t1 VNB.t4 1016.27
R99 VNB.t6 VNB.t5 993.177
R100 D_N.n0 D_N.t0 279.202
R101 D_N D_N.n0 158.847
R102 D_N.n0 D_N.t1 146.117
R103 a_27_424.t1 a_27_424.n1 411.289
R104 a_27_424.n1 a_27_424.t0 318.139
R105 a_27_424.n1 a_27_424.n0 267.759
R106 a_27_424.n0 a_27_424.t2 221.731
R107 a_27_424.n0 a_27_424.t3 190.935
C0 C_N VGND 0.015629f
C1 VPB D_N 0.067953f
C2 VGND VPB 0.011088f
C3 VPWR C_N 0.014793f
C4 A VGND 0.016765f
C5 VPWR VPB 0.139785f
C6 A VPWR 0.02051f
C7 X VGND 0.093068f
C8 X D_N 0.002125f
C9 C_N VPB 0.05639f
C10 A C_N 0.039056f
C11 VPWR X 0.015787f
C12 B VGND 0.14362f
C13 A VPB 0.042558f
C14 B VPWR 0.014953f
C15 X C_N 4.87e-20
C16 X VPB 0.004109f
C17 B C_N 0.003157f
C18 B VPB 0.029463f
C19 B A 0.06868f
C20 VGND D_N 0.010152f
C21 VPWR VGND 0.079507f
C22 VPWR D_N 0.014417f
C23 VGND VNB 0.64081f
C24 C_N VNB 0.192963f
C25 X VNB 0.009228f
C26 VPWR VNB 0.474822f
C27 A VNB 0.096095f
C28 B VNB 0.140466f
C29 D_N VNB 0.154947f
C30 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__or4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4bb_4 VNB VPB VPWR VGND D_N C_N A X B
X0 a_193_277.t5 a_27_94.t2 a_791_392.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X1 a_1060_392.t1 a_678_368.t2 a_791_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X2 VPWR.t2 D_N.t0 a_27_94.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2186 pd=1.52 as=0.295 ps=2.59 w=1 l=0.15
X3 VPWR.t7 a_193_277.t6 X.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2212 pd=1.515 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_1273_392.t2 A.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X5 X.t6 a_193_277.t7 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2186 ps=1.52 w=1.12 l=0.15
X6 a_678_368.t0 C_N.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2102 ps=1.505 w=1 l=0.15
X7 VPWR.t5 a_193_277.t8 X.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.3248 ps=1.7 w=1.12 l=0.15
X8 X.t4 a_193_277.t9 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=1.7 as=0.2212 ps=1.515 w=1.12 l=0.15
X9 VPWR.t0 A.t1 a_1273_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X10 VGND.t7 a_193_277.t10 X.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.24235 ps=1.395 w=0.74 l=0.15
X11 VGND.t0 a_678_368.t3 a_193_277.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.18315 pd=1.235 as=0.53465 ps=2.185 w=0.74 l=0.15
X12 a_1273_392.t0 B.t0 a_1060_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X13 a_678_368.t1 C_N.t1 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1719 pd=1.85 as=0.12945 ps=1.1 w=0.64 l=0.15
X14 a_1060_392.t3 B.t1 a_1273_392.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X15 VGND.t6 a_193_277.t11 X.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.19035 pd=1.37 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 X.t1 a_193_277.t12 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.24235 pd=1.395 as=0.19035 ps=1.37 w=0.74 l=0.15
X17 VGND.t1 D_N.t1 a_27_94.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1485 pd=1.165 as=0.1824 ps=1.85 w=0.64 l=0.15
X18 VGND.t3 A.t2 a_193_277.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.4625 pd=2.73 as=0.17205 ps=1.205 w=0.74 l=0.15
X19 a_791_392.t1 a_678_368.t4 a_1060_392.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X20 a_193_277.t0 B.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.17205 pd=1.205 as=0.18315 ps=1.235 w=0.74 l=0.15
X21 X.t0 a_193_277.t13 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1485 ps=1.165 w=0.74 l=0.15
X22 a_193_277.t3 a_27_94.t3 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.53465 pd=2.185 as=0.327 ps=3.11 w=0.74 l=0.15
X23 a_791_392.t2 a_27_94.t4 a_193_277.t4 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
R0 a_27_94.t0 a_27_94.n2 829.89
R1 a_27_94.t0 a_27_94.n3 735.255
R2 a_27_94.n2 a_27_94.n1 719.862
R3 a_27_94.n0 a_27_94.t4 302.659
R4 a_27_94.n1 a_27_94.t2 295.894
R5 a_27_94.n3 a_27_94.t1 205.857
R6 a_27_94.n0 a_27_94.t3 142.994
R7 a_27_94.n1 a_27_94.n0 69.3409
R8 a_27_94.n3 a_27_94.n2 12.8005
R9 a_791_392.n0 a_791_392.t3 847.016
R10 a_791_392.n0 a_791_392.t1 691.715
R11 a_791_392.n1 a_791_392.n0 585
R12 a_791_392.t0 a_791_392.n1 29.5505
R13 a_791_392.n1 a_791_392.t2 29.5505
R14 a_193_277.n12 a_193_277.n11 585
R15 a_193_277.n1 a_193_277.t7 260.332
R16 a_193_277.n5 a_193_277.t8 257.603
R17 a_193_277.n2 a_193_277.t9 257.603
R18 a_193_277.n0 a_193_277.t6 257.603
R19 a_193_277.n11 a_193_277.n7 172.906
R20 a_193_277.n10 a_193_277.n9 172.578
R21 a_193_277.n6 a_193_277.t10 172.206
R22 a_193_277.n1 a_193_277.t13 159.06
R23 a_193_277.n0 a_193_277.t11 159.06
R24 a_193_277.n3 a_193_277.t12 159.06
R25 a_193_277.n11 a_193_277.n10 157.582
R26 a_193_277.n7 a_193_277.n6 152
R27 a_193_277.n7 a_193_277.n4 84.5208
R28 a_193_277.n2 a_193_277.n0 79.6035
R29 a_193_277.n8 a_193_277.t3 75.0495
R30 a_193_277.n5 a_193_277.n4 66.4552
R31 a_193_277.n8 a_193_277.t2 64.9907
R32 a_193_277.n0 a_193_277.n1 63.5369
R33 a_193_277.n9 a_193_277.t1 52.7032
R34 a_193_277.n12 a_193_277.t4 29.5505
R35 a_193_277.t5 a_193_277.n12 29.5505
R36 a_193_277.n4 a_193_277.n3 27.6489
R37 a_193_277.n9 a_193_277.t0 22.7032
R38 a_193_277.n10 a_193_277.n8 10.6991
R39 a_193_277.n3 a_193_277.n2 5.84292
R40 a_193_277.n6 a_193_277.n5 3.65202
R41 VPB.t5 VPB.t11 515.861
R42 VPB.t3 VPB.t13 515.861
R43 VPB.t7 VPB.t8 372.849
R44 VPB.t0 VPB.t9 280.914
R45 VPB.t10 VPB.t7 278.361
R46 VPB.t8 VPB.t3 273.253
R47 VPB VPB.t0 257.93
R48 VPB.t1 VPB.t6 255.376
R49 VPB.t4 VPB.t5 255.376
R50 VPB.t2 VPB.t1 229.839
R51 VPB.t11 VPB.t2 229.839
R52 VPB.t12 VPB.t4 229.839
R53 VPB.t13 VPB.t12 229.839
R54 VPB.t9 VPB.t10 229.839
R55 a_678_368.t0 a_678_368.n2 887.222
R56 a_678_368.n0 a_678_368.t3 345.726
R57 a_678_368.n2 a_678_368.t1 315.267
R58 a_678_368.n1 a_678_368.t2 295.293
R59 a_678_368.n0 a_678_368.t4 263.762
R60 a_678_368.n2 a_678_368.n1 98.3116
R61 a_678_368.n1 a_678_368.n0 34.7778
R62 a_1060_392.n1 a_1060_392.n0 678.899
R63 a_1060_392.t1 a_1060_392.n1 39.4005
R64 a_1060_392.n0 a_1060_392.t2 29.5505
R65 a_1060_392.n0 a_1060_392.t3 29.5505
R66 a_1060_392.n1 a_1060_392.t0 29.5505
R67 D_N.n0 D_N.t0 230.919
R68 D_N.n0 D_N.t1 203.339
R69 D_N D_N.n0 154.03
R70 VPWR.n7 VPWR.n6 604.976
R71 VPWR.n14 VPWR.n1 604.107
R72 VPWR.n12 VPWR.n3 600.511
R73 VPWR.n8 VPWR.n5 322.005
R74 VPWR.n1 VPWR.t2 47.2805
R75 VPWR.n6 VPWR.t1 46.2955
R76 VPWR.n5 VPWR.t0 39.4005
R77 VPWR.n11 VPWR.n4 36.1417
R78 VPWR.n3 VPWR.t4 35.1791
R79 VPWR.n3 VPWR.t7 34.2996
R80 VPWR.n5 VPWR.t3 29.5505
R81 VPWR.n1 VPWR.t6 28.5142
R82 VPWR.n13 VPWR.n12 27.4829
R83 VPWR.n6 VPWR.t5 27.0196
R84 VPWR.n14 VPWR.n13 15.4358
R85 VPWR.n7 VPWR.n4 15.0593
R86 VPWR.n12 VPWR.n11 12.8005
R87 VPWR.n9 VPWR.n4 9.3005
R88 VPWR.n11 VPWR.n10 9.3005
R89 VPWR.n12 VPWR.n2 9.3005
R90 VPWR.n13 VPWR.n0 9.3005
R91 VPWR.n15 VPWR.n14 7.53404
R92 VPWR.n8 VPWR.n7 7.52486
R93 VPWR VPWR.n15 0.161409
R94 VPWR.n9 VPWR.n8 0.151452
R95 VPWR.n15 VPWR.n0 0.146411
R96 VPWR.n10 VPWR.n9 0.122949
R97 VPWR.n10 VPWR.n2 0.122949
R98 VPWR.n2 VPWR.n0 0.122949
R99 X.n2 X.n0 654.163
R100 X.n2 X.n1 585
R101 X.n5 X.n4 146.976
R102 X.n5 X.n3 91.112
R103 X.n0 X.t5 68.5987
R104 X.n4 X.t3 49.9505
R105 X.n4 X.t1 47.9644
R106 X.n0 X.t4 33.4201
R107 X.n1 X.t7 26.3844
R108 X.n1 X.t6 26.3844
R109 X.n3 X.t2 22.7032
R110 X.n3 X.t0 22.7032
R111 X X.n5 14.9485
R112 X X.n2 2.45529
R113 A.n1 A.t0 274.473
R114 A.n3 A.t1 274.473
R115 A.n1 A 188.227
R116 A.n3 A.t2 160.814
R117 A A.n4 157.017
R118 A.n2 A.n0 152
R119 A.n4 A.n2 49.6611
R120 A.n2 A.n1 15.3369
R121 A A.n0 9.85996
R122 A.n4 A.n3 8.03383
R123 A A.n0 6.74645
R124 a_1273_392.n1 a_1273_392.t3 692.458
R125 a_1273_392.t2 a_1273_392.n1 279.692
R126 a_1273_392.n1 a_1273_392.n0 189.115
R127 a_1273_392.n0 a_1273_392.t1 29.5505
R128 a_1273_392.n0 a_1273_392.t0 29.5505
R129 C_N.n0 C_N.t0 224.097
R130 C_N.n0 C_N.t1 196.516
R131 C_N C_N.n0 154.447
R132 VGND.n17 VGND.t9 251.048
R133 VGND.n22 VGND.n5 206.333
R134 VGND.n2 VGND.n1 203.621
R135 VGND.n30 VGND.n29 122.329
R136 VGND.n10 VGND.n9 114.883
R137 VGND.n8 VGND.t3 81.2404
R138 VGND.n9 VGND.t2 46.2167
R139 VGND.n5 VGND.t8 41.2505
R140 VGND.n29 VGND.t1 39.3755
R141 VGND.n29 VGND.t4 36.7236
R142 VGND.n11 VGND.n7 36.1417
R143 VGND.n15 VGND.n7 36.1417
R144 VGND.n24 VGND.n23 36.1417
R145 VGND.n1 VGND.t5 35.6762
R146 VGND.n1 VGND.t6 35.6762
R147 VGND.n9 VGND.t0 34.0546
R148 VGND.n16 VGND.n15 33.9171
R149 VGND.n11 VGND.n10 33.8829
R150 VGND.n28 VGND.n27 33.6699
R151 VGND.n18 VGND.n4 32.9284
R152 VGND.n22 VGND.n4 24.4711
R153 VGND.n23 VGND.n22 22.9652
R154 VGND.n30 VGND.n28 21.4593
R155 VGND.n5 VGND.t7 21.3263
R156 VGND.n24 VGND.n2 19.326
R157 VGND.n12 VGND.n11 9.3005
R158 VGND.n13 VGND.n7 9.3005
R159 VGND.n15 VGND.n14 9.3005
R160 VGND.n16 VGND.n6 9.3005
R161 VGND.n19 VGND.n18 9.3005
R162 VGND.n20 VGND.n4 9.3005
R163 VGND.n22 VGND.n21 9.3005
R164 VGND.n23 VGND.n3 9.3005
R165 VGND.n25 VGND.n24 9.3005
R166 VGND.n27 VGND.n26 9.3005
R167 VGND.n28 VGND.n0 9.3005
R168 VGND.n31 VGND.n30 7.43488
R169 VGND.n17 VGND.n16 6.46515
R170 VGND.n10 VGND.n8 6.33154
R171 VGND.n18 VGND.n17 5.94797
R172 VGND.n27 VGND.n2 2.97424
R173 VGND.n12 VGND.n8 0.267709
R174 VGND VGND.n31 0.160103
R175 VGND.n31 VGND.n0 0.1477
R176 VGND.n13 VGND.n12 0.122949
R177 VGND.n14 VGND.n13 0.122949
R178 VGND.n14 VGND.n6 0.122949
R179 VGND.n19 VGND.n6 0.122949
R180 VGND.n20 VGND.n19 0.122949
R181 VGND.n21 VGND.n20 0.122949
R182 VGND.n21 VGND.n3 0.122949
R183 VGND.n25 VGND.n3 0.122949
R184 VGND.n26 VGND.n25 0.122949
R185 VGND.n26 VGND.n0 0.122949
R186 VNB.t9 VNB.t0 3683.99
R187 VNB.t8 VNB.t9 3071.92
R188 VNB.t5 VNB.t7 1859.32
R189 VNB.t0 VNB.t2 1489.76
R190 VNB.t2 VNB.t3 1420.47
R191 VNB.t6 VNB.t5 1362.73
R192 VNB.t1 VNB.t4 1328.08
R193 VNB.t7 VNB.t8 1177.95
R194 VNB VNB.t1 1143.31
R195 VNB.t4 VNB.t6 993.177
R196 B.n0 B.t0 243.556
R197 B.n0 B.t2 228.148
R198 B.n1 B.t1 223.839
R199 B.n2 B.n1 152
R200 B.n1 B.n0 24.1005
R201 B.n2 B 16.0975
R202 B B.n2 2.52171
C0 VPB A 0.09572f
C1 D_N VPWR 0.015199f
C2 VPB X 0.003047f
C3 A VGND 0.093375f
C4 X VGND 0.253562f
C5 X C_N 4.47e-19
C6 VPB B 0.083125f
C7 VPB VPWR 0.222749f
C8 B VGND 0.0162f
C9 VPWR VGND 0.13926f
C10 VPWR C_N 0.012386f
C11 VPB D_N 0.041188f
C12 D_N VGND 0.038093f
C13 B A 0.061451f
C14 D_N C_N 0.001302f
C15 VPWR A 0.035455f
C16 VPWR X 0.04773f
C17 VPB VGND 0.014676f
C18 VPB C_N 0.051333f
C19 D_N X 0.031231f
C20 VPWR B 0.011465f
C21 C_N VGND 0.014663f
C22 VGND VNB 1.04412f
C23 A VNB 0.265209f
C24 B VNB 0.167137f
C25 C_N VNB 0.128822f
C26 X VNB 0.013675f
C27 VPWR VNB 0.794987f
C28 D_N VNB 0.140054f
C29 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfbbn_1 VNB VPB VPWR SET_B VGND D SCE SCD Q_N CLK_N RESET_B
+ Q
X0 a_212_464.t0 SCE.t0 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1056 ps=0.97 w=0.64 l=0.15
X1 a_1876_119.t1 a_977_243.t3 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.066 pd=0.79 as=0.11275 ps=0.96 w=0.55 l=0.15
X2 a_2392_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.17705 ps=1.38 w=0.74 l=0.15
X3 a_2133_410.t0 a_1954_119.t4 a_2509_392.t1 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X4 a_1081_497# a_977_243.t4 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.1239 ps=1.43 w=0.42 l=0.15
X5 a_977_243.t2 SET_B.t0 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=2.26 as=0.126 ps=1.14 w=0.84 l=0.15
X6 a_977_243.t0 a_1159_497.t2 a_1434_78.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1045 pd=0.93 as=0.2602 ps=2.24 w=0.55 l=0.15
X7 VGND.t5 RESET_B.t0 a_1579_258.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1828 pd=1.34 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 Q_N.t0 a_2133_410.t3 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1828 ps=1.34 w=0.74 l=0.15
X9 VPWR.t7 a_1579_258.t2 a_1528_424.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1134 ps=1.11 w=0.84 l=0.15
X10 a_119_119.t1 SCD.t0 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X11 a_2509_392.t0 a_1579_258.t3 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.269075 ps=1.705 w=1 l=0.15
X12 a_2133_410.t2 a_1579_258.t4 a_2392_74# VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1406 pd=1.12 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VGND.t2 SET_B.t1 a_1434_78.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.11275 pd=0.96 as=0.125125 ps=1.005 w=0.55 l=0.15
X14 a_1528_424.t1 a_1159_497.t3 a_977_243.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.3906 ps=2.61 w=0.84 l=0.15
X15 VPWR.t3 SET_B.t2 a_2133_410.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.269075 pd=1.705 as=0.295 ps=2.59 w=1 l=0.15
X16 Q.t0 a_3078_384.t2 VPWR.t14 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.203 ps=1.505 w=1.12 l=0.15
X17 VPWR.t9 SCD.t1 a_27_464.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1888 ps=1.87 w=0.64 l=0.15
X18 a_353_93.t0 SCE.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1449 ps=1.11 w=0.42 l=0.15
X19 a_353_93.t1 SCE.t2 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1888 ps=1.87 w=0.64 l=0.15
X20 VPWR.t6 RESET_B.t1 a_1579_258.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2748 pd=1.78 as=0.3625 ps=3.71 w=0.64 l=0.15
X21 VPWR.t13 a_2133_410.t4 a_3078_384.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X22 a_1954_119.t3 a_867_82.t2 a_1903_424.t0 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.1008 ps=1.08 w=0.84 l=0.15
X23 a_197_119.t0 a_867_82.t3 a_1159_497.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 VGND.t9 a_353_93.t2 a_305_119.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1449 pd=1.11 as=0.0504 ps=0.66 w=0.42 l=0.15
X25 a_197_119.t1 SCE.t3 a_119_119.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 VPWR.t0 a_2133_410.t5 a_2088_508.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.22775 pd=2.07 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 a_197_119.t4 a_662_82.t2 a_1159_497.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2208 pd=1.97 as=0.1133 ps=1.025 w=0.64 l=0.15
X28 a_305_119.t0 D.t0 a_197_119.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X29 a_2164_119.t0 a_867_82.t4 a_1954_119.t2 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.24035 ps=1.45 w=0.42 l=0.15
X30 VGND.t4 CLK_N.t0 a_662_82.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.19615 pd=1.41 as=0.2109 ps=2.05 w=0.74 l=0.15
X31 a_867_82.t1 a_662_82.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X32 a_1954_119.t0 a_662_82.t4 a_1876_119.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.24035 pd=1.45 as=0.066 ps=0.79 w=0.55 l=0.15
X33 a_27_464.t0 a_353_93.t3 a_197_119.t5 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1856 pd=1.86 as=0.096 ps=0.94 w=0.64 l=0.15
X34 VPWR.t12 CLK_N.t1 a_662_82.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X35 a_2088_508.t1 a_662_82.t5 a_1954_119.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.1428 ps=1.225 w=0.42 l=0.15
X36 a_197_119.t2 D.t1 a_212_464.t1 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X37 Q_N.t1 a_2133_410.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2748 ps=1.78 w=1.12 l=0.15
X38 VGND.t0 a_2133_410.t7 a_3078_384.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X39 a_867_82.t0 a_662_82.t6 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3219 pd=2.35 as=0.19615 ps=1.41 w=0.74 l=0.15
R0 SCE.t3 SCE.t1 922.227
R1 SCE.t1 SCE.t2 729.428
R2 SCE.n0 SCE.t0 271.394
R3 SCE.n0 SCE.t3 174.197
R4 SCE SCE.n0 67.4187
R5 VPWR.n35 VPWR.t0 759.761
R6 VPWR.n56 VPWR.t11 687.87
R7 VPWR.n15 VPWR.n14 649.534
R8 VPWR.n44 VPWR.n43 617.378
R9 VPWR.n23 VPWR.n22 585
R10 VPWR.n21 VPWR.n20 585
R11 VPWR.n63 VPWR.t5 381.726
R12 VPWR.n5 VPWR.n4 323.406
R13 VPWR.n69 VPWR.n1 315.932
R14 VPWR.n19 VPWR.n18 242.351
R15 VPWR.n22 VPWR.n21 110.812
R16 VPWR.n1 VPWR.t4 55.4067
R17 VPWR.n18 VPWR.t13 55.1136
R18 VPWR.n14 VPWR.t8 46.2955
R19 VPWR.n14 VPWR.t3 46.2955
R20 VPWR.n22 VPWR.t6 46.1724
R21 VPWR.n1 VPWR.t9 46.1724
R22 VPWR.n67 VPWR.n2 36.1417
R23 VPWR.n68 VPWR.n67 36.1417
R24 VPWR.n62 VPWR.n61 36.1417
R25 VPWR.n45 VPWR.n42 36.1417
R26 VPWR.n49 VPWR.n9 36.1417
R27 VPWR.n50 VPWR.n49 36.1417
R28 VPWR.n51 VPWR.n50 36.1417
R29 VPWR.n51 VPWR.n7 36.1417
R30 VPWR.n55 VPWR.n7 36.1417
R31 VPWR.n36 VPWR.n12 36.1417
R32 VPWR.n40 VPWR.n12 36.1417
R33 VPWR.n34 VPWR.n33 36.1417
R34 VPWR.n28 VPWR.n17 36.1417
R35 VPWR.n29 VPWR.n28 36.1417
R36 VPWR.n43 VPWR.t10 35.1791
R37 VPWR.n43 VPWR.t7 35.1791
R38 VPWR.n57 VPWR.n56 34.6358
R39 VPWR.n41 VPWR.n40 34.6358
R40 VPWR.n30 VPWR.n29 32.1866
R41 VPWR.n63 VPWR.n62 30.1181
R42 VPWR.n57 VPWR.n5 28.6123
R43 VPWR.n21 VPWR.t1 28.3632
R44 VPWR.n18 VPWR.t14 28.0072
R45 VPWR.n24 VPWR.n17 26.4622
R46 VPWR.n4 VPWR.t2 26.3844
R47 VPWR.n4 VPWR.t12 26.3844
R48 VPWR.n61 VPWR.n5 24.8476
R49 VPWR.n63 VPWR.n2 23.3417
R50 VPWR.n69 VPWR.n68 22.9652
R51 VPWR.n33 VPWR.n15 22.4407
R52 VPWR.n44 VPWR.n9 21.8358
R53 VPWR.n56 VPWR.n55 18.824
R54 VPWR.n45 VPWR.n44 14.3064
R55 VPWR.n42 VPWR.n41 12.8005
R56 VPWR.n36 VPWR.n35 12.276
R57 VPWR.n25 VPWR.n24 9.3005
R58 VPWR.n26 VPWR.n17 9.3005
R59 VPWR.n28 VPWR.n27 9.3005
R60 VPWR.n29 VPWR.n16 9.3005
R61 VPWR.n31 VPWR.n30 9.3005
R62 VPWR.n33 VPWR.n32 9.3005
R63 VPWR.n34 VPWR.n13 9.3005
R64 VPWR.n37 VPWR.n36 9.3005
R65 VPWR.n38 VPWR.n12 9.3005
R66 VPWR.n40 VPWR.n39 9.3005
R67 VPWR.n41 VPWR.n11 9.3005
R68 VPWR.n42 VPWR.n10 9.3005
R69 VPWR.n46 VPWR.n45 9.3005
R70 VPWR.n47 VPWR.n9 9.3005
R71 VPWR.n49 VPWR.n48 9.3005
R72 VPWR.n50 VPWR.n8 9.3005
R73 VPWR.n52 VPWR.n51 9.3005
R74 VPWR.n53 VPWR.n7 9.3005
R75 VPWR.n55 VPWR.n54 9.3005
R76 VPWR.n56 VPWR.n6 9.3005
R77 VPWR.n58 VPWR.n57 9.3005
R78 VPWR.n59 VPWR.n5 9.3005
R79 VPWR.n61 VPWR.n60 9.3005
R80 VPWR.n62 VPWR.n3 9.3005
R81 VPWR.n64 VPWR.n63 9.3005
R82 VPWR.n65 VPWR.n2 9.3005
R83 VPWR.n67 VPWR.n66 9.3005
R84 VPWR.n68 VPWR.n0 9.3005
R85 VPWR.n20 VPWR.n19 9.19461
R86 VPWR.n35 VPWR.n34 8.51127
R87 VPWR.n70 VPWR.n69 7.27223
R88 VPWR.n23 VPWR.n20 5.32767
R89 VPWR.n30 VPWR.n15 2.30162
R90 VPWR.n25 VPWR.n19 0.208615
R91 VPWR VPWR.n70 0.157962
R92 VPWR.n70 VPWR.n0 0.149814
R93 VPWR.n26 VPWR.n25 0.122949
R94 VPWR.n27 VPWR.n26 0.122949
R95 VPWR.n27 VPWR.n16 0.122949
R96 VPWR.n31 VPWR.n16 0.122949
R97 VPWR.n32 VPWR.n31 0.122949
R98 VPWR.n32 VPWR.n13 0.122949
R99 VPWR.n37 VPWR.n13 0.122949
R100 VPWR.n38 VPWR.n37 0.122949
R101 VPWR.n39 VPWR.n38 0.122949
R102 VPWR.n39 VPWR.n11 0.122949
R103 VPWR.n11 VPWR.n10 0.122949
R104 VPWR.n46 VPWR.n10 0.122949
R105 VPWR.n47 VPWR.n46 0.122949
R106 VPWR.n48 VPWR.n47 0.122949
R107 VPWR.n48 VPWR.n8 0.122949
R108 VPWR.n52 VPWR.n8 0.122949
R109 VPWR.n53 VPWR.n52 0.122949
R110 VPWR.n54 VPWR.n53 0.122949
R111 VPWR.n54 VPWR.n6 0.122949
R112 VPWR.n58 VPWR.n6 0.122949
R113 VPWR.n59 VPWR.n58 0.122949
R114 VPWR.n60 VPWR.n59 0.122949
R115 VPWR.n60 VPWR.n3 0.122949
R116 VPWR.n64 VPWR.n3 0.122949
R117 VPWR.n65 VPWR.n64 0.122949
R118 VPWR.n66 VPWR.n65 0.122949
R119 VPWR.n66 VPWR.n0 0.122949
R120 VPWR.n24 VPWR.n23 0.0744884
R121 a_212_464.t0 a_212_464.t1 83.1099
R122 VPB.n0 VPB 7814.52
R123 VPB VPB.n1 6471.57
R124 VPB.t20 VPB.t14 712.5
R125 VPB.t11 VPB.t2 669.087
R126 VPB.t5 VPB.t0 559.274
R127 VPB.t15 VPB.t3 515.861
R128 VPB.t16 VPB.t6 515.861
R129 VPB.t6 VPB.t13 513.307
R130 VPB.t2 VPB.t15 472.447
R131 VPB.t8 VPB.t1 390.61
R132 VPB.t10 VPB.t5 316.668
R133 VPB.t17 VPB.t21 273.253
R134 VPB.t4 VPB.t20 273.253
R135 VPB.n1 VPB.t19 270.7
R136 VPB.t1 VPB.n0 265.228
R137 VPB.t12 VPB 257.93
R138 VPB.n1 VPB.t8 250.762
R139 VPB.t7 VPB.t12 245.161
R140 VPB.n0 VPB.t17 234.946
R141 VPB.t14 VPB.t9 229.839
R142 VPB.t3 VPB.t16 229.839
R143 VPB.t13 VPB.t18 229.839
R144 VPB.t19 VPB.t10 214.517
R145 VPB.t9 VPB.t11 214.517
R146 VPB.t18 VPB.t7 214.517
R147 VPB.t0 VPB.t4 199.195
R148 a_977_243.t1 a_977_243.n6 686.678
R149 a_977_243.n5 a_977_243.n4 543.199
R150 a_977_243.n6 a_977_243.n5 345.432
R151 a_977_243.n3 a_977_243.t0 338.704
R152 a_977_243.n2 a_977_243.t2 333.947
R153 a_977_243.n1 a_977_243.t3 268.313
R154 a_977_243.n2 a_977_243.n1 206.55
R155 a_977_243.n1 a_977_243.n0 205.922
R156 a_977_243.n5 a_977_243.t4 163.637
R157 a_977_243.n3 a_977_243.n2 48.9417
R158 a_977_243.n6 a_977_243.n3 43.5205
R159 VGND.n65 VGND.t6 256.224
R160 VGND.n51 VGND.n50 220.173
R161 VGND.n36 VGND.n10 217.776
R162 VGND.n59 VGND.n58 214.868
R163 VGND.n18 VGND.n17 206.636
R164 VGND.n16 VGND.t0 177.649
R165 VGND.n58 VGND.t3 157.143
R166 VGND.n17 VGND.t5 120.811
R167 VGND.n10 VGND.t8 58.9096
R168 VGND.n58 VGND.t9 40.0005
R169 VGND.n20 VGND.n19 36.1417
R170 VGND.n20 VGND.n14 36.1417
R171 VGND.n24 VGND.n14 36.1417
R172 VGND.n25 VGND.n24 36.1417
R173 VGND.n26 VGND.n25 36.1417
R174 VGND.n30 VGND.n12 36.1417
R175 VGND.n31 VGND.n30 36.1417
R176 VGND.n32 VGND.n31 36.1417
R177 VGND.n32 VGND.n9 36.1417
R178 VGND.n38 VGND.n37 36.1417
R179 VGND.n38 VGND.n7 36.1417
R180 VGND.n42 VGND.n7 36.1417
R181 VGND.n43 VGND.n42 36.1417
R182 VGND.n44 VGND.n43 36.1417
R183 VGND.n49 VGND.n48 36.1417
R184 VGND.n56 VGND.n3 36.1417
R185 VGND.n57 VGND.n56 36.1417
R186 VGND.n63 VGND.n1 36.1417
R187 VGND.n64 VGND.n63 36.1417
R188 VGND.n50 VGND.t1 35.6762
R189 VGND.n50 VGND.t4 35.6762
R190 VGND.n52 VGND.n49 33.6699
R191 VGND.n59 VGND.n57 31.624
R192 VGND.n10 VGND.t2 30.546
R193 VGND.n37 VGND.n36 29.7417
R194 VGND.n17 VGND.t7 28.3794
R195 VGND.n44 VGND.n5 27.8593
R196 VGND.n48 VGND.n5 19.577
R197 VGND.n26 VGND.n12 19.3336
R198 VGND.n51 VGND.n3 19.326
R199 VGND.n19 VGND.n18 19.2005
R200 VGND.n65 VGND.n64 18.824
R201 VGND.n36 VGND.n9 17.6946
R202 VGND.n59 VGND.n1 15.8123
R203 VGND.n66 VGND.n65 9.3005
R204 VGND.n19 VGND.n15 9.3005
R205 VGND.n21 VGND.n20 9.3005
R206 VGND.n22 VGND.n14 9.3005
R207 VGND.n24 VGND.n23 9.3005
R208 VGND.n25 VGND.n13 9.3005
R209 VGND.n27 VGND.n26 9.3005
R210 VGND.n28 VGND.n12 9.3005
R211 VGND.n30 VGND.n29 9.3005
R212 VGND.n31 VGND.n11 9.3005
R213 VGND.n33 VGND.n32 9.3005
R214 VGND.n34 VGND.n9 9.3005
R215 VGND.n36 VGND.n35 9.3005
R216 VGND.n37 VGND.n8 9.3005
R217 VGND.n39 VGND.n38 9.3005
R218 VGND.n40 VGND.n7 9.3005
R219 VGND.n42 VGND.n41 9.3005
R220 VGND.n43 VGND.n6 9.3005
R221 VGND.n45 VGND.n44 9.3005
R222 VGND.n46 VGND.n5 9.3005
R223 VGND.n48 VGND.n47 9.3005
R224 VGND.n49 VGND.n4 9.3005
R225 VGND.n53 VGND.n52 9.3005
R226 VGND.n54 VGND.n3 9.3005
R227 VGND.n56 VGND.n55 9.3005
R228 VGND.n57 VGND.n2 9.3005
R229 VGND.n60 VGND.n59 9.3005
R230 VGND.n61 VGND.n1 9.3005
R231 VGND.n63 VGND.n62 9.3005
R232 VGND.n64 VGND.n0 9.3005
R233 VGND.n18 VGND.n16 7.33086
R234 VGND.n52 VGND.n51 2.97424
R235 VGND.n16 VGND.n15 0.216247
R236 VGND.n21 VGND.n15 0.122949
R237 VGND.n22 VGND.n21 0.122949
R238 VGND.n23 VGND.n22 0.122949
R239 VGND.n23 VGND.n13 0.122949
R240 VGND.n27 VGND.n13 0.122949
R241 VGND.n28 VGND.n27 0.122949
R242 VGND.n29 VGND.n28 0.122949
R243 VGND.n29 VGND.n11 0.122949
R244 VGND.n33 VGND.n11 0.122949
R245 VGND.n34 VGND.n33 0.122949
R246 VGND.n35 VGND.n34 0.122949
R247 VGND.n35 VGND.n8 0.122949
R248 VGND.n39 VGND.n8 0.122949
R249 VGND.n40 VGND.n39 0.122949
R250 VGND.n41 VGND.n40 0.122949
R251 VGND.n41 VGND.n6 0.122949
R252 VGND.n45 VGND.n6 0.122949
R253 VGND.n46 VGND.n45 0.122949
R254 VGND.n47 VGND.n46 0.122949
R255 VGND.n47 VGND.n4 0.122949
R256 VGND.n53 VGND.n4 0.122949
R257 VGND.n54 VGND.n53 0.122949
R258 VGND.n55 VGND.n54 0.122949
R259 VGND.n55 VGND.n2 0.122949
R260 VGND.n60 VGND.n2 0.122949
R261 VGND.n61 VGND.n60 0.122949
R262 VGND.n62 VGND.n61 0.122949
R263 VGND.n62 VGND.n0 0.122949
R264 VGND.n66 VGND.n0 0.122949
R265 VGND VGND.n66 0.0617245
R266 a_1876_119.t0 a_1876_119.t1 52.3641
R267 VNB VNB.n0 32895.8
R268 VNB.t10 VNB.t2 5104.46
R269 VNB.t16 VNB.t11 3626.25
R270 VNB.t9 VNB.t10 2633.07
R271 VNB.t3 VNB.t9 2621.52
R272 VNB.n0 VNB.t16 2552.23
R273 VNB.t12 VNB.t0 2426.74
R274 VNB.t11 VNB.t1 2425.2
R275 VNB.t6 VNB.t5 2286.61
R276 VNB.t5 VNB.t15 1940.16
R277 VNB.t7 VNB.t12 1838.44
R278 VNB.n0 VNB.t7 1507.52
R279 VNB.t2 VNB.t6 1362.73
R280 VNB.t13 VNB.t3 1293.44
R281 VNB.t14 VNB.t4 1247.24
R282 VNB.t8 VNB 1201.05
R283 VNB.t1 VNB.t13 900.788
R284 VNB.t15 VNB.t14 900.788
R285 VNB.t4 VNB.t8 900.788
R286 SET_B.n2 SET_B.t1 268.313
R287 SET_B.n1 SET_B.n0 258.673
R288 SET_B.n2 SET_B.t0 252.345
R289 SET_B.n1 SET_B.t2 231.629
R290 SET_B SET_B.n2 193.344
R291 SET_B SET_B.n1 176.862
R292 a_1954_119.t3 a_1954_119.n3 434.173
R293 a_1954_119.n3 a_1954_119.n1 296.832
R294 a_1954_119.n1 a_1954_119.n0 241.147
R295 a_1954_119.n1 a_1954_119.t4 207.529
R296 a_1954_119.n3 a_1954_119.n2 179.239
R297 a_1954_119.t3 a_1954_119.t1 111.264
R298 a_1954_119.n2 a_1954_119.t2 104.082
R299 a_1954_119.n2 a_1954_119.t0 75.2845
R300 a_2509_392.t0 a_2509_392.t1 53.1905
R301 a_2133_410.t0 a_2133_410.n3 825.947
R302 a_2133_410.n2 a_2133_410.t1 815.39
R303 a_2133_410.t0 a_2133_410.n8 744.648
R304 a_2133_410.n1 a_2133_410.n0 506.392
R305 a_2133_410.n7 a_2133_410.t2 443.003
R306 a_2133_410.n6 a_2133_410.t6 264.298
R307 a_2133_410.n4 a_2133_410.t4 232.7
R308 a_2133_410.n4 a_2133_410.t7 213.151
R309 a_2133_410.n2 a_2133_410.n1 212.44
R310 a_2133_410.n5 a_2133_410.t3 199.666
R311 a_2133_410.n7 a_2133_410.n6 152
R312 a_2133_410.n8 a_2133_410.n7 151.18
R313 a_2133_410.n5 a_2133_410.n4 147.279
R314 a_2133_410.n1 a_2133_410.t5 138.441
R315 a_2133_410.n3 a_2133_410.n2 93.376
R316 a_2133_410.n8 a_2133_410.n3 16.2914
R317 a_2133_410.n6 a_2133_410.n5 4.38232
R318 a_1159_497.n2 a_1159_497.n1 682.091
R319 a_1159_497.n0 a_1159_497.t3 347.652
R320 a_1159_497.n1 a_1159_497.t1 296.543
R321 a_1159_497.n1 a_1159_497.n0 169.002
R322 a_1159_497.n0 a_1159_497.t2 140.929
R323 a_1159_497.n3 a_1159_497.n2 73.4581
R324 a_1159_497.n2 a_1159_497.t0 34.2614
R325 a_1434_78.t0 a_1434_78.t1 624.962
R326 RESET_B.n0 RESET_B.t1 423.163
R327 RESET_B RESET_B.n0 159.345
R328 RESET_B.n0 RESET_B.t0 121.109
R329 a_1579_258.t1 a_1579_258.n4 1395.21
R330 a_1579_258.n3 a_1579_258.n1 536.135
R331 a_1579_258.n2 a_1579_258.t3 296.747
R332 a_1579_258.n1 a_1579_258.t2 287.731
R333 a_1579_258.n4 a_1579_258.t0 251.73
R334 a_1579_258.n2 a_1579_258.t4 178.34
R335 a_1579_258.n3 a_1579_258.n2 152
R336 a_1579_258.n1 a_1579_258.n0 149.826
R337 a_1579_258.n4 a_1579_258.n3 92.7467
R338 Q_N.n1 Q_N 589.157
R339 Q_N.n1 Q_N.n0 585
R340 Q_N.n2 Q_N.n1 585
R341 Q_N Q_N.t0 205.9
R342 Q_N.n1 Q_N.t1 26.3844
R343 Q_N Q_N.n2 11.1382
R344 Q_N Q_N.n0 9.64206
R345 Q_N Q_N.n0 2.66024
R346 Q_N.n2 Q_N 1.16414
R347 a_1528_424.t0 a_1528_424.t1 63.3219
R348 SCD.n0 SCD.t1 266.25
R349 SCD.n0 SCD.t0 169.072
R350 SCD SCD.n0 68.9655
R351 a_119_119.t0 a_119_119.t1 68.5719
R352 a_662_82.n1 a_662_82.t4 1372.09
R353 a_662_82.t4 a_662_82.t5 752.723
R354 a_662_82.t6 a_662_82.n1 740.673
R355 a_662_82.n0 a_662_82.t2 562.255
R356 a_662_82.n3 a_662_82.t0 327.75
R357 a_662_82.t1 a_662_82.n3 285.207
R358 a_662_82.n2 a_662_82.t3 253.587
R359 a_662_82.n2 a_662_82.t6 204.048
R360 a_662_82.n1 a_662_82.n0 176.733
R361 a_662_82.n3 a_662_82.n2 152
R362 a_3078_384.t1 a_3078_384.n2 417.993
R363 a_3078_384.n1 a_3078_384.t2 285.719
R364 a_3078_384.n2 a_3078_384.t0 242.31
R365 a_3078_384.n1 a_3078_384.n0 178.34
R366 a_3078_384.n2 a_3078_384.n1 176.825
R367 Q.n1 Q 589.444
R368 Q.n1 Q.n0 585
R369 Q.n2 Q.n1 585
R370 Q.n1 Q.t0 26.3844
R371 Q Q.n2 11.9116
R372 Q Q.n0 10.3116
R373 Q Q.n0 2.84494
R374 Q.n2 Q 1.24494
R375 a_27_464.t0 a_27_464.t1 898.692
R376 a_353_93.t1 a_353_93.n1 400.618
R377 a_353_93.n0 a_353_93.t3 295.627
R378 a_353_93.n0 a_353_93.t2 261.887
R379 a_353_93.n1 a_353_93.t0 254.635
R380 a_353_93.n1 a_353_93.n0 231.603
R381 a_867_82.n1 a_867_82.t3 434.137
R382 a_867_82.n1 a_867_82.n0 399.779
R383 a_867_82.n2 a_867_82.t2 367.358
R384 a_867_82.n2 a_867_82.t4 360.327
R385 a_867_82.n4 a_867_82.t0 284.536
R386 a_867_82.t1 a_867_82.n4 248.799
R387 a_867_82.n4 a_867_82.n3 50.4529
R388 a_867_82.n3 a_867_82.n2 22.3563
R389 a_867_82.n3 a_867_82.n1 2.52444
R390 a_197_119.n0 a_197_119.t4 862.105
R391 a_197_119.n3 a_197_119.n2 690.88
R392 a_197_119.n2 a_197_119.n0 515.686
R393 a_197_119.n2 a_197_119.n1 256.228
R394 a_197_119.n0 a_197_119.t0 246.429
R395 a_197_119.n1 a_197_119.t3 71.4291
R396 a_197_119.n3 a_197_119.t5 46.1724
R397 a_197_119.t2 a_197_119.n3 46.1724
R398 a_197_119.n1 a_197_119.t1 40.0005
R399 a_305_119.t0 a_305_119.t1 68.5719
R400 a_2088_508.t0 a_2088_508.t1 112.572
R401 D.n0 D.t1 279.83
R402 D.n0 D.t0 233.821
R403 D D.n0 154.522
R404 CLK_N.n0 CLK_N.t1 243.038
R405 CLK_N.n0 CLK_N.t0 199.392
R406 CLK_N CLK_N.n0 155.572
C0 D VPWR 0.006812f
C1 SET_B RESET_B 4.28e-19
C2 SCD SET_B 1.22e-20
C3 SCE CLK_N 0.043834f
C4 SCE SET_B 7.12e-20
C5 VPB VGND 0.028242f
C6 VGND a_2392_74# 0.164929f
C7 D SET_B 2.42e-20
C8 SCD SCE 0.146879f
C9 VPB VPWR 0.48333f
C10 VPB Q_N 0.018358f
C11 VPWR VGND 0.16365f
C12 VGND Q_N 0.070651f
C13 VPWR a_2392_74# 0.002163f
C14 VPWR Q_N 0.086288f
C15 VPB Q 0.014843f
C16 VGND Q 0.099051f
C17 VPB CLK_N 0.044092f
C18 VGND CLK_N 0.010022f
C19 SCE D 0.147216f
C20 VPWR Q 0.123984f
C21 VPB SET_B 0.165119f
C22 VPWR CLK_N 0.019917f
C23 VGND SET_B 0.069211f
C24 a_2392_74# SET_B 0.008212f
C25 VPWR a_1081_497# 0.001237f
C26 VPWR SET_B 0.163249f
C27 VPB RESET_B 0.130737f
C28 VGND RESET_B 0.007965f
C29 Q_N SET_B 1.99e-19
C30 a_2392_74# RESET_B 2.24e-19
C31 SCD VPB 0.075623f
C32 SCD VGND 0.048989f
C33 VPWR RESET_B 0.021231f
C34 Q_N RESET_B 0.002259f
C35 Q SET_B 6.36e-20
C36 SCD VPWR 0.019291f
C37 SCE VPB 0.166463f
C38 SCE VGND 0.085604f
C39 CLK_N SET_B 1.46e-20
C40 Q RESET_B 2.99e-19
C41 VGND a_1151_119# 0.001241f
C42 SCE VPWR 0.034375f
C43 D VPB 0.069028f
C44 D VGND 0.008699f
C45 Q VNB 0.113871f
C46 Q_N VNB 0.016951f
C47 VGND VNB 1.9026f
C48 RESET_B VNB 0.133097f
C49 SET_B VNB 0.217915f
C50 CLK_N VNB 0.119128f
C51 D VNB 0.106132f
C52 SCE VNB 0.506354f
C53 SCD VNB 0.189435f
C54 VPWR VNB 1.47044f
C55 VPB VNB 3.85939f
C56 a_2392_74# VNB 0.011608f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfbbn_2 VNB VPB VPWR SET_B VGND SCD SCE D CLK_N Q_N Q RESET_B
X0 a_1997_82.t2 a_868_368.t2 a_1986_424.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.1008 ps=1.08 w=0.84 l=0.15
X1 a_1185_125.t0 a_1007_366.t3 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.24385 ps=2.14 w=0.42 l=0.15
X2 a_2452_74.t2 SET_B.t0 VGND.t11 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1369 pd=1.11 as=0.173525 ps=1.395 w=0.74 l=0.15
X3 a_1070_464.t0 a_1007_366.t4 VPWR.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1239 ps=1.43 w=0.42 l=0.15
X4 a_363_119.t1 D.t0 a_197_119.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1428 ps=1.1 w=0.42 l=0.15
X5 VGND.t5 a_2216_410# Q_N.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2294 pd=2.1 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VGND.t6 a_2216_410# a_3272_94.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.16175 pd=1.19 as=0.1824 ps=1.85 w=0.64 l=0.15
X7 a_119_119.t1 SCD.t0 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 VGND.t4 SET_B.t1 a_1473_73.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.125125 ps=1.005 w=0.55 l=0.15
X9 a_2247_82.t1 a_868_368.t3 a_1997_82.t1 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.24725 ps=1.65 w=0.42 l=0.15
X10 VGND.t3 CLK_N.t0 a_688_98.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.30025 pd=1.74 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 a_868_368.t1 a_688_98.t2 VGND.t15 VNB.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.30025 ps=1.74 w=0.74 l=0.15
X12 VPWR.t4 a_3272_94.t2 Q.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_2452_74.t0 a_1997_82.t4 a_2216_410# VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.30055 pd=2.42 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t8 SCD.t1 a_27_464.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.1888 ps=1.87 w=0.64 l=0.15
X15 a_1986_424.t1 a_1007_366.t5 VPWR.t2 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.1008 pd=1.08 as=0.2478 ps=2.27 w=0.84 l=0.15
X16 VPWR.t7 a_2216_410# a_2171_508.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.0504 ps=0.66 w=0.42 l=0.15
X17 a_341_410.t1 SCE.t0 VPWR.t15 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1888 ps=1.87 w=0.64 l=0.15
X18 VPWR.t11 SET_B.t2 a_2216_410# VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.295 ps=2.59 w=1 l=0.15
X19 VGND.t12 a_3272_94.t3 Q.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t3 a_1643_257.t2 a_1592_424.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.23 as=0.1134 ps=1.11 w=0.84 l=0.15
X21 a_2171_508.t1 a_688_98.t3 a_1997_82.t3 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.1428 ps=1.225 w=0.42 l=0.15
X22 a_1997_82.t0 a_688_98.t4 a_1902_125.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.24725 pd=1.65 as=0.108175 ps=1.09 w=0.55 l=0.15
X23 a_2556_392# a_1643_257.t3 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X24 a_1592_424.t1 a_1154_464.t4 a_1007_366.t2 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.7476 ps=3.46 w=0.84 l=0.15
X25 a_1007_366.t0 SET_B.t3 VPWR.t10 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1638 ps=1.23 w=0.84 l=0.15
X26 VPWR.t0 RESET_B.t0 a_1643_257.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.58575 pd=2.345 as=0.1888 ps=1.87 w=0.64 l=0.15
X27 VPWR a_2216_410# Q_N VPB sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X28 a_2216_410# a_1643_257.t4 a_2452_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1369 ps=1.11 w=0.74 l=0.15
X29 a_197_119.t0 SCE.t1 a_119_119.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1428 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X30 Q_N.t2 a_2216_410# VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.58575 ps=2.345 w=1.12 l=0.15
X31 VGND.t8 a_2216_410# a_2247_82.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.173525 pd=1.395 as=0.0504 ps=0.66 w=0.42 l=0.15
X32 a_27_464.t1 a_341_410.t2 a_197_119.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.096 ps=0.94 w=0.64 l=0.15
X33 a_1473_73.t1 a_1643_257.t5 a_1007_366.t1 VNB.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.125125 pd=1.005 as=0.077 ps=0.83 w=0.55 l=0.15
X34 a_197_119.t4 D.t1 a_206_464.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0768 ps=0.88 w=0.64 l=0.15
X35 a_1154_464.t3 a_688_98.t5 a_1185_125.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 a_1902_125.t0 a_1007_366.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.108175 pd=1.09 as=0.09625 ps=0.9 w=0.55 l=0.15
X37 Q.t0 a_3272_94.t4 VGND.t13 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.16175 ps=1.19 w=0.74 l=0.15
X38 a_197_119.t2 a_688_98.t6 a_1154_464.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2208 pd=1.97 as=0.1133 ps=1.025 w=0.64 l=0.15
X39 VPWR.t6 a_2216_410# a_3272_94.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2038 pd=1.495 as=0.29 ps=2.58 w=1 l=0.15
X40 VGND.t10 RESET_B.t1 a_1643_257.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.188875 pd=1.83 as=0.1176 ps=1.4 w=0.42 l=0.15
X41 a_868_368.t0 a_688_98.t7 VPWR.t14 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X42 a_197_119.t5 a_868_368.t4 a_1154_464.t0 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.55 as=0.06405 ps=0.725 w=0.42 l=0.15
X43 a_206_464.t0 SCE.t2 VPWR.t13 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.0768 pd=0.88 as=0.096 ps=0.94 w=0.64 l=0.15
X44 VPWR.t12 CLK_N.t1 a_688_98.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X45 a_1154_464.t1 a_868_368.t5 a_1070_464.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1133 pd=1.025 as=0.0567 ps=0.69 w=0.42 l=0.15
X46 VGND.t0 a_341_410.t3 a_363_119.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.0504 ps=0.66 w=0.42 l=0.15
X47 a_341_410.t0 SCE.t3 VGND.t14 VNB.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1113 ps=0.95 w=0.42 l=0.15
X48 Q_N.t0 a_2216_410# VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.188875 ps=1.83 w=0.74 l=0.15
R0 a_868_368.n1 a_868_368.t4 421.892
R1 a_868_368.n0 a_868_368.t2 419.022
R2 a_868_368.n0 a_868_368.t3 414.721
R3 a_868_368.n2 a_868_368.t5 376.13
R4 a_868_368.t0 a_868_368.n3 279.914
R5 a_868_368.n3 a_868_368.t1 123.457
R6 a_868_368.n3 a_868_368.n2 61.9299
R7 a_868_368.n1 a_868_368.n0 27.5927
R8 a_868_368.n2 a_868_368.n1 4.65505
R9 a_1986_424.t0 a_1986_424.t1 56.2862
R10 a_1997_82.t2 a_1997_82.n3 430.704
R11 a_1997_82.n3 a_1997_82.n2 265.889
R12 a_1997_82.n2 a_1997_82.t4 258.673
R13 a_1997_82.n2 a_1997_82.n1 231.629
R14 a_1997_82.n3 a_1997_82.n0 145.655
R15 a_1997_82.t2 a_1997_82.t3 111.26
R16 a_1997_82.n0 a_1997_82.t0 110.177
R17 a_1997_82.n0 a_1997_82.t1 107.067
R18 VPB.t11 VPB.t22 845.297
R19 VPB.t6 VPB.t5 738.038
R20 VPB.t14 VPB.t0 730.376
R21 VPB.t0 VPB.t6 602.688
R22 VPB.t7 VPB.t10 523.521
R23 VPB.t2 VPB.t16 515.861
R24 VPB.t19 VPB.t15 515.861
R25 VPB.t20 VPB.t17 515.861
R26 VPB.t9 VPB.t20 515.861
R27 VPB.t5 VPB.t4 497.985
R28 VPB.t3 VPB.t2 275.807
R29 VPB.t13 VPB.t21 273.253
R30 VPB.t12 VPB.t11 273.253
R31 VPB.t10 VPB.t14 260.485
R32 VPB VPB.t8 257.93
R33 VPB.t17 VPB.t19 229.839
R34 VPB.t1 VPB.t9 229.839
R35 VPB.t8 VPB.t18 229.839
R36 VPB.t22 VPB.t3 214.517
R37 VPB.t15 VPB.t12 214.517
R38 VPB.t21 VPB.t7 199.195
R39 VPB.t16 VPB.t13 199.195
R40 VPB.t18 VPB.t1 199.195
R41 a_1007_366.n0 a_1007_366.t3 478.788
R42 a_1007_366.t0 a_1007_366.n4 391.717
R43 a_1007_366.n1 a_1007_366.t2 347.955
R44 a_1007_366.n1 a_1007_366.n0 345.156
R45 a_1007_366.n2 a_1007_366.t1 300.262
R46 a_1007_366.n3 a_1007_366.t6 268.899
R47 a_1007_366.n3 a_1007_366.t5 206.166
R48 a_1007_366.n4 a_1007_366.n3 198.649
R49 a_1007_366.n0 a_1007_366.t4 138.441
R50 a_1007_366.n4 a_1007_366.n2 71.1534
R51 a_1007_366.n2 a_1007_366.n1 59.8737
R52 VGND.n16 VGND.t10 333.315
R53 VGND.n5 VGND.t1 321.108
R54 VGND.n65 VGND.n64 269.916
R55 VGND.n79 VGND.t9 254.673
R56 VGND.n72 VGND.n71 223.912
R57 VGND.n10 VGND.n9 214.868
R58 VGND.n39 VGND.n38 205.663
R59 VGND.n22 VGND.t12 179.662
R60 VGND.n25 VGND.t5 160.254
R61 VGND.n17 VGND.n16 122.245
R62 VGND.n21 VGND.n20 115.93
R63 VGND.n71 VGND.t14 111.43
R64 VGND.n38 VGND.t8 80.0005
R65 VGND.n64 VGND.t15 76.2167
R66 VGND.n16 VGND.t7 49.211
R67 VGND.n9 VGND.t4 45.8187
R68 VGND.n20 VGND.t6 45.0005
R69 VGND.n71 VGND.t0 40.0005
R70 VGND.n27 VGND.n26 36.1417
R71 VGND.n31 VGND.n30 36.1417
R72 VGND.n32 VGND.n31 36.1417
R73 VGND.n32 VGND.n14 36.1417
R74 VGND.n36 VGND.n14 36.1417
R75 VGND.n37 VGND.n36 36.1417
R76 VGND.n44 VGND.n12 36.1417
R77 VGND.n45 VGND.n44 36.1417
R78 VGND.n46 VGND.n45 36.1417
R79 VGND.n51 VGND.n50 36.1417
R80 VGND.n52 VGND.n51 36.1417
R81 VGND.n52 VGND.n7 36.1417
R82 VGND.n56 VGND.n7 36.1417
R83 VGND.n57 VGND.n56 36.1417
R84 VGND.n58 VGND.n57 36.1417
R85 VGND.n63 VGND.n62 36.1417
R86 VGND.n69 VGND.n3 36.1417
R87 VGND.n70 VGND.n69 36.1417
R88 VGND.n73 VGND.n1 36.1417
R89 VGND.n77 VGND.n1 36.1417
R90 VGND.n78 VGND.n77 36.1417
R91 VGND.n64 VGND.t3 35.6762
R92 VGND.n46 VGND.n10 34.2593
R93 VGND.n25 VGND.n19 33.8829
R94 VGND.n40 VGND.n12 32.1065
R95 VGND.n62 VGND.n5 30.8711
R96 VGND.n9 VGND.t2 30.546
R97 VGND.n38 VGND.t11 30.3649
R98 VGND.n20 VGND.t13 30.2643
R99 VGND.n65 VGND.n63 28.6123
R100 VGND.n65 VGND.n3 24.8476
R101 VGND.n21 VGND.n19 23.3417
R102 VGND.n58 VGND.n5 21.0829
R103 VGND.n79 VGND.n78 18.824
R104 VGND.n39 VGND.n37 18.6522
R105 VGND.n72 VGND.n70 15.8123
R106 VGND.n30 VGND.n17 13.9299
R107 VGND.n26 VGND.n25 13.5534
R108 VGND.n50 VGND.n10 13.177
R109 VGND.n80 VGND.n79 9.3005
R110 VGND.n78 VGND.n0 9.3005
R111 VGND.n77 VGND.n76 9.3005
R112 VGND.n75 VGND.n1 9.3005
R113 VGND.n74 VGND.n73 9.3005
R114 VGND.n70 VGND.n2 9.3005
R115 VGND.n69 VGND.n68 9.3005
R116 VGND.n67 VGND.n3 9.3005
R117 VGND.n66 VGND.n65 9.3005
R118 VGND.n63 VGND.n4 9.3005
R119 VGND.n62 VGND.n61 9.3005
R120 VGND.n60 VGND.n5 9.3005
R121 VGND.n59 VGND.n58 9.3005
R122 VGND.n57 VGND.n6 9.3005
R123 VGND.n56 VGND.n55 9.3005
R124 VGND.n54 VGND.n7 9.3005
R125 VGND.n53 VGND.n52 9.3005
R126 VGND.n51 VGND.n8 9.3005
R127 VGND.n50 VGND.n49 9.3005
R128 VGND.n48 VGND.n10 9.3005
R129 VGND.n47 VGND.n46 9.3005
R130 VGND.n45 VGND.n11 9.3005
R131 VGND.n44 VGND.n43 9.3005
R132 VGND.n42 VGND.n12 9.3005
R133 VGND.n41 VGND.n40 9.3005
R134 VGND.n37 VGND.n13 9.3005
R135 VGND.n36 VGND.n35 9.3005
R136 VGND.n34 VGND.n14 9.3005
R137 VGND.n33 VGND.n32 9.3005
R138 VGND.n31 VGND.n15 9.3005
R139 VGND.n30 VGND.n29 9.3005
R140 VGND.n23 VGND.n19 9.3005
R141 VGND.n25 VGND.n24 9.3005
R142 VGND.n26 VGND.n18 9.3005
R143 VGND.n28 VGND.n27 9.3005
R144 VGND.n22 VGND.n21 6.7255
R145 VGND.n40 VGND.n39 2.61021
R146 VGND.n73 VGND.n72 1.50638
R147 VGND.n27 VGND.n17 0.753441
R148 VGND.n23 VGND.n22 0.585846
R149 VGND.n24 VGND.n23 0.122949
R150 VGND.n24 VGND.n18 0.122949
R151 VGND.n28 VGND.n18 0.122949
R152 VGND.n29 VGND.n28 0.122949
R153 VGND.n29 VGND.n15 0.122949
R154 VGND.n33 VGND.n15 0.122949
R155 VGND.n34 VGND.n33 0.122949
R156 VGND.n35 VGND.n34 0.122949
R157 VGND.n35 VGND.n13 0.122949
R158 VGND.n41 VGND.n13 0.122949
R159 VGND.n42 VGND.n41 0.122949
R160 VGND.n43 VGND.n42 0.122949
R161 VGND.n43 VGND.n11 0.122949
R162 VGND.n47 VGND.n11 0.122949
R163 VGND.n48 VGND.n47 0.122949
R164 VGND.n49 VGND.n48 0.122949
R165 VGND.n49 VGND.n8 0.122949
R166 VGND.n53 VGND.n8 0.122949
R167 VGND.n54 VGND.n53 0.122949
R168 VGND.n55 VGND.n54 0.122949
R169 VGND.n55 VGND.n6 0.122949
R170 VGND.n59 VGND.n6 0.122949
R171 VGND.n60 VGND.n59 0.122949
R172 VGND.n61 VGND.n60 0.122949
R173 VGND.n61 VGND.n4 0.122949
R174 VGND.n66 VGND.n4 0.122949
R175 VGND.n67 VGND.n66 0.122949
R176 VGND.n68 VGND.n67 0.122949
R177 VGND.n68 VGND.n2 0.122949
R178 VGND.n74 VGND.n2 0.122949
R179 VGND.n75 VGND.n74 0.122949
R180 VGND.n76 VGND.n75 0.122949
R181 VGND.n76 VGND.n0 0.122949
R182 VGND.n80 VGND.n0 0.122949
R183 VGND VGND.n80 0.0617245
R184 a_1185_125.t0 a_1185_125.t1 60.0005
R185 VNB.t20 VNB.t23 3845.67
R186 VNB.t14 VNB.t21 2887.14
R187 VNB.t24 VNB.t5 2794.75
R188 VNB.t1 VNB.t16 2459.84
R189 VNB.t11 VNB.t10 2448.29
R190 VNB.t16 VNB.t8 2379
R191 VNB.t22 VNB.t6 2286.61
R192 VNB.t6 VNB.t24 1940.16
R193 VNB.t2 VNB.t12 1917.06
R194 VNB.t0 VNB.t22 1570.6
R195 VNB.t9 VNB.t17 1466.67
R196 VNB.t23 VNB.t7 1397.38
R197 VNB.t10 VNB.t19 1385.83
R198 VNB.t17 VNB.t3 1201.05
R199 VNB VNB.t13 1201.05
R200 VNB.t7 VNB.t4 1154.86
R201 VNB.t4 VNB.t14 1097.11
R202 VNB.t15 VNB.t20 1050.92
R203 VNB.t19 VNB.t18 993.177
R204 VNB.t8 VNB.t11 993.177
R205 VNB.t3 VNB.t1 993.177
R206 VNB.t21 VNB.t9 900.788
R207 VNB.t12 VNB.t0 900.788
R208 VNB.t13 VNB.t2 900.788
R209 VNB.t5 VNB.t15 831.496
R210 SET_B.n0 SET_B.t2 298.572
R211 SET_B.n1 SET_B.t3 251.81
R212 SET_B.n1 SET_B.t1 198.523
R213 SET_B SET_B.n1 179.434
R214 SET_B.n0 SET_B.t0 178.34
R215 SET_B SET_B.n0 171.034
R216 a_2452_74.t0 a_2452_74.n0 541.014
R217 a_2452_74.n0 a_2452_74.t1 30.0005
R218 a_2452_74.n0 a_2452_74.t2 30.0005
R219 VPWR.n34 VPWR.n31 867.872
R220 VPWR.n35 VPWR.n34 867.872
R221 VPWR.n66 VPWR.t1 695.038
R222 VPWR.n14 VPWR.t7 676.303
R223 VPWR.n55 VPWR.n11 612.152
R224 VPWR.n42 VPWR.n16 605.946
R225 VPWR.n79 VPWR.n1 605.17
R226 VPWR.n73 VPWR.t15 374.271
R227 VPWR.n12 VPWR.t2 351.106
R228 VPWR.n5 VPWR.n4 316.211
R229 VPWR.n33 VPWR.n32 306.829
R230 VPWR.n23 VPWR.t6 268.163
R231 VPWR.n22 VPWR.t4 266.168
R232 VPWR.n34 VPWR.t0 114.466
R233 VPWR.n34 VPWR.n33 57.1611
R234 VPWR.n11 VPWR.t10 56.2862
R235 VPWR.n1 VPWR.t13 46.1724
R236 VPWR.n1 VPWR.t8 46.1724
R237 VPWR.n33 VPWR.t5 45.6634
R238 VPWR.n16 VPWR.t11 39.4005
R239 VPWR.n77 VPWR.n2 36.1417
R240 VPWR.n78 VPWR.n77 36.1417
R241 VPWR.n72 VPWR.n71 36.1417
R242 VPWR.n59 VPWR.n9 36.1417
R243 VPWR.n60 VPWR.n59 36.1417
R244 VPWR.n61 VPWR.n60 36.1417
R245 VPWR.n61 VPWR.n7 36.1417
R246 VPWR.n65 VPWR.n7 36.1417
R247 VPWR.n54 VPWR.n53 36.1417
R248 VPWR.n49 VPWR.n48 36.1417
R249 VPWR.n50 VPWR.n49 36.1417
R250 VPWR.n44 VPWR.n43 36.1417
R251 VPWR.n37 VPWR.n36 36.1417
R252 VPWR.n37 VPWR.n17 36.1417
R253 VPWR.n41 VPWR.n17 36.1417
R254 VPWR.n11 VPWR.t3 35.1791
R255 VPWR.n55 VPWR.n9 33.5064
R256 VPWR.n30 VPWR.n20 33.4998
R257 VPWR.n48 VPWR.n14 32.377
R258 VPWR.n16 VPWR.t9 31.5205
R259 VPWR.n67 VPWR.n66 30.4946
R260 VPWR.n25 VPWR.n24 30.4946
R261 VPWR.n73 VPWR.n72 28.2358
R262 VPWR.n67 VPWR.n5 26.7299
R263 VPWR.n4 VPWR.t14 26.3844
R264 VPWR.n4 VPWR.t12 26.3844
R265 VPWR.n24 VPWR.n23 25.224
R266 VPWR.n79 VPWR.n78 22.9652
R267 VPWR.n66 VPWR.n65 22.9652
R268 VPWR.n71 VPWR.n5 20.7064
R269 VPWR.n73 VPWR.n2 19.2005
R270 VPWR.n25 VPWR.n20 16.9417
R271 VPWR.n44 VPWR.n14 15.0593
R272 VPWR.n55 VPWR.n54 13.9299
R273 VPWR.n36 VPWR.n35 12.7411
R274 VPWR.n24 VPWR.n21 9.3005
R275 VPWR.n26 VPWR.n25 9.3005
R276 VPWR.n27 VPWR.n20 9.3005
R277 VPWR.n30 VPWR.n29 9.3005
R278 VPWR.n28 VPWR.n19 9.3005
R279 VPWR.n36 VPWR.n18 9.3005
R280 VPWR.n38 VPWR.n37 9.3005
R281 VPWR.n39 VPWR.n17 9.3005
R282 VPWR.n41 VPWR.n40 9.3005
R283 VPWR.n43 VPWR.n15 9.3005
R284 VPWR.n45 VPWR.n44 9.3005
R285 VPWR.n46 VPWR.n14 9.3005
R286 VPWR.n48 VPWR.n47 9.3005
R287 VPWR.n49 VPWR.n13 9.3005
R288 VPWR.n51 VPWR.n50 9.3005
R289 VPWR.n53 VPWR.n52 9.3005
R290 VPWR.n54 VPWR.n10 9.3005
R291 VPWR.n56 VPWR.n55 9.3005
R292 VPWR.n57 VPWR.n9 9.3005
R293 VPWR.n59 VPWR.n58 9.3005
R294 VPWR.n60 VPWR.n8 9.3005
R295 VPWR.n62 VPWR.n61 9.3005
R296 VPWR.n63 VPWR.n7 9.3005
R297 VPWR.n65 VPWR.n64 9.3005
R298 VPWR.n66 VPWR.n6 9.3005
R299 VPWR.n68 VPWR.n67 9.3005
R300 VPWR.n69 VPWR.n5 9.3005
R301 VPWR.n71 VPWR.n70 9.3005
R302 VPWR.n72 VPWR.n3 9.3005
R303 VPWR.n74 VPWR.n73 9.3005
R304 VPWR.n75 VPWR.n2 9.3005
R305 VPWR.n77 VPWR.n76 9.3005
R306 VPWR.n78 VPWR.n0 9.3005
R307 VPWR.n32 VPWR.n19 7.97243
R308 VPWR.n53 VPWR.n12 7.90638
R309 VPWR.n80 VPWR.n79 7.27223
R310 VPWR.n23 VPWR.n22 6.59649
R311 VPWR.n42 VPWR.n41 6.4005
R312 VPWR.n43 VPWR.n42 4.89462
R313 VPWR.n35 VPWR.n19 4.37945
R314 VPWR.n50 VPWR.n12 3.38874
R315 VPWR.n31 VPWR.n30 2.58296
R316 VPWR.n22 VPWR.n21 0.612104
R317 VPWR.n32 VPWR.n31 0.225061
R318 VPWR VPWR.n80 0.157962
R319 VPWR.n80 VPWR.n0 0.149814
R320 VPWR.n26 VPWR.n21 0.122949
R321 VPWR.n27 VPWR.n26 0.122949
R322 VPWR.n29 VPWR.n27 0.122949
R323 VPWR.n29 VPWR.n28 0.122949
R324 VPWR.n28 VPWR.n18 0.122949
R325 VPWR.n38 VPWR.n18 0.122949
R326 VPWR.n39 VPWR.n38 0.122949
R327 VPWR.n40 VPWR.n39 0.122949
R328 VPWR.n40 VPWR.n15 0.122949
R329 VPWR.n45 VPWR.n15 0.122949
R330 VPWR.n46 VPWR.n45 0.122949
R331 VPWR.n47 VPWR.n46 0.122949
R332 VPWR.n47 VPWR.n13 0.122949
R333 VPWR.n51 VPWR.n13 0.122949
R334 VPWR.n52 VPWR.n51 0.122949
R335 VPWR.n52 VPWR.n10 0.122949
R336 VPWR.n56 VPWR.n10 0.122949
R337 VPWR.n57 VPWR.n56 0.122949
R338 VPWR.n58 VPWR.n57 0.122949
R339 VPWR.n58 VPWR.n8 0.122949
R340 VPWR.n62 VPWR.n8 0.122949
R341 VPWR.n63 VPWR.n62 0.122949
R342 VPWR.n64 VPWR.n63 0.122949
R343 VPWR.n64 VPWR.n6 0.122949
R344 VPWR.n68 VPWR.n6 0.122949
R345 VPWR.n69 VPWR.n68 0.122949
R346 VPWR.n70 VPWR.n69 0.122949
R347 VPWR.n70 VPWR.n3 0.122949
R348 VPWR.n74 VPWR.n3 0.122949
R349 VPWR.n75 VPWR.n74 0.122949
R350 VPWR.n76 VPWR.n75 0.122949
R351 VPWR.n76 VPWR.n0 0.122949
R352 a_1070_464.t0 a_1070_464.t1 126.644
R353 D.n0 D.t1 268.767
R354 D.n0 D.t0 227.395
R355 D D.n0 154.133
R356 a_197_119.n0 a_197_119.t2 869.496
R357 a_197_119.n3 a_197_119.n2 696.903
R358 a_197_119.n2 a_197_119.n0 522.313
R359 a_197_119.n0 a_197_119.t5 245
R360 a_197_119.n2 a_197_119.n1 120.769
R361 a_197_119.n1 a_197_119.t0 85.8513
R362 a_197_119.n1 a_197_119.t3 82.3036
R363 a_197_119.t1 a_197_119.n3 46.1724
R364 a_197_119.n3 a_197_119.t4 46.1724
R365 a_363_119.t0 a_363_119.t1 68.5719
R366 Q_N.n1 Q_N.t2 249.188
R367 Q_N Q_N.n0 126.07
R368 Q_N.n0 Q_N.t1 22.7032
R369 Q_N.n0 Q_N.t0 22.7032
R370 Q_N Q_N.n1 6.12224
R371 Q_N.n1 Q_N 4.3525
R372 a_3272_94.n1 a_3272_94.t2 261.62
R373 a_3272_94.n3 a_3272_94.n0 261.62
R374 a_3272_94.t1 a_3272_94.n4 255.603
R375 a_3272_94.n4 a_3272_94.n3 183.81
R376 a_3272_94.n1 a_3272_94.t3 156.431
R377 a_3272_94.n2 a_3272_94.t4 154.24
R378 a_3272_94.n4 a_3272_94.t0 146.541
R379 a_3272_94.n2 a_3272_94.n1 60.6157
R380 a_3272_94.n3 a_3272_94.n2 5.11262
R381 SCD.n0 SCD.t1 197.399
R382 SCD.n2 SCD.n1 152
R383 SCD.n1 SCD.t0 124.035
R384 SCD SCD.n0 70.4022
R385 SCD.n1 SCD.n0 62.2601
R386 SCD SCD.n2 8.73462
R387 SCD.n2 SCD 2.40991
R388 a_119_119.t0 a_119_119.t1 68.5719
R389 a_1473_73.t0 a_1473_73.t1 99.2732
R390 a_2247_82.t0 a_2247_82.t1 68.5719
R391 CLK_N.n0 CLK_N.t1 250.2
R392 CLK_N.n0 CLK_N.t0 180.845
R393 CLK_N CLK_N.n0 158.4
R394 a_688_98.n0 a_688_98.t4 1327.11
R395 a_688_98.t4 a_688_98.t3 866.529
R396 a_688_98.t2 a_688_98.n0 698.9
R397 a_688_98.t5 a_688_98.t6 570.889
R398 a_688_98.n2 a_688_98.t0 340.637
R399 a_688_98.t1 a_688_98.n2 297.565
R400 a_688_98.n1 a_688_98.t7 231.677
R401 a_688_98.n1 a_688_98.t2 206.822
R402 a_688_98.n0 a_688_98.t5 186.374
R403 a_688_98.n2 a_688_98.n1 152
R404 Q Q.t2 232.097
R405 Q Q.n0 165.554
R406 Q.n0 Q.t1 22.7032
R407 Q.n0 Q.t0 22.7032
R408 a_27_464.t0 a_27_464.t1 864.181
R409 a_2171_508.t0 a_2171_508.t1 112.572
R410 SCE.t1 SCE.t3 964
R411 SCE.t3 SCE.t0 766.38
R412 SCE.n0 SCE.t2 271.527
R413 SCE SCE.n0 153.256
R414 SCE.n2 SCE.n1 152
R415 SCE.n1 SCE.t1 126.927
R416 SCE.n1 SCE.n0 49.6611
R417 SCE SCE.n2 7.27893
R418 SCE.n2 SCE 2.00834
R419 a_341_410.t1 a_341_410.n1 392.473
R420 a_341_410.n1 a_341_410.n0 328.733
R421 a_341_410.n0 a_341_410.t2 314.908
R422 a_341_410.n0 a_341_410.t3 274.74
R423 a_341_410.n1 a_341_410.t0 261.961
R424 a_1154_464.n4 a_1154_464.n3 685.501
R425 a_1154_464.n2 a_1154_464.t4 342.488
R426 a_1154_464.n3 a_1154_464.n0 245.944
R427 a_1154_464.n3 a_1154_464.n2 234.875
R428 a_1154_464.n2 a_1154_464.n1 143.798
R429 a_1154_464.n4 a_1154_464.t1 110.227
R430 a_1154_464.n0 a_1154_464.t3 47.1434
R431 a_1154_464.t2 a_1154_464.n4 46.1724
R432 a_1154_464.n0 a_1154_464.t0 40.0005
R433 a_1643_257.t0 a_1643_257.n3 690.153
R434 a_1643_257.n2 a_1643_257.n1 459.644
R435 a_1643_257.n0 a_1643_257.t3 298.572
R436 a_1643_257.n3 a_1643_257.t1 236.442
R437 a_1643_257.n1 a_1643_257.t2 229.44
R438 a_1643_257.n0 a_1643_257.t4 178.34
R439 a_1643_257.n1 a_1643_257.t5 168.529
R440 a_1643_257.n2 a_1643_257.n0 158.595
R441 a_1643_257.n3 a_1643_257.n2 62.0269
R442 a_1592_424.t0 a_1592_424.t1 63.3219
R443 a_1902_125.n0 a_1902_125.t1 54.1389
R444 a_1902_125.n1 a_1902_125.n0 50.4005
R445 a_1902_125.n0 a_1902_125.t0 17.5273
R446 RESET_B.n0 RESET_B.t0 173.788
R447 RESET_B RESET_B.n0 155.492
R448 RESET_B.n0 RESET_B.t1 151.028
R449 a_206_464.t0 a_206_464.t1 73.8755
C0 VGND RESET_B 0.004499f
C1 a_2556_392# a_2216_410# 0.015829f
C2 VGND CLK_N 0.009571f
C3 VPB a_2216_410# 0.367793f
C4 VPB Q_N 0.007503f
C5 VPWR a_2216_410# 0.520106f
C6 SET_B a_2216_410# 0.088776f
C7 VPB Q 0.006611f
C8 VPWR Q_N 0.191556f
C9 SET_B Q_N 1.28e-19
C10 VGND a_2216_410# 0.186265f
C11 VPWR Q 0.230711f
C12 RESET_B a_2216_410# 0.092363f
C13 SET_B Q 2.35e-20
C14 VGND Q_N 0.169575f
C15 VGND Q 0.160688f
C16 RESET_B Q_N 5.39e-19
C17 VPWR a_2556_392# 0.009205f
C18 RESET_B Q 8.13e-20
C19 VPB VPWR 0.545173f
C20 SET_B VPB 0.120336f
C21 VPB SCE 0.175372f
C22 VPB SCD 0.084478f
C23 VGND a_2556_392# 0.001297f
C24 SET_B VPWR 0.120812f
C25 VGND VPB 0.03157f
C26 Q_N a_2216_410# 0.115519f
C27 VPWR SCE 0.038727f
C28 VPB D 0.072242f
C29 VPWR SCD 0.017197f
C30 SET_B SCE 3.31e-20
C31 VGND VPWR 0.222133f
C32 RESET_B VPB 0.064251f
C33 Q a_2216_410# 0.001982f
C34 VPWR D 0.007011f
C35 SCD SCE 0.151885f
C36 VPB CLK_N 0.03553f
C37 SET_B VGND 0.073235f
C38 VGND SCE 0.0865f
C39 SET_B D 3.91e-20
C40 VGND SCD 0.04941f
C41 RESET_B VPWR 0.006627f
C42 SCE D 0.135725f
C43 VPWR CLK_N 0.019415f
C44 SCD D 0.001024f
C45 SET_B RESET_B 4.01e-19
C46 VGND D 0.008053f
C47 SET_B CLK_N 5.34e-20
C48 SCE CLK_N 0.042193f
C49 Q VNB 0.03091f
C50 Q_N VNB 0.01212f
C51 RESET_B VNB 0.102666f
C52 VGND VNB 2.10142f
C53 SET_B VNB 0.222804f
C54 CLK_N VNB 0.102503f
C55 D VNB 0.112703f
C56 SCE VNB 0.532319f
C57 SCD VNB 0.205879f
C58 VPWR VNB 1.63319f
C59 VPB VNB 4.15598f
C60 a_2216_410# VNB 0.613006f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfbbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfbbp_1 VNB VPB VPWR VGND Q_N RESET_B D SCE SCD Q CLK SET_B
X0 a_1580_379.t1 a_1092_96.t4 a_1250_231.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.1638 ps=1.23 w=0.84 l=0.15
X1 Q_N.t1 a_2037_442# VGND.t10 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10825 ps=1.065 w=0.74 l=0.15
X2 a_877_98.t0 a_622_98.t2 VPWR.t10 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_218_464.t0 SCE.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.1152 ps=1 w=0.64 l=0.15
X4 VPWR.t9 CLK.t0 a_622_98.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 a_2037_442# a_1878_420.t4 a_2271_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_2271_74.t0 a_1625_93.t1 a_2037_442# VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1443 ps=1.13 w=0.74 l=0.15
X7 a_1092_96.t3 a_622_98.t3 a_197_119.t3 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 a_119_119.t0 SCD.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 a_1418_125# SET_B.t0 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.229275 pd=1.45 as=0.17465 ps=1.35 w=0.55 l=0.15
X10 a_341_93.t1 SCE.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1155 ps=0.97 w=0.42 l=0.15
X11 VPWR.t15 RESET_B.t0 a_1625_93.t0 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.1828 pd=1.485 as=0.1792 ps=1.84 w=0.64 l=0.15
X12 Q.t1 a_2881_74.t1 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X13 a_2061_74.t0 a_622_98.t4 a_1878_420.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.117225 ps=1.17 w=0.42 l=0.15
X14 VPWR.t12 a_2037_442# a_1986_504.t1 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.267925 pd=1.88 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VPWR.t2 SCD.t1 a_27_464.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1152 pd=1 as=0.1888 ps=1.87 w=0.64 l=0.15
X16 Q_N.t0 a_2037_442# VPWR.t11 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1828 ps=1.485 w=1.12 l=0.15
X17 VPWR.t13 a_2037_442# a_2881_74.t0 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.1883 pd=1.48 as=0.2478 ps=2.27 w=0.84 l=0.15
X18 VGND.t7 a_341_93.t2 a_299_119.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 a_1878_420.t1 a_877_98.t2 a_1880_119.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.117225 pd=1.17 as=0.05775 ps=0.76 w=0.55 l=0.15
X20 a_2037_442# SET_B.t1 VPWR.t14 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.267925 ps=1.88 w=1 l=0.15
X21 a_341_93.t0 SCE.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1888 ps=1.87 w=0.64 l=0.15
X22 a_197_119.t0 SCE.t3 a_119_119.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 a_1880_119.t0 a_1250_231.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.05775 pd=0.76 as=0.15675 ps=1.67 w=0.55 l=0.15
X24 a_1250_231.t2 a_1092_96.t5 a_1418_125# VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.229275 ps=1.45 w=0.55 l=0.15
X25 Q.t0 a_2881_74.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1883 ps=1.48 w=1.12 l=0.15
X26 a_1986_504.t0 a_877_98.t3 a_1878_420.t0 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1449 ps=1.23 w=0.42 l=0.15
X27 a_299_119.t1 D.t0 a_197_119.t5 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X28 VGND.t9 a_2037_442# a_2061_74.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X29 VPWR.t4 a_1250_231.t4 a_1221_419.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2358 pd=1.525 as=0.0567 ps=0.69 w=0.42 l=0.15
X30 a_1221_419.t1 a_622_98.t5 a_1092_96.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1163 ps=1.055 w=0.42 l=0.15
X31 VGND.t8 CLK.t1 a_622_98.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.30025 pd=1.74 as=0.2109 ps=2.05 w=0.74 l=0.15
X32 a_877_98.t1 a_622_98.t6 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2516 pd=2.16 as=0.30025 ps=1.74 w=0.74 l=0.15
X33 a_1192_96# a_877_98.t4 a_1092_96.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.080925 pd=0.89 as=0.0735 ps=0.77 w=0.42 l=0.15
X34 a_27_464.t1 a_341_93.t3 a_197_119.t2 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.096 ps=0.94 w=0.64 l=0.15
X35 a_1250_231.t0 SET_B.t2 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.23 as=0.2358 ps=1.525 w=0.84 l=0.15
X36 a_197_119.t4 D.t1 a_218_464.t1 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X37 a_1092_96.t2 a_877_98.t5 a_197_119.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1163 pd=1.055 as=0.1888 ps=1.87 w=0.64 l=0.15
X38 VPWR.t7 a_1625_93.t2 a_1580_379.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.2 as=0.1134 ps=1.11 w=0.84 l=0.15
X39 a_1878_420.t3 a_622_98.t7 a_1766_379.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1449 pd=1.23 as=0.1845 ps=1.455 w=0.84 l=0.15
X40 VPWR.t8 a_1625_93.t3 a_2384_392.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.28 pd=2.56 as=0.12 ps=1.24 w=1 l=0.15
X41 a_2271_74.t1 SET_B.t3 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1212 ps=1.1 w=0.74 l=0.15
X42 a_1766_379.t0 a_1250_231.t5 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1845 pd=1.455 as=0.1512 ps=1.2 w=0.84 l=0.15
R0 a_1092_96.n3 a_1092_96.n2 624.085
R1 a_1092_96.n2 a_1092_96.n1 309.856
R2 a_1092_96.n2 a_1092_96.n0 266.017
R3 a_1092_96.n1 a_1092_96.t4 246.089
R4 a_1092_96.n1 a_1092_96.t5 147.814
R5 a_1092_96.n3 a_1092_96.t0 86.7743
R6 a_1092_96.n5 a_1092_96.n4 81.7741
R7 a_1092_96.n0 a_1092_96.t3 60.0005
R8 a_1092_96.n4 a_1092_96.n3 46.9053
R9 a_1092_96.n0 a_1092_96.t1 40.0005
R10 a_1092_96.n4 a_1092_96.t2 33.4995
R11 a_1250_231.n5 a_1250_231.n4 387.769
R12 a_1250_231.n2 a_1250_231.n1 284.308
R13 a_1250_231.n1 a_1250_231.t4 258.942
R14 a_1250_231.n3 a_1250_231.t3 240.311
R15 a_1250_231.n3 a_1250_231.t5 223.288
R16 a_1250_231.n2 a_1250_231.t2 215.546
R17 a_1250_231.n4 a_1250_231.n3 152
R18 a_1250_231.n1 a_1250_231.n0 126.927
R19 a_1250_231.n4 a_1250_231.n2 94.4562
R20 a_1250_231.t0 a_1250_231.n5 56.2862
R21 a_1250_231.n5 a_1250_231.t1 35.1791
R22 a_1580_379.t0 a_1580_379.t1 63.3219
R23 VPB.t20 VPB.t15 566.936
R24 VPB.t17 VPB.t16 564.383
R25 VPB.t18 VPB.t21 520.968
R26 VPB.t1 VPB.t13 515.861
R27 VPB.t12 VPB.t1 515.861
R28 VPB.t10 VPB.t22 500.538
R29 VPB.t21 VPB.t10 480.108
R30 VPB.t4 VPB.t5 426.478
R31 VPB.t15 VPB.t7 288.575
R32 VPB.t3 VPB.t8 286.022
R33 VPB.t8 VPB.t14 275.807
R34 VPB.t5 VPB.t11 275.807
R35 VPB.t22 VPB.t17 263.038
R36 VPB.t16 VPB.t6 260.485
R37 VPB.t9 VPB.t3 260.485
R38 VPB.t2 VPB.t0 260.485
R39 VPB VPB.t2 257.93
R40 VPB.t13 VPB.t20 229.839
R41 VPB.t19 VPB.t12 229.839
R42 VPB.t14 VPB.t18 214.517
R43 VPB.t11 VPB.t9 214.517
R44 VPB.t7 VPB.t4 214.517
R45 VPB.t0 VPB.t19 214.517
R46 VGND.n43 VGND.t5 316.443
R47 VGND.n9 VGND.t2 258.81
R48 VGND.n67 VGND.t1 254.673
R49 VGND.n52 VGND.n51 253.276
R50 VGND.n15 VGND.t10 252.929
R51 VGND.n60 VGND.n59 225.704
R52 VGND.n25 VGND.n22 202.409
R53 VGND.n25 VGND.n24 185
R54 VGND.n14 VGND.t3 156.862
R55 VGND.n59 VGND.t0 117.144
R56 VGND.n51 VGND.t8 76.2167
R57 VGND.n23 VGND.t9 61.4291
R58 VGND.t6 VGND.n22 52.5005
R59 VGND.n24 VGND.t6 40.0005
R60 VGND.n59 VGND.t7 40.0005
R61 VGND.n16 VGND.n13 36.1417
R62 VGND.n20 VGND.n13 36.1417
R63 VGND.n21 VGND.n20 36.1417
R64 VGND.n27 VGND.n21 36.1417
R65 VGND.n31 VGND.n11 36.1417
R66 VGND.n32 VGND.n31 36.1417
R67 VGND.n33 VGND.n32 36.1417
R68 VGND.n37 VGND.n36 36.1417
R69 VGND.n38 VGND.n37 36.1417
R70 VGND.n38 VGND.n7 36.1417
R71 VGND.n42 VGND.n7 36.1417
R72 VGND.n45 VGND.n44 36.1417
R73 VGND.n45 VGND.n5 36.1417
R74 VGND.n49 VGND.n5 36.1417
R75 VGND.n50 VGND.n49 36.1417
R76 VGND.n57 VGND.n3 36.1417
R77 VGND.n58 VGND.n57 36.1417
R78 VGND.n61 VGND.n58 36.1417
R79 VGND.n65 VGND.n1 36.1417
R80 VGND.n66 VGND.n65 36.1417
R81 VGND.n51 VGND.t4 35.6762
R82 VGND.n53 VGND.n50 30.8384
R83 VGND.n26 VGND.n25 25.8565
R84 VGND.n52 VGND.n3 22.4971
R85 VGND.n67 VGND.n66 18.824
R86 VGND.n15 VGND.n14 14.3664
R87 VGND.n60 VGND.n1 11.2946
R88 VGND.n36 VGND.n9 10.9181
R89 VGND.n27 VGND.n26 9.78874
R90 VGND.n68 VGND.n67 9.3005
R91 VGND.n17 VGND.n16 9.3005
R92 VGND.n18 VGND.n13 9.3005
R93 VGND.n20 VGND.n19 9.3005
R94 VGND.n21 VGND.n12 9.3005
R95 VGND.n28 VGND.n27 9.3005
R96 VGND.n29 VGND.n11 9.3005
R97 VGND.n31 VGND.n30 9.3005
R98 VGND.n32 VGND.n10 9.3005
R99 VGND.n34 VGND.n33 9.3005
R100 VGND.n36 VGND.n35 9.3005
R101 VGND.n37 VGND.n8 9.3005
R102 VGND.n39 VGND.n38 9.3005
R103 VGND.n40 VGND.n7 9.3005
R104 VGND.n42 VGND.n41 9.3005
R105 VGND.n44 VGND.n6 9.3005
R106 VGND.n46 VGND.n45 9.3005
R107 VGND.n47 VGND.n5 9.3005
R108 VGND.n49 VGND.n48 9.3005
R109 VGND.n50 VGND.n4 9.3005
R110 VGND.n54 VGND.n53 9.3005
R111 VGND.n55 VGND.n3 9.3005
R112 VGND.n57 VGND.n56 9.3005
R113 VGND.n58 VGND.n2 9.3005
R114 VGND.n62 VGND.n61 9.3005
R115 VGND.n63 VGND.n1 9.3005
R116 VGND.n65 VGND.n64 9.3005
R117 VGND.n66 VGND.n0 9.3005
R118 VGND.n26 VGND.n11 7.52991
R119 VGND.n16 VGND.n15 7.15344
R120 VGND.n33 VGND.n9 6.4005
R121 VGND.n61 VGND.n60 6.02403
R122 VGND.n43 VGND.n42 5.64756
R123 VGND.n23 VGND.n22 1.8755
R124 VGND.n53 VGND.n52 1.44746
R125 VGND.n24 VGND.n23 1.42907
R126 VGND.n44 VGND.n43 0.753441
R127 VGND.n17 VGND.n14 0.20927
R128 VGND.n18 VGND.n17 0.122949
R129 VGND.n19 VGND.n18 0.122949
R130 VGND.n19 VGND.n12 0.122949
R131 VGND.n28 VGND.n12 0.122949
R132 VGND.n29 VGND.n28 0.122949
R133 VGND.n30 VGND.n29 0.122949
R134 VGND.n30 VGND.n10 0.122949
R135 VGND.n34 VGND.n10 0.122949
R136 VGND.n35 VGND.n34 0.122949
R137 VGND.n35 VGND.n8 0.122949
R138 VGND.n39 VGND.n8 0.122949
R139 VGND.n40 VGND.n39 0.122949
R140 VGND.n41 VGND.n40 0.122949
R141 VGND.n41 VGND.n6 0.122949
R142 VGND.n46 VGND.n6 0.122949
R143 VGND.n47 VGND.n46 0.122949
R144 VGND.n48 VGND.n47 0.122949
R145 VGND.n48 VGND.n4 0.122949
R146 VGND.n54 VGND.n4 0.122949
R147 VGND.n55 VGND.n54 0.122949
R148 VGND.n56 VGND.n55 0.122949
R149 VGND.n56 VGND.n2 0.122949
R150 VGND.n62 VGND.n2 0.122949
R151 VGND.n63 VGND.n62 0.122949
R152 VGND.n64 VGND.n63 0.122949
R153 VGND.n64 VGND.n0 0.122949
R154 VGND.n68 VGND.n0 0.122949
R155 VGND VGND.n68 0.0617245
R156 Q_N Q_N.n0 585.79
R157 Q_N.n2 Q_N.n0 585
R158 Q_N.n1 Q_N.n0 585
R159 Q_N.n1 Q_N.t1 192.772
R160 Q_N.n0 Q_N.t0 26.3844
R161 Q_N.n2 Q_N 11.0622
R162 Q_N Q_N.n1 2.05482
R163 Q_N Q_N.n2 0.632599
R164 VNB VNB.n0 30909.7
R165 VNB.t17 VNB.t6 3961.22
R166 VNB.t4 VNB.t11 3591.6
R167 VNB.t9 VNB.t15 2609.97
R168 VNB.n0 VNB.t17 2535.18
R169 VNB.t18 VNB.t8 2482.94
R170 VNB.t13 VNB.t0 2286.61
R171 VNB.t8 VNB.t13 1940.16
R172 VNB.t11 VNB.t9 1743.83
R173 VNB.t0 VNB.t12 1616.8
R174 VNB.t7 VNB.t14 1258.79
R175 VNB.t5 VNB.t2 1247.24
R176 VNB.t16 VNB.t7 1247.24
R177 VNB.t3 VNB 1201.05
R178 VNB.t10 VNB.t16 1177.95
R179 VNB.t19 VNB.t1 1177.95
R180 VNB.t15 VNB.t18 1154.86
R181 VNB.n0 VNB.t5 993.177
R182 VNB.t2 VNB.t10 993.177
R183 VNB.t1 VNB.t3 900.788
R184 VNB.t14 VNB.t4 831.496
R185 VNB.t12 VNB.t19 831.496
R186 a_622_98.n0 a_622_98.t7 1192.95
R187 a_622_98.n1 a_622_98.n0 851.534
R188 a_622_98.t7 a_622_98.t4 795.054
R189 a_622_98.n1 a_622_98.t3 555.908
R190 a_622_98.n4 a_622_98.t1 306.55
R191 a_622_98.n3 a_622_98.t2 253.587
R192 a_622_98.n0 a_622_98.t5 241.536
R193 a_622_98.t0 a_622_98.n4 233.004
R194 a_622_98.n4 a_622_98.n3 197.827
R195 a_622_98.n2 a_622_98.t6 165.196
R196 a_622_98.n2 a_622_98.n1 99.6138
R197 a_622_98.n3 a_622_98.n2 13.146
R198 VPWR.n24 VPWR.t8 741.731
R199 VPWR.n61 VPWR.t1 660.869
R200 VPWR.n18 VPWR.n17 615.674
R201 VPWR.n40 VPWR.n11 610.601
R202 VPWR.n67 VPWR.n1 606.721
R203 VPWR.n33 VPWR.n32 585
R204 VPWR.n31 VPWR.n30 585
R205 VPWR.n54 VPWR.n53 333.466
R206 VPWR.n20 VPWR.n19 330.565
R207 VPWR.n46 VPWR.n8 324.853
R208 VPWR.n32 VPWR.n31 172.375
R209 VPWR.n8 VPWR.t5 130.096
R210 VPWR.n32 VPWR.t12 114.171
R211 VPWR.n8 VPWR.t4 86.8476
R212 VPWR.n31 VPWR.t14 71.3682
R213 VPWR.n17 VPWR.t15 69.2583
R214 VPWR.n1 VPWR.t2 61.563
R215 VPWR.n1 VPWR.t0 49.2505
R216 VPWR.n19 VPWR.t13 48.0779
R217 VPWR.n11 VPWR.t3 42.2148
R218 VPWR.n11 VPWR.t7 42.2148
R219 VPWR.n65 VPWR.n2 36.1417
R220 VPWR.n66 VPWR.n65 36.1417
R221 VPWR.n47 VPWR.n6 36.1417
R222 VPWR.n51 VPWR.n6 36.1417
R223 VPWR.n52 VPWR.n51 36.1417
R224 VPWR.n55 VPWR.n52 36.1417
R225 VPWR.n59 VPWR.n4 36.1417
R226 VPWR.n60 VPWR.n59 36.1417
R227 VPWR.n44 VPWR.n9 36.1417
R228 VPWR.n45 VPWR.n44 36.1417
R229 VPWR.n34 VPWR.n12 36.1417
R230 VPWR.n38 VPWR.n12 36.1417
R231 VPWR.n39 VPWR.n38 36.1417
R232 VPWR.n25 VPWR.n15 36.1417
R233 VPWR.n29 VPWR.n15 36.1417
R234 VPWR.n23 VPWR.n22 36.1417
R235 VPWR.n55 VPWR.n54 32.377
R236 VPWR.n19 VPWR.t6 32.1717
R237 VPWR.n40 VPWR.n9 29.7417
R238 VPWR.n61 VPWR.n60 27.4829
R239 VPWR.n53 VPWR.t10 26.3844
R240 VPWR.n53 VPWR.t9 26.3844
R241 VPWR.n61 VPWR.n2 25.977
R242 VPWR.n17 VPWR.t11 24.6255
R243 VPWR.n67 VPWR.n66 19.2005
R244 VPWR.n40 VPWR.n39 14.6829
R245 VPWR.n30 VPWR.n29 12.5861
R246 VPWR.n34 VPWR.n33 11.4567
R247 VPWR.n22 VPWR.n18 10.5417
R248 VPWR.n22 VPWR.n21 9.3005
R249 VPWR.n23 VPWR.n16 9.3005
R250 VPWR.n26 VPWR.n25 9.3005
R251 VPWR.n27 VPWR.n15 9.3005
R252 VPWR.n29 VPWR.n28 9.3005
R253 VPWR.n14 VPWR.n13 9.3005
R254 VPWR.n35 VPWR.n34 9.3005
R255 VPWR.n36 VPWR.n12 9.3005
R256 VPWR.n38 VPWR.n37 9.3005
R257 VPWR.n39 VPWR.n10 9.3005
R258 VPWR.n41 VPWR.n40 9.3005
R259 VPWR.n42 VPWR.n9 9.3005
R260 VPWR.n44 VPWR.n43 9.3005
R261 VPWR.n45 VPWR.n7 9.3005
R262 VPWR.n48 VPWR.n47 9.3005
R263 VPWR.n49 VPWR.n6 9.3005
R264 VPWR.n51 VPWR.n50 9.3005
R265 VPWR.n52 VPWR.n5 9.3005
R266 VPWR.n56 VPWR.n55 9.3005
R267 VPWR.n57 VPWR.n4 9.3005
R268 VPWR.n59 VPWR.n58 9.3005
R269 VPWR.n60 VPWR.n3 9.3005
R270 VPWR.n62 VPWR.n61 9.3005
R271 VPWR.n63 VPWR.n2 9.3005
R272 VPWR.n65 VPWR.n64 9.3005
R273 VPWR.n66 VPWR.n0 9.3005
R274 VPWR.n47 VPWR.n46 8.65932
R275 VPWR.n20 VPWR.n18 8.34873
R276 VPWR.n68 VPWR.n67 7.43488
R277 VPWR.n24 VPWR.n23 7.15344
R278 VPWR.n25 VPWR.n24 4.14168
R279 VPWR.n54 VPWR.n4 3.76521
R280 VPWR.n33 VPWR.n14 3.39123
R281 VPWR.n30 VPWR.n14 3.13692
R282 VPWR.n46 VPWR.n45 2.63579
R283 VPWR.n21 VPWR.n20 0.203618
R284 VPWR VPWR.n68 0.160103
R285 VPWR.n68 VPWR.n0 0.1477
R286 VPWR.n21 VPWR.n16 0.122949
R287 VPWR.n26 VPWR.n16 0.122949
R288 VPWR.n27 VPWR.n26 0.122949
R289 VPWR.n28 VPWR.n27 0.122949
R290 VPWR.n28 VPWR.n13 0.122949
R291 VPWR.n35 VPWR.n13 0.122949
R292 VPWR.n36 VPWR.n35 0.122949
R293 VPWR.n37 VPWR.n36 0.122949
R294 VPWR.n37 VPWR.n10 0.122949
R295 VPWR.n41 VPWR.n10 0.122949
R296 VPWR.n42 VPWR.n41 0.122949
R297 VPWR.n43 VPWR.n42 0.122949
R298 VPWR.n43 VPWR.n7 0.122949
R299 VPWR.n48 VPWR.n7 0.122949
R300 VPWR.n49 VPWR.n48 0.122949
R301 VPWR.n50 VPWR.n49 0.122949
R302 VPWR.n50 VPWR.n5 0.122949
R303 VPWR.n56 VPWR.n5 0.122949
R304 VPWR.n57 VPWR.n56 0.122949
R305 VPWR.n58 VPWR.n57 0.122949
R306 VPWR.n58 VPWR.n3 0.122949
R307 VPWR.n62 VPWR.n3 0.122949
R308 VPWR.n63 VPWR.n62 0.122949
R309 VPWR.n64 VPWR.n63 0.122949
R310 VPWR.n64 VPWR.n0 0.122949
R311 a_877_98.t4 a_877_98.t2 1558.47
R312 a_877_98.t2 a_877_98.t3 594.735
R313 a_877_98.n0 a_877_98.t4 344.466
R314 a_877_98.n1 a_877_98.t1 299.425
R315 a_877_98.t0 a_877_98.n1 242.393
R316 a_877_98.n0 a_877_98.t5 238.958
R317 a_877_98.n1 a_877_98.n0 171.589
R318 SCE.t3 SCE.t1 857.961
R319 SCE.t1 SCE.t2 623.654
R320 SCE.n0 SCE.t3 332.58
R321 SCE.n0 SCE.t0 191.194
R322 SCE SCE.n0 161.333
R323 a_218_464.t0 a_218_464.t1 83.1099
R324 a_1878_420.t3 a_1878_420.n4 778.717
R325 a_1878_420.t3 a_1878_420.n4 594.891
R326 a_1878_420.n1 a_1878_420.n0 298.572
R327 a_1878_420.n3 a_1878_420.n1 278.933
R328 a_1878_420.n3 a_1878_420.n2 220.52
R329 a_1878_420.n1 a_1878_420.t4 178.34
R330 a_1878_420.n2 a_1878_420.t2 115.715
R331 a_1878_420.t3 a_1878_420.t0 112.572
R332 a_1878_420.n4 a_1878_420.n3 50.6204
R333 a_1878_420.n2 a_1878_420.t1 30.546
R334 CLK.n0 CLK.t0 274.269
R335 CLK.n0 CLK.t1 172.499
R336 CLK CLK.n0 163.442
R337 a_2271_74.t0 a_2271_74.n0 291.813
R338 a_2271_74.n0 a_2271_74.t2 22.7032
R339 a_2271_74.n0 a_2271_74.t1 22.7032
R340 a_1625_93.t0 a_1625_93.n3 726.87
R341 a_1625_93.n2 a_1625_93.t3 277.459
R342 a_1625_93.n1 a_1625_93.t2 246.089
R343 a_1625_93.n3 a_1625_93.n2 204.583
R344 a_1625_93.n3 a_1625_93.n1 181.018
R345 a_1625_93.n2 a_1625_93.t1 154.24
R346 a_1625_93.n1 a_1625_93.n0 147.814
R347 a_197_119.n2 a_197_119.n0 676.889
R348 a_197_119.t1 a_197_119.n3 489.534
R349 a_197_119.n3 a_197_119.n2 305.38
R350 a_197_119.n2 a_197_119.n1 251.978
R351 a_197_119.n3 a_197_119.t3 225
R352 a_197_119.n1 a_197_119.t0 62.8576
R353 a_197_119.n0 a_197_119.t2 46.1724
R354 a_197_119.n0 a_197_119.t4 46.1724
R355 a_197_119.n1 a_197_119.t5 40.0005
R356 SCD.n0 SCD.t1 197.399
R357 SCD.n2 SCD.n1 152
R358 SCD.n1 SCD.t0 124.035
R359 SCD SCD.n0 70.4022
R360 SCD.n1 SCD.n0 62.2601
R361 SCD SCD.n2 8.73462
R362 SCD.n2 SCD 2.40991
R363 a_119_119.t0 a_119_119.t1 68.5719
R364 SET_B.n2 SET_B.n0 702.876
R365 SET_B.n1 SET_B.t3 258.673
R366 SET_B.n1 SET_B.t1 231.629
R367 SET_B.n0 SET_B.t2 209.476
R368 SET_B.n0 SET_B.t0 169.31
R369 SET_B.n2 SET_B.n1 157.781
R370 SET_B SET_B.n2 7.22631
R371 a_341_93.t0 a_341_93.n1 382.072
R372 a_341_93.n0 a_341_93.t2 380.781
R373 a_341_93.n1 a_341_93.t1 300.305
R374 a_341_93.n1 a_341_93.n0 191.489
R375 a_341_93.n0 a_341_93.t3 177.411
R376 RESET_B.n1 RESET_B.t0 181.821
R377 RESET_B RESET_B.n1 159.594
R378 RESET_B.n1 RESET_B.n0 126.927
R379 a_2881_74.t0 a_2881_74.n0 725.207
R380 a_2881_74.n0 a_2881_74.t2 295.579
R381 a_2881_74.n0 a_2881_74.t1 219.53
R382 Q.n3 Q 589.707
R383 Q.n3 Q.n0 585
R384 Q.n4 Q.n3 585
R385 Q.n2 Q.t1 279.738
R386 Q.t1 Q.n1 279.738
R387 Q.n3 Q.t0 26.3844
R388 Q Q.n4 12.6123
R389 Q.n1 Q 12.2358
R390 Q Q.n0 10.9181
R391 Q Q.n2 9.22403
R392 Q.n2 Q 4.70638
R393 Q Q.n0 3.01226
R394 Q.n1 Q 1.69462
R395 Q.n4 Q 1.31815
R396 a_2061_74.t0 a_2061_74.t1 111.43
R397 a_1986_504.t0 a_1986_504.t1 126.644
R398 a_27_464.t0 a_27_464.t1 1142.3
R399 a_299_119.t0 a_299_119.t1 60.0005
R400 a_1880_119.t0 a_1880_119.t1 45.8187
R401 D.n0 D.t1 249.856
R402 D.n0 D.t0 249.856
R403 D D.n0 156.542
R404 a_1221_419.t0 a_1221_419.t1 126.644
R405 a_1766_379.t0 a_1766_379.t1 110.376
C0 a_2037_442# SET_B 0.244235f
C1 a_2037_442# Q_N 0.155559f
C2 VPB SCD 0.082221f
C3 VPWR SCD 0.016409f
C4 CLK SCE 0.023923f
C5 VGND SCE 0.080294f
C6 VPB SCE 0.151553f
C7 VPWR SCE 0.032097f
C8 VGND D 0.0096f
C9 VPB D 0.068174f
C10 VPWR D 0.006736f
C11 VGND CLK 0.012211f
C12 a_2037_442# Q 0.003517f
C13 VPB CLK 0.049106f
C14 CLK VPWR 0.016841f
C15 VPB VGND 0.030383f
C16 VGND VPWR 0.189049f
C17 VGND RESET_B 0.021436f
C18 VPB VPWR 0.444602f
C19 VPB RESET_B 0.042454f
C20 RESET_B VPWR 0.005225f
C21 VGND SET_B 0.019142f
C22 VGND Q_N 0.108948f
C23 VPB SET_B 0.147543f
C24 VPWR SET_B 0.571798f
C25 VPB Q_N 0.016676f
C26 RESET_B SET_B 7.89e-20
C27 Q_N VPWR 0.072512f
C28 a_1192_96# VGND 0.004215f
C29 RESET_B Q_N 0.003341f
C30 a_1192_96# VPWR 6e-19
C31 a_1418_125# VGND 0.183922f
C32 SCD SCE 0.139793f
C33 a_1418_125# VPWR 0.001631f
C34 SCD D 0.00121f
C35 a_1418_125# SET_B 0.001723f
C36 a_2037_442# VGND 0.069619f
C37 VGND Q 0.089872f
C38 SCE D 0.133084f
C39 VPB a_2037_442# 0.3341f
C40 a_2037_442# VPWR 0.322136f
C41 VPB Q 0.014595f
C42 VPWR Q 0.109475f
C43 a_2037_442# RESET_B 0.089506f
C44 RESET_B Q 1.4e-19
C45 VGND SCD 0.049409f
C46 Q VNB 0.112393f
C47 Q_N VNB 0.019167f
C48 RESET_B VNB 0.1089f
C49 VGND VNB 1.82907f
C50 SET_B VNB 0.205362f
C51 VPWR VNB 1.40313f
C52 CLK VNB 0.132776f
C53 D VNB 0.103131f
C54 SCE VNB 0.467367f
C55 SCD VNB 0.209246f
C56 VPB VNB 3.63926f
C57 a_1418_125# VNB 0.013437f
C58 a_2037_442# VNB 0.444454f
.ends

* NGSPICE file created from sky130_fd_sc_hs__sdfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrbp_1 VNB VPB VPWR RESET_B VGND Q_N SCE CLK SCD D Q
X0 a_1369_71.t1 a_1221_97.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.24015 ps=1.585 w=0.64 l=0.15
X1 VPWR.t1 CLK.t0 a_850_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_512_464.t1 a_27_74.t2 a_413_90.t5 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.1248 pd=1.03 as=0.096 ps=0.94 w=0.64 l=0.15
X3 a_1023_74.t1 a_850_74.t2 VPWR.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_1966_74.t1 a_850_74.t3 a_1747_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.22595 ps=1.585 w=0.42 l=0.15
X5 a_413_90.t1 D.t0 a_338_464.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.096 pd=0.94 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 VPWR.t2 a_1369_71.t3 a_1328_463.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.126225 pd=1.105 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 VPWR.t7 SCD.t0 a_512_464.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.06 as=0.1248 ps=1.03 w=0.64 l=0.15
X8 VGND.t3 CLK.t1 a_850_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_2124_74.t0 RESET_B.t0 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_1328_463.t1 a_850_74.t4 a_1221_97.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X11 VGND.t5 SCE.t0 a_27_74.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X12 Q.t1 a_2513_424.t2 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1939 ps=1.49 w=1.12 l=0.15
X13 a_413_90.t2 D.t1 a_312_90.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.107525 pd=0.965 as=0.07455 ps=0.775 w=0.42 l=0.15
X14 a_1221_97.t2 RESET_B.t1 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.126225 ps=1.105 w=0.42 l=0.15
X15 a_1969_489.t0 a_1023_74.t2 a_1747_74.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.207425 ps=1.755 w=0.42 l=0.15
X16 a_2008_48.t0 RESET_B.t2 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.11785 ps=1.01 w=0.42 l=0.15
X17 a_225_90.t0 SCD.t1 a_545_97.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.085825 pd=0.855 as=0.0504 ps=0.66 w=0.42 l=0.15
X18 a_2008_48.t1 a_1747_74.t3 a_2124_74.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 VPWR.t8 a_1747_74.t4 a_2513_424.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1939 pd=1.49 as=0.231 ps=2.23 w=0.84 l=0.15
X20 VGND.t2 a_2008_48.t2 a_1966_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 a_338_464.t1 SCE.t1 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0864 pd=0.91 as=0.112 ps=0.99 w=0.64 l=0.15
X22 a_1321_97# a_1023_74.t3 a_1221_97.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X23 a_1221_97.t1 a_1023_74.t4 a_413_90.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X24 a_413_90.t6 RESET_B.t3 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1344 ps=1.06 w=0.64 l=0.15
X25 a_312_90.t1 a_27_74.t3 a_225_90.t2 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.07455 pd=0.775 as=0.1197 ps=1.41 w=0.42 l=0.15
X26 a_1747_74.t0 a_850_74.t5 a_1369_71.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.207425 pd=1.755 as=0.15 ps=1.3 w=1 l=0.15
X27 a_1369_71.t0 a_1221_97.t6 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.285 ps=2.57 w=1 l=0.15
X28 VGND.t9 a_1747_74.t5 a_2513_424.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.118675 pd=1.08 as=0.14575 ps=1.63 w=0.55 l=0.15
X29 a_1221_97.t4 a_850_74.t6 a_413_90.t4 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X30 VPWR.t5 SCE.t2 a_27_74.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.112 pd=0.99 as=0.5792 ps=3.09 w=0.64 l=0.15
X31 a_545_97.t1 SCE.t3 a_413_90.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.107525 ps=0.965 w=0.42 l=0.15
X32 VGND.t6 RESET_B.t4 a_1399_97.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.24015 pd=1.585 as=0.0504 ps=0.66 w=0.42 l=0.15
X33 VGND.t7 RESET_B.t5 a_225_90.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1365 pd=1.49 as=0.085825 ps=0.855 w=0.42 l=0.15
X34 a_1023_74.t0 a_850_74.t7 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X35 Q.t0 a_2513_424.t3 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.118675 ps=1.08 w=0.74 l=0.15
R0 a_1221_97.n1 a_1221_97.t2 669.625
R1 a_1221_97.n3 a_1221_97.n2 611.165
R2 a_1221_97.n4 a_1221_97.n3 313.697
R3 a_1221_97.n0 a_1221_97.t6 284.983
R4 a_1221_97.n1 a_1221_97.n0 239.508
R5 a_1221_97.n0 a_1221_97.t5 200.13
R6 a_1221_97.n2 a_1221_97.t3 70.3576
R7 a_1221_97.n2 a_1221_97.t1 70.3576
R8 a_1221_97.n4 a_1221_97.t4 60.0005
R9 a_1221_97.n3 a_1221_97.n1 48.5652
R10 a_1221_97.t0 a_1221_97.n4 40.0005
R11 VGND.n3 VGND.t7 259.12
R12 VGND.n46 VGND.t5 247.498
R13 VGND.n8 VGND.n7 210.602
R14 VGND.n14 VGND.n13 207.498
R15 VGND.n33 VGND.n32 206.333
R16 VGND.n12 VGND.n11 143.933
R17 VGND.n7 VGND.t0 117.376
R18 VGND.n7 VGND.t6 53.9524
R19 VGND.n11 VGND.t9 44.1118
R20 VGND.n13 VGND.t8 40.0005
R21 VGND.n13 VGND.t2 40.0005
R22 VGND.n15 VGND.n10 36.1417
R23 VGND.n19 VGND.n10 36.1417
R24 VGND.n20 VGND.n19 36.1417
R25 VGND.n21 VGND.n20 36.1417
R26 VGND.n25 VGND.n8 36.1417
R27 VGND.n26 VGND.n25 36.1417
R28 VGND.n27 VGND.n26 36.1417
R29 VGND.n27 VGND.n5 36.1417
R30 VGND.n31 VGND.n5 36.1417
R31 VGND.n35 VGND.n34 36.1417
R32 VGND.n39 VGND.n38 36.1417
R33 VGND.n40 VGND.n39 36.1417
R34 VGND.n40 VGND.n1 36.1417
R35 VGND.n44 VGND.n1 36.1417
R36 VGND.n45 VGND.n44 36.1417
R37 VGND.n15 VGND.n14 24.4711
R38 VGND.n46 VGND.n45 24.4711
R39 VGND.n32 VGND.t1 22.7032
R40 VGND.n32 VGND.t3 22.7032
R41 VGND.n11 VGND.t4 22.2507
R42 VGND.n21 VGND.n8 11.2946
R43 VGND.n16 VGND.n15 9.3005
R44 VGND.n17 VGND.n10 9.3005
R45 VGND.n19 VGND.n18 9.3005
R46 VGND.n20 VGND.n9 9.3005
R47 VGND.n22 VGND.n21 9.3005
R48 VGND.n23 VGND.n8 9.3005
R49 VGND.n25 VGND.n24 9.3005
R50 VGND.n26 VGND.n6 9.3005
R51 VGND.n28 VGND.n27 9.3005
R52 VGND.n29 VGND.n5 9.3005
R53 VGND.n31 VGND.n30 9.3005
R54 VGND.n34 VGND.n4 9.3005
R55 VGND.n36 VGND.n35 9.3005
R56 VGND.n38 VGND.n37 9.3005
R57 VGND.n39 VGND.n2 9.3005
R58 VGND.n41 VGND.n40 9.3005
R59 VGND.n42 VGND.n1 9.3005
R60 VGND.n44 VGND.n43 9.3005
R61 VGND.n45 VGND.n0 9.3005
R62 VGND.n34 VGND.n33 7.52991
R63 VGND.n47 VGND.n46 7.19894
R64 VGND.n14 VGND.n12 7.10595
R65 VGND.n35 VGND.n3 6.02403
R66 VGND.n38 VGND.n3 5.27109
R67 VGND.n33 VGND.n31 3.76521
R68 VGND.n16 VGND.n12 0.158857
R69 VGND VGND.n47 0.156997
R70 VGND.n47 VGND.n0 0.150766
R71 VGND.n17 VGND.n16 0.122949
R72 VGND.n18 VGND.n17 0.122949
R73 VGND.n18 VGND.n9 0.122949
R74 VGND.n22 VGND.n9 0.122949
R75 VGND.n23 VGND.n22 0.122949
R76 VGND.n24 VGND.n23 0.122949
R77 VGND.n24 VGND.n6 0.122949
R78 VGND.n28 VGND.n6 0.122949
R79 VGND.n29 VGND.n28 0.122949
R80 VGND.n30 VGND.n29 0.122949
R81 VGND.n30 VGND.n4 0.122949
R82 VGND.n36 VGND.n4 0.122949
R83 VGND.n37 VGND.n36 0.122949
R84 VGND.n37 VGND.n2 0.122949
R85 VGND.n41 VGND.n2 0.122949
R86 VGND.n42 VGND.n41 0.122949
R87 VGND.n43 VGND.n42 0.122949
R88 VGND.n43 VGND.n0 0.122949
R89 a_1369_71.n2 a_1369_71.n1 264.137
R90 a_1369_71.n3 a_1369_71.n2 258.861
R91 a_1369_71.n1 a_1369_71.n0 254.053
R92 a_1369_71.n1 a_1369_71.t3 237.986
R93 a_1369_71.n2 a_1369_71.t1 219.395
R94 a_1369_71.n3 a_1369_71.t2 29.5505
R95 a_1369_71.t0 a_1369_71.n3 29.5505
R96 VNB.n0 VNB 21976.9
R97 VNB.n1 VNB 19567.8
R98 VNB VNB.n2 9558.62
R99 VNB.t16 VNB.t14 4677.17
R100 VNB.t0 VNB.n0 3141.11
R101 VNB.t2 VNB.t15 2310.88
R102 VNB.t17 VNB.t10 2286.61
R103 VNB.t1 VNB.t11 1820.69
R104 VNB.t11 VNB.n1 1622.28
R105 VNB.t6 VNB.t4 1524.41
R106 VNB.t12 VNB.t9 1247.24
R107 VNB.n2 VNB.t5 1202.12
R108 VNB.n2 VNB.t12 1189.5
R109 VNB.t15 VNB.t1 1167.11
R110 VNB.t4 VNB.t17 1166.4
R111 VNB.t10 VNB 1143.31
R112 VNB.t14 VNB.t7 1131.76
R113 VNB.t5 VNB.t2 1003.71
R114 VNB.t3 VNB.t13 993.177
R115 VNB.t9 VNB.t6 900.788
R116 VNB.t13 VNB.t16 831.496
R117 VNB.t8 VNB.t3 831.496
R118 VNB.n0 VNB.t8 554.332
R119 VNB.n1 VNB.t0 550
R120 CLK.n0 CLK.t0 261.647
R121 CLK.n0 CLK.t1 154.24
R122 CLK CLK.n0 114.379
R123 a_850_74.n0 a_850_74.t5 998.812
R124 a_850_74.t0 a_850_74.n4 892.058
R125 a_850_74.n1 a_850_74.n0 838.681
R126 a_850_74.t5 a_850_74.t3 727.821
R127 a_850_74.n1 a_850_74.t6 294.021
R128 a_850_74.n3 a_850_74.t2 258.942
R129 a_850_74.n4 a_850_74.t1 198.273
R130 a_850_74.n0 a_850_74.t4 182.625
R131 a_850_74.n2 a_850_74.t7 153.948
R132 a_850_74.n4 a_850_74.n3 152
R133 a_850_74.n2 a_850_74.n1 99.6138
R134 a_850_74.n3 a_850_74.n2 29.9429
R135 VPWR.n14 VPWR.t9 718.654
R136 VPWR.n26 VPWR.n11 670.255
R137 VPWR.n7 VPWR.n6 606.139
R138 VPWR.n4 VPWR.n3 603.312
R139 VPWR.n1 VPWR.n0 315.151
R140 VPWR.n12 VPWR.t0 272.253
R141 VPWR.n16 VPWR.n15 242.188
R142 VPWR.n11 VPWR.t6 105.537
R143 VPWR.n11 VPWR.t2 105.537
R144 VPWR.n3 VPWR.t10 78.4927
R145 VPWR.n0 VPWR.t5 61.563
R146 VPWR.n3 VPWR.t7 50.7896
R147 VPWR.n15 VPWR.t8 46.4003
R148 VPWR.n0 VPWR.t4 46.1724
R149 VPWR.n43 VPWR.n42 36.1417
R150 VPWR.n44 VPWR.n43 36.1417
R151 VPWR.n37 VPWR.n36 36.1417
R152 VPWR.n38 VPWR.n37 36.1417
R153 VPWR.n27 VPWR.n9 36.1417
R154 VPWR.n31 VPWR.n9 36.1417
R155 VPWR.n32 VPWR.n31 36.1417
R156 VPWR.n33 VPWR.n32 36.1417
R157 VPWR.n25 VPWR.n24 36.1417
R158 VPWR.n19 VPWR.n18 36.1417
R159 VPWR.n20 VPWR.n19 36.1417
R160 VPWR.n15 VPWR.t11 35.6466
R161 VPWR.n18 VPWR.n14 35.0123
R162 VPWR.n42 VPWR.n4 33.5064
R163 VPWR.n20 VPWR.n12 29.7417
R164 VPWR.n6 VPWR.t3 26.3844
R165 VPWR.n6 VPWR.t1 26.3844
R166 VPWR.n24 VPWR.n12 23.7181
R167 VPWR.n38 VPWR.n4 11.6711
R168 VPWR.n36 VPWR.n7 10.9181
R169 VPWR.n27 VPWR.n26 9.78874
R170 VPWR.n46 VPWR.n1 9.53521
R171 VPWR.n44 VPWR.n1 9.41227
R172 VPWR.n18 VPWR.n17 9.3005
R173 VPWR.n19 VPWR.n13 9.3005
R174 VPWR.n21 VPWR.n20 9.3005
R175 VPWR.n22 VPWR.n12 9.3005
R176 VPWR.n24 VPWR.n23 9.3005
R177 VPWR.n25 VPWR.n10 9.3005
R178 VPWR.n28 VPWR.n27 9.3005
R179 VPWR.n29 VPWR.n9 9.3005
R180 VPWR.n31 VPWR.n30 9.3005
R181 VPWR.n32 VPWR.n8 9.3005
R182 VPWR.n34 VPWR.n33 9.3005
R183 VPWR.n36 VPWR.n35 9.3005
R184 VPWR.n37 VPWR.n5 9.3005
R185 VPWR.n39 VPWR.n38 9.3005
R186 VPWR.n40 VPWR.n4 9.3005
R187 VPWR.n42 VPWR.n41 9.3005
R188 VPWR.n43 VPWR.n2 9.3005
R189 VPWR.n45 VPWR.n44 9.3005
R190 VPWR.n16 VPWR.n14 6.19542
R191 VPWR.n26 VPWR.n25 1.50638
R192 VPWR.n33 VPWR.n7 0.376971
R193 VPWR VPWR.n46 0.282382
R194 VPWR.n17 VPWR.n16 0.175971
R195 VPWR.n46 VPWR.n45 0.148529
R196 VPWR.n17 VPWR.n13 0.122949
R197 VPWR.n21 VPWR.n13 0.122949
R198 VPWR.n22 VPWR.n21 0.122949
R199 VPWR.n23 VPWR.n22 0.122949
R200 VPWR.n23 VPWR.n10 0.122949
R201 VPWR.n28 VPWR.n10 0.122949
R202 VPWR.n29 VPWR.n28 0.122949
R203 VPWR.n30 VPWR.n29 0.122949
R204 VPWR.n30 VPWR.n8 0.122949
R205 VPWR.n34 VPWR.n8 0.122949
R206 VPWR.n35 VPWR.n34 0.122949
R207 VPWR.n35 VPWR.n5 0.122949
R208 VPWR.n39 VPWR.n5 0.122949
R209 VPWR.n40 VPWR.n39 0.122949
R210 VPWR.n41 VPWR.n40 0.122949
R211 VPWR.n41 VPWR.n2 0.122949
R212 VPWR.n45 VPWR.n2 0.122949
R213 VPB.n0 VPB 4859.81
R214 VPB VPB.n1 2069.28
R215 VPB.t14 VPB.t13 1082.8
R216 VPB.t10 VPB 569.49
R217 VPB.t1 VPB.t14 523.521
R218 VPB.t8 VPB.t2 515.427
R219 VPB.t11 VPB.t0 500.267
R220 VPB.t5 VPB.t11 303.192
R221 VPB.t15 VPB.t12 291.13
R222 VPB.n1 VPB.t3 277.926
R223 VPB.t12 VPB.t17 275.807
R224 VPB.t13 VPB.t16 265.591
R225 VPB.t6 VPB.n0 262.767
R226 VPB.n1 VPB.t15 255.376
R227 VPB.t9 VPB.t10 255.376
R228 VPB.t17 VPB.t4 229.839
R229 VPB.t0 VPB.t6 227.394
R230 VPB.t2 VPB.t7 227.394
R231 VPB.t3 VPB.t8 227.394
R232 VPB.t4 VPB.t9 214.517
R233 VPB.t7 VPB.t5 197.075
R234 VPB.n0 VPB.t1 130.243
R235 a_27_74.n4 a_27_74.n2 585
R236 a_27_74.n4 a_27_74.n3 585
R237 a_27_74.n3 a_27_74.t2 432.123
R238 a_27_74.n1 a_27_74.t3 346.248
R239 a_27_74.t1 a_27_74.n0 327.411
R240 a_27_74.n1 a_27_74.t0 245.481
R241 a_27_74.n2 a_27_74.n1 58.3767
R242 a_27_74.t1 a_27_74.n4 38.0944
R243 a_27_74.n2 a_27_74.n0 4.19131
R244 a_27_74.n3 a_27_74.n0 4.19131
R245 a_413_90.n0 a_413_90.t0 659.966
R246 a_413_90.n0 a_413_90.t4 403.32
R247 a_413_90.n3 a_413_90.n2 375.387
R248 a_413_90.n2 a_413_90.n1 366.747
R249 a_413_90.n2 a_413_90.t6 356.743
R250 a_413_90.n2 a_413_90.n0 131.185
R251 a_413_90.n1 a_413_90.t2 102.388
R252 a_413_90.n3 a_413_90.t5 46.1724
R253 a_413_90.t1 a_413_90.n3 46.1724
R254 a_413_90.n1 a_413_90.t3 27.0479
R255 a_512_464.t0 a_512_464.t1 120.047
R256 a_1023_74.t1 a_1023_74.n4 893.843
R257 a_1023_74.n2 a_1023_74.n1 446.021
R258 a_1023_74.n0 a_1023_74.t3 395.533
R259 a_1023_74.n3 a_1023_74.n2 362.329
R260 a_1023_74.n2 a_1023_74.t2 353.471
R261 a_1023_74.n0 a_1023_74.t4 205.387
R262 a_1023_74.n4 a_1023_74.n0 168.874
R263 a_1023_74.n3 a_1023_74.t0 134.338
R264 a_1023_74.n4 a_1023_74.n3 69.7496
R265 a_1747_74.n10 a_1747_74.n0 585
R266 a_1747_74.n9 a_1747_74.t1 326.538
R267 a_1747_74.n11 a_1747_74.n10 321.277
R268 a_1747_74.n7 a_1747_74.n1 290.272
R269 a_1747_74.n4 a_1747_74.t4 255.46
R270 a_1747_74.n4 a_1747_74.t5 230.339
R271 a_1747_74.n6 a_1747_74.n2 225.47
R272 a_1747_74.n8 a_1747_74.t3 206.712
R273 a_1747_74.n9 a_1747_74.n8 199.632
R274 a_1747_74.n5 a_1747_74.n3 159.06
R275 a_1747_74.n5 a_1747_74.n4 135.837
R276 a_1747_74.n10 a_1747_74.n9 92.578
R277 a_1747_74.n12 a_1747_74.n11 86.5611
R278 a_1747_74.n0 a_1747_74.t2 70.3576
R279 a_1747_74.n12 a_1747_74.n0 68.0124
R280 a_1747_74.n7 a_1747_74.n6 61.5894
R281 a_1747_74.n11 a_1747_74.t0 28.8409
R282 a_1747_74.n8 a_1747_74.n7 10.5176
R283 a_1747_74.n6 a_1747_74.n5 4.28494
R284 a_1966_74.t0 a_1966_74.t1 60.0005
R285 D.n0 D.t0 399.702
R286 D D.n0 160.704
R287 D.n0 D.t1 125.23
R288 a_338_464.t0 a_338_464.t1 83.1099
R289 a_1328_463.t0 a_1328_463.t1 112.572
R290 SCD.n1 SCD.t1 263.493
R291 SCD.n2 SCD.t0 187.178
R292 SCD.n1 SCD.n0 152
R293 SCD.n3 SCD.n2 152
R294 SCD.n2 SCD.n1 49.6611
R295 SCD.n3 SCD.n0 13.1884
R296 SCD.n0 SCD 0.970197
R297 SCD SCD.n3 0.194439
R298 RESET_B.n0 RESET_B.t0 414.521
R299 RESET_B.n2 RESET_B.t4 408.094
R300 RESET_B.n1 RESET_B.t5 378.151
R301 RESET_B.n3 RESET_B.n1 221.522
R302 RESET_B.n0 RESET_B.t2 217.589
R303 RESET_B.n3 RESET_B.n2 200.874
R304 RESET_B RESET_B.n0 167.919
R305 RESET_B.n1 RESET_B.t3 152.367
R306 RESET_B.n2 RESET_B.t1 122.364
R307 RESET_B RESET_B.n3 2.42441
R308 a_2124_74.t0 a_2124_74.t1 60.0005
R309 a_2008_48.n2 a_2008_48.t0 655.357
R310 a_2008_48.t1 a_2008_48.n2 418.49
R311 a_2008_48.n1 a_2008_48.t2 353.272
R312 a_2008_48.n1 a_2008_48.n0 213.493
R313 a_2008_48.n2 a_2008_48.n1 209.631
R314 SCE SCE.t3 414.675
R315 SCE.n5 SCE.t0 351.861
R316 SCE.n2 SCE.t1 248.767
R317 SCE.n3 SCE.t2 224.667
R318 SCE.n2 SCE.n1 152
R319 SCE.n4 SCE.n0 152
R320 SCE.n6 SCE.n5 152
R321 SCE.n5 SCE.n4 49.6611
R322 SCE.n3 SCE.n2 48.9308
R323 SCE.n6 SCE.n0 11.1595
R324 SCE.n1 SCE 10.9954
R325 SCE.n1 SCE 4.75947
R326 SCE SCE.n6 4.43127
R327 SCE.n4 SCE.n3 0.730803
R328 SCE SCE.n0 0.164603
R329 a_2513_424.t1 a_2513_424.n1 425.601
R330 a_2513_424.n0 a_2513_424.t2 264.298
R331 a_2513_424.n1 a_2513_424.t0 244.964
R332 a_2513_424.n0 a_2513_424.t3 204.048
R333 a_2513_424.n1 a_2513_424.n0 177.988
R334 Q.n1 Q 590.715
R335 Q.n1 Q.n0 585
R336 Q.n2 Q.n1 585
R337 Q.t0 Q.n3 279.738
R338 Q.n4 Q.t0 279.738
R339 Q.n3 Q 63.6826
R340 Q.n1 Q.t1 26.3844
R341 Q.n2 Q 15.3148
R342 Q.n0 Q 13.2576
R343 Q.n4 Q 11.3978
R344 Q.n3 Q 4.38406
R345 Q.n0 Q 3.65764
R346 Q Q.n2 1.6005
R347 Q Q.n4 1.57858
R348 a_312_90.t0 a_312_90.t1 101.43
R349 a_545_97.t0 a_545_97.t1 68.5719
R350 a_225_90.n0 a_225_90.t2 570.499
R351 a_225_90.n0 a_225_90.t1 31.4169
R352 a_225_90.n1 a_225_90.n0 30.4005
R353 a_225_90.n1 a_225_90.t0 26.5777
R354 a_225_90.n2 a_225_90.n1 9.6005
R355 Q_N.n1 Q_N.n0 1170.52
R356 Q_N Q_N.n2 14.2067
R357 Q_N.n2 Q_N 13.9734
R358 Q_N.n1 Q_N 10.2793
R359 Q_N.n0 Q_N 7.98149
R360 Q_N.n0 Q_N 6.2937
R361 Q_N Q_N.n1 4.07323
R362 Q_N.n2 Q_N 0.106323
C0 VPWR Q 0.116797f
C1 RESET_B SCE 3.11e-19
C2 SCD D 0.005619f
C3 VPWR VPB 0.400242f
C4 VPWR SCE 0.037063f
C5 RESET_B D 9.57e-19
C6 CLK VGND 0.022293f
C7 VPWR D 0.013171f
C8 Q VPB 0.014019f
C9 RESET_B CLK 0.063718f
C10 SCD VGND 0.00606f
C11 VGND Q_N 0.048348f
C12 RESET_B VGND 0.201925f
C13 VPWR CLK 0.010474f
C14 VPB SCE 0.187816f
C15 SCD RESET_B 0.085032f
C16 VPWR VGND 0.112211f
C17 RESET_B Q_N 7.99e-19
C18 VPB D 0.054885f
C19 SCD VPWR 0.014629f
C20 VPWR Q_N 0.116593f
C21 SCE D 0.161492f
C22 RESET_B VPWR 0.350099f
C23 CLK VPB 0.050696f
C24 Q VGND 0.103685f
C25 a_1321_97# VGND 4.68e-19
C26 VGND VPB 0.024704f
C27 CLK SCE 2.82e-19
C28 SCD VPB 0.074598f
C29 Q_N VPB 0.011934f
C30 VGND SCE 0.027606f
C31 RESET_B Q 1.95e-19
C32 RESET_B a_1321_97# 2.54e-19
C33 SCD SCE 0.077107f
C34 RESET_B VPB 0.358063f
C35 VGND D 0.010157f
C36 Q VNB 0.112219f
C37 Q_N VNB 0.010543f
C38 VGND VNB 1.59395f
C39 CLK VNB 0.160769f
C40 VPWR VNB 1.23448f
C41 RESET_B VNB 0.4347f
C42 SCD VNB 0.115736f
C43 D VNB 0.145853f
C44 SCE VNB 0.366736f
C45 VPB VNB 3.22017f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o22a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o22a_2 VNB VPB VPWR VGND X B2 B1 A2 A1
X0 a_82_48.t0 B2.t0 a_383_384.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X1 VPWR.t2 a_82_48.t4 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.35 pd=1.785 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_383_384.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.35 ps=1.785 w=1 l=0.15
X3 a_575_384.t1 A2.t0 a_82_48.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.18 ps=1.36 w=1 l=0.15
X4 VPWR.t3 A1.t0 a_575_384.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.195 ps=1.39 w=1 l=0.15
X5 VGND.t3 A2.t1 a_307_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X6 VGND.t1 a_82_48.t5 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.19325 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 X.t2 a_82_48.t6 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X8 X.t3 a_82_48.t7 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2035 ps=2.03 w=0.74 l=0.15
X9 a_307_74.t0 B2.t1 a_82_48.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1147 ps=1.05 w=0.74 l=0.15
X10 a_307_74.t1 A1.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 a_82_48.t2 B1.t1 a_307_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.195 ps=2.03 w=0.74 l=0.15
R0 B2.n0 B2.t1 245.821
R1 B2.n0 B2.t0 231.629
R2 B2 B2.n0 161.51
R3 a_383_384.t0 a_383_384.t1 59.1005
R4 a_82_48.n5 a_82_48.n4 320.082
R5 a_82_48.n2 a_82_48.t4 252.636
R6 a_82_48.n4 a_82_48.n0 248.66
R7 a_82_48.n1 a_82_48.t6 240.197
R8 a_82_48.n1 a_82_48.t7 226.942
R9 a_82_48.n3 a_82_48.t5 197.05
R10 a_82_48.n4 a_82_48.n3 152
R11 a_82_48.n2 a_82_48.n1 53.2213
R12 a_82_48.n5 a_82_48.t3 41.3705
R13 a_82_48.t0 a_82_48.n5 29.5505
R14 a_82_48.n0 a_82_48.t1 25.1356
R15 a_82_48.n0 a_82_48.t2 25.1356
R16 a_82_48.n3 a_82_48.n2 4.66502
R17 VPB.t3 VPB.t0 416.264
R18 VPB VPB.t2 293.683
R19 VPB.t4 VPB.t5 275.807
R20 VPB.t1 VPB.t4 260.485
R21 VPB.t0 VPB.t1 229.839
R22 VPB.t2 VPB.t3 229.839
R23 X.n2 X.n0 271.49
R24 X.n2 X.n1 95.4914
R25 X.n0 X.t1 26.3844
R26 X.n0 X.t2 26.3844
R27 X.n1 X.t0 22.7032
R28 X.n1 X.t3 22.7032
R29 X X.n2 1.80288
R30 VPWR.n1 VPWR.t3 260.738
R31 VPWR.n5 VPWR.t1 258.875
R32 VPWR.n3 VPWR.n2 142.531
R33 VPWR.n2 VPWR.t0 61.4512
R34 VPWR.n2 VPWR.t2 56.9872
R35 VPWR.n4 VPWR.n3 31.2476
R36 VPWR.n5 VPWR.n4 19.2005
R37 VPWR.n4 VPWR.n0 9.3005
R38 VPWR.n6 VPWR.n5 9.3005
R39 VPWR.n3 VPWR.n1 4.06016
R40 VPWR.n1 VPWR.n0 0.216549
R41 VPWR.n6 VPWR.n0 0.122949
R42 VPWR VPWR.n6 0.0617245
R43 B1.n0 B1.t1 240.885
R44 B1.n0 B1.t0 226.692
R45 B1 B1.n0 156.207
R46 A2.n0 A2.t1 245.821
R47 A2.n0 A2.t0 231.629
R48 A2 A2.n0 157.851
R49 a_575_384.t0 a_575_384.t1 76.8305
R50 A1.n0 A1.t0 258.738
R51 A1.n0 A1.t1 196.345
R52 A1 A1.n0 156.462
R53 a_307_74.n0 a_307_74.t2 274.51
R54 a_307_74.n0 a_307_74.t1 212.136
R55 a_307_74.n1 a_307_74.n0 88.3339
R56 a_307_74.t0 a_307_74.n1 34.0546
R57 a_307_74.n1 a_307_74.t3 22.7032
R58 VGND.n3 VGND.t1 231.476
R59 VGND.n2 VGND.n1 215.543
R60 VGND.n5 VGND.t0 170.655
R61 VGND.n1 VGND.t3 34.0546
R62 VGND.n5 VGND.n4 26.7299
R63 VGND.n1 VGND.t2 22.7032
R64 VGND.n4 VGND.n3 18.4476
R65 VGND.n6 VGND.n5 9.3005
R66 VGND.n4 VGND.n0 9.3005
R67 VGND.n3 VGND.n2 7.38408
R68 VGND.n2 VGND.n0 0.163687
R69 VGND.n6 VGND.n0 0.122949
R70 VGND VGND.n6 0.0617245
R71 VNB.t2 VNB.t4 2240.42
R72 VNB.t5 VNB.t3 1154.86
R73 VNB.t0 VNB.t5 1154.86
R74 VNB VNB.t1 1120.21
R75 VNB.t4 VNB.t0 1062.47
R76 VNB.t1 VNB.t2 993.177
C0 VPB VPWR 0.129089f
C1 X B2 2.88e-19
C2 A2 VGND 0.015836f
C3 A2 VPB 0.041177f
C4 VPWR A1 0.054362f
C5 B2 VPWR 0.012826f
C6 VPB VGND 0.009375f
C7 X B1 0.001026f
C8 B2 A2 0.084504f
C9 A1 VGND 0.018001f
C10 A2 A1 0.092903f
C11 B2 VGND 0.007988f
C12 B1 VPWR 0.020946f
C13 VPB A1 0.04978f
C14 B2 VPB 0.038068f
C15 B2 A1 2.44e-19
C16 B1 VGND 0.00792f
C17 X VPWR 0.195371f
C18 B1 VPB 0.048132f
C19 X VGND 0.125724f
C20 B1 A1 1.32e-19
C21 B1 B2 0.096072f
C22 X VPB 0.00592f
C23 VPWR VGND 0.074593f
C24 A2 VPWR 0.024877f
C25 VGND VNB 0.530047f
C26 A1 VNB 0.173096f
C27 A2 VNB 0.1041f
C28 B2 VNB 0.102658f
C29 B1 VNB 0.116184f
C30 X VNB 0.03051f
C31 VPWR VNB 0.465638f
C32 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21ba_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21ba_2 VNB VPB VPWR VGND A1 X A2 B1_N
X0 VPWR.t1 B1_N.t0 a_27_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2086 pd=1.515 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VGND.t3 A2.t0 a_487_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1797 pd=1.34 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VGND.t0 a_177_48.t3 X.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_582_368.t1 A2.t1 a_177_48.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X4 a_177_48.t0 a_27_74.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.4044 ps=1.855 w=1 l=0.15
X5 VPWR.t0 A1.t0 a_582_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.18 ps=1.36 w=1 l=0.15
X6 a_487_74.t1 a_27_74.t3 a_177_48.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2035 ps=2.03 w=0.74 l=0.15
X7 VGND.t2 B1_N.t1 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.113125 pd=1.065 as=0.15125 ps=1.65 w=0.55 l=0.15
X8 X.t0 a_177_48.t4 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.113125 ps=1.065 w=0.74 l=0.15
X9 a_487_74.t0 A1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1797 ps=1.34 w=0.74 l=0.15
X10 VPWR.t4 a_177_48.t5 X.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4044 pd=1.855 as=0.168 ps=1.42 w=1.12 l=0.15
X11 X.t2 a_177_48.t6 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2086 ps=1.515 w=1.12 l=0.15
R0 B1_N.n0 B1_N.t1 227.395
R1 B1_N.n0 B1_N.t0 212.131
R2 B1_N B1_N.n0 155.601
R3 a_27_74.t0 a_27_74.n1 340.853
R4 a_27_74.n1 a_27_74.t1 324.497
R5 a_27_74.n1 a_27_74.n0 313.762
R6 a_27_74.n0 a_27_74.t2 211.179
R7 a_27_74.n0 a_27_74.t3 196.013
R8 VPWR.n10 VPWR.n1 649.676
R9 VPWR.n3 VPWR.n2 589.49
R10 VPWR.n5 VPWR.n4 585
R11 VPWR.n6 VPWR.t0 263.921
R12 VPWR.n4 VPWR.n3 58.1488
R13 VPWR.n1 VPWR.t1 56.2862
R14 VPWR.n4 VPWR.t2 47.2805
R15 VPWR.n1 VPWR.t3 30.268
R16 VPWR.n9 VPWR.n8 29.2457
R17 VPWR.n3 VPWR.t4 21.4094
R18 VPWR.n10 VPWR.n9 16.5652
R19 VPWR.n8 VPWR.n7 9.3005
R20 VPWR.n9 VPWR.n0 9.3005
R21 VPWR.n6 VPWR.n5 8.80459
R22 VPWR.n11 VPWR.n10 7.53404
R23 VPWR.n5 VPWR.n2 5.21248
R24 VPWR.n8 VPWR.n2 0.766967
R25 VPWR.n7 VPWR.n6 0.224492
R26 VPWR VPWR.n11 0.161409
R27 VPWR.n11 VPWR.n0 0.146411
R28 VPWR.n7 VPWR.n0 0.122949
R29 VPB.t5 VPB.t3 452.017
R30 VPB.t2 VPB.t4 278.361
R31 VPB.t0 VPB.t1 260.485
R32 VPB VPB.t2 257.93
R33 VPB.t3 VPB.t0 229.839
R34 VPB.t4 VPB.t5 229.839
R35 A2.n0 A2.t1 266.44
R36 A2.n0 A2.t0 178.34
R37 A2 A2.n0 156.351
R38 a_487_74.t0 a_487_74.n0 381.606
R39 a_487_74.n0 a_487_74.t2 22.7032
R40 a_487_74.n0 a_487_74.t1 22.7032
R41 VGND.n3 VGND.t0 240.471
R42 VGND.n2 VGND.n1 219.627
R43 VGND.n6 VGND.n5 216.232
R44 VGND.n1 VGND.t1 34.0546
R45 VGND.n1 VGND.t3 34.0546
R46 VGND.n5 VGND.t4 33.8208
R47 VGND.n6 VGND.n4 31.2476
R48 VGND.n5 VGND.t2 30.546
R49 VGND.n4 VGND.n3 24.0946
R50 VGND.n4 VGND.n0 9.3005
R51 VGND.n3 VGND.n2 7.34285
R52 VGND.n7 VGND.n6 7.16028
R53 VGND.n2 VGND.n0 0.219268
R54 VGND VGND.n7 0.156488
R55 VGND.n7 VGND.n0 0.151269
R56 VNB.t0 VNB.t3 2240.42
R57 VNB.t4 VNB.t1 1316.54
R58 VNB VNB.t2 1120.21
R59 VNB.t2 VNB.t5 1097.11
R60 VNB.t3 VNB.t4 993.177
R61 VNB.t5 VNB.t0 993.177
R62 a_177_48.n3 a_177_48.n2 272.697
R63 a_177_48.n0 a_177_48.t5 261.747
R64 a_177_48.n1 a_177_48.t6 248.231
R65 a_177_48.n1 a_177_48.t4 211.418
R66 a_177_48.n0 a_177_48.t3 201.737
R67 a_177_48.n2 a_177_48.n0 196.424
R68 a_177_48.n2 a_177_48.t1 153.784
R69 a_177_48.n0 a_177_48.n1 50.751
R70 a_177_48.n3 a_177_48.t2 29.5505
R71 a_177_48.t0 a_177_48.n3 29.5505
R72 X.n1 X.n0 652.569
R73 X.n2 X.n1 185
R74 X.n3 X.n2 185
R75 X.n0 X.t3 26.3844
R76 X.n0 X.t2 26.3844
R77 X.n2 X.t1 22.7032
R78 X.n2 X.t0 22.7032
R79 X.n3 X 12.6066
R80 X.n1 X 4.84898
R81 X X.n3 1.74595
R82 a_582_368.t0 a_582_368.t1 70.9205
R83 A1.n0 A1.t0 260.012
R84 A1.n0 A1.t1 171.913
R85 A1 A1.n0 158.788
C0 VPB X 0.003827f
C1 A1 VPWR 0.047742f
C2 VGND A2 0.016534f
C3 VGND VPB 0.008411f
C4 VPB B1_N 0.048029f
C5 A1 A2 0.085865f
C6 VGND X 0.110817f
C7 A1 VPB 0.04068f
C8 VPWR A2 0.021572f
C9 B1_N X 0.001625f
C10 VPB VPWR 0.132132f
C11 VGND B1_N 0.016968f
C12 VPWR X 0.017627f
C13 A1 VGND 0.013108f
C14 VPB A2 0.032624f
C15 VGND VPWR 0.065639f
C16 VPWR B1_N 0.0099f
C17 VGND VNB 0.49597f
C18 A1 VNB 0.166018f
C19 A2 VNB 0.107226f
C20 X VNB 0.008189f
C21 B1_N VNB 0.191431f
C22 VPWR VNB 0.433021f
C23 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21ba_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21ba_1 VNB VPB VPWR VGND B1_N A2 A1 X
X0 a_116_392.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X1 VGND.t1 B1_N.t0 a_281_244.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.14495 pd=1.16 as=0.275 ps=2.1 w=0.55 l=0.15
X2 VPWR.t2 B1_N.t1 a_281_244.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.3108 ps=2.42 w=0.84 l=0.15
X3 VGND.t0 A1.t1 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.1824 ps=1.85 w=0.64 l=0.15
X4 a_200_392.t2 a_281_244.t2 a_27_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2176 pd=1.96 as=0.0944 ps=0.935 w=0.64 l=0.15
X5 a_200_392.t0 A2.t0 a_116_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t1 a_281_244.t3 a_200_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.21 ps=1.42 w=1 l=0.15
X7 a_27_74.t1 A2.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0944 pd=0.935 as=0.1344 ps=1.06 w=0.64 l=0.15
X8 X.t0 a_200_392.t3 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.231 ps=1.555 w=1.12 l=0.15
X9 X.t1 a_200_392.t4 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.14495 ps=1.16 w=0.74 l=0.15
R0 A1.n0 A1.t0 232.321
R1 A1.n1 A1.t1 164.111
R2 A1 A1.n0 153.656
R3 A1.n2 A1.n1 152
R4 A1.n1 A1.n0 46.8234
R5 A1 A1.n2 8.58403
R6 A1.n2 A1 2.5605
R7 VPWR.n1 VPWR.t1 820.029
R8 VPWR.n3 VPWR.n2 669.462
R9 VPWR.n7 VPWR.t0 251.702
R10 VPWR.n2 VPWR.t2 60.9767
R11 VPWR.n6 VPWR.n5 36.1417
R12 VPWR.n2 VPWR.t3 32.6589
R13 VPWR.n5 VPWR.n1 26.7299
R14 VPWR.n7 VPWR.n6 20.7064
R15 VPWR.n5 VPWR.n4 9.3005
R16 VPWR.n6 VPWR.n0 9.3005
R17 VPWR.n8 VPWR.n7 9.3005
R18 VPWR.n3 VPWR.n1 6.89086
R19 VPWR.n4 VPWR.n3 0.244332
R20 VPWR.n4 VPWR.n0 0.122949
R21 VPWR.n8 VPWR.n0 0.122949
R22 VPWR VPWR.n8 0.0617245
R23 a_116_392.t0 a_116_392.t1 53.1905
R24 VPB.t1 VPB.t3 640.995
R25 VPB.t3 VPB.t4 298.791
R26 VPB.t2 VPB.t1 291.13
R27 VPB VPB.t0 257.93
R28 VPB.t0 VPB.t2 214.517
R29 B1_N.n0 B1_N.t1 240.732
R30 B1_N B1_N.n0 158.788
R31 B1_N.n0 B1_N.t0 147.814
R32 a_281_244.t0 a_281_244.n1 763.032
R33 a_281_244.n0 a_281_244.t3 287.676
R34 a_281_244.n1 a_281_244.n0 253.387
R35 a_281_244.n1 a_281_244.t1 250.751
R36 a_281_244.n0 a_281_244.t2 170.308
R37 VGND.n2 VGND.n0 211.155
R38 VGND.n2 VGND.n1 125.219
R39 VGND.n1 VGND.t1 51.509
R40 VGND.n0 VGND.t3 39.3755
R41 VGND.n0 VGND.t0 39.3755
R42 VGND.n1 VGND.t2 28.7381
R43 VGND VGND.n2 0.200367
R44 VNB.t4 VNB.t1 2910.24
R45 VNB.t1 VNB.t2 1316.54
R46 VNB.t0 VNB.t3 1316.54
R47 VNB VNB.t0 1143.31
R48 VNB.t3 VNB.t4 1027.82
R49 a_27_74.t0 a_27_74.n0 279.127
R50 a_27_74.n0 a_27_74.t2 29.063
R51 a_27_74.n0 a_27_74.t1 26.2505
R52 a_200_392.n1 a_200_392.n0 312.43
R53 a_200_392.n0 a_200_392.t3 258.233
R54 a_200_392.n0 a_200_392.t4 209.764
R55 a_200_392.n1 a_200_392.t2 209.514
R56 a_200_392.n2 a_200_392.n1 208.197
R57 a_200_392.t0 a_200_392.n2 43.3405
R58 a_200_392.n2 a_200_392.t1 39.4005
R59 A2.n0 A2.t0 231.629
R60 A2.n1 A2.t1 165.488
R61 A2 A2.n0 153.468
R62 A2.n2 A2.n1 152
R63 A2.n1 A2.n0 49.6611
R64 A2 A2.n2 7.6005
R65 A2.n2 A2 2.26717
R66 X.n1 X 589.444
R67 X.n1 X.n0 585
R68 X.n2 X.n1 585
R69 X X.t1 206.069
R70 X.n1 X.t0 26.3844
R71 X X.n2 11.9116
R72 X X.n0 10.3116
R73 X X.n0 2.84494
R74 X.n2 X 1.24494
C0 A1 VPWR 0.054993f
C1 VPB B1_N 0.042034f
C2 VPWR X 0.070036f
C3 A2 VGND 0.015789f
C4 VPB VPWR 0.137003f
C5 VPWR B1_N 0.00907f
C6 A1 A2 0.108315f
C7 A1 VGND 0.014873f
C8 X VGND 0.096634f
C9 VPB A2 0.042513f
C10 VPB VGND 0.010684f
C11 B1_N VGND 0.016853f
C12 VPB A1 0.047319f
C13 VPB X 0.014492f
C14 A2 VPWR 0.022234f
C15 B1_N X 0.006303f
C16 VPWR VGND 0.063349f
C17 VGND VNB 0.501821f
C18 X VNB 0.113859f
C19 B1_N VNB 0.121771f
C20 VPWR VNB 0.426054f
C21 A2 VNB 0.117312f
C22 A1 VNB 0.184577f
C23 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21ai_4 VNB VPB VPWR VGND Y A1 A2 B1
X0 a_116_368.t6 A1.t0 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t7 B1.t0 a_27_74.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t3 A2.t0 a_116_368.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 Y.t6 B1.t1 a_27_74.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t3 A2.t1 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VGND.t7 A1.t1 a_27_74.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_27_74.t9 B1.t2 Y.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_27_74.t0 A2.t2 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_27_74.t8 B1.t3 Y.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VGND.t1 A2.t3 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11285 ps=1.045 w=0.74 l=0.15
X10 VPWR.t0 B1.t4 Y.t9 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.4256 pd=3 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t8 B1.t5 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_27_74.t4 A1.t2 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.10915 ps=1.035 w=0.74 l=0.15
X13 VPWR.t4 A1.t3 a_116_368.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_27_74.t2 A2.t4 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_116_368.t4 A1.t4 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VPWR.t2 A1.t5 a_116_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_27_74.t7 A1.t6 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 Y.t0 A2.t5 a_116_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_116_368.t1 A2.t6 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X20 a_116_368.t2 A2.t7 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X21 VGND.t4 A1.t7 a_27_74.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A1.n3 A1.t3 242.875
R1 A1.n5 A1.t4 234.841
R2 A1.n8 A1.t5 234.841
R3 A1.n1 A1.t0 234.841
R4 A1.n1 A1.t1 187.834
R5 A1.n9 A1.t6 186.374
R6 A1.n6 A1.t7 186.374
R7 A1.n3 A1.t2 186.374
R8 A1.n11 A1.n2 165.189
R9 A1.n4 A1 152.975
R10 A1.n11 A1.n10 152
R11 A1.n7 A1.n0 152
R12 A1.n8 A1.n7 48.9308
R13 A1.n9 A1.n2 46.0096
R14 A1.n5 A1.n4 32.8641
R15 A1.n4 A1.n3 24.8308
R16 A1.n2 A1.n1 15.3369
R17 A1.n7 A1.n6 9.49444
R18 A1 A1.n0 8.48746
R19 A1.n6 A1.n5 7.30353
R20 A1 A1.n11 6.07165
R21 A1 A1.n0 4.87007
R22 A1.n10 A1.n9 3.65202
R23 A1.n10 A1.n8 0.730803
R24 VPWR.n5 VPWR.t0 820.899
R25 VPWR.n4 VPWR.n3 611.88
R26 VPWR.n9 VPWR.n1 331.5
R27 VPWR.n11 VPWR.t5 259.171
R28 VPWR.n8 VPWR.n2 36.1417
R29 VPWR.n10 VPWR.n9 34.6358
R30 VPWR.n11 VPWR.n10 26.7299
R31 VPWR.n1 VPWR.t3 26.3844
R32 VPWR.n1 VPWR.t2 26.3844
R33 VPWR.n3 VPWR.t1 26.3844
R34 VPWR.n3 VPWR.t4 26.3844
R35 VPWR.n4 VPWR.n2 23.7181
R36 VPWR.n6 VPWR.n2 9.3005
R37 VPWR.n8 VPWR.n7 9.3005
R38 VPWR.n10 VPWR.n0 9.3005
R39 VPWR.n12 VPWR.n11 9.3005
R40 VPWR.n5 VPWR.n4 7.01265
R41 VPWR.n9 VPWR.n8 1.50638
R42 VPWR.n6 VPWR.n5 0.535129
R43 VPWR.n7 VPWR.n6 0.122949
R44 VPWR.n7 VPWR.n0 0.122949
R45 VPWR.n12 VPWR.n0 0.122949
R46 VPWR VPWR.n12 0.0617245
R47 a_116_368.n2 a_116_368.t7 315.435
R48 a_116_368.n1 a_116_368.n0 305.901
R49 a_116_368.n1 a_116_368.t2 301.389
R50 a_116_368.n5 a_116_368.n4 255.745
R51 a_116_368.n4 a_116_368.n3 195.787
R52 a_116_368.n4 a_116_368.n2 138.744
R53 a_116_368.n2 a_116_368.n1 72.7942
R54 a_116_368.n3 a_116_368.t5 26.3844
R55 a_116_368.n3 a_116_368.t4 26.3844
R56 a_116_368.n0 a_116_368.t0 26.3844
R57 a_116_368.n0 a_116_368.t1 26.3844
R58 a_116_368.n5 a_116_368.t3 26.3844
R59 a_116_368.t6 a_116_368.n5 26.3844
R60 VPB.t3 VPB.t9 559.274
R61 VPB VPB.t8 257.93
R62 VPB.t9 VPB.t1 255.376
R63 VPB.t0 VPB.t2 229.839
R64 VPB.t1 VPB.t0 229.839
R65 VPB.t4 VPB.t3 229.839
R66 VPB.t7 VPB.t4 229.839
R67 VPB.t6 VPB.t7 229.839
R68 VPB.t5 VPB.t6 229.839
R69 VPB.t8 VPB.t5 229.839
R70 B1.n1 B1.t2 266.971
R71 B1.n0 B1.t4 261.62
R72 B1.n5 B1.t5 261.62
R73 B1.n3 B1.n2 163.762
R74 B1.n5 B1.t1 152.898
R75 B1.n4 B1.n3 152
R76 B1.n7 B1.n6 152
R77 B1.n4 B1.t3 142.994
R78 B1.n1 B1.t0 142.994
R79 B1.n6 B1.n4 44.8991
R80 B1.n2 B1.n0 32.3539
R81 B1.n4 B1.n0 12.5457
R82 B1.n2 B1.n1 11.8854
R83 B1 B1.n7 8.47618
R84 B1.n7 B1 8.13023
R85 B1.n3 B1 3.63293
R86 B1.n6 B1.n5 1.98132
R87 a_27_74.n2 a_27_74.t5 211.385
R88 a_27_74.t0 a_27_74.n9 210.411
R89 a_27_74.n6 a_27_74.n5 185
R90 a_27_74.n9 a_27_74.n0 103.65
R91 a_27_74.n2 a_27_74.n1 98.8814
R92 a_27_74.n4 a_27_74.n3 86.4329
R93 a_27_74.n8 a_27_74.n7 84.741
R94 a_27_74.n9 a_27_74.n8 83.6621
R95 a_27_74.n8 a_27_74.n6 81.5983
R96 a_27_74.n6 a_27_74.n4 74.8264
R97 a_27_74.n4 a_27_74.n2 73.2298
R98 a_27_74.n7 a_27_74.t9 26.7573
R99 a_27_74.n7 a_27_74.t1 22.7032
R100 a_27_74.n5 a_27_74.t11 22.7032
R101 a_27_74.n5 a_27_74.t8 22.7032
R102 a_27_74.n3 a_27_74.t10 22.7032
R103 a_27_74.n3 a_27_74.t4 22.7032
R104 a_27_74.n1 a_27_74.t6 22.7032
R105 a_27_74.n1 a_27_74.t7 22.7032
R106 a_27_74.n0 a_27_74.t3 22.7032
R107 a_27_74.n0 a_27_74.t2 22.7032
R108 Y.n4 Y.n0 619.347
R109 Y.n3 Y.n1 342.868
R110 Y.n3 Y.n2 299.95
R111 Y.n7 Y.n5 243.353
R112 Y.n7 Y.n6 190.614
R113 Y Y.n7 45.4874
R114 Y.n2 Y.t3 35.1791
R115 Y.n0 Y.t9 26.3844
R116 Y.n0 Y.t8 26.3844
R117 Y.n1 Y.t2 26.3844
R118 Y.n1 Y.t0 26.3844
R119 Y.n2 Y.t1 26.3844
R120 Y.n6 Y.t5 22.7032
R121 Y.n6 Y.t7 22.7032
R122 Y.n5 Y.t4 22.7032
R123 Y.n5 Y.t6 22.7032
R124 Y.n4 Y.n3 20.637
R125 Y Y.n4 13.1373
R126 VNB VNB.t7 1143.31
R127 VNB.t9 VNB.t1 1050.92
R128 VNB.t4 VNB.t6 1027.82
R129 VNB.t3 VNB.t0 993.177
R130 VNB.t2 VNB.t3 993.177
R131 VNB.t1 VNB.t2 993.177
R132 VNB.t11 VNB.t9 993.177
R133 VNB.t8 VNB.t11 993.177
R134 VNB.t10 VNB.t8 993.177
R135 VNB.t6 VNB.t10 993.177
R136 VNB.t5 VNB.t4 993.177
R137 VNB.t7 VNB.t5 993.177
R138 A2.n3 A2.t0 230.861
R139 A2.n0 A2.t7 214.758
R140 A2.n1 A2.t5 214.758
R141 A2.n5 A2.t6 214.758
R142 A2.n0 A2.t2 197.941
R143 A2.n3 A2.t3 196.013
R144 A2.n6 A2.t4 196.013
R145 A2.n11 A2.t1 196.013
R146 A2.n13 A2.n12 152
R147 A2.n10 A2.n9 152
R148 A2.n8 A2.n7 152
R149 A2.n4 A2.n2 152
R150 A2.n7 A2.n1 42.4165
R151 A2.n12 A2.n11 40.4885
R152 A2.n5 A2.n4 28.2778
R153 A2.n4 A2.n3 19.9232
R154 A2.n12 A2.n0 12.8538
R155 A2.n8 A2.n2 10.1214
R156 A2.n9 A2 9.97259
R157 A2 A2.n13 8.48422
R158 A2.n7 A2.n6 8.35517
R159 A2.n6 A2.n5 7.06983
R160 A2.n13 A2 5.80515
R161 A2.n9 A2 4.31678
R162 A2.n2 A2 4.0191
R163 A2.n11 A2.n10 3.21383
R164 A2.n10 A2.n1 1.28583
R165 A2 A2.n8 0.149337
R166 VGND.n7 VGND.n6 213.62
R167 VGND.n18 VGND.n17 209.048
R168 VGND.n5 VGND.n4 208.079
R169 VGND.n15 VGND.n2 206.333
R170 VGND.n10 VGND.n9 36.1417
R171 VGND.n11 VGND.n10 36.1417
R172 VGND.n11 VGND.n1 36.1417
R173 VGND.n9 VGND.n5 32.0005
R174 VGND.n15 VGND.n1 32.0005
R175 VGND.n2 VGND.t6 25.1356
R176 VGND.n18 VGND.n16 24.4711
R177 VGND.n6 VGND.t2 22.7032
R178 VGND.n6 VGND.t3 22.7032
R179 VGND.n4 VGND.t0 22.7032
R180 VGND.n4 VGND.t1 22.7032
R181 VGND.n2 VGND.t4 22.7032
R182 VGND.n17 VGND.t5 22.7032
R183 VGND.n17 VGND.t7 22.7032
R184 VGND.n16 VGND.n15 15.4358
R185 VGND.n9 VGND.n8 9.3005
R186 VGND.n10 VGND.n3 9.3005
R187 VGND.n12 VGND.n11 9.3005
R188 VGND.n13 VGND.n1 9.3005
R189 VGND.n15 VGND.n14 9.3005
R190 VGND.n16 VGND.n0 9.3005
R191 VGND.n19 VGND.n18 7.19894
R192 VGND.n7 VGND.n5 6.08503
R193 VGND.n8 VGND.n7 0.64127
R194 VGND VGND.n19 0.156997
R195 VGND.n19 VGND.n0 0.150766
R196 VGND.n8 VGND.n3 0.122949
R197 VGND.n12 VGND.n3 0.122949
R198 VGND.n13 VGND.n12 0.122949
R199 VGND.n14 VGND.n13 0.122949
R200 VGND.n14 VGND.n0 0.122949
C0 B1 Y 0.224308f
C1 A2 VPWR 0.025913f
C2 Y VPB 0.016122f
C3 VPWR A1 0.065913f
C4 B1 VGND 0.022177f
C5 VPB VGND 0.008916f
C6 B1 VPWR 0.037388f
C7 VPWR VPB 0.157412f
C8 Y VGND 0.022687f
C9 B1 A2 0.030476f
C10 A2 VPB 0.145527f
C11 B1 A1 0.082555f
C12 VPB A1 0.138768f
C13 VPWR Y 0.04867f
C14 VPWR VGND 0.092871f
C15 B1 VPB 0.090327f
C16 A2 Y 0.199409f
C17 Y A1 0.006032f
C18 A2 VGND 0.072549f
C19 A1 VGND 0.067837f
C20 VGND VNB 0.679414f
C21 Y VNB 0.027128f
C22 VPWR VNB 0.585288f
C23 A2 VNB 0.449649f
C24 B1 VNB 0.342522f
C25 A1 VNB 0.437536f
C26 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21ai_2 VNB VPB VPWR VGND B1 A2 A1 Y
X0 Y.t1 B1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_116_368.t1 A1.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t0 A1.t1 a_116_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3 a_27_74.t1 B1.t1 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.11655 ps=1.055 w=0.74 l=0.15
X4 a_27_74.t5 A1.t2 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.12395 ps=1.075 w=0.74 l=0.15
X5 VGND.t2 A1.t3 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_116_368.t3 A2.t0 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X7 VGND.t1 A2.t1 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.12395 pd=1.075 as=0.10915 ps=1.035 w=0.74 l=0.15
X8 Y.t3 B1.t2 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.12025 ps=1.065 w=0.74 l=0.15
X9 Y.t4 A2.t2 a_116_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_27_74.t2 A2.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 VPWR.t1 B1.t3 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B1.n0 B1.t0 245.805
R1 B1.n1 B1.t3 244.214
R2 B1.n0 B1.t2 204.337
R3 B1.n2 B1.t1 182.81
R4 B1 B1.n2 165.135
R5 B1.n1 B1.n0 87.6133
R6 B1.n2 B1.n1 11.8622
R7 VPWR.n3 VPWR.n2 611.88
R8 VPWR.n9 VPWR.t3 349.788
R9 VPWR.n4 VPWR.t1 266.168
R10 VPWR.n7 VPWR.n1 36.1417
R11 VPWR.n8 VPWR.n7 36.1417
R12 VPWR.n3 VPWR.n1 31.2476
R13 VPWR.n9 VPWR.n8 26.7299
R14 VPWR.n2 VPWR.t2 26.3844
R15 VPWR.n2 VPWR.t0 26.3844
R16 VPWR.n5 VPWR.n1 9.3005
R17 VPWR.n7 VPWR.n6 9.3005
R18 VPWR.n8 VPWR.n0 9.3005
R19 VPWR.n10 VPWR.n9 9.3005
R20 VPWR.n4 VPWR.n3 6.59649
R21 VPWR.n5 VPWR.n4 0.612104
R22 VPWR.n6 VPWR.n5 0.122949
R23 VPWR.n6 VPWR.n0 0.122949
R24 VPWR.n10 VPWR.n0 0.122949
R25 VPWR VPWR.n10 0.0617245
R26 Y.n1 Y.n0 674.828
R27 Y.n5 Y.n4 585
R28 Y.n4 Y.n3 290.577
R29 Y Y.n2 245.529
R30 Y.n0 Y.t4 35.1791
R31 Y.n2 Y.t3 27.5681
R32 Y.n4 Y.t0 26.3844
R33 Y.n4 Y.t1 26.3844
R34 Y.n0 Y.t5 26.3844
R35 Y.n2 Y.t2 23.514
R36 Y Y.n5 15.882
R37 Y.n3 Y.n1 7.94658
R38 Y.n3 Y 6.82988
R39 Y Y.n1 2.60791
R40 Y.n5 Y 1.65976
R41 VPB VPB.t3 257.93
R42 VPB.t5 VPB.t0 255.376
R43 VPB.t4 VPB.t5 255.376
R44 VPB.t2 VPB.t1 229.839
R45 VPB.t0 VPB.t2 229.839
R46 VPB.t3 VPB.t4 229.839
R47 A1 A1.n0 270.712
R48 A1.n1 A1.t1 250.909
R49 A1.n0 A1.t0 250.909
R50 A1.n1 A1.t2 220.113
R51 A1.n0 A1.t3 220.113
R52 A1 A1.n1 153.601
R53 a_116_368.n1 a_116_368.n0 945.361
R54 a_116_368.n0 a_116_368.t3 35.1791
R55 a_116_368.n0 a_116_368.t0 26.3844
R56 a_116_368.n1 a_116_368.t2 26.3844
R57 a_116_368.t1 a_116_368.n1 26.3844
R58 a_27_74.t1 a_27_74.n3 203.608
R59 a_27_74.n1 a_27_74.t4 200.344
R60 a_27_74.n1 a_27_74.n0 104.579
R61 a_27_74.n3 a_27_74.n2 87.0786
R62 a_27_74.n3 a_27_74.n1 68.7017
R63 a_27_74.n2 a_27_74.t0 30.0005
R64 a_27_74.n0 a_27_74.t3 25.1356
R65 a_27_74.n2 a_27_74.t5 22.7032
R66 a_27_74.n0 a_27_74.t2 22.7032
R67 VNB.t4 VNB.t2 1154.86
R68 VNB VNB.t4 1143.31
R69 VNB.t3 VNB.t5 1120.21
R70 VNB.t5 VNB.t0 1097.11
R71 VNB.t0 VNB.t1 1074.02
R72 VNB.t2 VNB.t3 1027.82
R73 VGND.n2 VGND.n0 216.446
R74 VGND.n2 VGND.n1 216.231
R75 VGND.n1 VGND.t2 34.0546
R76 VGND.n0 VGND.t1 31.6221
R77 VGND.n0 VGND.t3 22.7032
R78 VGND.n1 VGND.t0 22.7032
R79 VGND VGND.n2 0.536269
R80 A2.n1 A2.t2 232.65
R81 A2.n0 A2.t0 228.47
R82 A2.n0 A2.t1 196.013
R83 A2.n1 A2.t3 196.013
R84 A2 A2.n2 67.8006
R85 A2.n2 A2.n0 34.8513
R86 A2.n2 A2.n1 23.3684
C0 VPB VPWR 0.103867f
C1 A1 B1 0.067148f
C2 A2 VGND 0.034189f
C3 B1 VPWR 0.055317f
C4 Y VGND 0.009385f
C5 VPB B1 0.073204f
C6 A2 Y 0.017153f
C7 A1 VGND 0.035131f
C8 A1 A2 0.240997f
C9 VPWR VGND 0.055642f
C10 A2 VPWR 0.011478f
C11 A1 Y 0.170243f
C12 VPB VGND 0.005895f
C13 VPB A2 0.065864f
C14 B1 VGND 0.016517f
C15 VPWR Y 0.204785f
C16 A1 VPWR 0.056487f
C17 VPB Y 0.006831f
C18 VPB A1 0.076065f
C19 B1 Y 0.104983f
C20 VGND VNB 0.426767f
C21 Y VNB 0.025526f
C22 VPWR VNB 0.415511f
C23 B1 VNB 0.26721f
C24 A2 VNB 0.196758f
C25 A1 VNB 0.270875f
C26 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21bai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21bai_4 VNB VPB VPWR VGND Y A1 A2 B1_N
X0 a_27_74.t8 A2.t0 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1889 ps=1.36 w=0.74 l=0.15
X1 VGND.t0 A1.t0 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t7 a_828_48.t3 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 VPWR.t5 A1.t1 a_28_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4 a_28_368.t7 A2.t1 Y.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X5 VGND.t8 A1.t2 a_27_74.t9 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 Y.t9 a_828_48.t4 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X7 VGND.t5 A2.t2 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1889 pd=1.36 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_27_74.t10 a_828_48.t5 Y.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 Y.t2 A2.t3 a_28_368.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VPWR.t0 B1_N.t0 a_828_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X11 a_28_368.t5 A2.t4 Y.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VGND.t7 B1_N.t1 a_828_48.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 a_828_48.t1 B1_N.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2478 ps=2.27 w=0.84 l=0.15
X14 a_27_74.t6 A2.t5 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 Y.t0 A2.t6 a_28_368.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_28_368.t2 A1.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 VPWR.t3 A1.t4 a_28_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 Y.t5 a_828_48.t6 a_27_74.t11 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X19 VPWR.t6 a_828_48.t7 Y.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.3304 ps=2.83 w=1.12 l=0.15
X20 a_27_74.t2 A1.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 a_28_368.t0 A1.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_27_74.t1 a_828_48.t8 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X23 a_27_74.t3 A1.t7 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X24 VGND.t3 A2.t7 a_27_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A2.n2 A2.t6 292.223
R1 A2.n8 A2.t3 226.809
R2 A2.n4 A2.t4 226.809
R3 A2.n2 A2.t7 213.228
R4 A2.n1 A2.t1 206.865
R5 A2.n1 A2.t0 197.465
R6 A2.n7 A2.t2 196.013
R7 A2.n3 A2.t5 196.013
R8 A2.n10 A2.n9 152
R9 A2.n7 A2.n0 152
R10 A2.n6 A2.n5 152
R11 A2.n3 A2.n2 81.6484
R12 A2.n7 A2.n6 49.6611
R13 A2.n9 A2.n8 37.246
R14 A2.n9 A2.n1 35.0616
R15 A2.n8 A2.n7 12.4157
R16 A2.n10 A2.n0 10.1214
R17 A2.n4 A2.n3 9.49444
R18 A2.n5 A2 7.44236
R19 A2.n5 A2 6.84701
R20 A2.n6 A2.n4 3.65202
R21 A2 A2.n0 2.67957
R22 A2 A2.n10 1.48887
R23 VGND.n6 VGND.n5 212.477
R24 VGND.n9 VGND.n8 211.183
R25 VGND.n13 VGND.n2 211.183
R26 VGND.n16 VGND.n15 211.183
R27 VGND.n4 VGND.t7 177.669
R28 VGND.n9 VGND.n7 35.7652
R29 VGND.n5 VGND.t6 35.6762
R30 VGND.n5 VGND.t5 35.6762
R31 VGND.n15 VGND.t2 30.8113
R32 VGND.n13 VGND.n1 28.2358
R33 VGND.n16 VGND.n14 24.4711
R34 VGND.n8 VGND.t4 22.7032
R35 VGND.n8 VGND.t3 22.7032
R36 VGND.n2 VGND.t1 22.7032
R37 VGND.n2 VGND.t0 22.7032
R38 VGND.n15 VGND.t8 22.7032
R39 VGND.n14 VGND.n13 19.2005
R40 VGND.n9 VGND.n1 11.6711
R41 VGND.n7 VGND.n6 10.1652
R42 VGND.n14 VGND.n0 9.3005
R43 VGND.n13 VGND.n12 9.3005
R44 VGND.n11 VGND.n1 9.3005
R45 VGND.n10 VGND.n9 9.3005
R46 VGND.n7 VGND.n3 9.3005
R47 VGND.n6 VGND.n4 8.7798
R48 VGND.n17 VGND.n16 7.19894
R49 VGND VGND.n17 0.156997
R50 VGND.n17 VGND.n0 0.150766
R51 VGND.n4 VGND.n3 0.149535
R52 VGND.n10 VGND.n3 0.122949
R53 VGND.n11 VGND.n10 0.122949
R54 VGND.n12 VGND.n11 0.122949
R55 VGND.n12 VGND.n0 0.122949
R56 a_27_74.n2 a_27_74.t9 214.175
R57 a_27_74.n7 a_27_74.t1 190.583
R58 a_27_74.n7 a_27_74.n6 185
R59 a_27_74.n9 a_27_74.n8 185
R60 a_27_74.n2 a_27_74.n1 103.65
R61 a_27_74.n3 a_27_74.n0 103.65
R62 a_27_74.n5 a_27_74.n4 92.8625
R63 a_27_74.n5 a_27_74.n3 70.0708
R64 a_27_74.n3 a_27_74.n2 64.7534
R65 a_27_74.n8 a_27_74.n7 63.9487
R66 a_27_74.n8 a_27_74.n5 63.557
R67 a_27_74.n6 a_27_74.t10 34.0546
R68 a_27_74.n9 a_27_74.t11 34.0546
R69 a_27_74.n4 a_27_74.t7 22.7032
R70 a_27_74.n4 a_27_74.t6 22.7032
R71 a_27_74.n1 a_27_74.t0 22.7032
R72 a_27_74.n1 a_27_74.t3 22.7032
R73 a_27_74.n0 a_27_74.t5 22.7032
R74 a_27_74.n0 a_27_74.t2 22.7032
R75 a_27_74.n6 a_27_74.t4 22.7032
R76 a_27_74.t8 a_27_74.n9 22.7032
R77 VNB.t1 VNB.t9 2448.29
R78 VNB.t7 VNB.t8 1362.73
R79 VNB.t4 VNB.t1 1154.86
R80 VNB.t11 VNB.t4 1154.86
R81 VNB.t8 VNB.t12 1154.86
R82 VNB VNB.t10 1143.31
R83 VNB.t10 VNB.t3 1108.66
R84 VNB.t12 VNB.t11 993.177
R85 VNB.t6 VNB.t7 993.177
R86 VNB.t5 VNB.t6 993.177
R87 VNB.t2 VNB.t5 993.177
R88 VNB.t0 VNB.t2 993.177
R89 VNB.t3 VNB.t0 993.177
R90 A1.n0 A1.t3 283.041
R91 A1.n1 A1.t4 226.809
R92 A1.n8 A1.t6 226.809
R93 A1.n3 A1.t1 226.809
R94 A1.n3 A1.t2 198.204
R95 A1.n0 A1.t5 196.013
R96 A1.n9 A1.t7 196.013
R97 A1.n2 A1.t0 196.013
R98 A1.n11 A1.n10 152
R99 A1.n7 A1.n6 152
R100 A1.n5 A1.n4 152
R101 A1.n1 A1.n0 120.793
R102 A1.n7 A1.n4 49.6611
R103 A1.n10 A1.n9 42.3581
R104 A1.n10 A1.n2 20.449
R105 A1.n5 A1 12.8005
R106 A1.n4 A1.n3 10.955
R107 A1 A1.n11 9.82376
R108 A1.n6 A1 8.63306
R109 A1.n6 A1 5.65631
R110 A1.n8 A1.n7 5.11262
R111 A1.n11 A1 4.46562
R112 A1.n9 A1.n8 2.19141
R113 A1 A1.n5 1.48887
R114 A1.n2 A1.n1 0.730803
R115 a_828_48.n12 a_828_48.n11 363.481
R116 a_828_48.n3 a_828_48.t6 242.754
R117 a_828_48.n8 a_828_48.t4 226.809
R118 a_828_48.n1 a_828_48.t7 226.809
R119 a_828_48.n9 a_828_48.t8 209.16
R120 a_828_48.n2 a_828_48.t5 196.013
R121 a_828_48.n6 a_828_48.t3 196.013
R122 a_828_48.n11 a_828_48.t2 188.274
R123 a_828_48.n4 a_828_48.n3 165.189
R124 a_828_48.n5 a_828_48.n4 152
R125 a_828_48.n7 a_828_48.n0 152
R126 a_828_48.n10 a_828_48.n9 152
R127 a_828_48.n9 a_828_48.n8 46.7399
R128 a_828_48.n6 a_828_48.n5 39.4369
R129 a_828_48.t0 a_828_48.n12 35.1791
R130 a_828_48.n12 a_828_48.t1 35.1791
R131 a_828_48.n2 a_828_48.n1 18.2581
R132 a_828_48.n3 a_828_48.n2 16.0672
R133 a_828_48.n5 a_828_48.n1 15.3369
R134 a_828_48.n10 a_828_48.n0 13.1884
R135 a_828_48.n4 a_828_48.n0 13.1884
R136 a_828_48.n11 a_828_48.n10 12.6066
R137 a_828_48.n7 a_828_48.n6 10.2247
R138 a_828_48.n8 a_828_48.n7 2.92171
R139 Y.n2 Y.n0 351.899
R140 Y.n2 Y.n1 297.598
R141 Y.n3 Y.t9 280.557
R142 Y.n7 Y.n5 248.173
R143 Y.n3 Y.t8 229.291
R144 Y.n7 Y.n6 185
R145 Y.n1 Y.t2 35.1791
R146 Y.n5 Y.t7 34.0546
R147 Y.n0 Y.t1 26.3844
R148 Y.n0 Y.t0 26.3844
R149 Y.n1 Y.t3 26.3844
R150 Y Y.n4 25.3222
R151 Y.n4 Y.n2 23.7181
R152 Y.n6 Y.t6 22.7032
R153 Y.n6 Y.t5 22.7032
R154 Y.n5 Y.t4 22.7032
R155 Y Y.n7 15.2813
R156 Y.n4 Y.n3 14.1995
R157 a_28_368.n4 a_28_368.t7 389.12
R158 a_28_368.n5 a_28_368.n4 302.74
R159 a_28_368.n1 a_28_368.t3 281.322
R160 a_28_368.n1 a_28_368.n0 205.998
R161 a_28_368.n3 a_28_368.n2 183.916
R162 a_28_368.n4 a_28_368.n3 88.7484
R163 a_28_368.n3 a_28_368.n1 84.7995
R164 a_28_368.n2 a_28_368.t4 26.3844
R165 a_28_368.n2 a_28_368.t2 26.3844
R166 a_28_368.n0 a_28_368.t1 26.3844
R167 a_28_368.n0 a_28_368.t0 26.3844
R168 a_28_368.t6 a_28_368.n5 26.3844
R169 a_28_368.n5 a_28_368.t5 26.3844
R170 VPWR.n8 VPWR.t0 416.245
R171 VPWR.n9 VPWR.t1 358.584
R172 VPWR.n12 VPWR.n11 333.288
R173 VPWR.n26 VPWR.n1 323.406
R174 VPWR.n24 VPWR.n3 315.928
R175 VPWR.n13 VPWR.n10 36.1417
R176 VPWR.n17 VPWR.n6 36.1417
R177 VPWR.n18 VPWR.n17 36.1417
R178 VPWR.n19 VPWR.n18 36.1417
R179 VPWR.n19 VPWR.n4 36.1417
R180 VPWR.n23 VPWR.n4 36.1417
R181 VPWR.n12 VPWR.n6 32.7534
R182 VPWR.n11 VPWR.t7 29.0228
R183 VPWR.n26 VPWR.n25 28.6123
R184 VPWR.n24 VPWR.n23 27.1064
R185 VPWR.n1 VPWR.t2 26.3844
R186 VPWR.n1 VPWR.t5 26.3844
R187 VPWR.n3 VPWR.t4 26.3844
R188 VPWR.n3 VPWR.t3 26.3844
R189 VPWR.n11 VPWR.t6 26.3844
R190 VPWR.n10 VPWR.n9 25.224
R191 VPWR.n25 VPWR.n24 20.3299
R192 VPWR.n10 VPWR.n7 9.3005
R193 VPWR.n14 VPWR.n13 9.3005
R194 VPWR.n15 VPWR.n6 9.3005
R195 VPWR.n17 VPWR.n16 9.3005
R196 VPWR.n18 VPWR.n5 9.3005
R197 VPWR.n20 VPWR.n19 9.3005
R198 VPWR.n21 VPWR.n4 9.3005
R199 VPWR.n23 VPWR.n22 9.3005
R200 VPWR.n24 VPWR.n2 9.3005
R201 VPWR.n25 VPWR.n0 9.3005
R202 VPWR.n27 VPWR.n26 7.28976
R203 VPWR.n9 VPWR.n8 6.88165
R204 VPWR.n13 VPWR.n12 3.38874
R205 VPWR.n8 VPWR.n7 0.610715
R206 VPWR VPWR.n27 0.158192
R207 VPWR.n27 VPWR.n0 0.149586
R208 VPWR.n14 VPWR.n7 0.122949
R209 VPWR.n15 VPWR.n14 0.122949
R210 VPWR.n16 VPWR.n15 0.122949
R211 VPWR.n16 VPWR.n5 0.122949
R212 VPWR.n20 VPWR.n5 0.122949
R213 VPWR.n21 VPWR.n20 0.122949
R214 VPWR.n22 VPWR.n21 0.122949
R215 VPWR.n22 VPWR.n2 0.122949
R216 VPWR.n2 VPWR.n0 0.122949
R217 VPB.t9 VPB.t10 541.399
R218 VPB.t11 VPB.t1 515.861
R219 VPB VPB.t5 260.485
R220 VPB.t8 VPB.t9 255.376
R221 VPB.t10 VPB.t11 237.5
R222 VPB.t1 VPB.t0 229.839
R223 VPB.t7 VPB.t8 229.839
R224 VPB.t6 VPB.t7 229.839
R225 VPB.t4 VPB.t6 229.839
R226 VPB.t3 VPB.t4 229.839
R227 VPB.t2 VPB.t3 229.839
R228 VPB.t5 VPB.t2 229.839
R229 B1_N.n1 B1_N.t2 269.457
R230 B1_N.n0 B1_N.t0 230.022
R231 B1_N.n0 B1_N.t1 181.407
R232 B1_N.n2 B1_N.n1 152
R233 B1_N.n1 B1_N.n0 24.1005
R234 B1_N B1_N.n2 13.3823
R235 B1_N.n2 B1_N 5.23686
C0 B1_N VPB 0.116055f
C1 Y A2 0.199259f
C2 VGND A1 0.074568f
C3 VPWR VGND 0.115776f
C4 A1 A2 0.075138f
C5 VPWR A2 0.024676f
C6 Y A1 3.01e-19
C7 VGND VPB 0.013078f
C8 VPWR Y 0.299927f
C9 B1_N VGND 0.051982f
C10 VPB A2 0.140777f
C11 VPWR A1 0.078812f
C12 Y VPB 0.034166f
C13 B1_N Y 0.002952f
C14 VPB A1 0.136284f
C15 VPWR VPB 0.205126f
C16 B1_N VPWR 0.059005f
C17 VGND A2 0.058462f
C18 Y VGND 0.028205f
C19 VGND VNB 0.880137f
C20 Y VNB 0.024501f
C21 VPWR VNB 0.696098f
C22 B1_N VNB 0.196951f
C23 A2 VNB 0.409484f
C24 A1 VNB 0.44936f
C25 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21bai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21bai_2 VNB VPB VPWR VGND A1 A2 B1_N Y
X0 VGND.t4 A2.t0 a_225_74.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VGND.t0 B1_N.t0 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1824 ps=1.85 w=0.64 l=0.15
X2 a_225_74.t3 A1.t0 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 VGND.t1 A1.t1 a_225_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1406 pd=1.12 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 Y.t1 a_27_74.t2 a_225_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_225_74.t4 A2.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1406 ps=1.12 w=0.74 l=0.15
X6 VPWR.t4 B1_N.t1 a_27_74.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3364 pd=1.74 as=0.305 ps=2.61 w=1 l=0.15
X7 a_225_74.t1 a_27_74.t3 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t3 a_27_74.t4 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_507_368.t3 A2.t2 Y.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t2 a_27_74.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3364 ps=1.74 w=1.12 l=0.15
X11 Y.t4 A2.t3 a_507_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_507_368.t1 A1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2184 ps=1.51 w=1.12 l=0.15
X13 VPWR.t0 A1.t3 a_507_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1708 ps=1.425 w=1.12 l=0.15
R0 A2.n1 A2.t3 231.921
R1 A2.n0 A2.t2 226.809
R2 A2.n0 A2.t0 198.204
R3 A2.n1 A2.t1 196.013
R4 A2 A2.n2 154.006
R5 A2.n2 A2.n0 48.2005
R6 A2.n2 A2.n1 12.4157
R7 a_225_74.t0 a_225_74.n3 280.997
R8 a_225_74.n1 a_225_74.t3 202.476
R9 a_225_74.n1 a_225_74.n0 107.79
R10 a_225_74.n3 a_225_74.n2 88.3339
R11 a_225_74.n3 a_225_74.n1 69.0952
R12 a_225_74.n2 a_225_74.t1 34.0546
R13 a_225_74.n2 a_225_74.t2 22.7032
R14 a_225_74.n0 a_225_74.t5 22.7032
R15 a_225_74.n0 a_225_74.t4 22.7032
R16 VGND.n10 VGND.t0 237.433
R17 VGND.n5 VGND.n2 215.594
R18 VGND.n4 VGND.n3 211.183
R19 VGND.n8 VGND.n1 36.1417
R20 VGND.n9 VGND.n8 36.1417
R21 VGND.n3 VGND.t1 34.0546
R22 VGND.n4 VGND.n1 28.2358
R23 VGND.n3 VGND.t3 27.5681
R24 VGND.n10 VGND.n9 24.4711
R25 VGND.n2 VGND.t2 22.7032
R26 VGND.n2 VGND.t4 22.7032
R27 VGND.n6 VGND.n1 9.3005
R28 VGND.n8 VGND.n7 9.3005
R29 VGND.n9 VGND.n0 9.3005
R30 VGND.n11 VGND.n10 7.19894
R31 VGND.n5 VGND.n4 6.39688
R32 VGND.n6 VGND.n5 0.607862
R33 VGND VGND.n11 0.156997
R34 VGND.n11 VGND.n0 0.150766
R35 VGND.n7 VGND.n6 0.122949
R36 VGND.n7 VGND.n0 0.122949
R37 VNB.t2 VNB.t0 2286.61
R38 VNB.t3 VNB.t5 1224.15
R39 VNB.t1 VNB.t3 1154.86
R40 VNB VNB.t2 1143.31
R41 VNB.t6 VNB.t4 993.177
R42 VNB.t5 VNB.t6 993.177
R43 VNB.t0 VNB.t1 993.177
R44 B1_N.n0 B1_N.t0 233.576
R45 B1_N.n0 B1_N.t1 229.023
R46 B1_N B1_N.n0 154.22
R47 a_27_74.t0 a_27_74.n3 293.498
R48 a_27_74.n2 a_27_74.t5 261.62
R49 a_27_74.n3 a_27_74.n2 253.487
R50 a_27_74.n0 a_27_74.t4 247.881
R51 a_27_74.n0 a_27_74.t3 154.976
R52 a_27_74.n1 a_27_74.t2 154.24
R53 a_27_74.n3 a_27_74.t1 145.45
R54 a_27_74.n1 a_27_74.n0 66.3208
R55 a_27_74.n2 a_27_74.n1 2.19141
R56 A1.n2 A1.n0 261.738
R57 A1.n1 A1.t3 258.942
R58 A1.n0 A1.t2 250.909
R59 A1.n0 A1.t1 220.113
R60 A1.n1 A1.t0 210.474
R61 A1.n2 A1.n1 163.249
R62 A1 A1.n2 3.89615
R63 A1.n2 A1 3.29747
R64 Y.n2 Y.n0 689.341
R65 Y Y.n3 205.602
R66 Y.n2 Y.n1 194.364
R67 Y.n0 Y.t5 26.3844
R68 Y.n0 Y.t4 26.3844
R69 Y.n1 Y.t3 26.3844
R70 Y.n1 Y.t2 26.3844
R71 Y.n3 Y.t0 22.7032
R72 Y.n3 Y.t1 22.7032
R73 Y Y.n2 11.0417
R74 VPWR.n4 VPWR.n3 602.817
R75 VPWR.n2 VPWR.t0 266.877
R76 VPWR.n1 VPWR.n0 223.696
R77 VPWR.n0 VPWR.t4 77.8155
R78 VPWR.n3 VPWR.t1 38.6969
R79 VPWR.n0 VPWR.t2 36.5101
R80 VPWR.n3 VPWR.t3 29.9023
R81 VPWR.n5 VPWR.n1 25.977
R82 VPWR.n5 VPWR.n4 22.5887
R83 VPWR.n6 VPWR.n5 9.3005
R84 VPWR.n4 VPWR.n2 7.03002
R85 VPWR.n7 VPWR.n1 7.02605
R86 VPWR VPWR.n7 0.272696
R87 VPWR.n6 VPWR.n2 0.172977
R88 VPWR.n7 VPWR.n6 0.158067
R89 VPB.t4 VPB.t2 393.281
R90 VPB VPB.t4 357.527
R91 VPB.t3 VPB.t1 275.807
R92 VPB.t6 VPB.t0 232.393
R93 VPB.t5 VPB.t6 229.839
R94 VPB.t1 VPB.t5 229.839
R95 VPB.t2 VPB.t3 229.839
R96 a_507_368.n1 a_507_368.n0 938.424
R97 a_507_368.n0 a_507_368.t0 27.2639
R98 a_507_368.n0 a_507_368.t3 26.3844
R99 a_507_368.n1 a_507_368.t2 26.3844
R100 a_507_368.t1 a_507_368.n1 26.3844
C0 A2 Y 0.013408f
C1 VPB VPWR 0.127493f
C2 A1 VGND 0.03429f
C3 A2 VPWR 0.012451f
C4 VPB A2 0.059481f
C5 Y VGND 0.011656f
C6 B1_N VGND 0.018645f
C7 A1 Y 0.136365f
C8 VPWR VGND 0.072935f
C9 B1_N Y 0.00772f
C10 VPB VGND 0.007533f
C11 A1 VPWR 0.076431f
C12 VPB A1 0.07388f
C13 A2 VGND 0.034432f
C14 VPWR Y 0.215682f
C15 B1_N VPWR 0.019542f
C16 A1 A2 0.233027f
C17 VPB Y 0.007694f
C18 VPB B1_N 0.047123f
C19 VGND VNB 0.537587f
C20 Y VNB 0.017874f
C21 VPWR VNB 0.471698f
C22 A2 VNB 0.188504f
C23 A1 VNB 0.262649f
C24 B1_N VNB 0.157241f
C25 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21bai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21bai_1 VNB VPB VPWR VGND B1_N Y A2 A1
X0 VGND.t0 A2.t0 a_308_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1221 ps=1.07 w=0.74 l=0.15
X1 a_395_368.t0 A2.t1 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t2 A1.t0 a_395_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.1848 ps=1.45 w=1.12 l=0.15
X3 Y.t2 a_27_74.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3626 ps=1.895 w=1.12 l=0.15
X4 a_308_74.t0 a_27_74.t3 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.2072 ps=2.04 w=0.74 l=0.15
X5 VPWR.t0 B1_N.t0 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3626 pd=1.895 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 VGND.t1 B1_N.t1 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.15125 pd=1.65 as=0.154 ps=1.66 w=0.55 l=0.15
X7 a_308_74.t2 A1.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1073 ps=1.03 w=0.74 l=0.15
R0 A2.n0 A2.t1 264.298
R1 A2.n0 A2.t0 204.048
R2 A2 A2.n0 158.207
R3 A2.n1 A2 17.8092
R4 A2.n1 A2 3.29747
R5 A2 A2.n1 2.78311
R6 a_308_74.n0 a_308_74.t2 308.784
R7 a_308_74.t0 a_308_74.n0 30.8113
R8 a_308_74.n0 a_308_74.t1 22.7032
R9 VGND.n1 VGND.t1 246.365
R10 VGND.n1 VGND.n0 210.522
R11 VGND.n0 VGND.t2 23.514
R12 VGND.n0 VGND.t0 23.514
R13 VGND VGND.n1 0.242184
R14 VNB.t2 VNB.t0 2251.97
R15 VNB VNB.t2 1131.76
R16 VNB.t0 VNB.t1 1108.66
R17 VNB.t1 VNB.t3 1016.27
R18 Y.n1 Y 589.385
R19 Y.n1 Y.n0 585
R20 Y.n2 Y.n1 585
R21 Y Y.t0 209.661
R22 Y.n1 Y.t1 26.3844
R23 Y.n1 Y.t2 26.3844
R24 Y Y.n2 11.7484
R25 Y Y.n0 10.1704
R26 Y Y.n0 2.80598
R27 Y.n2 Y 1.2279
R28 a_395_368.t0 a_395_368.t1 58.0451
R29 VPB.t0 VPB.t2 472.447
R30 VPB VPB.t0 268.146
R31 VPB.t1 VPB.t3 245.161
R32 VPB.t2 VPB.t1 229.839
R33 A1.n0 A1.t0 256.596
R34 A1.n0 A1.t1 196.345
R35 A1 A1.n0 156.462
R36 VPWR.n2 VPWR.n0 585
R37 VPWR.n1 VPWR.n0 585
R38 VPWR.n4 VPWR.n3 273.839
R39 VPWR.n5 VPWR.t2 265.103
R40 VPWR.n1 VPWR.t1 50.9336
R41 VPWR.n2 VPWR.t0 46.9053
R42 VPWR.n3 VPWR.n2 37.3262
R43 VPWR.n3 VPWR.n1 37.3262
R44 VPWR.n5 VPWR.n4 13.4759
R45 VPWR.n4 VPWR.n0 6.87811
R46 VPWR VPWR.n5 0.283677
R47 a_27_74.t0 a_27_74.n1 455.497
R48 a_27_74.n0 a_27_74.t2 308.481
R49 a_27_74.n1 a_27_74.t1 286.015
R50 a_27_74.n1 a_27_74.n0 248.4
R51 a_27_74.n0 a_27_74.t3 200.03
R52 B1_N.n0 B1_N.t1 282.774
R53 B1_N.n0 B1_N.t0 254.924
R54 B1_N B1_N.n0 161.504
C0 A2 A1 0.116967f
C1 VPWR Y 0.117379f
C2 Y VPB 0.007754f
C3 VPWR B1_N 0.018982f
C4 VPB B1_N 0.073658f
C5 VGND A2 0.017769f
C6 A1 Y 8.18e-19
C7 VPWR VPB 0.092744f
C8 VGND Y 0.087869f
C9 VGND B1_N 0.018527f
C10 A2 Y 0.128233f
C11 A1 VPWR 0.046388f
C12 A2 B1_N 2.04e-19
C13 A1 VPB 0.043355f
C14 VGND VPWR 0.04895f
C15 VGND VPB 0.006895f
C16 A2 VPWR 0.101136f
C17 A2 VPB 0.035511f
C18 Y B1_N 0.003147f
C19 VGND A1 0.01712f
C20 VGND VNB 0.39416f
C21 Y VNB 0.021294f
C22 VPWR VNB 0.343284f
C23 A1 VNB 0.167514f
C24 A2 VNB 0.108983f
C25 B1_N VNB 0.186246f
C26 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21ba_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21ba_4 VNB VPB VPWR VGND A1 A2 B1_N X
X0 VPWR.t4 a_193_48.t6 X.t5 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.371 pd=1.915 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t5 B1_N.t0 a_27_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 X.t2 a_193_48.t7 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_193_48.t3 a_27_368.t2 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.371 ps=1.915 w=0.84 l=0.15
X4 VPWR.t2 a_193_48.t8 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_193_48.t1 A2.t0 a_892_392.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X6 VPWR.t6 A1.t0 a_892_392.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X7 X.t0 a_193_48.t9 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X8 a_892_392.t3 A1.t1 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2039 ps=1.435 w=1 l=0.15
X9 a_892_392.t0 A2.t1 a_193_48.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X10 a_618_94.t1 a_27_368.t3 a_193_48.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.123625 pd=1.145 as=0.0896 ps=0.92 w=0.64 l=0.15
X11 VGND.t3 a_193_48.t10 X.t7 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_618_94.t4 A2.t2 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
X13 VGND.t2 a_193_48.t11 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1073 ps=1.03 w=0.74 l=0.15
X14 VGND.t7 B1_N.t1 a_27_368.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.13505 pd=1.105 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 a_193_48.t5 a_27_368.t4 a_618_94.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X16 X.t4 a_193_48.t12 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t4 A1.t2 a_618_94.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.123625 ps=1.145 w=0.64 l=0.15
X18 VGND.t5 A2.t3 a_618_94.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X19 VPWR.t0 a_27_368.t5 a_193_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2039 pd=1.435 as=0.126 ps=1.14 w=0.84 l=0.15
X20 X.t3 a_193_48.t13 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.13505 ps=1.105 w=0.74 l=0.15
R0 a_193_48.n14 a_193_48.n13 345.587
R1 a_193_48.n13 a_193_48.n12 306.5
R2 a_193_48.n11 a_193_48.n1 306.349
R3 a_193_48.n3 a_193_48.t9 261.62
R4 a_193_48.n0 a_193_48.t6 252.369
R5 a_193_48.n8 a_193_48.t7 242.875
R6 a_193_48.n5 a_193_48.t8 242.875
R7 a_193_48.n3 a_193_48.t13 179.514
R8 a_193_48.n4 a_193_48.t11 176.733
R9 a_193_48.n7 a_193_48.t12 176.733
R10 a_193_48.n0 a_193_48.t10 176.733
R11 a_193_48.n6 a_193_48.n2 165.189
R12 a_193_48.n9 a_193_48.n2 152
R13 a_193_48.n10 a_193_48.n0 152
R14 a_193_48.n13 a_193_48.n11 97.7916
R15 a_193_48.n4 a_193_48.n3 75.8397
R16 a_193_48.n0 a_193_48.n9 51.1217
R17 a_193_48.n7 a_193_48.n6 37.9763
R18 a_193_48.n12 a_193_48.t0 35.1791
R19 a_193_48.n12 a_193_48.t3 35.1791
R20 a_193_48.n14 a_193_48.t2 29.5505
R21 a_193_48.t1 a_193_48.n14 29.5505
R22 a_193_48.n1 a_193_48.t4 26.2505
R23 a_193_48.n1 a_193_48.t5 26.2505
R24 a_193_48.n11 a_193_48.n10 21.9157
R25 a_193_48.n6 a_193_48.n5 21.1793
R26 a_193_48.n10 a_193_48.n2 13.1884
R27 a_193_48.n8 a_193_48.n7 6.57323
R28 a_193_48.n9 a_193_48.n8 5.11262
R29 a_193_48.n5 a_193_48.n4 3.65202
R30 X.n2 X.n0 613.801
R31 X.n2 X.n1 585
R32 X.n5 X.n3 148.589
R33 X.n5 X.n4 104.451
R34 X X.n5 39.626
R35 X.n1 X.t1 26.3844
R36 X.n1 X.t0 26.3844
R37 X.n0 X.t5 26.3844
R38 X.n0 X.t2 26.3844
R39 X.n4 X.t6 24.3248
R40 X.n4 X.t3 22.7032
R41 X.n3 X.t7 22.7032
R42 X.n3 X.t4 22.7032
R43 X.n6 X 13.357
R44 X X.n6 2.7205
R45 X.n6 X.n2 2.5605
R46 VPWR.n7 VPWR.n6 611.958
R47 VPWR.n19 VPWR.n3 604.976
R48 VPWR.n21 VPWR.n1 602.347
R49 VPWR.n12 VPWR.n4 585
R50 VPWR.n14 VPWR.n13 585
R51 VPWR.n8 VPWR.t6 268.305
R52 VPWR.n13 VPWR.n12 96.1553
R53 VPWR.n13 VPWR.t8 55.1136
R54 VPWR.n6 VPWR.t0 55.1136
R55 VPWR.n6 VPWR.t7 43.3808
R56 VPWR.n1 VPWR.t5 39.5764
R57 VPWR.n11 VPWR.n10 31.33
R58 VPWR.n12 VPWR.t4 31.284
R59 VPWR.n1 VPWR.t1 30.7817
R60 VPWR.n20 VPWR.n19 27.4829
R61 VPWR.n3 VPWR.t3 26.3844
R62 VPWR.n3 VPWR.t2 26.3844
R63 VPWR.n18 VPWR.n4 26.0484
R64 VPWR.n10 VPWR.n7 25.977
R65 VPWR.n19 VPWR.n18 19.9534
R66 VPWR.n21 VPWR.n20 15.4358
R67 VPWR.n10 VPWR.n9 9.3005
R68 VPWR.n11 VPWR.n5 9.3005
R69 VPWR.n16 VPWR.n15 9.3005
R70 VPWR.n18 VPWR.n17 9.3005
R71 VPWR.n19 VPWR.n2 9.3005
R72 VPWR.n20 VPWR.n0 9.3005
R73 VPWR.n15 VPWR.n14 7.47495
R74 VPWR.n22 VPWR.n21 7.43488
R75 VPWR.n8 VPWR.n7 7.00784
R76 VPWR.n14 VPWR.n11 1.49539
R77 VPWR.n15 VPWR.n4 0.187361
R78 VPWR.n9 VPWR.n8 0.173461
R79 VPWR VPWR.n22 0.160103
R80 VPWR.n22 VPWR.n0 0.1477
R81 VPWR.n9 VPWR.n5 0.122949
R82 VPWR.n16 VPWR.n5 0.122949
R83 VPWR.n17 VPWR.n16 0.122949
R84 VPWR.n17 VPWR.n2 0.122949
R85 VPWR.n2 VPWR.n0 0.122949
R86 VPB.t4 VPB.t10 482.661
R87 VPB.t0 VPB.t7 298.791
R88 VPB.t5 VPB.t1 280.914
R89 VPB VPB.t5 257.93
R90 VPB.t9 VPB.t6 229.839
R91 VPB.t8 VPB.t9 229.839
R92 VPB.t7 VPB.t8 229.839
R93 VPB.t10 VPB.t0 229.839
R94 VPB.t3 VPB.t4 229.839
R95 VPB.t2 VPB.t3 229.839
R96 VPB.t1 VPB.t2 229.839
R97 B1_N.n0 B1_N.t0 285.01
R98 B1_N.n0 B1_N.t1 177.631
R99 B1_N B1_N.n0 157.464
R100 a_27_368.n3 a_27_368.n2 410.945
R101 a_27_368.n0 a_27_368.t3 286.368
R102 a_27_368.n1 a_27_368.t4 269.921
R103 a_27_368.t0 a_27_368.n3 218.899
R104 a_27_368.n3 a_27_368.t1 218.751
R105 a_27_368.n0 a_27_368.t5 181.821
R106 a_27_368.n2 a_27_368.t2 181.821
R107 a_27_368.n1 a_27_368.n0 51.1217
R108 a_27_368.n2 a_27_368.n1 14.6066
R109 A2.n1 A2.t0 219.457
R110 A2.n0 A2.t1 212.883
R111 A2.n0 A2.t3 166.136
R112 A2.n1 A2.t2 162.274
R113 A2.n3 A2.n2 152
R114 A2.n2 A2.n0 40.1672
R115 A2.n2 A2.n1 18.9884
R116 A2.n3 A2 16.4853
R117 A2 A2.n3 2.13383
R118 a_892_392.n1 a_892_392.n0 850.86
R119 a_892_392.n0 a_892_392.t2 29.5505
R120 a_892_392.n0 a_892_392.t0 29.5505
R121 a_892_392.t1 a_892_392.n1 29.5505
R122 a_892_392.n1 a_892_392.t3 29.5505
R123 A1.t2 A1.n0 880.453
R124 A1.n0 A1.t0 457.632
R125 A1.n1 A1.t1 236.983
R126 A1.n1 A1.t2 186.374
R127 A1 A1.n1 157.237
R128 VGND.n7 VGND.t5 305.219
R129 VGND.n6 VGND.n5 224.424
R130 VGND.n16 VGND.n2 213.929
R131 VGND.n12 VGND.t3 170.673
R132 VGND.n19 VGND.n18 115.692
R133 VGND.n5 VGND.t4 39.3755
R134 VGND.n10 VGND.n4 36.1417
R135 VGND.n11 VGND.n10 36.1417
R136 VGND.n12 VGND.n11 36.1417
R137 VGND.n18 VGND.t7 34.0546
R138 VGND.n6 VGND.n4 31.624
R139 VGND.n16 VGND.n1 28.6123
R140 VGND.n5 VGND.t6 26.2505
R141 VGND.n18 VGND.t0 25.1356
R142 VGND.n17 VGND.n16 24.8476
R143 VGND.n2 VGND.t1 22.7032
R144 VGND.n2 VGND.t2 22.7032
R145 VGND.n12 VGND.n1 17.3181
R146 VGND.n19 VGND.n17 16.9417
R147 VGND.n17 VGND.n0 9.3005
R148 VGND.n16 VGND.n15 9.3005
R149 VGND.n14 VGND.n1 9.3005
R150 VGND.n8 VGND.n4 9.3005
R151 VGND.n10 VGND.n9 9.3005
R152 VGND.n11 VGND.n3 9.3005
R153 VGND.n13 VGND.n12 9.3005
R154 VGND.n20 VGND.n19 7.52053
R155 VGND.n7 VGND.n6 6.60377
R156 VGND.n8 VGND.n7 0.571275
R157 VGND VGND.n20 0.161231
R158 VGND.n20 VGND.n0 0.146587
R159 VGND.n9 VGND.n8 0.122949
R160 VGND.n9 VGND.n3 0.122949
R161 VGND.n13 VGND.n3 0.122949
R162 VGND.n14 VGND.n13 0.122949
R163 VGND.n15 VGND.n14 0.122949
R164 VGND.n15 VGND.n0 0.122949
R165 a_618_94.n1 a_618_94.t0 279.132
R166 a_618_94.n2 a_618_94.n1 185
R167 a_618_94.n1 a_618_94.n0 149.118
R168 a_618_94.t1 a_618_94.n2 43.2736
R169 a_618_94.n0 a_618_94.t3 26.2505
R170 a_618_94.n0 a_618_94.t4 26.2505
R171 a_618_94.n2 a_618_94.t2 25.954
R172 VNB.t5 VNB.t0 2563.78
R173 VNB VNB.t9 1212.6
R174 VNB.t9 VNB.t2 1189.5
R175 VNB.t6 VNB.t8 1154.86
R176 VNB.t1 VNB.t6 1154.86
R177 VNB.t2 VNB.t4 1016.27
R178 VNB.t8 VNB.t7 993.177
R179 VNB.t0 VNB.t1 993.177
R180 VNB.t3 VNB.t5 993.177
R181 VNB.t4 VNB.t3 993.177
C0 VPWR VGND 0.10433f
C1 A1 VPB 0.079975f
C2 A2 VPWR 0.037356f
C3 VPWR X 0.041229f
C4 A2 VGND 0.022946f
C5 X VGND 0.282064f
C6 B1_N VPB 0.035159f
C7 A1 VPWR 0.032124f
C8 A1 VGND 0.085219f
C9 B1_N VPWR 0.016706f
C10 A1 A2 0.18268f
C11 VPWR VPB 0.16928f
C12 A1 X 9e-20
C13 B1_N VGND 0.039974f
C14 VGND VPB 0.010523f
C15 A2 VPB 0.076707f
C16 B1_N X 0.024534f
C17 X VPB 0.010304f
C18 VGND VNB 0.762916f
C19 X VNB 0.017431f
C20 VPWR VNB 0.619415f
C21 A2 VNB 0.173878f
C22 A1 VNB 0.406799f
C23 B1_N VNB 0.139518f
C24 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o22a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o22a_1 VNB VPB VPWR VGND X B1 A2 B2 A1
X0 VPWR.t2 a_83_260.t4 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.6459 pd=2.38 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_299_139.t3 B2.t0 a_83_260.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1024 ps=0.96 w=0.64 l=0.15
X2 a_299_139.t2 A1.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.18205 pd=1.85 as=0.144725 ps=1.125 w=0.64 l=0.15
X3 VGND.t1 a_83_260.t5 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 VGND.t0 A2.t0 a_299_139.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.144725 pd=1.125 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 a_572_392.t0 A2.t1 a_83_260.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.15 ps=1.3 w=1 l=0.15
X6 a_83_260.t0 B1.t0 a_299_139.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1705 ps=1.85 w=0.64 l=0.15
X7 a_83_260.t3 B2.t1 a_398_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t1 A1.t1 a_572_392.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.195 ps=1.39 w=1 l=0.15
X9 a_398_392.t1 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.6459 ps=2.38 w=1 l=0.15
R0 a_83_260.n3 a_83_260.n2 277.051
R1 a_83_260.n0 a_83_260.t4 240.197
R2 a_83_260.n2 a_83_260.n0 185.857
R3 a_83_260.n2 a_83_260.n1 185
R4 a_83_260.n0 a_83_260.t5 181.407
R5 a_83_260.n1 a_83_260.t1 30.0005
R6 a_83_260.n1 a_83_260.t0 30.0005
R7 a_83_260.t2 a_83_260.n3 29.5505
R8 a_83_260.n3 a_83_260.t3 29.5505
R9 X.n1 X 589.444
R10 X.n1 X.n0 585
R11 X.n2 X.n1 585
R12 X X.t0 208.948
R13 X.n1 X.t1 26.3844
R14 X X.n2 11.9116
R15 X X.n0 10.3116
R16 X X.n0 2.84494
R17 X.n2 X 1.24494
R18 VPWR.n4 VPWR.t1 258.868
R19 VPWR.n10 VPWR.n9 195
R20 VPWR.n3 VPWR.n2 195
R21 VPWR.n8 VPWR.n7 195
R22 VPWR.n9 VPWR.n8 98.5005
R23 VPWR.n8 VPWR.n2 88.6505
R24 VPWR.n4 VPWR.n3 32.3988
R25 VPWR.n2 VPWR.t0 30.5355
R26 VPWR.n9 VPWR.t2 28.6759
R27 VPWR.n6 VPWR.n5 9.3005
R28 VPWR.n1 VPWR.n0 9.3005
R29 VPWR.n11 VPWR.n10 7.60576
R30 VPWR.n10 VPWR.n1 4.16274
R31 VPWR.n7 VPWR.n6 3.98372
R32 VPWR.n7 VPWR.n1 0.313787
R33 VPWR.n5 VPWR.n4 0.218694
R34 VPWR VPWR.n11 0.160585
R35 VPWR.n11 VPWR.n0 0.147224
R36 VPWR.n5 VPWR.n0 0.122949
R37 VPWR.n6 VPWR.n3 0.0452552
R38 VPB VPB.t0 140.7
R39 VPB.t0 VPB.t1 13.5076
R40 B2.t0 B2.t1 438.889
R41 B2.n0 B2.t0 357.329
R42 B2 B2.n0 6.69141
R43 B2.n0 B2 3.10353
R44 a_299_139.n2 a_299_139.n1 249
R45 a_299_139.n1 a_299_139.t2 200.894
R46 a_299_139.n1 a_299_139.n0 185
R47 a_299_139.n2 a_299_139.t0 70.2297
R48 a_299_139.n0 a_299_139.t1 26.2505
R49 a_299_139.n0 a_299_139.t3 26.2505
R50 VNB.n0 VNB 3692.86
R51 VNB VNB.n1 2658.33
R52 VNB.n1 VNB.t0 1592.71
R53 VNB.n1 VNB.t4 1535.96
R54 VNB.n0 VNB.t2 1388.1
R55 VNB.t4 VNB 1143.31
R56 VNB.t0 VNB.t3 1077.08
R57 VNB.t1 VNB.n0 996.875
R58 VNB.t3 VNB.t1 985.418
R59 A1.n0 A1.t1 231.629
R60 A1.n0 A1.t0 184.768
R61 A1 A1.n0 156.462
R62 VGND.n1 VGND.n0 221.28
R63 VGND.n1 VGND.t1 144.397
R64 VGND.n0 VGND.t0 41.336
R65 VGND.n0 VGND.t2 32.4623
R66 VGND VGND.n1 0.191665
R67 A2.n0 A2.t1 231.629
R68 A2.n0 A2.t0 170.308
R69 A2 A2.n0 162.667
R70 a_572_392.t0 a_572_392.t1 76.8305
R71 B1.n0 B1.t1 216.292
R72 B1.n0 B1.t0 146.208
R73 B1 B1.n0 92.5936
R74 a_398_392.t0 a_398_392.t1 53.1905
C0 B1 VGND 0.006699f
C1 B2 VPWR 0.014574f
C2 X VGND 0.083988f
C3 B1 B2 0.058845f
C4 VPB A2 0.04116f
C5 VPB VGND 0.00852f
C6 B1 VPWR 0.075457f
C7 B2 X 1.53e-19
C8 A2 A1 0.064333f
C9 X VPWR 0.124773f
C10 A1 VGND 0.011719f
C11 VPB B2 0.028808f
C12 B2 A1 9e-19
C13 VPB VPWR 0.117869f
C14 B1 X 0.004097f
C15 A1 VPWR 0.055229f
C16 A2 VGND 0.0117f
C17 VPB B1 0.070685f
C18 VPB X 0.017547f
C19 B2 A2 0.05686f
C20 B2 VGND 0.21297f
C21 A2 VPWR 0.019911f
C22 VPWR VGND 0.064851f
C23 VPB A1 0.047668f
C24 VGND VNB 0.520547f
C25 VPWR VNB 0.418676f
C26 X VNB 0.116529f
C27 A1 VNB 0.135823f
C28 A2 VNB 0.091983f
C29 B2 VNB 0.162706f
C30 B1 VNB 0.127114f
C31 VPB VNB 0.93825f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o31a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o31a_1 VNB VPB VPWR VGND B1 A2 A1 A3 X
X0 VGND.t3 a_84_48.t3 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VGND.t1 A2.t0 a_230_94.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.21 as=0.1136 ps=0.995 w=0.64 l=0.15
X2 VPWR.t2 a_84_48.t4 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2907 pd=1.66 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_84_48.t0 B1.t0 a_230_94.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.1104 ps=0.985 w=0.64 l=0.15
X4 a_340_368.t0 A2.t1 a_256_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X5 a_84_48.t2 A3.t0 a_340_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1874 pd=1.39 as=0.18 ps=1.36 w=1 l=0.15
X6 a_256_368.t1 A1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2907 ps=1.66 w=1 l=0.15
X7 a_230_94.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1136 pd=0.995 as=0.15535 ps=1.17 w=0.64 l=0.15
X8 VPWR.t0 B1.t1 a_84_48.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.399 pd=2.63 as=0.1874 ps=1.39 w=0.84 l=0.15
X9 a_230_94.t3 A3.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1104 pd=0.985 as=0.1824 ps=1.21 w=0.64 l=0.15
R0 a_84_48.n3 a_84_48.n2 292.108
R1 a_84_48.n1 a_84_48.n0 7.73055
R2 a_84_48.n2 a_84_48.t4 258.582
R3 a_84_48.n3 a_84_48.t0 251.575
R4 a_84_48.n2 a_84_48.t3 210.114
R5 a_84_48.n0 a_84_48.t1 56.2862
R6 a_84_48.n4 a_84_48.n1 46.2119
R7 a_84_48.n0 a_84_48.t2 29.5767
R8 a_84_48.n1 a_84_48.n3 196.948
R9 X.n1 X 589.324
R10 X.n1 X.n0 585
R11 X.n2 X.n1 585
R12 X X.t0 206.076
R13 X.n1 X.t1 26.3844
R14 X X.n2 11.5897
R15 X X.n0 10.0329
R16 X X.n0 2.76807
R17 X.n2 X 1.21131
R18 VGND.n2 VGND.n1 212.499
R19 VGND.n2 VGND.n0 122.294
R20 VGND.n1 VGND.t1 54.3755
R21 VGND.n1 VGND.t2 52.5005
R22 VGND.n0 VGND.t0 41.2505
R23 VGND.n0 VGND.t3 30.6984
R24 VGND VGND.n2 0.33901
R25 VNB.t2 VNB.t3 1662.99
R26 VNB.t4 VNB.t0 1339.63
R27 VNB.t0 VNB.t2 1166.4
R28 VNB.t3 VNB.t1 1143.31
R29 VNB VNB.t4 1143.31
R30 A2.n0 A2.t1 245.018
R31 A2.n0 A2.t0 187.981
R32 A2 A2.n0 156.462
R33 a_230_94.n1 a_230_94.n0 269.567
R34 a_230_94.n1 a_230_94.t1 40.313
R35 a_230_94.n0 a_230_94.t3 38.438
R36 a_230_94.n0 a_230_94.t2 26.2505
R37 a_230_94.t0 a_230_94.n1 26.2505
R38 VPWR.n1 VPWR.t0 709.237
R39 VPWR.n1 VPWR.n0 307.974
R40 VPWR.n0 VPWR.t1 53.5134
R41 VPWR.n0 VPWR.t2 48.3439
R42 VPWR VPWR.n1 0.223188
R43 VPB.t4 VPB.t3 352.42
R44 VPB.t2 VPB.t1 275.807
R45 VPB VPB.t4 263.038
R46 VPB.t0 VPB.t2 260.485
R47 VPB.t3 VPB.t0 214.517
R48 B1.n0 B1.t1 205.922
R49 B1.n0 B1.t0 204.048
R50 B1 B1.n0 157.805
R51 a_256_368.t0 a_256_368.t1 53.1905
R52 a_340_368.t0 a_340_368.t1 70.9205
R53 A3.n0 A3.t0 231.629
R54 A3.n0 A3.t1 204.048
R55 A3 A3.n0 156.019
R56 A1.n0 A1.t0 231.629
R57 A1.n0 A1.t1 204.048
R58 A1 A1.n0 154.377
C0 A1 VPB 0.03636f
C1 B1 VGND 0.012931f
C2 X A1 0.001814f
C3 VPB VGND 0.007876f
C4 VPWR B1 0.013273f
C5 X VGND 0.105028f
C6 VPWR VPB 0.11349f
C7 A3 VGND 0.013744f
C8 X VPWR 0.101561f
C9 VPB B1 0.042634f
C10 A1 A2 0.093016f
C11 X B1 1.38e-19
C12 VPWR A3 0.007992f
C13 A2 VGND 0.013457f
C14 X VPB 0.014306f
C15 A3 B1 0.085324f
C16 VPB A3 0.036808f
C17 VPWR A2 0.010158f
C18 X A3 2.31e-19
C19 A1 VGND 0.020187f
C20 A2 B1 1.1e-19
C21 A2 VPB 0.032129f
C22 X A2 8.58e-19
C23 VPWR A1 0.014794f
C24 A2 A3 0.080056f
C25 VPWR VGND 0.056475f
C26 VGND VNB 0.447943f
C27 B1 VNB 0.133864f
C28 A3 VNB 0.106732f
C29 A2 VNB 0.107651f
C30 A1 VNB 0.108627f
C31 VPWR VNB 0.375924f
C32 X VNB 0.115257f
C33 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o22ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o22ai_4 VNB VPB VPWR VGND B1 B2 Y A2 A1
X0 VPWR.t6 A1.t0 a_117_368.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_117_368.t1 A2.t0 Y.t8 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_27_74.t3 B1.t0 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1258 ps=1.08 w=0.74 l=0.15
X3 Y.t13 B2.t0 a_877_368.t5 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t3 A2.t1 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1406 pd=1.12 as=0.1184 ps=1.06 w=0.74 l=0.15
X5 Y.t7 A2.t2 a_117_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_27_74.t6 A2.t3 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 a_117_368.t2 A2.t4 Y.t6 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8 a_877_368.t4 B2.t1 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.1736 ps=1.43 w=1.12 l=0.15
X9 Y.t14 B2.t2 a_877_368.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X10 a_117_368.t5 A1.t1 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X11 a_27_74.t5 A2.t5 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X12 a_27_74.t12 B2.t3 Y.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 Y.t2 B1.t1 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1073 ps=1.03 w=0.74 l=0.15
X14 VGND.t7 A1.t2 a_27_74.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 VGND.t0 A2.t6 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VPWR.t0 B1.t2 a_877_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 Y.t5 A2.t7 a_117_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_877_368.t1 B1.t3 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X19 a_877_368.t0 B1.t4 VPWR.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X20 VGND.t6 A1.t3 a_27_74.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 Y.t10 B2.t4 a_27_74.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_117_368.t4 A1.t4 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X23 Y.t3 B1.t5 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1073 ps=1.03 w=0.74 l=0.15
X24 a_27_74.t9 A1.t5 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1406 ps=1.12 w=0.74 l=0.15
X25 a_27_74.t0 B1.t6 Y.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2991 pd=2.41 as=0.1295 ps=1.09 w=0.74 l=0.15
X26 a_27_74.t8 A1.t6 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X27 a_27_74.t14 B2.t5 Y.t11 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VPWR.t3 A1.t7 a_117_368.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X29 Y.t12 B2.t6 a_27_74.t15 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
R0 A1.n0 A1.t0 250.909
R1 A1.n2 A1.t4 239.953
R2 A1.n5 A1.t7 234.841
R3 A1.n3 A1.t1 234.841
R4 A1.n0 A1.t5 220.113
R5 A1 A1.n0 204.26
R6 A1.n3 A1.t2 188.565
R7 A1.n6 A1.t6 186.374
R8 A1.n2 A1.t3 186.374
R9 A1.n4 A1.n1 165.189
R10 A1.n9 A1.n8 152
R11 A1.n7 A1.n1 152
R12 A1 A1.n9 89.0789
R13 A1.n8 A1.n7 49.6611
R14 A1.n5 A1.n4 37.246
R15 A1.n4 A1.n3 28.4823
R16 A1.n9 A1.n1 13.1884
R17 A1.n7 A1.n6 7.30353
R18 A1.n8 A1.n2 5.84292
R19 A1.n6 A1.n5 5.11262
R20 a_117_368.n4 a_117_368.n0 621
R21 a_117_368.n5 a_117_368.n4 585
R22 a_117_368.n3 a_117_368.n2 286.889
R23 a_117_368.n3 a_117_368.n1 263.615
R24 a_117_368.n4 a_117_368.n3 42.8178
R25 a_117_368.n0 a_117_368.t6 26.3844
R26 a_117_368.n0 a_117_368.t1 26.3844
R27 a_117_368.n2 a_117_368.t3 26.3844
R28 a_117_368.n2 a_117_368.t4 26.3844
R29 a_117_368.n1 a_117_368.t7 26.3844
R30 a_117_368.n1 a_117_368.t5 26.3844
R31 a_117_368.t0 a_117_368.n5 26.3844
R32 a_117_368.n5 a_117_368.t2 26.3844
R33 VPWR.n8 VPWR.n7 620.29
R34 VPWR.n6 VPWR.n5 606.333
R35 VPWR.n17 VPWR.n2 315.349
R36 VPWR.n19 VPWR.t5 259.171
R37 VPWR.n11 VPWR.n10 36.1417
R38 VPWR.n12 VPWR.n11 36.1417
R39 VPWR.n12 VPWR.n3 36.1417
R40 VPWR.n16 VPWR.n3 36.1417
R41 VPWR.n2 VPWR.t4 35.1791
R42 VPWR.n5 VPWR.t1 35.1791
R43 VPWR.n5 VPWR.t6 35.1791
R44 VPWR.n2 VPWR.t3 26.3844
R45 VPWR.n7 VPWR.t2 26.3844
R46 VPWR.n7 VPWR.t0 26.3844
R47 VPWR.n19 VPWR.n18 26.3534
R48 VPWR.n17 VPWR.n16 24.8476
R49 VPWR.n18 VPWR.n17 22.5887
R50 VPWR.n10 VPWR.n6 20.3299
R51 VPWR.n10 VPWR.n9 9.3005
R52 VPWR.n11 VPWR.n4 9.3005
R53 VPWR.n13 VPWR.n12 9.3005
R54 VPWR.n14 VPWR.n3 9.3005
R55 VPWR.n16 VPWR.n15 9.3005
R56 VPWR.n17 VPWR.n1 9.3005
R57 VPWR.n18 VPWR.n0 9.3005
R58 VPWR.n20 VPWR.n19 9.3005
R59 VPWR.n8 VPWR.n6 6.95043
R60 VPWR.n9 VPWR.n8 0.498883
R61 VPWR.n9 VPWR.n4 0.122949
R62 VPWR.n13 VPWR.n4 0.122949
R63 VPWR.n14 VPWR.n13 0.122949
R64 VPWR.n15 VPWR.n14 0.122949
R65 VPWR.n15 VPWR.n1 0.122949
R66 VPWR.n1 VPWR.n0 0.122949
R67 VPWR.n20 VPWR.n0 0.122949
R68 VPWR VPWR.n20 0.0617245
R69 VPB.t13 VPB.t12 459.678
R70 VPB.t11 VPB.t6 280.914
R71 VPB VPB.t10 260.485
R72 VPB.t7 VPB.t13 255.376
R73 VPB.t4 VPB.t3 255.376
R74 VPB.t8 VPB.t9 255.376
R75 VPB.t12 VPB.t1 234.946
R76 VPB.t5 VPB.t7 229.839
R77 VPB.t6 VPB.t5 229.839
R78 VPB.t2 VPB.t11 229.839
R79 VPB.t0 VPB.t2 229.839
R80 VPB.t3 VPB.t0 229.839
R81 VPB.t9 VPB.t4 229.839
R82 VPB.t10 VPB.t8 229.839
R83 A2.n2 A2.t0 261.62
R84 A2.n3 A2.t2 261.62
R85 A2.n7 A2.t4 261.62
R86 A2.n10 A2.t7 261.62
R87 A2.n2 A2.t1 156.431
R88 A2.n10 A2.t5 154.24
R89 A2.n9 A2.t6 154.24
R90 A2.n1 A2.t3 154.24
R91 A2 A2.n4 153.212
R92 A2 A2.n11 152.865
R93 A2.n6 A2.n5 152
R94 A2.n8 A2.n0 152
R95 A2.n7 A2.n6 46.7399
R96 A2.n11 A2.n9 44.549
R97 A2.n4 A2.n2 35.055
R98 A2.n4 A2.n3 30.6732
R99 A2.n6 A2.n1 18.2581
R100 A2.n11 A2.n10 18.2581
R101 A2 A2.n0 10.8978
R102 A2.n5 A2 10.5519
R103 A2.n5 A2 6.05455
R104 A2 A2.n0 5.70861
R105 A2.n9 A2.n8 5.11262
R106 A2.n8 A2.n7 2.92171
R107 A2.n3 A2.n1 0.730803
R108 Y.n2 Y.n0 645.254
R109 Y.n2 Y.n1 585
R110 Y.n3 Y.t14 386.277
R111 Y.n5 Y.n4 299.95
R112 Y.n3 Y.n2 228.274
R113 Y.n7 Y.n5 192.099
R114 Y.n7 Y.n6 185
R115 Y.n9 Y.n8 185
R116 Y.n11 Y.n10 185
R117 Y.n13 Y.n12 185
R118 Y.n11 Y.n9 64.099
R119 Y.n9 Y.n7 63.4445
R120 Y.n5 Y.n3 43.2763
R121 Y.n0 Y.t5 35.1791
R122 Y.n8 Y.t10 34.0546
R123 Y.n6 Y.t12 34.0546
R124 Y.n12 Y.t2 32.4329
R125 Y Y.n11 28.1962
R126 Y.n4 Y.t0 28.1434
R127 Y.n1 Y.t8 26.3844
R128 Y.n1 Y.t7 26.3844
R129 Y.n0 Y.t6 26.3844
R130 Y.n4 Y.t13 26.3844
R131 Y.n12 Y.t1 22.7032
R132 Y.n10 Y.t11 22.7032
R133 Y.n10 Y.t3 22.7032
R134 Y.n8 Y.t9 22.7032
R135 Y.n6 Y.t4 22.7032
R136 Y.n13 Y 12.9689
R137 Y Y.n13 3.2005
R138 B1.n2 B1.n1 300.05
R139 B1.n1 B1.n0 285.719
R140 B1.n4 B1.t4 240.197
R141 B1.n7 B1.t2 240.197
R142 B1.n5 B1.t3 240.197
R143 B1.n5 B1.t1 182.138
R144 B1.n4 B1.t5 182.138
R145 B1.n8 B1.t0 179.947
R146 B1.n1 B1.t6 178.34
R147 B1.n6 B1.n3 165.189
R148 B1.n11 B1.n10 152
R149 B1.n9 B1.n3 152
R150 B1.n10 B1.n9 49.6611
R151 B1.n7 B1.n6 44.549
R152 B1.n6 B1.n5 21.1793
R153 B1.n11 B1.n3 13.1884
R154 B1 B1.n11 11.6369
R155 B1.n10 B1.n4 10.955
R156 B1.n2 B1 5.18145
R157 B1.n8 B1.n7 3.65202
R158 B1 B1.n2 3.29747
R159 B1.n9 B1.n8 1.46111
R160 a_27_74.n1 a_27_74.t0 356.046
R161 a_27_74.n5 a_27_74.t11 205.264
R162 a_27_74.n1 a_27_74.n0 185
R163 a_27_74.n3 a_27_74.n2 185
R164 a_27_74.n13 a_27_74.n12 185
R165 a_27_74.n7 a_27_74.n6 97.4677
R166 a_27_74.n9 a_27_74.n8 97.4677
R167 a_27_74.n5 a_27_74.n4 96.9594
R168 a_27_74.n11 a_27_74.n10 89.0748
R169 a_27_74.n3 a_27_74.n1 63.4445
R170 a_27_74.n11 a_27_74.n9 58.105
R171 a_27_74.n7 a_27_74.n5 52.2744
R172 a_27_74.n9 a_27_74.n7 51.2005
R173 a_27_74.n12 a_27_74.n11 41.7992
R174 a_27_74.n12 a_27_74.n3 34.0682
R175 a_27_74.n0 a_27_74.t12 34.0546
R176 a_27_74.n8 a_27_74.t7 29.1897
R177 a_27_74.n10 a_27_74.t2 24.3248
R178 a_27_74.n13 a_27_74.t1 23.514
R179 a_27_74.t3 a_27_74.n13 23.514
R180 a_27_74.n2 a_27_74.t13 22.7032
R181 a_27_74.n2 a_27_74.t14 22.7032
R182 a_27_74.n10 a_27_74.t9 22.7032
R183 a_27_74.n4 a_27_74.t10 22.7032
R184 a_27_74.n4 a_27_74.t8 22.7032
R185 a_27_74.n6 a_27_74.t4 22.7032
R186 a_27_74.n6 a_27_74.t5 22.7032
R187 a_27_74.n8 a_27_74.t6 22.7032
R188 a_27_74.n0 a_27_74.t15 22.7032
R189 VNB.t7 VNB.t9 1224.15
R190 VNB.t15 VNB.t0 1154.86
R191 VNB.t12 VNB.t15 1154.86
R192 VNB.t13 VNB.t12 1154.86
R193 VNB.t4 VNB.t6 1154.86
R194 VNB.t10 VNB.t5 1154.86
R195 VNB.t11 VNB.t8 1154.86
R196 VNB VNB.t11 1143.31
R197 VNB.t2 VNB.t3 1131.76
R198 VNB.t6 VNB.t7 1085.56
R199 VNB.t3 VNB.t1 1016.27
R200 VNB.t9 VNB.t2 1016.27
R201 VNB.t14 VNB.t13 993.177
R202 VNB.t1 VNB.t14 993.177
R203 VNB.t5 VNB.t4 993.177
R204 VNB.t8 VNB.t10 993.177
R205 B2.n0 B2.t1 226.809
R206 B2.n10 B2.t0 226.809
R207 B2.n3 B2.n2 226.809
R208 B2.n5 B2.t2 226.809
R209 B2.n5 B2.t5 204.048
R210 B2.n0 B2.t6 198.204
R211 B2.n4 B2.t4 196.013
R212 B2.n9 B2.t3 196.013
R213 B2.n7 B2.n6 169.409
R214 B2 B2.n1 156.207
R215 B2.n8 B2.n7 152
R216 B2.n12 B2.n11 152
R217 B2.n11 B2.n1 49.6611
R218 B2.n9 B2.n8 40.1672
R219 B2.n6 B2.n5 37.9763
R220 B2.n8 B2.n3 21.9096
R221 B2.n6 B2.n4 16.7975
R222 B2.n1 B2.n0 11.6853
R223 B2.n4 B2.n3 10.955
R224 B2.n12 B2 9.32621
R225 B2 B2.n12 8.22907
R226 B2.n11 B2.n10 5.84292
R227 B2.n7 B2 3.91364
R228 B2.n10 B2.n9 3.65202
R229 a_877_368.n0 a_877_368.t4 395.264
R230 a_877_368.n3 a_877_368.n2 362.32
R231 a_877_368.n0 a_877_368.t5 332.284
R232 a_877_368.n2 a_877_368.n1 286.729
R233 a_877_368.n2 a_877_368.n0 81.8693
R234 a_877_368.n1 a_877_368.t0 35.1791
R235 a_877_368.n1 a_877_368.t3 26.3844
R236 a_877_368.t2 a_877_368.n3 26.3844
R237 a_877_368.n3 a_877_368.t1 26.3844
R238 VGND.n6 VGND.n3 211.893
R239 VGND.n12 VGND.n11 209.048
R240 VGND.n5 VGND.n4 206.333
R241 VGND.n9 VGND.n2 206.333
R242 VGND.n3 VGND.t5 34.0546
R243 VGND.n4 VGND.t0 34.0546
R244 VGND.n2 VGND.t6 34.0546
R245 VGND.n11 VGND.t7 34.0546
R246 VGND.n3 VGND.t3 27.5681
R247 VGND.n10 VGND.n9 25.977
R248 VGND.n5 VGND.n1 23.7181
R249 VGND.n4 VGND.t2 22.7032
R250 VGND.n2 VGND.t1 22.7032
R251 VGND.n11 VGND.t4 22.7032
R252 VGND.n9 VGND.n1 21.4593
R253 VGND.n12 VGND.n10 19.2005
R254 VGND.n7 VGND.n1 9.3005
R255 VGND.n9 VGND.n8 9.3005
R256 VGND.n10 VGND.n0 9.3005
R257 VGND.n13 VGND.n12 7.43488
R258 VGND.n6 VGND.n5 6.70158
R259 VGND.n7 VGND.n6 0.570057
R260 VGND VGND.n13 0.160103
R261 VGND.n13 VGND.n0 0.1477
R262 VGND.n8 VGND.n7 0.122949
R263 VGND.n8 VGND.n0 0.122949
C0 B2 VPWR 0.023639f
C1 Y VGND 0.046132f
C2 VPB VPWR 0.215441f
C3 A1 B2 0.001913f
C4 B1 Y 0.523326f
C5 A2 VGND 0.063782f
C6 VPB A1 0.150732f
C7 A2 B1 0.003119f
C8 VPWR VGND 0.129096f
C9 VPB B2 0.138223f
C10 A2 Y 0.031489f
C11 B1 VPWR 0.064686f
C12 A1 VGND 0.066985f
C13 A1 B1 0.072575f
C14 B2 VGND 0.022452f
C15 VPWR Y 0.142626f
C16 A2 VPWR 0.025158f
C17 VPB VGND 0.010587f
C18 A1 Y 0.168355f
C19 B1 B2 0.303445f
C20 VPB B1 0.132058f
C21 A1 A2 0.303792f
C22 B2 Y 0.225421f
C23 A1 VPWR 0.081345f
C24 VPB Y 0.018689f
C25 B1 VGND 0.029471f
C26 VPB A2 0.126352f
C27 VGND VNB 0.91208f
C28 Y VNB 0.081469f
C29 VPWR VNB 0.808777f
C30 B2 VNB 0.399902f
C31 B1 VNB 0.450543f
C32 A2 VNB 0.41542f
C33 A1 VNB 0.460234f
C34 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o22ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o22ai_2 VNB VPB VPWR VGND B2 B1 A2 A1 Y
X0 a_27_74.t4 B1.t0 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1406 ps=1.12 w=0.74 l=0.15
X1 a_510_368.t2 A1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t0 A1.t1 a_510_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_510_368.t3 A2.t0 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_27_74.t0 A1.t2 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 VPWR.t3 B1.t1 a_28_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 Y.t0 A2.t1 a_510_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 a_27_74.t6 B2.t0 Y.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2812 pd=1.5 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 a_27_74.t2 A2.t2 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1184 ps=1.06 w=0.74 l=0.15
X9 Y.t1 B1.t2 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1406 pd=1.12 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 VGND.t2 A2.t3 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2812 ps=1.5 w=0.74 l=0.15
X11 VGND.t0 A1.t3 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_28_368.t3 B2.t1 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X13 Y.t6 B2.t2 a_28_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y.t3 B2.t3 a_27_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1184 ps=1.06 w=0.74 l=0.15
X15 a_28_368.t0 B1.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
R0 B1.n0 B1.t3 226.809
R1 B1.n1 B1.t1 226.809
R2 B1.n1 B1.t2 198.204
R3 B1.n0 B1.t0 198.204
R4 B1.n5 B1.n4 152
R5 B1.n3 B1.n2 152
R6 B1.n4 B1.n3 49.6611
R7 B1.n2 B1 12.8005
R8 B1.n4 B1.n0 12.4157
R9 B1.n3 B1.n1 10.955
R10 B1.n5 B1 8.63306
R11 B1 B1.n5 5.65631
R12 B1.n2 B1 1.48887
R13 Y.n2 Y.n0 364.027
R14 Y.n2 Y.n1 329.945
R15 Y.n5 Y.n3 248.441
R16 Y.n5 Y.n4 197.994
R17 Y Y.n2 37.5657
R18 Y.n3 Y.t1 34.0546
R19 Y.n4 Y.t3 34.0546
R20 Y.n3 Y.t2 27.5681
R21 Y.n1 Y.t7 26.3844
R22 Y.n1 Y.t6 26.3844
R23 Y.n0 Y.t5 26.3844
R24 Y.n0 Y.t0 26.3844
R25 Y.n4 Y.t4 22.7032
R26 Y Y.n5 13.9299
R27 a_27_74.n1 a_27_74.t0 205.819
R28 a_27_74.n6 a_27_74.t3 201.337
R29 a_27_74.n7 a_27_74.n6 197.994
R30 a_27_74.n5 a_27_74.n4 185
R31 a_27_74.n1 a_27_74.n0 102.019
R32 a_27_74.n3 a_27_74.n2 91.6858
R33 a_27_74.n4 a_27_74.n3 77.8383
R34 a_27_74.n2 a_27_74.n1 59.6989
R35 a_27_74.n6 a_27_74.n5 52.5262
R36 a_27_74.t4 a_27_74.n7 29.1897
R37 a_27_74.n3 a_27_74.t7 22.7032
R38 a_27_74.n4 a_27_74.t6 22.7032
R39 a_27_74.n0 a_27_74.t1 22.7032
R40 a_27_74.n0 a_27_74.t2 22.7032
R41 a_27_74.n7 a_27_74.t5 22.7032
R42 a_27_74.n5 a_27_74.n2 11.3748
R43 VNB.t6 VNB.t7 2101.84
R44 VNB.t3 VNB.t4 1224.15
R45 VNB.t1 VNB.t0 1154.86
R46 VNB.t5 VNB.t6 1154.86
R47 VNB VNB.t3 1143.31
R48 VNB.t7 VNB.t2 1085.56
R49 VNB.t4 VNB.t5 1085.56
R50 VNB.t2 VNB.t1 993.177
R51 A1.n3 A1.t0 226.809
R52 A1.n1 A1.t1 226.809
R53 A1.n1 A1.t3 198.204
R54 A1.n4 A1.t2 196.013
R55 A1.n5 A1.n4 168.067
R56 A1.n2 A1.n0 152
R57 A1.n2 A1.n1 37.246
R58 A1.n3 A1.n2 28.4823
R59 A1.n5 A1.n0 10.1214
R60 A1.n4 A1.n3 5.11262
R61 A1.n0 A1 2.3819
R62 A1 A1.n5 1.78655
R63 VPWR.n2 VPWR.n0 330.219
R64 VPWR.n2 VPWR.n1 321.772
R65 VPWR.n1 VPWR.t2 35.1791
R66 VPWR.n1 VPWR.t3 26.3844
R67 VPWR.n0 VPWR.t1 26.3844
R68 VPWR.n0 VPWR.t0 26.3844
R69 VPWR VPWR.n2 0.192514
R70 a_510_368.n1 a_510_368.t0 417.757
R71 a_510_368.t2 a_510_368.n1 312.199
R72 a_510_368.n1 a_510_368.n0 183.911
R73 a_510_368.n0 a_510_368.t1 26.3844
R74 a_510_368.n0 a_510_368.t3 26.3844
R75 VPB.t7 VPB.t0 515.861
R76 VPB VPB.t4 260.485
R77 VPB.t4 VPB.t3 255.376
R78 VPB.t1 VPB.t2 229.839
R79 VPB.t5 VPB.t1 229.839
R80 VPB.t0 VPB.t5 229.839
R81 VPB.t6 VPB.t7 229.839
R82 VPB.t3 VPB.t6 229.839
R83 A2.n1 A2.t0 240.197
R84 A2.n2 A2.t1 240.197
R85 A2.n1 A2.t2 180.678
R86 A2.n0 A2.t3 179.947
R87 A2.n4 A2.n0 176.143
R88 A2.n4 A2.n3 152
R89 A2.n3 A2.n2 36.5157
R90 A2.n3 A2.n1 29.2126
R91 A2 A2.n4 16.0005
R92 A2.n2 A2.n0 2.19141
R93 VGND.n2 VGND.n0 216.948
R94 VGND.n2 VGND.n1 214.714
R95 VGND.n0 VGND.t0 34.0546
R96 VGND.n1 VGND.t3 29.1897
R97 VGND.n0 VGND.t1 22.7032
R98 VGND.n1 VGND.t2 22.7032
R99 VGND VGND.n2 1.10625
R100 a_28_368.n1 a_28_368.t3 392.853
R101 a_28_368.t1 a_28_368.n1 304.238
R102 a_28_368.n1 a_28_368.n0 189.115
R103 a_28_368.n0 a_28_368.t2 26.3844
R104 a_28_368.n0 a_28_368.t0 26.3844
R105 B2.n1 B2.t2 231.921
R106 B2.n0 B2.t1 226.809
R107 B2.n0 B2.t0 212.448
R108 B2.n1 B2.t3 196.013
R109 B2 B2.n2 154.522
R110 B2.n2 B2.n0 37.9763
R111 B2.n2 B2.n1 22.6399
C0 VPB B1 0.070874f
C1 A1 VPB 0.076334f
C2 B2 A2 0.021659f
C3 Y B2 0.156325f
C4 VGND B1 0.014309f
C5 VPWR A2 0.012963f
C6 A1 VGND 0.035976f
C7 VPWR Y 0.025466f
C8 VGND VPB 0.008337f
C9 Y B1 0.081507f
C10 VPWR B2 0.01203f
C11 A1 A2 0.095472f
C12 A1 Y 0.001283f
C13 B1 B2 0.094846f
C14 VPB A2 0.074236f
C15 Y VPB 0.018184f
C16 VPWR B1 0.041015f
C17 A1 VPWR 0.037169f
C18 VGND A2 0.036306f
C19 Y VGND 0.023245f
C20 VPB B2 0.067198f
C21 VPWR VPB 0.122665f
C22 VGND B2 0.01209f
C23 Y A2 0.104337f
C24 VPWR VGND 0.074901f
C25 VGND VNB 0.565559f
C26 Y VNB 0.037599f
C27 VPWR VNB 0.464578f
C28 A1 VNB 0.260763f
C29 A2 VNB 0.224097f
C30 B2 VNB 0.206303f
C31 B1 VNB 0.252182f
C32 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o22ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o22ai_1 VNB VPB VPWR VGND B2 B1 Y A2 A1
X0 VGND.t1 A2.t0 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 Y.t0 B2.t0 a_142_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X2 a_27_74.t1 B2.t1 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.21275 ps=1.315 w=0.74 l=0.15
X3 Y.t3 B1.t0 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.21275 pd=1.315 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 a_27_74.t0 A1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 a_142_368.t0 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.4648 ps=3.07 w=1.12 l=0.15
X6 a_340_368.t1 A2.t1 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X7 VPWR.t1 A1.t1 a_340_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
R0 A2.n0 A2.t1 250.909
R1 A2.n0 A2.t0 220.113
R2 A2 A2.n0 155.126
R3 a_27_74.n1 a_27_74.t3 224.279
R4 a_27_74.t0 a_27_74.n1 209.089
R5 a_27_74.n1 a_27_74.n0 88.3339
R6 a_27_74.n0 a_27_74.t1 34.0546
R7 a_27_74.n0 a_27_74.t2 22.7032
R8 VGND VGND.n0 215.262
R9 VGND.n0 VGND.t0 34.0546
R10 VGND.n0 VGND.t1 34.0546
R11 VNB.t3 VNB.t1 1674.54
R12 VNB.t2 VNB.t0 1316.54
R13 VNB.t1 VNB.t2 1154.86
R14 VNB VNB.t3 1143.31
R15 B2.n0 B2.t0 250.909
R16 B2.n0 B2.t1 220.113
R17 B2 B2.n0 154.377
R18 a_142_368.t0 a_142_368.t1 47.4916
R19 Y Y.n0 586.731
R20 Y.n3 Y.n0 585
R21 Y.n2 Y.n0 585
R22 Y.n2 Y.n1 257.274
R23 Y.n1 Y.t1 47.0275
R24 Y.n1 Y.t3 46.2167
R25 Y.n0 Y.t2 37.8175
R26 Y.n0 Y.t0 36.0585
R27 Y Y.n3 3.11401
R28 Y Y.n2 2.83726
R29 Y.n3 Y 2.00699
R30 VPB VPB.t0 324.329
R31 VPB.t2 VPB.t3 291.13
R32 VPB.t1 VPB.t2 291.13
R33 VPB.t0 VPB.t1 214.517
R34 B1.n0 B1.t1 287.793
R35 B1.n0 B1.t0 171.72
R36 B1 B1.n0 158.788
R37 A1.n1 A1.t1 251.151
R38 A1.n0 A1 200.207
R39 A1.n0 A1.t0 179.947
R40 A1.n2 A1.n1 152
R41 A1.n2 A1 7.6005
R42 A1 A1.n2 5.2005
R43 A1.n1 A1.n0 2.92171
R44 VPWR.n0 VPWR.t0 278.111
R45 VPWR.n0 VPWR.t1 256.252
R46 VPWR VPWR.n0 0.105349
R47 a_340_368.t0 a_340_368.t1 73.8755
C0 B2 VPWR 0.005328f
C1 A2 A1 0.083724f
C2 B1 B2 0.048808f
C3 VPB A2 0.035513f
C4 Y B2 0.101923f
C5 VGND VPWR 0.047512f
C6 B1 VGND 0.007823f
C7 B2 A1 1.37e-19
C8 VPB B2 0.032767f
C9 B1 VPWR 0.039f
C10 Y VGND 0.013685f
C11 Y VPWR 0.231996f
C12 VGND A1 0.01926f
C13 VPB VGND 0.007678f
C14 B1 Y 0.061303f
C15 B2 A2 0.081229f
C16 A1 VPWR 0.059166f
C17 VPB VPWR 0.10598f
C18 VPB B1 0.044948f
C19 VGND A2 0.012652f
C20 Y A1 0.004846f
C21 VPB Y 0.01142f
C22 A2 VPWR 0.018089f
C23 VPB A1 0.059774f
C24 Y A2 0.012028f
C25 VGND B2 0.006232f
C26 VGND VNB 0.37717f
C27 Y VNB 0.032912f
C28 VPWR VNB 0.387424f
C29 A1 VNB 0.19261f
C30 A2 VNB 0.105064f
C31 B2 VNB 0.108046f
C32 B1 VNB 0.180554f
C33 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o22a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o22a_4 VNB VPB VPWR VGND B1 X A1 A2 B2
X0 a_116_392.t1 A1.t0 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X1 VPWR.t6 A1.t1 a_116_392.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.175 ps=1.35 w=1 l=0.15
X2 a_516_392.t3 B2.t0 a_206_392.t4 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X3 VGND.t1 A2.t0 a_27_136.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 a_206_392.t6 B2.t1 a_27_136.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1136 ps=0.995 w=0.64 l=0.15
X5 X.t3 a_206_392.t8 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.2186 ps=1.52 w=1.12 l=0.15
X6 VPWR.t2 a_206_392.t9 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X7 X.t1 a_206_392.t10 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.322 ps=1.695 w=1.12 l=0.15
X8 a_27_136.t3 A1.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.12 pd=1.015 as=0.1248 ps=1.03 w=0.64 l=0.15
X9 a_27_136.t5 B2.t2 a_206_392.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1136 pd=0.995 as=0.0912 ps=0.925 w=0.64 l=0.15
X10 a_116_392.t2 A2.t1 a_206_392.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X11 X.t6 a_206_392.t11 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VPWR.t4 a_206_392.t12 X.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.322 pd=1.695 as=0.1876 ps=1.455 w=1.12 l=0.15
X13 a_206_392.t3 B2.t3 a_516_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X14 a_516_392.t1 B1.t0 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X15 a_27_136.t4 B1.t1 a_206_392.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 X.t5 a_206_392.t13 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2991 ps=2.41 w=0.74 l=0.15
X17 a_206_392.t1 A2.t2 a_116_392.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND.t2 A1.t3 a_27_136.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X19 VGND.t6 a_206_392.t14 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t0 B1.t2 a_516_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2186 pd=1.52 as=0.175 ps=1.35 w=1 l=0.15
X21 a_206_392.t7 B1.t3 a_27_136.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0912 pd=0.925 as=0.12 ps=1.015 w=0.64 l=0.15
X22 a_27_136.t0 A2.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
R0 A1.t2 A1.t3 915.801
R1 A1.t3 A1.t0 449.384
R2 A1.n0 A1.t1 236.983
R3 A1.n0 A1.t2 168.701
R4 A1 A1.n0 154.522
R5 VPWR.n8 VPWR.n7 316.87
R6 VPWR.n20 VPWR.n3 315.928
R7 VPWR.n9 VPWR.t2 265.644
R8 VPWR.n26 VPWR.t7 260.733
R9 VPWR.n13 VPWR.n6 223.389
R10 VPWR.n7 VPWR.t4 52.7684
R11 VPWR.n7 VPWR.t3 48.371
R12 VPWR.n6 VPWR.t0 46.2955
R13 VPWR.n3 VPWR.t5 39.4005
R14 VPWR.n3 VPWR.t6 39.4005
R15 VPWR.n24 VPWR.n1 36.1417
R16 VPWR.n25 VPWR.n24 36.1417
R17 VPWR.n14 VPWR.n4 36.1417
R18 VPWR.n18 VPWR.n4 36.1417
R19 VPWR.n19 VPWR.n18 36.1417
R20 VPWR.n12 VPWR.n11 36.1417
R21 VPWR.n6 VPWR.t1 29.4992
R22 VPWR.n20 VPWR.n1 28.9887
R23 VPWR.n26 VPWR.n25 26.7299
R24 VPWR.n20 VPWR.n19 18.4476
R25 VPWR.n11 VPWR.n8 12.0476
R26 VPWR.n13 VPWR.n12 9.78874
R27 VPWR.n11 VPWR.n10 9.3005
R28 VPWR.n12 VPWR.n5 9.3005
R29 VPWR.n15 VPWR.n14 9.3005
R30 VPWR.n16 VPWR.n4 9.3005
R31 VPWR.n18 VPWR.n17 9.3005
R32 VPWR.n19 VPWR.n2 9.3005
R33 VPWR.n21 VPWR.n20 9.3005
R34 VPWR.n22 VPWR.n1 9.3005
R35 VPWR.n24 VPWR.n23 9.3005
R36 VPWR.n25 VPWR.n0 9.3005
R37 VPWR.n27 VPWR.n26 9.3005
R38 VPWR.n9 VPWR.n8 7.21497
R39 VPWR.n14 VPWR.n13 1.50638
R40 VPWR.n10 VPWR.n9 0.543582
R41 VPWR.n10 VPWR.n5 0.122949
R42 VPWR.n15 VPWR.n5 0.122949
R43 VPWR.n16 VPWR.n15 0.122949
R44 VPWR.n17 VPWR.n16 0.122949
R45 VPWR.n17 VPWR.n2 0.122949
R46 VPWR.n21 VPWR.n2 0.122949
R47 VPWR.n22 VPWR.n21 0.122949
R48 VPWR.n23 VPWR.n22 0.122949
R49 VPWR.n23 VPWR.n0 0.122949
R50 VPWR.n27 VPWR.n0 0.122949
R51 VPWR VPWR.n27 0.0617245
R52 a_116_392.n1 a_116_392.n0 562.359
R53 a_116_392.n0 a_116_392.t2 39.4005
R54 a_116_392.n0 a_116_392.t0 29.5505
R55 a_116_392.n1 a_116_392.t3 29.5505
R56 a_116_392.t1 a_116_392.n1 29.5505
R57 VPB.t6 VPB.t5 370.296
R58 VPB.t0 VPB.t3 280.914
R59 VPB.t8 VPB.t7 280.914
R60 VPB VPB.t9 257.93
R61 VPB.t1 VPB.t0 255.376
R62 VPB.t2 VPB.t1 255.376
R63 VPB.t10 VPB.t8 255.376
R64 VPB.t11 VPB.t10 255.376
R65 VPB.t3 VPB.t6 247.715
R66 VPB.t5 VPB.t4 229.839
R67 VPB.t7 VPB.t2 229.839
R68 VPB.t9 VPB.t11 229.839
R69 B2.n0 B2.t0 213.614
R70 B2.n2 B2.t3 212.883
R71 B2 B2.n1 163.831
R72 B2.n4 B2.n3 152
R73 B2.n2 B2.t2 148.982
R74 B2.n0 B2.t1 140.88
R75 B2.n3 B2.n1 49.6611
R76 B2.n4 B2 17.2611
R77 B2.n1 B2.n0 16.0672
R78 B2.n3 B2.n2 6.57323
R79 B2 B2.n4 1.35808
R80 a_206_392.n19 a_206_392.n18 425.692
R81 a_206_392.n18 a_206_392.n17 299.95
R82 a_206_392.n4 a_206_392.n2 247.88
R83 a_206_392.n14 a_206_392.t8 237.762
R84 a_206_392.n7 a_206_392.t9 226.809
R85 a_206_392.n9 a_206_392.t10 226.809
R86 a_206_392.n13 a_206_392.t12 226.809
R87 a_206_392.n7 a_206_392.n6 205.796
R88 a_206_392.n1 a_206_392.t13 196.013
R89 a_206_392.n5 a_206_392.t14 196.013
R90 a_206_392.n8 a_206_392.t11 196.013
R91 a_206_392.n4 a_206_392.n3 185
R92 a_206_392.n11 a_206_392.n10 165.189
R93 a_206_392.n15 a_206_392.n14 152
R94 a_206_392.n1 a_206_392.n0 152
R95 a_206_392.n12 a_206_392.n11 152
R96 a_206_392.n18 a_206_392.n16 100.427
R97 a_206_392.n16 a_206_392.n4 92.453
R98 a_206_392.n8 a_206_392.n7 54.7732
R99 a_206_392.n14 a_206_392.n1 49.6611
R100 a_206_392.n13 a_206_392.n12 39.4369
R101 a_206_392.n17 a_206_392.t3 39.4005
R102 a_206_392.n19 a_206_392.t1 39.4005
R103 a_206_392.n10 a_206_392.n5 35.055
R104 a_206_392.n17 a_206_392.t4 29.5505
R105 a_206_392.t0 a_206_392.n19 29.5505
R106 a_206_392.n2 a_206_392.t7 27.188
R107 a_206_392.n3 a_206_392.t2 26.2505
R108 a_206_392.n3 a_206_392.t6 26.2505
R109 a_206_392.n2 a_206_392.t5 26.2505
R110 a_206_392.n10 a_206_392.n9 16.7975
R111 a_206_392.n12 a_206_392.n5 14.6066
R112 a_206_392.n11 a_206_392.n0 13.1884
R113 a_206_392.n15 a_206_392.n0 13.1884
R114 a_206_392.n9 a_206_392.n8 10.955
R115 a_206_392.n1 a_206_392.n13 10.2247
R116 a_206_392.n16 a_206_392.n15 3.10353
R117 a_516_392.n1 a_516_392.n0 655.923
R118 a_516_392.n0 a_516_392.t3 39.4005
R119 a_516_392.n0 a_516_392.t0 29.5505
R120 a_516_392.t2 a_516_392.n1 29.5505
R121 a_516_392.n1 a_516_392.t1 29.5505
R122 A2.n1 A2.t2 218.726
R123 A2.n0 A2.t1 216.254
R124 A2.n1 A2.t3 144.601
R125 A2.n0 A2.t0 142.994
R126 A2 A2.n2 68.5461
R127 A2.n2 A2.n0 33.4961
R128 A2.n2 A2.n1 23.3196
R129 a_27_136.n4 a_27_136.t4 316.649
R130 a_27_136.n1 a_27_136.t2 186.381
R131 a_27_136.n1 a_27_136.n0 185
R132 a_27_136.n3 a_27_136.n2 185
R133 a_27_136.n5 a_27_136.n4 185
R134 a_27_136.n4 a_27_136.n3 58.6952
R135 a_27_136.n3 a_27_136.n1 58.654
R136 a_27_136.n2 a_27_136.t7 38.438
R137 a_27_136.t6 a_27_136.n5 33.7505
R138 a_27_136.n5 a_27_136.t5 32.813
R139 a_27_136.n2 a_27_136.t3 31.8755
R140 a_27_136.n0 a_27_136.t1 26.2505
R141 a_27_136.n0 a_27_136.t0 26.2505
R142 VGND.n6 VGND.t4 307.947
R143 VGND.n16 VGND.n2 217.583
R144 VGND.n19 VGND.n18 217.583
R145 VGND.n7 VGND.n5 214.775
R146 VGND.n2 VGND.t1 39.3755
R147 VGND.n18 VGND.t2 39.3755
R148 VGND.n10 VGND.n4 36.1417
R149 VGND.n11 VGND.n10 36.1417
R150 VGND.n12 VGND.n11 36.1417
R151 VGND.n12 VGND.n1 36.1417
R152 VGND.n2 VGND.t3 33.7505
R153 VGND.n6 VGND.n4 29.3652
R154 VGND.n18 VGND.t0 26.2505
R155 VGND.n17 VGND.n16 25.977
R156 VGND.n5 VGND.t5 22.7032
R157 VGND.n5 VGND.t6 22.7032
R158 VGND.n16 VGND.n1 21.4593
R159 VGND.n19 VGND.n17 19.2005
R160 VGND.n8 VGND.n4 9.3005
R161 VGND.n10 VGND.n9 9.3005
R162 VGND.n11 VGND.n3 9.3005
R163 VGND.n13 VGND.n12 9.3005
R164 VGND.n14 VGND.n1 9.3005
R165 VGND.n16 VGND.n15 9.3005
R166 VGND.n17 VGND.n0 9.3005
R167 VGND.n20 VGND.n19 7.43488
R168 VGND.n7 VGND.n6 6.39061
R169 VGND.n8 VGND.n7 0.551106
R170 VGND VGND.n20 0.160103
R171 VGND.n20 VGND.n0 0.1477
R172 VGND.n9 VGND.n8 0.122949
R173 VGND.n9 VGND.n3 0.122949
R174 VGND.n13 VGND.n3 0.122949
R175 VGND.n14 VGND.n13 0.122949
R176 VGND.n15 VGND.n14 0.122949
R177 VGND.n15 VGND.n0 0.122949
R178 VNB.t7 VNB.t5 2471.39
R179 VNB.t1 VNB.t3 1247.24
R180 VNB.t3 VNB.t10 1212.6
R181 VNB.t8 VNB.t9 1166.4
R182 VNB.t2 VNB.t0 1154.86
R183 VNB VNB.t2 1143.31
R184 VNB.t10 VNB.t8 1004.72
R185 VNB.t4 VNB.t6 993.177
R186 VNB.t5 VNB.t4 993.177
R187 VNB.t9 VNB.t7 993.177
R188 VNB.t0 VNB.t1 993.177
R189 X.n2 X.n0 270.14
R190 X.n2 X.n1 206.517
R191 X.n4 X.t6 157.087
R192 X.n4 X.n3 156.532
R193 X.n5 X.n2 36.4269
R194 X.n0 X.t3 32.5407
R195 X.n1 X.t2 26.3844
R196 X.n1 X.t1 26.3844
R197 X.n0 X.t0 26.3844
R198 X.n3 X.t4 22.7032
R199 X.n3 X.t5 22.7032
R200 X X.n5 20.8701
R201 X.n5 X.n4 5.88158
R202 B1.n0 B1.t1 648.217
R203 B1.t3 B1.t0 442.904
R204 B1.t1 B1.t2 430.546
R205 B1.n1 B1.n0 163.582
R206 B1.n0 B1.t3 162.274
R207 B1 B1.n1 5.56572
R208 B1.n1 B1 3.45447
C0 B1 A1 0.082105f
C1 B2 VPB 0.080826f
C2 VGND A2 0.021678f
C3 B2 VGND 0.009262f
C4 B2 X 1.25e-19
C5 VPB A1 0.081076f
C6 B1 VPB 0.073465f
C7 VGND A1 0.089332f
C8 VPWR A2 0.01181f
C9 B1 VGND 0.151638f
C10 B2 VPWR 0.012655f
C11 B1 X 0.002543f
C12 VGND VPB 0.011241f
C13 X VPB 0.015267f
C14 VPWR A1 0.035756f
C15 B1 VPWR 0.039002f
C16 X VGND 0.276142f
C17 A1 A2 0.138091f
C18 B2 A1 0.021577f
C19 VPWR VPB 0.189417f
C20 B1 B2 0.137699f
C21 VPWR VGND 0.112018f
C22 VPWR X 0.446557f
C23 VPB A2 0.080002f
C24 VGND VNB 0.848287f
C25 X VNB 0.05157f
C26 VPWR VNB 0.706456f
C27 B2 VNB 0.159082f
C28 B1 VNB 0.387475f
C29 A2 VNB 0.166982f
C30 A1 VNB 0.39914f
C31 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o31ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o31ai_4 VNB VPB VPWR VGND Y B1 A3 A2 A1
X0 a_27_82.t13 A3.t0 VGND.t11 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3627 ps=1.75 w=0.74 l=0.15
X1 Y.t3 B1.t0 a_27_82.t14 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t4 B1.t1 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.5852 ps=2.165 w=1.12 l=0.15
X3 a_27_82.t8 A2.t0 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2183 ps=1.33 w=0.74 l=0.15
X4 a_28_368.t7 A2.t1 a_487_368.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=1.69 as=0.196 ps=1.47 w=1.12 l=0.15
X5 VPWR.t0 A1.t0 a_28_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 a_27_82.t9 A1.t1 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 a_487_368.t1 A3.t1 Y.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8 VGND.t4 A1.t2 a_27_82.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_487_368.t5 A2.t2 a_28_368.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t0 A2.t3 a_27_82.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2183 pd=1.33 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_28_368.t5 A2.t4 a_487_368.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_28_368.t2 A1.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X13 VGND.t5 A1.t4 a_27_82.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_27_82.t1 A2.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0.5852 pd=2.165 as=0.196 ps=1.47 w=1.12 l=0.15
X16 a_27_82.t15 B1.t2 Y.t2 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_27_82.t6 B1.t3 Y.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_487_368.t3 A2.t6 a_28_368.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=1.69 w=1.12 l=0.15
X19 VGND.t10 A3.t2 a_27_82.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.3627 pd=1.75 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VGND.t9 A3.t3 a_27_82.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.201 pd=1.42 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VPWR.t3 A1.t5 a_28_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_27_82.t3 A1.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X23 a_28_368.t1 A1.t7 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 VGND.t2 A2.t7 a_27_82.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X25 a_27_82.t10 A3.t4 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.201 ps=1.42 w=0.74 l=0.15
X26 Y.t0 B1.t4 a_27_82.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 a_487_368.t0 A3.t5 Y.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A3.n6 A3.t2 329.368
R1 A3.n2 A3.t5 253.587
R2 A3.n1 A3.n0 243.483
R3 A3.n11 A3.n4 226.809
R4 A3.n5 A3.t1 226.809
R5 A3.n1 A3.t4 224.934
R6 A3.n10 A3.t0 183.161
R7 A3.n3 A3.t3 183.161
R8 A3.n13 A3.n12 152
R9 A3.n9 A3.n8 152
R10 A3.n7 A3.n6 152
R11 A3.n2 A3.n1 117.555
R12 A3.n9 A3.n5 36.5157
R13 A3.n12 A3.n3 21.1793
R14 A3.n11 A3.n10 21.1793
R15 A3.n12 A3.n11 20.449
R16 A3.n6 A3.n5 13.146
R17 A3.n3 A3.n2 10.955
R18 A3.n8 A3.n7 10.1214
R19 A3.n10 A3.n9 8.03383
R20 A3.n13 A3 7.29352
R21 A3 A3.n13 6.99585
R22 A3.n8 A3 2.82841
R23 A3.n7 A3 1.34003
R24 VGND.n12 VGND.n11 280.455
R25 VGND.n13 VGND.n12 280.455
R26 VGND.n10 VGND.n9 225.596
R27 VGND.n5 VGND.n4 210.406
R28 VGND.n25 VGND.n2 207.109
R29 VGND.n28 VGND.n27 207.109
R30 VGND.n21 VGND.n20 203.444
R31 VGND.n12 VGND.t11 64.0546
R32 VGND.n12 VGND.t10 64.0546
R33 VGND.n20 VGND.t6 47.8383
R34 VGND.n20 VGND.t0 47.8383
R35 VGND.n9 VGND.t8 36.487
R36 VGND.n9 VGND.t9 36.487
R37 VGND.n15 VGND.n14 36.1417
R38 VGND.n19 VGND.n18 36.1417
R39 VGND.n2 VGND.t7 34.0546
R40 VGND.n27 VGND.t4 34.0546
R41 VGND.n11 VGND.n10 29.2129
R42 VGND.n25 VGND.n1 26.7299
R43 VGND.n21 VGND.n1 25.224
R44 VGND.n4 VGND.t1 22.7032
R45 VGND.n4 VGND.t2 22.7032
R46 VGND.n2 VGND.t5 22.7032
R47 VGND.n27 VGND.t3 22.7032
R48 VGND.n26 VGND.n25 20.7064
R49 VGND.n28 VGND.n26 19.2005
R50 VGND.n21 VGND.n19 12.0476
R51 VGND.n26 VGND.n0 9.3005
R52 VGND.n25 VGND.n24 9.3005
R53 VGND.n23 VGND.n1 9.3005
R54 VGND.n22 VGND.n21 9.3005
R55 VGND.n8 VGND.n7 9.3005
R56 VGND.n14 VGND.n6 9.3005
R57 VGND.n16 VGND.n15 9.3005
R58 VGND.n18 VGND.n17 9.3005
R59 VGND.n19 VGND.n3 9.3005
R60 VGND.n15 VGND.n5 7.90638
R61 VGND.n29 VGND.n28 7.43488
R62 VGND.n13 VGND.n7 6.3458
R63 VGND.n14 VGND.n13 5.49311
R64 VGND.n18 VGND.n5 3.38874
R65 VGND.n11 VGND.n7 1.31332
R66 VGND.n10 VGND.n8 1.30579
R67 VGND VGND.n29 0.160103
R68 VGND.n29 VGND.n0 0.1477
R69 VGND.n8 VGND.n6 0.122949
R70 VGND.n16 VGND.n6 0.122949
R71 VGND.n17 VGND.n16 0.122949
R72 VGND.n17 VGND.n3 0.122949
R73 VGND.n22 VGND.n3 0.122949
R74 VGND.n23 VGND.n22 0.122949
R75 VGND.n24 VGND.n23 0.122949
R76 VGND.n24 VGND.n0 0.122949
R77 a_27_82.n1 a_27_82.t15 199.03
R78 a_27_82.n5 a_27_82.n4 185
R79 a_27_82.n1 a_27_82.n0 185
R80 a_27_82.n3 a_27_82.n2 185
R81 a_27_82.n13 a_27_82.n12 185
R82 a_27_82.n5 a_27_82.t4 183.508
R83 a_27_82.n12 a_27_82.n11 101.576
R84 a_27_82.n9 a_27_82.n8 100.159
R85 a_27_82.n7 a_27_82.n6 98.414
R86 a_27_82.n11 a_27_82.n10 91.6106
R87 a_27_82.n9 a_27_82.n7 64.993
R88 a_27_82.n11 a_27_82.n9 63.8544
R89 a_27_82.n12 a_27_82.n3 63.2664
R90 a_27_82.n3 a_27_82.n1 51.6397
R91 a_27_82.n7 a_27_82.n5 37.662
R92 a_27_82.n8 a_27_82.t2 34.0546
R93 a_27_82.n10 a_27_82.t12 22.7032
R94 a_27_82.n10 a_27_82.t1 22.7032
R95 a_27_82.n6 a_27_82.t0 22.7032
R96 a_27_82.n6 a_27_82.t9 22.7032
R97 a_27_82.n4 a_27_82.t5 22.7032
R98 a_27_82.n4 a_27_82.t3 22.7032
R99 a_27_82.n8 a_27_82.t8 22.7032
R100 a_27_82.n2 a_27_82.t14 22.7032
R101 a_27_82.n2 a_27_82.t10 22.7032
R102 a_27_82.n0 a_27_82.t7 22.7032
R103 a_27_82.n0 a_27_82.t6 22.7032
R104 a_27_82.n13 a_27_82.t11 22.7032
R105 a_27_82.t13 a_27_82.n13 22.7032
R106 VNB.t12 VNB.t13 2171.13
R107 VNB.t0 VNB.t8 1709.19
R108 VNB.t11 VNB.t10 1385.83
R109 VNB.t8 VNB.t2 1154.86
R110 VNB.t5 VNB.t9 1154.86
R111 VNB.t4 VNB.t3 1154.86
R112 VNB VNB.t4 1143.31
R113 VNB.t7 VNB.t15 993.177
R114 VNB.t6 VNB.t7 993.177
R115 VNB.t14 VNB.t6 993.177
R116 VNB.t10 VNB.t14 993.177
R117 VNB.t13 VNB.t11 993.177
R118 VNB.t1 VNB.t12 993.177
R119 VNB.t2 VNB.t1 993.177
R120 VNB.t9 VNB.t0 993.177
R121 VNB.t3 VNB.t5 993.177
R122 B1.n0 B1.t1 295.091
R123 B1.n5 B1.n4 226.809
R124 B1.n0 B1.t2 201.948
R125 B1.n5 B1.t0 195.576
R126 B1.n7 B1.t3 183.161
R127 B1.n1 B1.t4 183.161
R128 B1 B1.n2 160.037
R129 B1.n8 B1.n7 152
R130 B1.n6 B1.n3 152
R131 B1.n1 B1.n0 92.895
R132 B1.n7 B1.n2 49.6611
R133 B1.n7 B1.n6 49.6611
R134 B1.n2 B1.n1 13.146
R135 B1.n8 B1.n3 10.1214
R136 B1 B1.n8 2.08422
R137 B1.n3 B1 2.08422
R138 B1.n6 B1.n5 0.730803
R139 Y.n4 Y.t6 386.01
R140 Y.n3 Y.t4 375.205
R141 Y.n3 Y.t5 374.149
R142 Y.n2 Y.n0 227.339
R143 Y.n5 Y.n2 211.042
R144 Y.n2 Y.n1 185
R145 Y.n4 Y.n3 47.8159
R146 Y.n1 Y.t1 22.7032
R147 Y.n1 Y.t3 22.7032
R148 Y.n0 Y.t2 22.7032
R149 Y.n0 Y.t0 22.7032
R150 Y Y.n5 12.4805
R151 Y.n5 Y.n4 4.38555
R152 VPWR.n15 VPWR.n14 361.099
R153 VPWR.n33 VPWR.n3 315.928
R154 VPWR.n35 VPWR.n1 315.926
R155 VPWR.n14 VPWR.n13 292.5
R156 VPWR.n12 VPWR.n11 292.5
R157 VPWR.n14 VPWR.n11 62.4425
R158 VPWR.n16 VPWR.n8 36.1417
R159 VPWR.n20 VPWR.n8 36.1417
R160 VPWR.n21 VPWR.n20 36.1417
R161 VPWR.n22 VPWR.n21 36.1417
R162 VPWR.n22 VPWR.n6 36.1417
R163 VPWR.n26 VPWR.n6 36.1417
R164 VPWR.n27 VPWR.n26 36.1417
R165 VPWR.n28 VPWR.n27 36.1417
R166 VPWR.n28 VPWR.n4 36.1417
R167 VPWR.n32 VPWR.n4 36.1417
R168 VPWR.n3 VPWR.t2 35.1791
R169 VPWR.n33 VPWR.n32 27.1064
R170 VPWR.n11 VPWR.t4 26.3844
R171 VPWR.n1 VPWR.t1 26.3844
R172 VPWR.n1 VPWR.t0 26.3844
R173 VPWR.n3 VPWR.t3 26.3844
R174 VPWR.n35 VPWR.n34 22.5887
R175 VPWR.n34 VPWR.n33 20.3299
R176 VPWR.n10 VPWR.n9 9.3005
R177 VPWR.n17 VPWR.n16 9.3005
R178 VPWR.n18 VPWR.n8 9.3005
R179 VPWR.n20 VPWR.n19 9.3005
R180 VPWR.n21 VPWR.n7 9.3005
R181 VPWR.n23 VPWR.n22 9.3005
R182 VPWR.n24 VPWR.n6 9.3005
R183 VPWR.n26 VPWR.n25 9.3005
R184 VPWR.n27 VPWR.n5 9.3005
R185 VPWR.n29 VPWR.n28 9.3005
R186 VPWR.n30 VPWR.n4 9.3005
R187 VPWR.n32 VPWR.n31 9.3005
R188 VPWR.n33 VPWR.n2 9.3005
R189 VPWR.n34 VPWR.n0 9.3005
R190 VPWR.n16 VPWR.n15 8.08542
R191 VPWR.n12 VPWR.n9 7.74056
R192 VPWR.n36 VPWR.n35 7.28976
R193 VPWR.n13 VPWR.n12 4.03961
R194 VPWR.n15 VPWR.n10 3.12939
R195 VPWR.n13 VPWR.n10 1.30894
R196 VPWR VPWR.n36 0.158192
R197 VPWR.n36 VPWR.n0 0.149586
R198 VPWR.n17 VPWR.n9 0.122949
R199 VPWR.n18 VPWR.n17 0.122949
R200 VPWR.n19 VPWR.n18 0.122949
R201 VPWR.n19 VPWR.n7 0.122949
R202 VPWR.n23 VPWR.n7 0.122949
R203 VPWR.n24 VPWR.n23 0.122949
R204 VPWR.n25 VPWR.n24 0.122949
R205 VPWR.n25 VPWR.n5 0.122949
R206 VPWR.n29 VPWR.n5 0.122949
R207 VPWR.n30 VPWR.n29 0.122949
R208 VPWR.n31 VPWR.n30 0.122949
R209 VPWR.n31 VPWR.n2 0.122949
R210 VPWR.n2 VPWR.n0 0.122949
R211 VPB.t7 VPB.t6 1095.56
R212 VPB.t2 VPB.t8 541.399
R213 VPB.t8 VPB.t7 459.678
R214 VPB.t10 VPB.t3 367.743
R215 VPB VPB.t0 260.485
R216 VPB.t9 VPB.t10 255.376
R217 VPB.t5 VPB.t4 255.376
R218 VPB.t3 VPB.t2 229.839
R219 VPB.t4 VPB.t9 229.839
R220 VPB.t1 VPB.t5 229.839
R221 VPB.t0 VPB.t1 229.839
R222 A2.n4 A2.t2 296.272
R223 A2.n1 A2.t5 263.594
R224 A2.n1 A2.t4 251.471
R225 A2.n3 A2.t6 226.809
R226 A2.n7 A2.t1 226.809
R227 A2.n4 A2.t3 204.425
R228 A2.n8 A2.t0 183.161
R229 A2.n2 A2.t7 183.161
R230 A2.n11 A2.n10 152
R231 A2.n9 A2.n0 152
R232 A2.n6 A2.n5 152
R233 A2.n2 A2.n1 97.715
R234 A2.n6 A2.n4 91.5805
R235 A2.n10 A2.n9 49.6611
R236 A2.n8 A2.n7 34.3247
R237 A2.n10 A2.n3 10.955
R238 A2.n9 A2.n8 10.2247
R239 A2.n11 A2.n0 10.1214
R240 A2.n5 A2 8.03771
R241 A2.n5 A2 6.25166
R242 A2.n7 A2.n6 5.11262
R243 A2 A2.n0 3.87027
R244 A2.n3 A2.n2 2.19141
R245 A2 A2.n11 0.298174
R246 a_487_368.n2 a_487_368.n1 585
R247 a_487_368.n3 a_487_368.t0 387.346
R248 a_487_368.n2 a_487_368.n0 371.772
R249 a_487_368.t1 a_487_368.n3 332.382
R250 a_487_368.n3 a_487_368.n2 94.6339
R251 a_487_368.n0 a_487_368.t5 35.1791
R252 a_487_368.n1 a_487_368.t4 26.3844
R253 a_487_368.n1 a_487_368.t3 26.3844
R254 a_487_368.n0 a_487_368.t2 26.3844
R255 a_28_368.n3 a_28_368.t5 695.759
R256 a_28_368.n1 a_28_368.t0 296.526
R257 a_28_368.n3 a_28_368.n2 290.351
R258 a_28_368.n1 a_28_368.n0 208.897
R259 a_28_368.n5 a_28_368.n4 203.127
R260 a_28_368.n2 a_28_368.t4 65.0809
R261 a_28_368.n4 a_28_368.n3 60.047
R262 a_28_368.n4 a_28_368.n1 59.1064
R263 a_28_368.n2 a_28_368.t7 35.1791
R264 a_28_368.n0 a_28_368.t3 26.3844
R265 a_28_368.n0 a_28_368.t1 26.3844
R266 a_28_368.t6 a_28_368.n5 26.3844
R267 a_28_368.n5 a_28_368.t2 26.3844
R268 A1.n0 A1.t3 295.091
R269 A1.n2 A1.t5 226.809
R270 A1.n8 A1.t7 226.809
R271 A1.n3 A1.t0 226.809
R272 A1.n0 A1.t1 203.244
R273 A1.n3 A1.t2 185.351
R274 A1.n9 A1.t6 183.161
R275 A1.n1 A1.t4 183.161
R276 A1.n11 A1.n10 152
R277 A1.n7 A1.n6 152
R278 A1.n5 A1.n4 152
R279 A1.n1 A1.n0 113.781
R280 A1.n7 A1.n4 49.6611
R281 A1.n10 A1.n9 39.4369
R282 A1.n10 A1.n2 21.1793
R283 A1.n5 A1 12.8005
R284 A1.n4 A1.n3 10.955
R285 A1 A1.n11 9.82376
R286 A1.n6 A1 8.63306
R287 A1.n6 A1 5.65631
R288 A1.n9 A1.n8 5.11262
R289 A1.n8 A1.n7 5.11262
R290 A1.n11 A1 4.46562
R291 A1.n2 A1.n1 2.19141
R292 A1 A1.n5 1.48887
C0 VPB Y 0.036941f
C1 B1 VPB 0.119142f
C2 A2 Y 0.045793f
C3 VPWR VGND 0.139344f
C4 VPB A1 0.139741f
C5 A2 A1 0.071268f
C6 A3 VPB 0.161801f
C7 Y VGND 0.046889f
C8 A2 A3 0.036999f
C9 B1 VGND 0.026607f
C10 VPWR Y 0.337398f
C11 B1 VPWR 0.046731f
C12 A2 VPB 0.159321f
C13 A1 VGND 0.066192f
C14 VPWR A1 0.082356f
C15 B1 Y 0.320078f
C16 A3 VGND 0.045666f
C17 A3 VPWR 0.025426f
C18 VPB VGND 0.010173f
C19 A1 Y 2.33e-19
C20 VPWR VPB 0.196517f
C21 A2 VGND 0.059873f
C22 A3 Y 0.371966f
C23 A2 VPWR 0.028562f
C24 A3 B1 0.094007f
C25 VGND VNB 0.993108f
C26 Y VNB 0.082519f
C27 VPWR VNB 0.778706f
C28 B1 VNB 0.383144f
C29 A3 VNB 0.457677f
C30 A2 VNB 0.430857f
C31 A1 VNB 0.448174f
C32 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o31ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o31ai_2 VNB VPB VPWR VGND A2 B1 A3 A1 Y
X0 VPWR.t1 B1.t0 Y.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1 VGND.t4 A3.t0 a_27_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.32 pd=1.645 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t3 A1.t0 a_28_368.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 Y.t5 A3.t1 a_297_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t2 A1.t1 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_27_74.t3 A2.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6 a_297_368.t1 A3.t2 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 a_27_74.t2 B1.t1 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=2.09 as=0.1221 ps=1.07 w=0.74 l=0.15
X8 Y.t0 B1.t2 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VGND.t5 A2.t1 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_28_368.t2 A2.t2 a_297_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_297_368.t3 A2.t3 a_28_368.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_27_74.t5 A3.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.32 ps=1.645 w=0.74 l=0.15
X13 a_27_74.t0 A1.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X14 a_28_368.t0 A1.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Y.t2 B1.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B1.n2 B1.t3 226.809
R1 B1.n1 B1.t0 226.809
R2 B1.n1 B1.t2 185.655
R3 B1.n2 B1.n0 184.595
R4 B1.n3 B1.t1 179.947
R5 B1 B1.n4 80.7407
R6 B1.n4 B1.n3 29.6098
R7 B1.n4 B1.n1 20.4067
R8 B1.n0 B1 5.4308
R9 B1 B1.n0 2.13383
R10 B1.n3 B1.n2 1.90313
R11 Y.n2 Y.n1 585
R12 Y.n4 Y.t4 393.301
R13 Y.n4 Y.n3 335.877
R14 Y.n1 Y.n0 290.661
R15 Y.n2 Y.t2 289.37
R16 Y Y.n4 70.3681
R17 Y.n1 Y.t5 35.1791
R18 Y.n3 Y.t1 30.8113
R19 Y.n1 Y.t3 26.3844
R20 Y.n3 Y.t0 22.7032
R21 Y Y.n5 18.0005
R22 Y Y.n2 15.4358
R23 Y.n5 Y 11.6005
R24 Y.n5 Y 10.9181
R25 Y.n0 Y 8.41828
R26 Y.n5 Y.n0 8.285
R27 VPWR.n2 VPWR.n0 341.183
R28 VPWR.n2 VPWR.n1 329.45
R29 VPWR.n1 VPWR.t2 26.3844
R30 VPWR.n1 VPWR.t3 26.3844
R31 VPWR.n0 VPWR.t0 26.3844
R32 VPWR.n0 VPWR.t1 26.3844
R33 VPWR VPWR.n2 0.187828
R34 VPB.t5 VPB.t2 528.63
R35 VPB VPB.t7 260.485
R36 VPB.t4 VPB.t1 255.376
R37 VPB.t1 VPB.t0 229.839
R38 VPB.t2 VPB.t4 229.839
R39 VPB.t6 VPB.t5 229.839
R40 VPB.t3 VPB.t6 229.839
R41 VPB.t7 VPB.t3 229.839
R42 A3.n1 A3.t0 308.772
R43 A3.n0 A3.t1 226.809
R44 A3.n1 A3.t2 226.809
R45 A3.n0 A3.t3 199.666
R46 A3 A3.n2 159.293
R47 A3.n2 A3.n1 56.2338
R48 A3.n2 A3.n0 9.49444
R49 a_27_74.t2 a_27_74.n5 207.849
R50 a_27_74.n1 a_27_74.t4 199.591
R51 a_27_74.n5 a_27_74.n4 185
R52 a_27_74.n1 a_27_74.n0 101.71
R53 a_27_74.n3 a_27_74.n2 92.7788
R54 a_27_74.n5 a_27_74.n3 85.6897
R55 a_27_74.n3 a_27_74.n1 59.3797
R56 a_27_74.n4 a_27_74.t1 22.7032
R57 a_27_74.n4 a_27_74.t5 22.7032
R58 a_27_74.n2 a_27_74.t6 22.7032
R59 a_27_74.n2 a_27_74.t3 22.7032
R60 a_27_74.n0 a_27_74.t7 22.7032
R61 a_27_74.n0 a_27_74.t0 22.7032
R62 VGND.n4 VGND.n3 210.601
R63 VGND.n7 VGND.n6 210.601
R64 VGND.n2 VGND.n1 198.657
R65 VGND.n1 VGND.t3 59.1897
R66 VGND.n1 VGND.t4 58.3789
R67 VGND.n3 VGND.t1 34.0546
R68 VGND.n3 VGND.t5 34.0546
R69 VGND.n6 VGND.t0 34.0546
R70 VGND.n6 VGND.t2 34.0546
R71 VGND.n5 VGND.n4 31.2476
R72 VGND.n7 VGND.n5 19.2005
R73 VGND.n5 VGND.n0 9.3005
R74 VGND.n8 VGND.n7 7.43488
R75 VGND.n4 VGND.n2 6.45226
R76 VGND.n2 VGND.n0 0.368054
R77 VGND VGND.n8 0.160103
R78 VGND.n8 VGND.n0 0.1477
R79 VNB.t6 VNB.t5 2021
R80 VNB.t7 VNB.t3 1316.54
R81 VNB.t4 VNB.t0 1316.54
R82 VNB VNB.t4 1143.31
R83 VNB.t1 VNB.t2 1108.66
R84 VNB.t5 VNB.t1 993.177
R85 VNB.t3 VNB.t6 993.177
R86 VNB.t0 VNB.t7 993.177
R87 A1.n0 A1.t3 226.809
R88 A1.n1 A1.t0 226.809
R89 A1.n1 A1.t1 198.204
R90 A1.n0 A1.t2 180.13
R91 A1.n3 A1.n2 152
R92 A1.n2 A1.n0 54.7732
R93 A1.n3 A1 12.8005
R94 A1.n2 A1.n1 10.955
R95 A1 A1.n3 1.48887
R96 a_28_368.n1 a_28_368.t2 418.31
R97 a_28_368.t1 a_28_368.n1 284.103
R98 a_28_368.n1 a_28_368.n0 205.487
R99 a_28_368.n0 a_28_368.t3 26.3844
R100 a_28_368.n0 a_28_368.t0 26.3844
R101 a_297_368.n1 a_297_368.n0 708.027
R102 a_297_368.n0 a_297_368.t0 26.3844
R103 a_297_368.n0 a_297_368.t3 26.3844
R104 a_297_368.t2 a_297_368.n1 26.3844
R105 a_297_368.n1 a_297_368.t1 26.3844
R106 A2.n0 A2.t0 244.536
R107 A2.n1 A2.t3 222.093
R108 A2.n0 A2.t2 214.758
R109 A2.n1 A2.t1 196.013
R110 A2.n3 A2.n2 152
R111 A2.n2 A2.n1 30.2058
R112 A2.n2 A2.n0 16.7098
R113 A2 A2.n3 10.2703
R114 A2.n3 A2 4.0191
C0 Y A3 0.182281f
C1 VGND A2 0.033245f
C2 B1 VPWR 0.0336f
C3 B1 VPB 0.082116f
C4 Y VGND 0.026491f
C5 Y A2 0.023049f
C6 VPWR A3 0.016837f
C7 VGND A1 0.034972f
C8 VPB A3 0.081314f
C9 A1 A2 0.088492f
C10 VPWR VGND 0.076963f
C11 B1 A3 0.08077f
C12 VGND VPB 0.009108f
C13 VPWR A2 0.017424f
C14 Y A1 5.82e-19
C15 VPB A2 0.073583f
C16 B1 VGND 0.01545f
C17 VPWR Y 0.24103f
C18 VPWR A1 0.03734f
C19 Y VPB 0.02664f
C20 VPB A1 0.069334f
C21 VGND A3 0.026402f
C22 A2 A3 0.041755f
C23 B1 Y 0.195122f
C24 VPWR VPB 0.121558f
C25 VGND VNB 0.56627f
C26 Y VNB 0.071226f
C27 VPWR VNB 0.46789f
C28 B1 VNB 0.283372f
C29 A3 VNB 0.23921f
C30 A2 VNB 0.21543f
C31 A1 VNB 0.256796f
C32 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o31ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o31ai_1 VNB VPB VPWR VGND A3 A2 B1 A1 Y
X0 VPWR.t0 B1.t0 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=1.81 w=1.12 l=0.15
X1 a_203_368.t1 A2.t0 a_119_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X2 Y.t2 A3.t0 a_203_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=1.81 as=0.2352 ps=1.54 w=1.12 l=0.15
X3 a_114_74.t1 A1.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 Y.t0 B1.t1 a_114_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2479 pd=2.15 as=0.111 ps=1.04 w=0.74 l=0.15
X5 a_119_368.t0 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 VGND.t2 A2.t1 a_114_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.3492 pd=1.7 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_114_74.t2 A3.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.3492 ps=1.7 w=0.74 l=0.15
R0 B1.n0 B1.t0 255.639
R1 B1.n0 B1.t1 195.389
R2 B1 B1.n0 156.462
R3 Y.n4 Y.n1 585
R4 Y.n4 Y.n3 585
R5 Y.n2 Y.n1 585
R6 Y.n3 Y.n2 585
R7 Y.n2 Y.t0 279.563
R8 Y Y.n0 278.12
R9 Y.n1 Y.n0 32.4005
R10 Y.n3 Y.n0 32.4005
R11 Y.n3 Y.t1 26.3844
R12 Y.n1 Y.t2 26.3844
R13 Y Y.n4 3.27323
R14 Y.n2 Y 2.98232
R15 Y.n4 Y 2.10959
R16 VPWR.n0 VPWR.t1 266.411
R17 VPWR.n0 VPWR.t0 256.139
R18 VPWR VPWR.n0 0.0973887
R19 VPB.t1 VPB.t0 429.033
R20 VPB.t3 VPB.t1 291.13
R21 VPB VPB.t2 265.591
R22 VPB.t2 VPB.t3 214.517
R23 A2.n0 A2.t0 264.298
R24 A2.n0 A2.t1 204.048
R25 A2 A2.n0 154.56
R26 a_119_368.t0 a_119_368.t1 47.4916
R27 a_203_368.t0 a_203_368.t1 73.8755
R28 A3.n0 A3.t0 288.957
R29 A3.n0 A3.t1 220.113
R30 A3 A3.n0 158.549
R31 A1.n0 A1.t1 279.529
R32 A1.n0 A1.t0 171.344
R33 A1 A1.n0 158.788
R34 VGND.n1 VGND.n0 170.821
R35 VGND.n1 VGND.t0 166.325
R36 VGND.n0 VGND.t1 65.6762
R37 VGND.n0 VGND.t2 65.6762
R38 VGND VGND.n1 0.341406
R39 a_114_74.n1 a_114_74.n0 367.865
R40 a_114_74.t0 a_114_74.n1 25.9464
R41 a_114_74.n0 a_114_74.t3 22.7032
R42 a_114_74.n0 a_114_74.t1 22.7032
R43 a_114_74.n1 a_114_74.t2 22.7032
R44 VNB.t3 VNB.t2 2217.32
R45 VNB VNB.t1 1143.31
R46 VNB.t2 VNB.t0 1039.37
R47 VNB.t1 VNB.t3 993.177
C0 A3 VGND 0.012977f
C1 A3 B1 0.092828f
C2 VPWR Y 0.18686f
C3 A2 VGND 0.017477f
C4 Y VPB 0.008945f
C5 VPWR A1 0.04152f
C6 VPB A1 0.040418f
C7 Y VGND 0.05789f
C8 B1 Y 0.0607f
C9 A1 VGND 0.053624f
C10 VPWR VPB 0.100149f
C11 A3 A2 0.03397f
C12 VPWR VGND 0.05035f
C13 B1 VPWR 0.054417f
C14 A3 Y 0.168304f
C15 VPB VGND 0.006107f
C16 B1 VPB 0.049114f
C17 Y A2 0.13541f
C18 A1 A2 0.100389f
C19 B1 VGND 0.012417f
C20 A3 VPWR 0.007033f
C21 A3 VPB 0.05223f
C22 VPWR A2 0.134832f
C23 Y A1 0.00356f
C24 VPB A2 0.038208f
C25 VGND VNB 0.40206f
C26 Y VNB 0.058332f
C27 VPWR VNB 0.387896f
C28 B1 VNB 0.171593f
C29 A3 VNB 0.13378f
C30 A2 VNB 0.122703f
C31 A1 VNB 0.168846f
C32 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o31a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o31a_4 VNB VPB VPWR VGND A2 A1 A3 B1 X
X0 a_86_260.t3 B1.t0 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2102 ps=1.505 w=1 l=0.15
X1 VPWR.t0 a_86_260.t6 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_492_125.t1 A1.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 X.t7 a_86_260.t7 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.10915 ps=1.035 w=0.74 l=0.15
X4 X.t2 a_86_260.t8 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t2 a_86_260.t9 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t0 A3.t0 a_492_125.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1408 ps=1.08 w=0.64 l=0.15
X7 a_86_260.t5 B1.t1 a_492_125.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1056 pd=0.97 as=0.1952 ps=1.89 w=0.64 l=0.15
X8 a_492_125.t4 B1.t2 a_86_260.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1408 pd=1.08 as=0.1056 ps=0.97 w=0.64 l=0.15
X9 a_968_392.t2 A1.t1 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.17 pd=1.34 as=0.175 ps=1.35 w=1 l=0.15
X10 a_492_125.t3 A3.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X11 VGND.t3 a_86_260.t10 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 X.t0 a_86_260.t11 VPWR.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X13 X.t5 a_86_260.t12 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 a_968_392.t3 A2.t0 a_699_392.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X15 a_699_392.t1 A3.t2 a_86_260.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X16 VPWR.t5 A1.t2 a_968_392.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X17 VGND.t6 A2.t1 a_492_125.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X18 a_86_260.t1 A3.t3 a_699_392.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X19 a_699_392.t2 A2.t2 a_968_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.17 ps=1.34 w=1 l=0.15
X20 VGND.t1 a_86_260.t13 X.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VPWR.t6 B1.t3 a_86_260.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
R0 B1.n0 B1.t0 373.526
R1 B1.n1 B1.t3 207.529
R2 B1.n2 B1.t2 205.215
R3 B1.n0 B1.t1 168.701
R4 B1.n3 B1.n2 152
R5 B1.n2 B1.n1 31.4035
R6 B1.n3 B1 12.2187
R7 B1.n1 B1.n0 2.19141
R8 B1 B1.n3 2.13383
R9 VPWR.n7 VPWR.t6 835.754
R10 VPWR.n6 VPWR.n5 611.84
R11 VPWR.n13 VPWR.n2 325.255
R12 VPWR.n15 VPWR.t3 259.171
R13 VPWR.n4 VPWR.n3 232.787
R14 VPWR.n3 VPWR.t7 46.2955
R15 VPWR.n5 VPWR.t4 39.4005
R16 VPWR.n13 VPWR.n12 30.1181
R17 VPWR.n5 VPWR.t5 29.5505
R18 VPWR.n8 VPWR.n4 28.6123
R19 VPWR.n3 VPWR.t0 27.0196
R20 VPWR.n2 VPWR.t1 26.3844
R21 VPWR.n2 VPWR.t2 26.3844
R22 VPWR.n15 VPWR.n14 25.6005
R23 VPWR.n12 VPWR.n4 24.8476
R24 VPWR.n14 VPWR.n13 23.3417
R25 VPWR.n8 VPWR.n7 20.7064
R26 VPWR.n9 VPWR.n8 9.3005
R27 VPWR.n10 VPWR.n4 9.3005
R28 VPWR.n12 VPWR.n11 9.3005
R29 VPWR.n13 VPWR.n1 9.3005
R30 VPWR.n14 VPWR.n0 9.3005
R31 VPWR.n16 VPWR.n15 9.3005
R32 VPWR.n7 VPWR.n6 7.29369
R33 VPWR.n9 VPWR.n6 0.157378
R34 VPWR.n10 VPWR.n9 0.122949
R35 VPWR.n11 VPWR.n10 0.122949
R36 VPWR.n11 VPWR.n1 0.122949
R37 VPWR.n1 VPWR.n0 0.122949
R38 VPWR.n16 VPWR.n0 0.122949
R39 VPWR VPWR.n16 0.0617245
R40 a_86_260.n14 a_86_260.n13 393.005
R41 a_86_260.n2 a_86_260.t11 265.301
R42 a_86_260.n10 a_86_260.t6 243.119
R43 a_86_260.n7 a_86_260.t8 240.197
R44 a_86_260.n4 a_86_260.t9 240.197
R45 a_86_260.n15 a_86_260.n14 193.002
R46 a_86_260.n2 a_86_260.t12 179.947
R47 a_86_260.n3 a_86_260.t10 179.947
R48 a_86_260.n6 a_86_260.t7 179.947
R49 a_86_260.n9 a_86_260.t13 179.947
R50 a_86_260.n5 a_86_260.n1 165.189
R51 a_86_260.n8 a_86_260.n1 152
R52 a_86_260.n11 a_86_260.n10 152
R53 a_86_260.n12 a_86_260.n0 124.353
R54 a_86_260.n3 a_86_260.n2 82.2509
R55 a_86_260.n9 a_86_260.n8 46.7399
R56 a_86_260.n14 a_86_260.n12 36.1334
R57 a_86_260.n0 a_86_260.t5 35.6255
R58 a_86_260.n6 a_86_260.n5 33.5944
R59 a_86_260.n13 a_86_260.t0 29.5505
R60 a_86_260.n13 a_86_260.t1 29.5505
R61 a_86_260.n15 a_86_260.t2 29.5505
R62 a_86_260.t3 a_86_260.n15 29.5505
R63 a_86_260.n5 a_86_260.n4 29.2126
R64 a_86_260.n12 a_86_260.n11 28.7035
R65 a_86_260.n0 a_86_260.t4 26.2505
R66 a_86_260.n11 a_86_260.n1 13.1884
R67 a_86_260.n8 a_86_260.n7 13.146
R68 a_86_260.n10 a_86_260.n9 2.92171
R69 a_86_260.n7 a_86_260.n6 2.92171
R70 a_86_260.n4 a_86_260.n3 2.19141
R71 VPB.t10 VPB.t7 515.861
R72 VPB.t3 VPB.t11 273.253
R73 VPB VPB.t0 265.591
R74 VPB.t9 VPB.t8 255.376
R75 VPB.t8 VPB.t4 250.269
R76 VPB.t5 VPB.t9 229.839
R77 VPB.t6 VPB.t5 229.839
R78 VPB.t7 VPB.t6 229.839
R79 VPB.t11 VPB.t10 229.839
R80 VPB.t2 VPB.t3 229.839
R81 VPB.t1 VPB.t2 229.839
R82 VPB.t0 VPB.t1 229.839
R83 X.n8 X 591.154
R84 X.n8 X.n0 585
R85 X.n9 X.n8 585
R86 X.n7 X.n1 256.164
R87 X.n3 X.n2 198.827
R88 X.n6 X.n5 185
R89 X.n5 X.n4 185
R90 X.n8 X.t1 26.3844
R91 X.n8 X.t0 26.3844
R92 X.n1 X.t3 26.3844
R93 X.n1 X.t2 26.3844
R94 X.n5 X.t6 22.7032
R95 X.n5 X.t5 22.7032
R96 X.n2 X.t4 22.7032
R97 X.n2 X.t7 22.7032
R98 X X.n9 16.4928
R99 X.n7 X 15.0159
R100 X X.n0 14.2774
R101 X X.n6 12.062
R102 X.n4 X.n3 11.0774
R103 X.n6 X 6.15435
R104 X.n3 X 4.92358
R105 X X.n0 3.93896
R106 X X.n7 3.2005
R107 X.n4 X 2.21588
R108 X.n9 X 1.72358
R109 A1.n3 A1.t1 212.275
R110 A1.n1 A1.t2 211.544
R111 A1.n1 A1.t0 166.071
R112 A1.n2 A1.n0 163.881
R113 A1 A1.n3 162.667
R114 A1.n2 A1.n1 70.8399
R115 A1.n3 A1.n2 1.46111
R116 VGND.n7 VGND.n6 224.68
R117 VGND.n18 VGND.n1 221.518
R118 VGND.n8 VGND.n5 220.573
R119 VGND.n20 VGND.t2 171.77
R120 VGND.n13 VGND.t1 164.077
R121 VGND.n11 VGND.n4 36.1417
R122 VGND.n12 VGND.n11 36.1417
R123 VGND.n17 VGND.n2 36.1417
R124 VGND.n19 VGND.n18 33.8829
R125 VGND.n13 VGND.n12 32.377
R126 VGND.n7 VGND.n4 27.1064
R127 VGND.n5 VGND.t5 26.2505
R128 VGND.n5 VGND.t6 26.2505
R129 VGND.n6 VGND.t7 26.2505
R130 VGND.n6 VGND.t0 26.2505
R131 VGND.n1 VGND.t4 25.1356
R132 VGND.n20 VGND.n19 24.4711
R133 VGND.n1 VGND.t3 22.7032
R134 VGND.n13 VGND.n2 15.0593
R135 VGND.n21 VGND.n20 9.3005
R136 VGND.n9 VGND.n4 9.3005
R137 VGND.n11 VGND.n10 9.3005
R138 VGND.n12 VGND.n3 9.3005
R139 VGND.n14 VGND.n13 9.3005
R140 VGND.n15 VGND.n2 9.3005
R141 VGND.n17 VGND.n16 9.3005
R142 VGND.n19 VGND.n0 9.3005
R143 VGND.n8 VGND.n7 6.83265
R144 VGND.n18 VGND.n17 2.25932
R145 VGND.n9 VGND.n8 0.566085
R146 VGND.n10 VGND.n9 0.122949
R147 VGND.n10 VGND.n3 0.122949
R148 VGND.n14 VGND.n3 0.122949
R149 VGND.n15 VGND.n14 0.122949
R150 VGND.n16 VGND.n15 0.122949
R151 VGND.n16 VGND.n0 0.122949
R152 VGND.n21 VGND.n0 0.122949
R153 VGND VGND.n21 0.0617245
R154 a_492_125.n1 a_492_125.t5 340.637
R155 a_492_125.t1 a_492_125.n3 191.446
R156 a_492_125.n3 a_492_125.n2 100.871
R157 a_492_125.n1 a_492_125.n0 89.2272
R158 a_492_125.n3 a_492_125.n1 55.5811
R159 a_492_125.n0 a_492_125.t0 41.2505
R160 a_492_125.n0 a_492_125.t4 41.2505
R161 a_492_125.n2 a_492_125.t2 26.2505
R162 a_492_125.n2 a_492_125.t3 26.2505
R163 VNB.t1 VNB.t9 2332.81
R164 VNB.t8 VNB.t0 1362.73
R165 VNB VNB.t2 1212.6
R166 VNB.t9 VNB.t8 1108.66
R167 VNB.t3 VNB.t4 1027.82
R168 VNB.t6 VNB.t5 993.177
R169 VNB.t7 VNB.t6 993.177
R170 VNB.t0 VNB.t7 993.177
R171 VNB.t4 VNB.t1 993.177
R172 VNB.t2 VNB.t3 993.177
R173 A3.n2 A3.t3 216.657
R174 A3.n0 A3.t2 211.544
R175 A3.n0 A3.t1 167.743
R176 A3.n3 A3.t0 163.881
R177 A3.n5 A3.n4 152
R178 A3.n2 A3.n1 152
R179 A3.n4 A3.n3 48.2005
R180 A3.n1 A3 14.9338
R181 A3.n4 A3.n0 10.955
R182 A3.n5 A3 9.50353
R183 A3 A3.n5 9.11565
R184 A3.n1 A3 3.68535
R185 A3.n3 A3.n2 1.46111
R186 a_968_392.n1 a_968_392.n0 647.33
R187 a_968_392.n1 a_968_392.t0 37.4305
R188 a_968_392.n0 a_968_392.t1 29.5505
R189 a_968_392.n0 a_968_392.t3 29.5505
R190 a_968_392.t2 a_968_392.n1 29.5505
R191 A2.n0 A2.t1 902.947
R192 A2.t1 A2.t0 457.632
R193 A2.n1 A2.t2 235.644
R194 A2.n1 A2.n0 187.981
R195 A2 A2.n1 156.462
R196 a_699_392.n0 a_699_392.t0 858.131
R197 a_699_392.n0 a_699_392.t2 365.029
R198 a_699_392.n1 a_699_392.n0 204.349
R199 a_699_392.n1 a_699_392.t3 29.5505
R200 a_699_392.t1 a_699_392.n1 29.5505
C0 VPWR B1 0.045861f
C1 X VPB 0.012206f
C2 A1 A3 0.030339f
C3 VGND A2 0.094623f
C4 A1 VPWR 0.02953f
C5 VPB A3 0.086038f
C6 X VGND 0.296895f
C7 VPWR VPB 0.19434f
C8 A1 B1 1.97e-19
C9 VGND A3 0.026867f
C10 X A2 4.86e-20
C11 VPB B1 0.115492f
C12 VPWR VGND 0.119615f
C13 A3 A2 0.069894f
C14 A1 VPB 0.08055f
C15 VGND B1 0.013588f
C16 VPWR A2 0.021279f
C17 VPWR X 0.415298f
C18 A1 VGND 0.02482f
C19 B1 A2 2.46e-19
C20 VGND VPB 0.01313f
C21 A1 A2 0.154526f
C22 VPWR A3 0.0229f
C23 X B1 0.001472f
C24 B1 A3 0.060601f
C25 VPB A2 0.079187f
C26 VGND VNB 0.866044f
C27 X VNB 0.038706f
C28 VPWR VNB 0.668885f
C29 A1 VNB 0.166432f
C30 A2 VNB 0.428229f
C31 A3 VNB 0.186012f
C32 B1 VNB 0.22501f
C33 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o31a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o31a_2 VNB VPB VPWR VGND B1 A3 A2 A1 X
X0 X.t1 a_55_264.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.475 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 X.t3 a_55_264.t4 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X2 VGND.t3 A2.t0 a_328_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.12765 ps=1.085 w=0.74 l=0.15
X3 a_430_392.t1 A2.t1 a_346_392.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X4 a_328_74.t0 A1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12765 pd=1.085 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 VPWR.t1 a_55_264.t5 X.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2634 pd=1.615 as=0.1988 ps=1.475 w=1.12 l=0.15
X6 a_346_392.t0 A1.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2634 ps=1.615 w=1 l=0.15
X7 a_328_74.t3 A3.t0 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.18315 pd=1.235 as=0.1554 ps=1.16 w=0.74 l=0.15
X8 a_55_264.t0 A3.t1 a_430_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.21 ps=1.42 w=1 l=0.15
X9 VPWR.t3 B1.t0 a_55_264.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.445 pd=2.89 as=0.195 ps=1.39 w=1 l=0.15
X10 VGND.t1 a_55_264.t6 X.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_55_264.t1 B1.t1 a_328_74.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.18315 ps=1.235 w=0.74 l=0.15
R0 a_55_264.n3 a_55_264.n2 395.635
R1 a_55_264.n0 a_55_264.t5 303.125
R2 a_55_264.n2 a_55_264.t3 256.63
R3 a_55_264.n3 a_55_264.t1 228.124
R4 a_55_264.n0 a_55_264.t6 206.458
R5 a_55_264.n1 a_55_264.t4 196.278
R6 a_55_264.n4 a_55_264.n3 194.917
R7 a_55_264.n1 a_55_264.n0 89.9738
R8 a_55_264.t0 a_55_264.n4 41.3705
R9 a_55_264.n4 a_55_264.t2 35.4605
R10 a_55_264.n2 a_55_264.n1 11.8854
R11 VPWR.n7 VPWR.t2 860.096
R12 VPWR.n2 VPWR.n1 585
R13 VPWR.n3 VPWR.t3 288.853
R14 VPWR.n1 VPWR.t0 49.2505
R15 VPWR.n1 VPWR.t1 46.4059
R16 VPWR.n6 VPWR.n5 28.5574
R17 VPWR.n7 VPWR.n6 20.7064
R18 VPWR.n3 VPWR.n2 18.5313
R19 VPWR.n5 VPWR.n4 9.3005
R20 VPWR.n6 VPWR.n0 9.3005
R21 VPWR.n8 VPWR.n7 9.3005
R22 VPWR.n5 VPWR.n2 2.20447
R23 VPWR.n4 VPWR.n3 0.161319
R24 VPWR.n4 VPWR.n0 0.122949
R25 VPWR.n8 VPWR.n0 0.122949
R26 VPWR VPWR.n8 0.0617245
R27 X.n2 X.n1 585
R28 X.n2 X.n0 159.095
R29 X.n1 X.t0 31.6612
R30 X.n1 X.t1 30.7817
R31 X.n0 X.t2 22.7032
R32 X.n0 X.t3 22.7032
R33 X X.n2 4.65505
R34 VPB.t2 VPB.t1 329.435
R35 VPB.t5 VPB.t0 291.13
R36 VPB.t0 VPB.t4 275.807
R37 VPB.t3 VPB.t2 257.93
R38 VPB VPB.t3 257.93
R39 VPB.t1 VPB.t5 214.517
R40 VGND.n2 VGND.n1 206.816
R41 VGND.n6 VGND.t2 154.727
R42 VGND.n4 VGND.n3 116.644
R43 VGND.n1 VGND.t4 39.7302
R44 VGND.n3 VGND.t0 34.0546
R45 VGND.n3 VGND.t1 34.0546
R46 VGND.n5 VGND.n4 29.7417
R47 VGND.n1 VGND.t3 28.3789
R48 VGND.n6 VGND.n5 20.7064
R49 VGND.n7 VGND.n6 9.3005
R50 VGND.n5 VGND.n0 9.3005
R51 VGND.n4 VGND.n2 6.44889
R52 VGND.n2 VGND.n0 0.477682
R53 VGND.n7 VGND.n0 0.122949
R54 VGND VGND.n7 0.0617245
R55 VNB.t5 VNB.t1 1489.76
R56 VNB.t4 VNB.t5 1316.54
R57 VNB.t2 VNB.t0 1316.54
R58 VNB VNB.t3 1304.99
R59 VNB.t0 VNB.t4 1143.31
R60 VNB.t3 VNB.t2 993.177
R61 A2.n0 A2.t0 258.673
R62 A2.n0 A2.t1 231.629
R63 A2.n1 A2.n0 152
R64 A2.n1 A2 12.2187
R65 A2 A2.n1 2.13383
R66 a_328_74.n1 a_328_74.n0 358.351
R67 a_328_74.n0 a_328_74.t2 40.541
R68 a_328_74.n0 a_328_74.t3 39.7302
R69 a_328_74.n1 a_328_74.t1 33.2437
R70 a_328_74.t0 a_328_74.n1 22.7032
R71 a_346_392.t0 a_346_392.t1 53.1905
R72 a_430_392.t0 a_430_392.t1 82.7405
R73 A1.n0 A1.t1 263.762
R74 A1.n0 A1.t0 220.113
R75 A1 A1.n0 154.19
R76 A3.n0 A3.t1 298.572
R77 A3.n0 A3.t0 178.34
R78 A3 A3.n0 158.222
R79 B1.n0 B1.t0 274.887
R80 B1 B1.n0 198.089
R81 B1.n0 B1.t1 179.947
C0 A3 VPWR 0.007584f
C1 A1 VGND 0.025288f
C2 VPB A1 0.046189f
C3 X VGND 0.167625f
C4 VPB X 0.003959f
C5 A1 VPWR 0.019115f
C6 A3 B1 0.050935f
C7 VPB VGND 0.009809f
C8 VPWR X 0.017665f
C9 VPWR VGND 0.070061f
C10 A2 A3 0.064593f
C11 VPB VPWR 0.119431f
C12 A1 A2 0.119257f
C13 B1 VGND 0.011215f
C14 VPB B1 0.061006f
C15 A1 A3 0.00389f
C16 A2 X 3.8e-19
C17 B1 VPWR 0.041681f
C18 A3 X 0.002563f
C19 A2 VGND 0.014941f
C20 VPB A2 0.043982f
C21 A3 VGND 0.011271f
C22 VPB A3 0.0397f
C23 A2 VPWR 0.011088f
C24 A1 X 0.034851f
C25 VGND VNB 0.52251f
C26 X VNB 0.018994f
C27 VPWR VNB 0.437997f
C28 B1 VNB 0.184639f
C29 A3 VNB 0.113974f
C30 A2 VNB 0.10431f
C31 A1 VNB 0.110133f
C32 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o32a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32a_1 VNB VPB VPWR VGND B1 A1 A2 A3 B2 X
X0 VPWR.t2 a_83_264.t4 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2757 pd=1.63 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_251_74.t2 A3.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1344 ps=1.06 w=0.64 l=0.15
X2 a_332_368.t0 A2.t0 a_248_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X3 a_83_264.t2 A3.t1 a_332_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_248_368.t1 A1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2757 ps=1.63 w=1 l=0.15
X5 VGND.t3 a_83_264.t5 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1469 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_548_368.t1 B2.t0 a_83_264.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2225 pd=1.445 as=0.195 ps=1.39 w=1 l=0.15
X7 VPWR.t0 B1.t0 a_548_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2225 ps=1.445 w=1 l=0.15
X8 a_251_74.t1 A1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1469 ps=1.16 w=0.64 l=0.15
X9 VGND.t0 A2.t1 a_251_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0896 ps=0.92 w=0.64 l=0.15
X10 a_83_264.t1 B2.t1 a_251_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1424 pd=1.085 as=0.112 ps=0.99 w=0.64 l=0.15
X11 a_251_74.t4 B1.t1 a_83_264.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2144 pd=1.95 as=0.1424 ps=1.085 w=0.64 l=0.15
R0 a_83_264.n2 a_83_264.n0 301.692
R1 a_83_264.n2 a_83_264.n1 293.774
R2 a_83_264.n1 a_83_264.t4 258.942
R3 a_83_264.n1 a_83_264.t5 210.474
R4 a_83_264.n3 a_83_264.n2 201.093
R5 a_83_264.n0 a_83_264.t3 42.188
R6 a_83_264.n0 a_83_264.t1 41.2505
R7 a_83_264.t0 a_83_264.n3 38.4155
R8 a_83_264.n3 a_83_264.t2 38.4155
R9 X.n0 X.t0 291.661
R10 X.t1 X.n0 279.738
R11 X.n1 X.t1 279.738
R12 X.n1 X 8.75839
R13 X.n0 X 3.36892
R14 X X.n1 1.21313
R15 VPWR.n1 VPWR.t0 422.94
R16 VPWR.n1 VPWR.n0 321.719
R17 VPWR.n0 VPWR.t1 61.0705
R18 VPWR.n0 VPWR.t2 35.4615
R19 VPWR VPWR.n1 0.198419
R20 VPB.t4 VPB.t2 337.098
R21 VPB.t0 VPB.t1 303.899
R22 VPB.t5 VPB.t0 275.807
R23 VPB.t3 VPB.t5 275.807
R24 VPB VPB.t4 257.93
R25 VPB.t2 VPB.t3 214.517
R26 A3.n0 A3.t0 236.18
R27 A3.n0 A3.t1 231.629
R28 A3 A3.n0 155.721
R29 VGND.n2 VGND.n1 216.838
R30 VGND.n2 VGND.n0 121.2
R31 VGND.n1 VGND.t2 39.3755
R32 VGND.n1 VGND.t0 39.3755
R33 VGND.n0 VGND.t1 39.3755
R34 VGND.n0 VGND.t3 35.7861
R35 VGND VGND.n2 0.501259
R36 a_251_74.n1 a_251_74.t4 201.054
R37 a_251_74.n2 a_251_74.n1 170.612
R38 a_251_74.n1 a_251_74.n0 89.2272
R39 a_251_74.n0 a_251_74.t3 39.3755
R40 a_251_74.n0 a_251_74.t2 26.2505
R41 a_251_74.t0 a_251_74.n2 26.2505
R42 a_251_74.n2 a_251_74.t1 26.2505
R43 VNB VNB.t4 1408.92
R44 VNB.t3 VNB.t5 1374.28
R45 VNB.t0 VNB.t2 1316.54
R46 VNB.t4 VNB.t1 1316.54
R47 VNB.t2 VNB.t3 1154.86
R48 VNB.t1 VNB.t0 993.177
R49 A2.n0 A2.t1 236.18
R50 A2.n0 A2.t0 231.629
R51 A2 A2.n0 153.935
R52 a_248_368.t0 a_248_368.t1 53.1905
R53 a_332_368.t0 a_332_368.t1 76.8305
R54 A1.n0 A1.t1 236.18
R55 A1.n0 A1.t0 231.629
R56 A1 A1.n0 154.311
R57 B2.n0 B2.t1 236.18
R58 B2.n0 B2.t0 231.629
R59 B2 B2.n0 157.507
R60 a_548_368.t0 a_548_368.t1 87.6655
R61 B1.n0 B1.t0 267.127
R62 B1.n0 B1.t1 171.53
R63 B1.n1 B1.n0 152
R64 B1 B1.n1 9.25588
R65 B1.n1 B1 5.31742
C0 A2 VGND 0.013877f
C1 A1 VPB 0.036139f
C2 B2 X 5.98e-20
C3 A3 VPWR 0.007574f
C4 VPB VGND 0.008793f
C5 A1 VGND 0.025465f
C6 X VPWR 0.100649f
C7 B2 VPB 0.03543f
C8 A3 X 2.37e-19
C9 A2 VPWR 0.010323f
C10 VPB B1 0.048161f
C11 A2 A3 0.086923f
C12 B2 VGND 0.006842f
C13 B1 VGND 0.010897f
C14 VPB VPWR 0.128487f
C15 A1 VPWR 0.013454f
C16 A3 VPB 0.034603f
C17 A2 X 4.58e-19
C18 VPWR VGND 0.062572f
C19 B2 B1 0.048213f
C20 A3 VGND 0.011999f
C21 VPB X 0.01375f
C22 A1 X 0.002178f
C23 A2 VPB 0.032849f
C24 B2 VPWR 0.009f
C25 A1 A2 0.10451f
C26 X VGND 0.109068f
C27 VPWR B1 0.043315f
C28 A3 B2 0.094984f
C29 VGND VNB 0.48596f
C30 B1 VNB 0.198284f
C31 B2 VNB 0.111347f
C32 A3 VNB 0.109659f
C33 A2 VNB 0.108019f
C34 A1 VNB 0.113473f
C35 VPWR VNB 0.430397f
C36 X VNB 0.119531f
C37 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o41ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41ai_2 VNB VPB VPWR VGND A1 Y B1 A4 A3 A2
X0 VGND.t5 A4.t0 a_132_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 a_132_74.t2 A3.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.10545 ps=1.025 w=0.74 l=0.15
X2 VGND.t3 A1.t0 a_132_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 VPWR.t3 B1.t0 Y.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_132_74.t6 B1.t1 Y.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_807_368.t3 A2.t0 a_607_368.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_807_368.t1 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_607_368.t2 A2.t1 a_807_368.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X8 VPWR.t0 A1.t2 a_807_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_132_74.t1 A2.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X10 a_314_368.t3 A3.t1 a_607_368.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t2 B1.t2 a_132_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 VGND.t7 A3.t2 a_132_74.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.12765 ps=1.085 w=0.74 l=0.15
X13 a_607_368.t1 A3.t3 a_314_368.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2436 ps=1.555 w=1.12 l=0.15
X14 Y.t4 B1.t3 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X15 VGND.t0 A2.t3 a_132_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1147 ps=1.05 w=0.74 l=0.15
X16 a_132_74.t4 A4.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.12765 pd=1.085 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 a_132_74.t8 A1.t3 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 a_314_368.t1 A4.t2 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=1.555 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t0 A4.t3 a_314_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
R0 A4.n2 A4.t2 248.017
R1 A4.n0 A4.t3 245.917
R2 A4.n1 A4.t1 213.365
R3 A4.n0 A4.t0 196.013
R4 A4 A4.n2 154.377
R5 A4.n1 A4.n0 58.7169
R6 A4.n2 A4.n1 3.8565
R7 a_132_74.n1 a_132_74.t7 194.131
R8 a_132_74.n5 a_132_74.t8 190.242
R9 a_132_74.n3 a_132_74.n2 104.579
R10 a_132_74.n7 a_132_74.n6 103.317
R11 a_132_74.n5 a_132_74.n4 101.71
R12 a_132_74.n1 a_132_74.n0 88.3339
R13 a_132_74.n3 a_132_74.n1 64.5775
R14 a_132_74.n6 a_132_74.n3 51.2005
R15 a_132_74.n6 a_132_74.n5 50.4476
R16 a_132_74.n0 a_132_74.t6 34.0546
R17 a_132_74.n2 a_132_74.t9 33.2437
R18 a_132_74.t0 a_132_74.n7 25.1356
R19 a_132_74.n7 a_132_74.t2 25.1356
R20 a_132_74.n4 a_132_74.t3 22.7032
R21 a_132_74.n4 a_132_74.t1 22.7032
R22 a_132_74.n0 a_132_74.t5 22.7032
R23 a_132_74.n2 a_132_74.t4 22.7032
R24 VGND.n6 VGND.n3 215.004
R25 VGND.n5 VGND.n4 209.436
R26 VGND.n9 VGND.n2 209.436
R27 VGND.n12 VGND.n11 209.436
R28 VGND.n3 VGND.t3 34.0546
R29 VGND.n4 VGND.t1 34.0546
R30 VGND.n4 VGND.t0 34.0546
R31 VGND.n11 VGND.t5 34.0546
R32 VGND.n5 VGND.n1 27.1064
R33 VGND.n10 VGND.n9 27.1064
R34 VGND.n2 VGND.t7 23.514
R35 VGND.n3 VGND.t6 22.7032
R36 VGND.n2 VGND.t2 22.7032
R37 VGND.n11 VGND.t4 22.7032
R38 VGND.n9 VGND.n1 20.3299
R39 VGND.n12 VGND.n10 18.0711
R40 VGND.n7 VGND.n1 9.3005
R41 VGND.n9 VGND.n8 9.3005
R42 VGND.n10 VGND.n0 9.3005
R43 VGND.n13 VGND.n12 7.40976
R44 VGND.n6 VGND.n5 6.59734
R45 VGND VGND.n13 0.523687
R46 VGND.n7 VGND.n6 0.501235
R47 VGND.n13 VGND.n0 0.153233
R48 VGND.n8 VGND.n7 0.122949
R49 VGND.n8 VGND.n0 0.122949
R50 VNB VNB.t7 2355.91
R51 VNB.t0 VNB.t1 1316.54
R52 VNB.t3 VNB.t8 1154.86
R53 VNB.t5 VNB.t4 1154.86
R54 VNB.t6 VNB.t5 1154.86
R55 VNB.t4 VNB.t9 1143.31
R56 VNB.t2 VNB.t0 1062.47
R57 VNB.t9 VNB.t2 1004.72
R58 VNB.t1 VNB.t3 993.177
R59 VNB.t7 VNB.t6 993.177
R60 A3.n0 A3.t1 229.812
R61 A3.n1 A3.t3 226.809
R62 A3.n1 A3.t2 198.204
R63 A3.n0 A3.t0 196.013
R64 A3 A3.n2 159.591
R65 A3.n2 A3.n1 48.2005
R66 A3.n2 A3.n0 13.146
R67 A1.n1 A1.t0 269.045
R68 A1.n4 A1.t1 226.809
R69 A1.n1 A1.t2 226.809
R70 A1.n5 A1.n4 162.712
R71 A1.n3 A1.n0 152
R72 A1.n2 A1.t3 142.994
R73 A1.n4 A1.n3 22.3965
R74 A1.n3 A1.n2 17.0409
R75 A1.n5 A1.n0 10.1214
R76 A1.n2 A1.n1 4.38232
R77 A1.n0 A1 2.3819
R78 A1 A1.n5 1.78655
R79 B1.n0 B1.t1 285.926
R80 B1.n3 B1.t3 262.363
R81 B1.n1 B1.t0 261.62
R82 B1 B1.n2 155.459
R83 B1.n0 B1.t2 151.053
R84 B1.n4 B1.n3 58.7236
R85 B1.n2 B1.n1 30.6732
R86 B1.n3 B1.n2 25.1486
R87 B1 B1.n4 11.9356
R88 B1.n1 B1.n0 11.8887
R89 B1.n4 B1 4.67077
R90 Y Y.n1 327.979
R91 Y Y.n3 246.738
R92 Y.n2 Y.n0 213.703
R93 Y.n3 Y.t5 26.3844
R94 Y.n3 Y.t4 26.3844
R95 Y.n1 Y.t1 26.3844
R96 Y.n1 Y.t0 26.3844
R97 Y.n0 Y.t3 22.7032
R98 Y.n0 Y.t2 22.7032
R99 Y.n2 Y 13.5534
R100 Y Y.n2 4.51815
R101 VPWR.n3 VPWR.t3 418.663
R102 VPWR.n2 VPWR.n1 339.101
R103 VPWR.n5 VPWR.t2 250.081
R104 VPWR.n1 VPWR.t1 26.3844
R105 VPWR.n1 VPWR.t0 26.3844
R106 VPWR.n4 VPWR.n3 21.4593
R107 VPWR.n5 VPWR.n4 21.4593
R108 VPWR.n4 VPWR.n0 9.3005
R109 VPWR.n6 VPWR.n5 9.3005
R110 VPWR.n3 VPWR.n2 7.26096
R111 VPWR.n2 VPWR.n0 0.155613
R112 VPWR.n6 VPWR.n0 0.122949
R113 VPWR VPWR.n6 0.0617245
R114 VPB.t8 VPB.t9 503.091
R115 VPB.t6 VPB.t3 500.538
R116 VPB.t4 VPB.t7 298.791
R117 VPB VPB.t5 252.823
R118 VPB.t0 VPB.t1 229.839
R119 VPB.t2 VPB.t0 229.839
R120 VPB.t9 VPB.t2 229.839
R121 VPB.t7 VPB.t8 229.839
R122 VPB.t3 VPB.t4 229.839
R123 VPB.t5 VPB.t6 229.839
R124 A2.n0 A2.t0 331.241
R125 A2.n2 A2.t3 227.585
R126 A2.n1 A2.t1 214.758
R127 A2.n0 A2.t2 196.013
R128 A2 A2.n2 96.1448
R129 A2.n2 A2.n1 34.4739
R130 A2.n1 A2.n0 1.9285
R131 a_607_368.n1 a_607_368.n0 713.544
R132 a_607_368.n0 a_607_368.t3 26.3844
R133 a_607_368.n0 a_607_368.t2 26.3844
R134 a_607_368.t0 a_607_368.n1 26.3844
R135 a_607_368.n1 a_607_368.t1 26.3844
R136 a_807_368.n1 a_807_368.t2 434.082
R137 a_807_368.t1 a_807_368.n1 274.788
R138 a_807_368.n1 a_807_368.n0 205.487
R139 a_807_368.n0 a_807_368.t0 26.3844
R140 a_807_368.n0 a_807_368.t3 26.3844
R141 a_314_368.n0 a_314_368.t0 468.45
R142 a_314_368.n0 a_314_368.t3 448.839
R143 a_314_368.n1 a_314_368.n0 189.115
R144 a_314_368.n1 a_314_368.t2 50.13
R145 a_314_368.t1 a_314_368.n1 26.3844
C0 B1 Y 0.136794f
C1 VPB VGND 0.01009f
C2 VPB A3 0.066452f
C3 A2 VPWR 0.018999f
C4 B1 VPWR 0.083342f
C5 Y VGND 0.013671f
C6 A3 Y 8.57e-19
C7 VPB Y 0.018745f
C8 VPWR VGND 0.099106f
C9 A2 A1 0.106784f
C10 A3 VPWR 0.015839f
C11 VPB VPWR 0.168445f
C12 B1 A4 0.029836f
C13 VPWR Y 0.23197f
C14 A1 VGND 0.045203f
C15 A4 VGND 0.033915f
C16 VPB A1 0.081133f
C17 A4 A3 0.086087f
C18 VPB A4 0.075637f
C19 A1 Y 2.56e-19
C20 A2 VGND 0.035648f
C21 B1 VGND 0.070201f
C22 A4 Y 0.070697f
C23 A3 A2 0.066772f
C24 VPB A2 0.097692f
C25 A1 VPWR 0.033237f
C26 VPB B1 0.092926f
C27 A4 VPWR 0.013042f
C28 A2 Y 1.83e-19
C29 A3 VGND 0.034957f
C30 VGND VNB 0.728952f
C31 Y VNB 0.032686f
C32 VPWR VNB 0.626143f
C33 A1 VNB 0.30881f
C34 A2 VNB 0.240444f
C35 A3 VNB 0.188365f
C36 A4 VNB 0.217715f
C37 B1 VNB 0.502672f
C38 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o41ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41ai_1 VNB VPB VPWR VGND A3 A2 B1 Y A4 A1
X0 a_157_74.t3 A1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X1 a_260_368.t1 A4.t0 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.196 ps=1.47 w=1.12 l=0.15
X2 VGND.t3 A4.t1 a_157_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.16095 pd=1.175 as=0.14615 ps=1.135 w=0.74 l=0.15
X3 a_157_74.t2 B1.t0 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.14615 pd=1.135 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 Y.t2 B1.t1 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.5768 ps=3.27 w=1.12 l=0.15
X5 a_358_368.t0 A3.t0 a_260_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1904 ps=1.46 w=1.12 l=0.15
X6 a_157_74.t0 A3.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.16095 ps=1.175 w=0.74 l=0.15
X7 a_472_368.t1 A2.t0 a_358_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X8 VGND.t1 A2.t1 a_157_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t1 A1.t1 a_472_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
R0 A1.n0 A1.t1 248.017
R1 A1.n0 A1.t0 217.221
R2 A1 A1.n0 153.958
R3 VGND.n2 VGND.n1 213.785
R4 VGND.n2 VGND.n0 213.316
R5 VGND.n0 VGND.t0 36.487
R6 VGND.n1 VGND.t2 34.0546
R7 VGND.n1 VGND.t1 34.0546
R8 VGND.n0 VGND.t3 34.0546
R9 VGND VGND.n2 0.687027
R10 a_157_74.n1 a_157_74.t3 199.591
R11 a_157_74.n1 a_157_74.n0 156.155
R12 a_157_74.n2 a_157_74.n1 101.71
R13 a_157_74.n0 a_157_74.t2 41.3519
R14 a_157_74.n0 a_157_74.t4 22.7032
R15 a_157_74.n2 a_157_74.t1 22.7032
R16 a_157_74.t0 a_157_74.n2 22.7032
R17 VNB VNB.t2 1639.9
R18 VNB.t4 VNB.t0 1351.18
R19 VNB.t1 VNB.t3 1316.54
R20 VNB.t2 VNB.t4 1258.79
R21 VNB.t0 VNB.t1 993.177
R22 A4.n0 A4.t0 250.909
R23 A4.n0 A4.t1 220.113
R24 A4 A4.n0 155.126
R25 Y.n1 Y.n0 289.245
R26 Y.n1 Y.t1 113.465
R27 Y.n0 Y.t2 35.1791
R28 Y.n0 Y.t0 26.3844
R29 Y Y.n1 4.36513
R30 a_260_368.t0 a_260_368.t1 59.8041
R31 VPB VPB.t3 370.296
R32 VPB.t2 VPB.t4 291.13
R33 VPB.t0 VPB.t2 291.13
R34 VPB.t3 VPB.t1 255.376
R35 VPB.t1 VPB.t0 250.269
R36 B1.n0 B1.t1 263.81
R37 B1 B1.n0 223.055
R38 B1.n0 B1.t0 154.24
R39 VPWR.n0 VPWR.t1 265.368
R40 VPWR.n0 VPWR.t0 248.638
R41 VPWR VPWR.n0 0.128232
R42 A3.n0 A3.t0 250.909
R43 A3.n0 A3.t1 220.113
R44 A3.n1 A3.n0 156.268
R45 A3.n1 A3 15.0266
R46 A3 A3.n1 5.56572
R47 A3.n1 A3 3.29747
R48 a_358_368.t0 a_358_368.t1 73.8755
R49 A2.n0 A2.t0 250.909
R50 A2.n0 A2.t1 220.113
R51 A2 A2.n0 176.887
R52 a_472_368.t0 a_472_368.t1 73.8755
C0 VGND A3 0.016515f
C1 Y A2 3.32e-19
C2 VPWR VPB 0.111718f
C3 VPB B1 0.050619f
C4 A1 VPWR 0.045391f
C5 Y VGND 0.072461f
C6 VGND A4 0.013343f
C7 Y A3 0.051063f
C8 VPWR A2 0.065191f
C9 A1 VPB 0.040953f
C10 A4 A3 0.091638f
C11 VPB A2 0.039248f
C12 VPWR VGND 0.056251f
C13 A1 A2 0.077155f
C14 VPWR A3 0.02743f
C15 Y A4 0.059083f
C16 VGND B1 0.007175f
C17 VGND VPB 0.00727f
C18 VPB A3 0.036283f
C19 A1 VGND 0.016488f
C20 VPWR Y 0.136813f
C21 Y B1 0.108828f
C22 VPWR A4 0.011272f
C23 B1 A4 0.051234f
C24 VGND A2 0.016633f
C25 Y VPB 0.007478f
C26 A3 A2 0.158932f
C27 VPB A4 0.033158f
C28 A1 Y 1.74e-19
C29 VPWR B1 0.046014f
C30 VGND VNB 0.432343f
C31 Y VNB 0.062248f
C32 VPWR VNB 0.438554f
C33 A1 VNB 0.158529f
C34 A2 VNB 0.109169f
C35 A3 VNB 0.104634f
C36 A4 VNB 0.105677f
C37 B1 VNB 0.191312f
C38 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o41a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41a_4 VNB VPB VPWR VGND B1 X A1 A2 A3 A4
X0 a_523_124.t2 A3.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 VGND.t7 A4.t0 a_523_124.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 VGND.t11 A1.t0 a_523_124.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.113125 pd=1.005 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 a_1213_368# A1.t1 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1904 ps=1.46 w=1.12 l=0.15
X4 VPWR.t2 a_110_48.t6 X.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.20015 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_851_368.t1 A4.t1 a_110_48.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X6 VGND.t10 a_110_48.t7 X.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 X.t6 a_110_48.t8 VPWR.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VGND.t1 A3.t1 a_523_124.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.19135 pd=1.26 as=0.1184 ps=1.01 w=0.64 l=0.15
X9 VPWR.t4 a_110_48.t9 X.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 X.t4 a_110_48.t10 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X11 X.t2 a_110_48.t11 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X12 VGND.t0 A2.t0 a_523_124.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0928 ps=0.93 w=0.64 l=0.15
X13 X.t1 a_110_48.t12 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X14 a_110_48.t3 B1.t0 a_523_124.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X15 a_523_124.t5 A4.t2 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.19135 ps=1.26 w=0.64 l=0.15
X16 a_110_48.t0 A4.t3 a_851_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X17 VPWR A1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VGND.t5 a_110_48.t13 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_523_124.t3 A2.t1 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.113125 ps=1.005 w=0.64 l=0.15
X20 VPWR.t0 B1.t1 a_110_48.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X21 a_851_368.t2 A3.t2 a_762_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X22 a_523_124.t6 A1.t2 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X23 a_110_48.t5 B1.t2 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.20015 ps=1.505 w=0.84 l=0.15
X24 a_1213_368# A2.t2 a_762_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 a_762_368.t1 A2.t3 a_1213_368# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X26 a_523_124.t8 B1.t3 a_110_48.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.01 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 A3.n1 A3.t0 661.178
R1 A3.t1 A3.t2 479.055
R2 A3.t0 A3.n0 451.474
R3 A3.n1 A3.t1 160.577
R4 A3 A3.n1 156.849
R5 VGND.n33 VGND.t4 240.582
R6 VGND.n20 VGND.n6 235.242
R7 VGND.n11 VGND.n10 227.853
R8 VGND.n13 VGND.n12 223.144
R9 VGND.n8 VGND.n7 213.898
R10 VGND.n31 VGND.n2 206.528
R11 VGND.n27 VGND.t10 160.755
R12 VGND.n6 VGND.t1 85.3772
R13 VGND.n10 VGND.t6 36.9402
R14 VGND.n15 VGND.n14 36.1417
R15 VGND.n19 VGND.n18 36.1417
R16 VGND.n21 VGND.n4 36.1417
R17 VGND.n25 VGND.n4 36.1417
R18 VGND.n26 VGND.n25 36.1417
R19 VGND.n2 VGND.t3 34.0546
R20 VGND.n32 VGND.n31 28.9887
R21 VGND.n21 VGND.n20 28.6123
R22 VGND.n27 VGND.n1 26.7299
R23 VGND.n12 VGND.t9 26.2505
R24 VGND.n12 VGND.t0 26.2505
R25 VGND.n7 VGND.t2 26.2505
R26 VGND.n7 VGND.t7 26.2505
R27 VGND.n10 VGND.t11 23.5002
R28 VGND.n2 VGND.t5 22.7032
R29 VGND.n6 VGND.t8 22.1719
R30 VGND.n13 VGND.n11 21.4625
R31 VGND.n27 VGND.n26 20.7064
R32 VGND.n31 VGND.n1 18.4476
R33 VGND.n33 VGND.n32 16.1887
R34 VGND.n34 VGND.n33 9.3005
R35 VGND.n32 VGND.n0 9.3005
R36 VGND.n31 VGND.n30 9.3005
R37 VGND.n29 VGND.n1 9.3005
R38 VGND.n28 VGND.n27 9.3005
R39 VGND.n14 VGND.n9 9.3005
R40 VGND.n16 VGND.n15 9.3005
R41 VGND.n18 VGND.n17 9.3005
R42 VGND.n19 VGND.n5 9.3005
R43 VGND.n22 VGND.n21 9.3005
R44 VGND.n23 VGND.n4 9.3005
R45 VGND.n25 VGND.n24 9.3005
R46 VGND.n26 VGND.n3 9.3005
R47 VGND.n18 VGND.n8 8.65932
R48 VGND.n20 VGND.n19 7.52991
R49 VGND.n15 VGND.n8 2.63579
R50 VGND.n14 VGND.n13 1.88285
R51 VGND.n11 VGND.n9 1.55938
R52 VGND.n16 VGND.n9 0.122949
R53 VGND.n17 VGND.n16 0.122949
R54 VGND.n17 VGND.n5 0.122949
R55 VGND.n22 VGND.n5 0.122949
R56 VGND.n23 VGND.n22 0.122949
R57 VGND.n24 VGND.n23 0.122949
R58 VGND.n24 VGND.n3 0.122949
R59 VGND.n28 VGND.n3 0.122949
R60 VGND.n29 VGND.n28 0.122949
R61 VGND.n30 VGND.n29 0.122949
R62 VGND.n30 VGND.n0 0.122949
R63 VGND.n34 VGND.n0 0.122949
R64 VGND VGND.n34 0.0617245
R65 a_523_124.n3 a_523_124.t7 344.699
R66 a_523_124.n1 a_523_124.t3 272.178
R67 a_523_124.n7 a_523_124.n6 103.587
R68 a_523_124.n5 a_523_124.n4 100.812
R69 a_523_124.n1 a_523_124.n0 100.754
R70 a_523_124.n5 a_523_124.n3 88.4419
R71 a_523_124.n3 a_523_124.n2 88.3446
R72 a_523_124.n6 a_523_124.n5 52.309
R73 a_523_124.n6 a_523_124.n1 45.9299
R74 a_523_124.n2 a_523_124.t1 43.1255
R75 a_523_124.n7 a_523_124.t0 27.188
R76 a_523_124.t2 a_523_124.n7 27.188
R77 a_523_124.n2 a_523_124.t8 26.2505
R78 a_523_124.n4 a_523_124.t4 26.2505
R79 a_523_124.n4 a_523_124.t5 26.2505
R80 a_523_124.n0 a_523_124.t9 26.2505
R81 a_523_124.n0 a_523_124.t6 26.2505
R82 VNB.t11 VNB.t10 2286.61
R83 VNB.t1 VNB.t8 1732.28
R84 VNB VNB.t4 1443.57
R85 VNB.t12 VNB.t1 1201.05
R86 VNB.t13 VNB.t6 1154.86
R87 VNB.t5 VNB.t3 1154.86
R88 VNB.t2 VNB.t0 1016.27
R89 VNB.t9 VNB.t13 993.177
R90 VNB.t0 VNB.t9 993.177
R91 VNB.t7 VNB.t2 993.177
R92 VNB.t8 VNB.t7 993.177
R93 VNB.t10 VNB.t12 993.177
R94 VNB.t3 VNB.t11 993.177
R95 VNB.t4 VNB.t5 993.177
R96 A4.n2 A4.t3 233.381
R97 A4.n0 A4.t1 226.809
R98 A4 A4.n1 154.163
R99 A4.n3 A4.n2 152
R100 A4.n0 A4.t0 140.364
R101 A4.n2 A4.t2 138.173
R102 A4.n2 A4.n1 49.6611
R103 A4.n1 A4.n0 10.955
R104 A4 A4.n3 10.0963
R105 A4.n3 A4 7.21177
R106 A1.n0 A1.t1 240.361
R107 A1.n2 A1.n1 226.809
R108 A1.n4 A1.n3 152
R109 A1.n2 A1.t2 143.286
R110 A1.n0 A1.t0 138.173
R111 A1.n3 A1.n0 49.6611
R112 A1 A1.n4 13.5116
R113 A1.n3 A1.n2 8.03383
R114 A1.n4 A1 3.55606
R115 VPWR.n7 VPWR.t1 856.317
R116 VPWR.n6 VPWR.t0 752.33
R117 VPWR.n18 VPWR.t5 361.084
R118 VPWR.n11 VPWR.n4 335.473
R119 VPWR.n2 VPWR.n1 334.702
R120 VPWR.n4 VPWR.t6 55.1136
R121 VPWR.n19 VPWR.n18 37.1593
R122 VPWR.n13 VPWR.n12 36.1417
R123 VPWR.n17 VPWR.n16 36.1417
R124 VPWR.n10 VPWR.n5 36.1417
R125 VPWR.n4 VPWR.t2 29.3574
R126 VPWR.n1 VPWR.t3 26.3844
R127 VPWR.n1 VPWR.t4 26.3844
R128 VPWR.n16 VPWR.n2 23.3417
R129 VPWR.n6 VPWR.n5 14.3064
R130 VPWR.n13 VPWR.n2 12.8005
R131 VPWR.n12 VPWR.n11 12.424
R132 VPWR.n7 VPWR.n6 10.6621
R133 VPWR.n8 VPWR.n5 9.3005
R134 VPWR.n10 VPWR.n9 9.3005
R135 VPWR.n12 VPWR.n3 9.3005
R136 VPWR.n14 VPWR.n13 9.3005
R137 VPWR.n16 VPWR.n15 9.3005
R138 VPWR.n17 VPWR.n0 9.3005
R139 VPWR.n18 VPWR.n17 8.28285
R140 VPWR.n11 VPWR.n10 4.89462
R141 VPWR.n8 VPWR.n7 0.149596
R142 VPWR.n9 VPWR.n8 0.122949
R143 VPWR.n9 VPWR.n3 0.122949
R144 VPWR.n14 VPWR.n3 0.122949
R145 VPWR.n15 VPWR.n14 0.122949
R146 VPWR.n15 VPWR.n0 0.122949
R147 VPWR.n19 VPWR.n0 0.122949
R148 VPWR VPWR.n19 0.0617245
R149 VPB.t3 VPB.t2 515.861
R150 VPB.t4 VPB.t6 480.108
R151 VPB.t1 VPB.t4 459.678
R152 VPB VPB.t10 426.478
R153 VPB.t7 VPB.t11 273.253
R154 VPB.t6 VPB.t5 255.376
R155 VPB.t0 VPB.t1 234.946
R156 VPB.t2 VPB.t0 229.839
R157 VPB.t11 VPB.t3 229.839
R158 VPB.t8 VPB.t7 229.839
R159 VPB.t9 VPB.t8 229.839
R160 VPB.t10 VPB.t9 229.839
R161 a_110_48.n19 a_110_48.n18 716.765
R162 a_110_48.n18 a_110_48.n0 299.291
R163 a_110_48.n15 a_110_48.t6 259.185
R164 a_110_48.n12 a_110_48.t8 248.231
R165 a_110_48.n3 a_110_48.t9 248.231
R166 a_110_48.n5 a_110_48.t10 248.231
R167 a_110_48.n4 a_110_48.t12 188.565
R168 a_110_48.n6 a_110_48.t13 170.308
R169 a_110_48.n11 a_110_48.t11 170.308
R170 a_110_48.n14 a_110_48.t7 170.308
R171 a_110_48.n8 a_110_48.n4 165.189
R172 a_110_48.n8 a_110_48.n7 152
R173 a_110_48.n10 a_110_48.n9 152
R174 a_110_48.n13 a_110_48.n2 152
R175 a_110_48.n16 a_110_48.n15 152
R176 a_110_48.n17 a_110_48.n1 107.853
R177 a_110_48.n0 a_110_48.t2 35.1791
R178 a_110_48.n0 a_110_48.t5 35.1791
R179 a_110_48.n17 a_110_48.n16 32.3884
R180 a_110_48.n6 a_110_48.n5 32.1338
R181 a_110_48.n14 a_110_48.n13 31.4035
R182 a_110_48.n7 a_110_48.n3 28.4823
R183 a_110_48.n19 a_110_48.t1 27.2639
R184 a_110_48.t0 a_110_48.n19 27.2639
R185 a_110_48.n12 a_110_48.n11 26.2914
R186 a_110_48.n1 a_110_48.t4 26.2505
R187 a_110_48.n1 a_110_48.t3 26.2505
R188 a_110_48.n10 a_110_48.n3 21.1793
R189 a_110_48.n15 a_110_48.n14 18.2581
R190 a_110_48.n11 a_110_48.n10 18.2581
R191 a_110_48.n18 a_110_48.n17 16.8732
R192 a_110_48.n16 a_110_48.n2 13.1884
R193 a_110_48.n9 a_110_48.n2 13.1884
R194 a_110_48.n9 a_110_48.n8 13.1884
R195 a_110_48.n5 a_110_48.n4 12.4157
R196 a_110_48.n13 a_110_48.n12 5.11262
R197 a_110_48.n7 a_110_48.n6 5.11262
R198 X.n2 X.n0 251.68
R199 X.n2 X.n1 208.763
R200 X.n5 X.n3 152.879
R201 X.n5 X.n4 101.678
R202 X.n6 X.n5 90.1898
R203 X.n6 X.n2 40.6593
R204 X.n0 X.t7 26.3844
R205 X.n0 X.t6 26.3844
R206 X.n1 X.t5 26.3844
R207 X.n1 X.t4 26.3844
R208 X.n3 X.t3 22.7032
R209 X.n3 X.t2 22.7032
R210 X.n4 X.t0 22.7032
R211 X.n4 X.t1 22.7032
R212 X X.n6 5.28746
R213 a_851_368.t1 a_851_368.n0 1469.23
R214 a_851_368.n0 a_851_368.t0 26.3844
R215 a_851_368.n0 a_851_368.t2 26.3844
R216 A2.n0 A2.t0 644.917
R217 A2.t0 A2.t2 451.474
R218 A2.t1 A2.t3 435.099
R219 A2 A2.n0 176.031
R220 A2.n0 A2.t1 159.381
R221 B1.n0 B1.t2 303.125
R222 B1.n1 B1.t1 181.821
R223 B1.n0 B1.t0 160.667
R224 B1.n2 B1.t3 160.667
R225 B1 B1.n2 160.478
R226 B1.n1 B1.n0 46.886
R227 B1.n2 B1.n1 34.3247
R228 a_762_368.t0 a_762_368.n0 461.668
R229 a_762_368.n0 a_762_368.t1 380.303
R230 a_762_368.n0 a_762_368.t2 221.444
C0 a_1213_368# VPB 0.004821f
C1 A3 A4 0.127718f
C2 X VGND 0.313739f
C3 A3 A2 0.068849f
C4 VPB X 0.038372f
C5 B1 VGND 0.013429f
C6 A3 VPWR 0.015108f
C7 A4 A2 0.001192f
C8 A3 A1 0.001258f
C9 VPB B1 0.109984f
C10 A4 VPWR 0.01087f
C11 A4 A1 0.007042f
C12 VPB VGND 0.015708f
C13 A2 VPWR 0.01508f
C14 A2 A1 0.125398f
C15 A3 X 8.02e-20
C16 A2 a_1213_368# 0.015104f
C17 A1 VPWR 0.023969f
C18 A3 B1 0.042754f
C19 a_1213_368# VPWR 0.169483f
C20 A1 a_1213_368# 0.028392f
C21 A3 VGND 0.155241f
C22 A4 B1 0.02226f
C23 A3 VPB 0.062438f
C24 VPWR X 0.504985f
C25 A4 VGND 0.01963f
C26 A4 VPB 0.063649f
C27 VPWR B1 0.03058f
C28 A1 B1 1.49e-21
C29 A2 VGND 0.177406f
C30 a_1213_368# B1 6.3e-20
C31 A2 VPB 0.060653f
C32 VPWR VGND 0.132481f
C33 A1 VGND 0.020959f
C34 VPB VPWR 0.235828f
C35 a_1213_368# VGND 0.003122f
C36 A1 VPB 0.067931f
C37 X B1 0.002403f
C38 VGND VNB 0.981787f
C39 B1 VNB 0.218958f
C40 X VNB 0.104277f
C41 VPWR VNB 0.77651f
C42 A1 VNB 0.175516f
C43 A2 VNB 0.440022f
C44 A4 VNB 0.164831f
C45 A3 VNB 0.402413f
C46 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o41a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41a_2 VNB VPB VPWR VGND A1 A2 A3 A4 B1 X
X0 X.t3 a_428_368.t3 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.5459 ps=2.18 w=1.12 l=0.15
X1 a_116_368.t1 A1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VGND.t5 a_428_368.t4 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_27_74.t4 A4.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.21645 ps=1.325 w=0.74 l=0.15
X4 VPWR.t1 B1.t0 a_428_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.5459 pd=2.18 as=0.2277 ps=1.54 w=1 l=0.15
X5 VGND.t1 A1.t1 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 X.t0 a_428_368.t5 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X7 VGND.t3 A3.t0 a_27_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.21645 pd=1.325 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_200_368.t1 A2.t0 a_116_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X9 a_314_368.t0 A3.t1 a_200_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X10 a_27_74.t2 A2.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X11 a_428_368.t0 B1.t1 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.10915 ps=1.035 w=0.74 l=0.15
X12 a_428_368.t1 A4.t1 a_314_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X13 VPWR.t2 a_428_368.t6 X.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 a_428_368.n0 a_428_368.n4 299.125
R1 a_428_368.n1 a_428_368.t6 248.596
R2 a_428_368.n2 a_428_368.t3 240.197
R3 a_428_368.n4 a_428_368.n3 186.325
R4 a_428_368.n4 a_428_368.t0 182.713
R5 a_428_368.n3 a_428_368.t5 179.947
R6 a_428_368.n1 a_428_368.t4 179.947
R7 a_428_368.n2 a_428_368.n1 56.9641
R8 a_428_368.n0 a_428_368.t2 53.1905
R9 a_428_368.n5 a_428_368.n0 40.0683
R10 a_428_368.n0 a_428_368.t1 27.0196
R11 a_428_368.n3 a_428_368.n2 5.84292
R12 VPWR.n13 VPWR.n12 292.5
R13 VPWR.n11 VPWR.n10 292.5
R14 VPWR.n5 VPWR.n4 292.5
R15 VPWR.n6 VPWR.t2 255.03
R16 VPWR.n21 VPWR.t0 248.744
R17 VPWR.n11 VPWR.n4 78.8005
R18 VPWR.n12 VPWR.n11 69.9355
R19 VPWR.n15 VPWR.n14 36.1417
R20 VPWR.n15 VPWR.n1 36.1417
R21 VPWR.n19 VPWR.n1 36.1417
R22 VPWR.n20 VPWR.n19 36.1417
R23 VPWR.n12 VPWR.t1 29.5505
R24 VPWR.n6 VPWR.n5 29.3505
R25 VPWR.n4 VPWR.t3 28.5357
R26 VPWR.n21 VPWR.n20 20.7064
R27 VPWR.n9 VPWR.n8 9.3005
R28 VPWR.n7 VPWR.n3 9.3005
R29 VPWR.n14 VPWR.n2 9.3005
R30 VPWR.n16 VPWR.n15 9.3005
R31 VPWR.n17 VPWR.n1 9.3005
R32 VPWR.n19 VPWR.n18 9.3005
R33 VPWR.n20 VPWR.n0 9.3005
R34 VPWR.n22 VPWR.n21 9.3005
R35 VPWR.n14 VPWR.n13 6.01901
R36 VPWR.n10 VPWR.n9 4.38094
R37 VPWR.n13 VPWR.n3 2.95872
R38 VPWR.n8 VPWR.n6 2.34593
R39 VPWR.n10 VPWR.n3 1.08139
R40 VPWR.n9 VPWR.n5 0.171167
R41 VPWR.n8 VPWR.n7 0.122949
R42 VPWR.n7 VPWR.n2 0.122949
R43 VPWR.n16 VPWR.n2 0.122949
R44 VPWR.n17 VPWR.n16 0.122949
R45 VPWR.n18 VPWR.n17 0.122949
R46 VPWR.n18 VPWR.n0 0.122949
R47 VPWR.n22 VPWR.n0 0.122949
R48 VPWR VPWR.n22 0.0617245
R49 X X.n0 255.624
R50 X X.n1 107.427
R51 X.n0 X.t2 26.3844
R52 X.n0 X.t3 26.3844
R53 X.n1 X.t1 22.7032
R54 X.n1 X.t0 22.7032
R55 VPB.t3 VPB.t6 618.011
R56 VPB.t2 VPB.t3 291.13
R57 VPB.t4 VPB.t2 291.13
R58 VPB.t0 VPB.t4 291.13
R59 VPB VPB.t1 257.93
R60 VPB.t6 VPB.t5 229.839
R61 VPB.t1 VPB.t0 214.517
R62 A1.n0 A1.t0 250.909
R63 A1.n0 A1.t1 220.113
R64 A1 A1.n0 160.186
R65 a_116_368.t0 a_116_368.t1 47.4916
R66 VGND.n5 VGND.t4 233.109
R67 VGND.n14 VGND.n13 208.079
R68 VGND.n11 VGND.n2 200.435
R69 VGND.n4 VGND.t5 150.393
R70 VGND.n2 VGND.t3 48.6491
R71 VGND.n2 VGND.t0 46.2167
R72 VGND.n7 VGND.n6 36.1417
R73 VGND.n7 VGND.n1 36.1417
R74 VGND.n13 VGND.t2 34.0546
R75 VGND.n13 VGND.t1 34.0546
R76 VGND.n12 VGND.n11 31.2476
R77 VGND.n14 VGND.n12 19.2005
R78 VGND.n6 VGND.n5 17.6946
R79 VGND.n12 VGND.n0 9.3005
R80 VGND.n11 VGND.n10 9.3005
R81 VGND.n9 VGND.n1 9.3005
R82 VGND.n8 VGND.n7 9.3005
R83 VGND.n6 VGND.n3 9.3005
R84 VGND.n15 VGND.n14 7.43488
R85 VGND.n5 VGND.n4 6.96039
R86 VGND.n11 VGND.n1 2.63579
R87 VGND.n4 VGND.n3 0.594857
R88 VGND VGND.n15 0.160103
R89 VGND.n15 VGND.n0 0.1477
R90 VGND.n8 VGND.n3 0.122949
R91 VGND.n9 VGND.n8 0.122949
R92 VGND.n10 VGND.n9 0.122949
R93 VGND.n10 VGND.n0 0.122949
R94 VNB.t0 VNB.t5 2609.97
R95 VNB.t4 VNB.t1 1697.64
R96 VNB.t2 VNB.t3 1316.54
R97 VNB VNB.t2 1143.31
R98 VNB.t1 VNB.t0 1027.82
R99 VNB.t5 VNB.t6 993.177
R100 VNB.t3 VNB.t4 993.177
R101 A4.n0 A4.t1 250.909
R102 A4.n0 A4.t0 220.113
R103 A4 A4.n0 153.935
R104 a_27_74.n1 a_27_74.t1 199.591
R105 a_27_74.n2 a_27_74.n1 165.71
R106 a_27_74.n1 a_27_74.n0 101.71
R107 a_27_74.n2 a_27_74.t4 25.1356
R108 a_27_74.n0 a_27_74.t3 22.7032
R109 a_27_74.n0 a_27_74.t2 22.7032
R110 a_27_74.t0 a_27_74.n2 22.7032
R111 B1.n0 B1.t0 231.629
R112 B1.n0 B1.t1 220.113
R113 B1.n1 B1.n0 152
R114 B1 B1.n1 9.67492
R115 B1.n1 B1 4.61445
R116 A3.n0 A3.t1 250.909
R117 A3.n0 A3.t0 220.113
R118 A3 A3.n0 154.133
R119 A3.n1 A3 15.0266
R120 A3 A3.n1 5.56572
R121 A3.n1 A3 3.28255
R122 A2.n0 A2.t0 250.909
R123 A2.n0 A2.t1 220.113
R124 A2 A2.n0 168.51
R125 a_200_368.t0 a_200_368.t1 73.8755
R126 a_314_368.t0 a_314_368.t1 73.8755
C0 VPB A1 0.036315f
C1 B1 VGND 0.013315f
C2 A3 VPWR 0.035875f
C3 A2 VGND 0.017443f
C4 A4 VPB 0.037442f
C5 B1 A2 8.36e-20
C6 X VGND 0.135213f
C7 VPWR VGND 0.093863f
C8 B1 X 3.23e-19
C9 A3 A4 0.086591f
C10 VPWR B1 0.018814f
C11 A1 VGND 0.015976f
C12 A3 VPB 0.038231f
C13 VPWR A2 0.094704f
C14 VPWR X 0.179106f
C15 A4 VGND 0.01538f
C16 A1 A2 0.089706f
C17 A4 B1 0.0798f
C18 VPB VGND 0.008399f
C19 VPWR A1 0.055186f
C20 B1 VPB 0.046167f
C21 A3 VGND 0.018121f
C22 VPB A2 0.037367f
C23 A4 VPWR 0.013172f
C24 A3 B1 5.47e-19
C25 VPB X 0.004934f
C26 VPWR VPB 0.14753f
C27 A3 A2 0.161362f
C28 VGND VNB 0.627261f
C29 X VNB 0.03546f
C30 B1 VNB 0.120136f
C31 VPWR VNB 0.547692f
C32 A4 VNB 0.106261f
C33 A3 VNB 0.106957f
C34 A2 VNB 0.109548f
C35 A1 VNB 0.15441f
C36 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o41a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41a_1 VNB VPB VPWR VGND A4 B1 A1 A3 A2 X
X0 VPWR.t2 a_83_270.t3 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4712 pd=2.07 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t4 a_83_270.t4 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VGND.t2 A4.t0 a_326_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.112 ps=0.99 w=0.64 l=0.15
X3 a_527_368.t0 A3.t0 a_443_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X4 a_83_270.t0 B1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.200825 pd=1.505 as=0.4712 ps=2.07 w=0.84 l=0.15
X5 a_326_74.t4 B1.t1 a_83_270.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X6 a_326_74.t2 A3.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1088 pd=0.98 as=0.1344 ps=1.06 w=0.64 l=0.15
X7 a_443_368.t1 A4.t1 a_83_270.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.200825 ps=1.505 w=1.12 l=0.15
X8 a_641_368.t1 A2.t0 a_527_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X9 a_326_74.t0 A1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1792 ps=1.2 w=0.64 l=0.15
X10 VGND.t3 A2.t1 a_326_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1792 pd=1.2 as=0.1088 ps=0.98 w=0.64 l=0.15
X11 VPWR.t1 A1.t1 a_641_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.4592 pd=3.06 as=0.2352 ps=1.54 w=1.12 l=0.15
R0 a_83_270.n2 a_83_270.n1 394.252
R1 a_83_270.n0 a_83_270.t3 248.303
R2 a_83_270.n0 a_83_270.t4 217.508
R3 a_83_270.n1 a_83_270.t2 192.887
R4 a_83_270.n1 a_83_270.n0 152
R5 a_83_270.n4 a_83_270.n3 56.0753
R6 a_83_270.n2 a_83_270.t0 55.1136
R7 a_83_270.n3 a_83_270.t1 25.7866
R8 a_83_270.n3 a_83_270.n2 3.16009
R9 X X.n0 589.85
R10 X.n1 X.n0 585
R11 X X.t0 241.826
R12 X.n0 X.t1 26.3844
R13 X X.n1 9.11565
R14 X.n1 X 5.23686
R15 VPWR.n3 VPWR.n1 588.029
R16 VPWR.n4 VPWR.n0 585
R17 VPWR.n5 VPWR.t1 343.63
R18 VPWR.n3 VPWR.n2 301.06
R19 VPWR.n2 VPWR.n0 80.6115
R20 VPWR.n1 VPWR.n0 38.6969
R21 VPWR.n1 VPWR.t0 36.3517
R22 VPWR.n2 VPWR.t2 24.1092
R23 VPWR.n5 VPWR.n4 10.4363
R24 VPWR.n4 VPWR.n3 3.02956
R25 VPWR VPWR.n5 0.267985
R26 VPB.t5 VPB.t1 561.828
R27 VPB.t4 VPB.t2 291.13
R28 VPB.t0 VPB.t4 291.13
R29 VPB.t1 VPB.t3 273.253
R30 VPB VPB.t5 257.93
R31 VPB.t3 VPB.t0 214.517
R32 VGND.n3 VGND.n2 204.976
R33 VGND.n5 VGND.n4 190.796
R34 VGND.n10 VGND.t4 133.686
R35 VGND.n4 VGND.t0 58.1255
R36 VGND.n4 VGND.t3 46.8755
R37 VGND.n2 VGND.t1 39.3755
R38 VGND.n2 VGND.t2 39.3755
R39 VGND.n8 VGND.n1 36.1417
R40 VGND.n9 VGND.n8 36.1417
R41 VGND.n10 VGND.n9 19.2005
R42 VGND.n5 VGND.n3 17.1625
R43 VGND.n6 VGND.n1 9.3005
R44 VGND.n8 VGND.n7 9.3005
R45 VGND.n9 VGND.n0 9.3005
R46 VGND.n11 VGND.n10 7.19894
R47 VGND.n3 VGND.n1 1.12991
R48 VGND.n6 VGND.n5 0.756849
R49 VGND VGND.n11 0.156997
R50 VGND.n11 VGND.n0 0.150766
R51 VGND.n7 VGND.n6 0.122949
R52 VGND.n7 VGND.n0 0.122949
R53 VNB.t5 VNB.t4 2448.29
R54 VNB.t3 VNB.t0 1639.9
R55 VNB.t2 VNB.t1 1316.54
R56 VNB.t4 VNB.t2 1154.86
R57 VNB VNB.t5 1143.31
R58 VNB.t1 VNB.t3 1131.76
R59 A4.n0 A4.t1 291.926
R60 A4.n0 A4.t0 184.768
R61 A4 A4.n0 159.112
R62 a_326_74.t0 a_326_74.n2 200.871
R63 a_326_74.n2 a_326_74.n0 149.234
R64 a_326_74.n2 a_326_74.n1 98.788
R65 a_326_74.n0 a_326_74.t4 39.3755
R66 a_326_74.n1 a_326_74.t3 37.5005
R67 a_326_74.n0 a_326_74.t1 26.2505
R68 a_326_74.n1 a_326_74.t2 26.2505
R69 A3.n0 A3.t0 285.719
R70 A3.n0 A3.t1 194.407
R71 A3 A3.n0 159.565
R72 a_443_368.t0 a_443_368.t1 47.4916
R73 a_527_368.t0 a_527_368.t1 73.8755
R74 B1.n0 B1.t1 265.142
R75 B1.n0 B1.t0 196.089
R76 B1 B1.n0 163.637
R77 A2.n0 A2.t0 264.298
R78 A2.n0 A2.t1 220.113
R79 A2 A2.n0 156.034
R80 a_641_368.t0 a_641_368.t1 73.8755
R81 A1.n0 A1.t1 250.909
R82 A1.n0 A1.t0 236.18
R83 A1 A1.n0 153.423
C0 X VPWR 0.097331f
C1 VPWR A4 0.012444f
C2 A4 A3 0.111152f
C3 B1 VGND 0.013152f
C4 VGND A2 0.014639f
C5 B1 A1 1.41e-19
C6 VGND VPB 0.007739f
C7 A2 A1 0.105452f
C8 A1 VPB 0.043303f
C9 VPWR VGND 0.07122f
C10 VGND A3 0.01256f
C11 B1 A2 2.59e-19
C12 VPWR A1 0.069452f
C13 B1 VPB 0.071939f
C14 A3 A1 1.58e-19
C15 A2 VPB 0.037935f
C16 X VGND 0.082573f
C17 VPWR B1 0.019213f
C18 VPWR A2 0.066211f
C19 B1 A3 0.001532f
C20 VGND A4 0.014043f
C21 VPWR VPB 0.122682f
C22 A3 A2 0.174138f
C23 A4 A1 2.94e-20
C24 A3 VPB 0.034984f
C25 X B1 6.71e-19
C26 B1 A4 0.071976f
C27 VPWR A3 0.035628f
C28 X VPB 0.012551f
C29 A4 A2 8.01e-20
C30 A4 VPB 0.035554f
C31 VGND A1 0.016381f
C32 VGND VNB 0.549442f
C33 B1 VNB 0.135537f
C34 VPWR VNB 0.455778f
C35 X VNB 0.109151f
C36 A1 VNB 0.181245f
C37 A2 VNB 0.121898f
C38 A3 VNB 0.116605f
C39 A4 VNB 0.122155f
C40 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o32ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32ai_4 VNB VPB VPWR VGND Y B2 B1 A3 A2 A1
X0 Y.t7 B2.t0 a_27_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_861_368.t7 A3.t0 Y.t15 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_27_74.t9 B1.t0 Y.t10 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 a_27_74.t4 A2.t0 VGND.t7 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1554 ps=1.16 w=0.74 l=0.15
X4 VGND.t3 A3.t1 a_27_74.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.12765 ps=1.085 w=0.74 l=0.15
X5 a_1330_368.t7 A2.t1 a_861_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X6 Y.t3 B2.t1 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 VGND.t2 A3.t2 a_27_74.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1773 pd=1.28 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 Y.t8 B1.t1 a_27_74.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.12395 ps=1.075 w=0.74 l=0.15
X9 VPWR.t5 B1.t2 a_27_368.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VPWR.t0 A1.t0 a_1330_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_27_368.t5 B1.t3 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 Y.t11 A3.t3 a_861_368.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X13 Y.t12 A3.t4 a_861_368.t5 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_861_368.t4 A3.t5 Y.t13 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Y.t2 B2.t2 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 VPWR.t3 B1.t4 a_27_368.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_27_368.t2 B2.t3 Y.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_861_368.t1 A2.t2 a_1330_368.t6 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_27_74.t1 B2.t4 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.12395 pd=1.075 as=0.10915 ps=1.035 w=0.74 l=0.15
X20 a_27_74.t11 A3.t6 VGND.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.12765 pd=1.085 as=0.1773 ps=1.28 w=0.74 l=0.15
X21 VPWR.t1 A1.t1 a_1330_368.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X22 Y.t5 B2.t5 a_27_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_27_368.t0 B2.t6 Y.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_27_74.t7 B1.t5 Y.t9 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X25 a_27_74.t14 A1.t2 VGND.t4 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X26 a_27_74.t5 A2.t3 VGND.t6 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X27 a_1330_368.t2 A1.t3 VPWR.t6 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X28 a_27_368.t7 B1.t6 VPWR.t2 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1736 ps=1.43 w=1.12 l=0.15
X29 a_27_74.t0 B2.t7 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 a_1330_368.t5 A2.t4 a_861_368.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X31 a_1330_368.t3 A1.t4 VPWR.t7 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X32 Y.t14 B1.t7 a_27_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X33 a_27_74.t10 A3.t7 VGND.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2626 pd=1.455 as=0.10545 ps=1.025 w=0.74 l=0.15
X34 VGND.t5 A1.t5 a_27_74.t15 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X35 a_861_368.t3 A2.t5 a_1330_368.t4 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
R0 B2.n0 B2.t3 226.809
R1 B2.n3 B2.t5 226.809
R2 B2.n10 B2.t6 226.809
R3 B2.n4 B2.t0 226.809
R4 B2.n0 B2.t4 198.204
R5 B2.n4 B2.t1 197.475
R6 B2.n9 B2.t7 196.013
R7 B2.n2 B2.t2 196.013
R8 B2 B2.n1 152.184
R9 B2.n12 B2.n11 152
R10 B2.n8 B2.n7 152
R11 B2.n6 B2.n5 152
R12 B2.n8 B2.n5 49.6611
R13 B2.n11 B2.n10 44.549
R14 B2.n1 B2.n0 37.246
R15 B2.n2 B2.n1 25.5611
R16 B2.n11 B2.n3 21.1793
R17 B2.n6 B2 15.5434
R18 B2 B2.n12 12.2519
R19 B2.n5 B2.n4 10.955
R20 B2.n7 B2 10.4234
R21 B2.n7 B2 7.13193
R22 B2.n12 B2 5.30336
R23 B2.n10 B2.n9 4.38232
R24 B2.n3 B2.n2 2.92171
R25 B2 B2.n6 2.01193
R26 B2.n9 B2.n8 0.730803
R27 a_27_368.n1 a_27_368.t7 369.108
R28 a_27_368.n5 a_27_368.n4 305.998
R29 a_27_368.n1 a_27_368.n0 299.053
R30 a_27_368.n3 a_27_368.n2 287.964
R31 a_27_368.n4 a_27_368.t3 278.474
R32 a_27_368.n4 a_27_368.n3 72.9988
R33 a_27_368.n3 a_27_368.n1 56.0877
R34 a_27_368.n2 a_27_368.t6 26.3844
R35 a_27_368.n2 a_27_368.t2 26.3844
R36 a_27_368.n0 a_27_368.t4 26.3844
R37 a_27_368.n0 a_27_368.t5 26.3844
R38 a_27_368.n5 a_27_368.t1 26.3844
R39 a_27_368.t0 a_27_368.n5 26.3844
R40 Y.n12 Y.n0 356.074
R41 Y.n11 Y.n10 299.95
R42 Y.n9 Y.n1 296.8
R43 Y.n14 Y.n13 292.93
R44 Y.n4 Y.n2 248.418
R45 Y.n12 Y.n11 221.365
R46 Y.n9 Y.n8 218.894
R47 Y.n4 Y.n3 201.129
R48 Y.n6 Y.n5 185
R49 Y.n8 Y.n7 185
R50 Y.n8 Y.n6 56.7994
R51 Y.n11 Y.n9 55.3417
R52 Y.n6 Y.n4 53.6235
R53 Y.n7 Y.t14 34.0546
R54 Y.n5 Y.t8 34.0546
R55 Y.n13 Y.t6 26.3844
R56 Y.n13 Y.t5 26.3844
R57 Y.n1 Y.t15 26.3844
R58 Y.n1 Y.t12 26.3844
R59 Y.n10 Y.t13 26.3844
R60 Y.n10 Y.t11 26.3844
R61 Y.n0 Y.t4 26.3844
R62 Y.n0 Y.t7 26.3844
R63 Y.n3 Y.t1 25.1356
R64 Y.n7 Y.t9 22.7032
R65 Y.n5 Y.t10 22.7032
R66 Y.n2 Y.t0 22.7032
R67 Y.n2 Y.t3 22.7032
R68 Y.n3 Y.t2 22.7032
R69 Y.n14 Y.n12 7.02071
R70 Y Y.n14 3.9826
R71 VPB.t12 VPB.t17 541.399
R72 VPB.t16 VPB.t13 515.861
R73 VPB.t6 VPB.t18 280.914
R74 VPB.t19 VPB.t11 280.914
R75 VPB VPB.t3 257.93
R76 VPB.t4 VPB.t12 255.376
R77 VPB.t5 VPB.t4 255.376
R78 VPB.t8 VPB.t16 234.946
R79 VPB.t18 VPB.t7 229.839
R80 VPB.t17 VPB.t6 229.839
R81 VPB.t11 VPB.t5 229.839
R82 VPB.t14 VPB.t19 229.839
R83 VPB.t15 VPB.t14 229.839
R84 VPB.t13 VPB.t15 229.839
R85 VPB.t9 VPB.t8 229.839
R86 VPB.t10 VPB.t9 229.839
R87 VPB.t2 VPB.t10 229.839
R88 VPB.t1 VPB.t2 229.839
R89 VPB.t0 VPB.t1 229.839
R90 VPB.t3 VPB.t0 229.839
R91 A3.n4 A3.t2 283.065
R92 A3.n1 A3.t0 254.231
R93 A3.n2 A3.t4 226.809
R94 A3.n9 A3.t5 226.809
R95 A3.n4 A3.t3 226.809
R96 A3.n7 A3.t6 196.013
R97 A3.n3 A3.t1 196.013
R98 A3.n1 A3.t7 196.013
R99 A3.n11 A3.n10 152
R100 A3.n8 A3.n0 152
R101 A3.n6 A3.n5 152
R102 A3.n10 A3.n9 44.549
R103 A3.n2 A3.n1 43.8187
R104 A3.n7 A3.n6 28.4823
R105 A3.n8 A3.n7 21.1793
R106 A3.n3 A3.n2 19.7187
R107 A3.n11 A3.n0 12.4348
R108 A3.n6 A3.n4 10.955
R109 A3.n5 A3 10.0576
R110 A3.n5 A3 7.49764
R111 A3.n9 A3.n8 5.11262
R112 A3 A3.n0 4.93764
R113 A3.n10 A3.n3 1.46111
R114 A3 A3.n11 0.183357
R115 a_861_368.t6 a_861_368.n5 393.745
R116 a_861_368.n2 a_861_368.t3 388.365
R117 a_861_368.n5 a_861_368.n0 305.901
R118 a_861_368.n2 a_861_368.n1 302.74
R119 a_861_368.n4 a_861_368.n3 209.739
R120 a_861_368.n5 a_861_368.n4 59.8593
R121 a_861_368.n4 a_861_368.n2 50.4476
R122 a_861_368.n1 a_861_368.t1 35.1791
R123 a_861_368.n3 a_861_368.t2 35.1791
R124 a_861_368.n3 a_861_368.t7 35.1791
R125 a_861_368.n1 a_861_368.t0 26.3844
R126 a_861_368.n0 a_861_368.t5 26.3844
R127 a_861_368.n0 a_861_368.t4 26.3844
R128 B1.n2 B1.t4 234.112
R129 B1.n13 B1.t6 226.809
R130 B1.n1 B1.t2 226.809
R131 B1.n7 B1.t3 226.809
R132 B1.n14 B1.t5 212.81
R133 B1.n2 B1.t1 196.013
R134 B1.n8 B1.t0 196.013
R135 B1.n0 B1.t7 196.013
R136 B1.n15 B1.n14 152
R137 B1.n12 B1.n11 152
R138 B1.n10 B1.n9 152
R139 B1.n6 B1.n5 152
R140 B1.n4 B1.n3 152
R141 B1.n6 B1.n3 49.6611
R142 B1.n13 B1.n12 38.7066
R143 B1.n9 B1.n8 29.9429
R144 B1.n1 B1.n0 21.9096
R145 B1.n9 B1.n1 21.1793
R146 B1.n8 B1.n7 14.6066
R147 B1.n11 B1.n10 12.4348
R148 B1.n5 B1 11.5205
R149 B1.n4 B1 11.1548
R150 B1.n14 B1.n13 10.955
R151 B1 B1.n15 9.32621
R152 B1.n15 B1 8.22907
R153 B1.n12 B1.n0 6.57323
R154 B1 B1.n4 6.4005
R155 B1.n5 B1 6.03479
R156 B1.n7 B1.n6 5.11262
R157 B1.n11 B1 4.20621
R158 B1.n3 B1.n2 3.65202
R159 B1.n10 B1 0.914786
R160 a_27_74.t3 a_27_74.n13 208.738
R161 a_27_74.n1 a_27_74.t14 200.438
R162 a_27_74.n7 a_27_74.n6 185
R163 a_27_74.n9 a_27_74.n8 185
R164 a_27_74.n11 a_27_74.n10 185
R165 a_27_74.n13 a_27_74.n12 185
R166 a_27_74.n2 a_27_74.t5 149.99
R167 a_27_74.n3 a_27_74.t10 106.09
R168 a_27_74.n1 a_27_74.n0 101.71
R169 a_27_74.n5 a_27_74.n4 95.685
R170 a_27_74.n9 a_27_74.n7 65.0659
R171 a_27_74.n3 a_27_74.n2 61.3469
R172 a_27_74.n7 a_27_74.n5 59.711
R173 a_27_74.n5 a_27_74.n3 56.9675
R174 a_27_74.n11 a_27_74.n9 56.7994
R175 a_27_74.n13 a_27_74.n11 51.5289
R176 a_27_74.n2 a_27_74.n1 50.4476
R177 a_27_74.n12 a_27_74.t0 34.0546
R178 a_27_74.n8 a_27_74.t9 34.0546
R179 a_27_74.n6 a_27_74.t7 34.0546
R180 a_27_74.n0 a_27_74.t15 34.0546
R181 a_27_74.n4 a_27_74.t13 33.2437
R182 a_27_74.n10 a_27_74.t1 31.6221
R183 a_27_74.n12 a_27_74.t2 22.7032
R184 a_27_74.n10 a_27_74.t8 22.7032
R185 a_27_74.n8 a_27_74.t6 22.7032
R186 a_27_74.n6 a_27_74.t12 22.7032
R187 a_27_74.n0 a_27_74.t4 22.7032
R188 a_27_74.n4 a_27_74.t11 22.7032
R189 VNB.t10 VNB.t5 3268.24
R190 VNB.t5 VNB.t4 2309.71
R191 VNB.t12 VNB.t11 1362.73
R192 VNB.t15 VNB.t14 1154.86
R193 VNB.t4 VNB.t15 1154.86
R194 VNB.t7 VNB.t12 1154.86
R195 VNB.t6 VNB.t7 1154.86
R196 VNB.t9 VNB.t6 1154.86
R197 VNB.t8 VNB.t9 1154.86
R198 VNB.t0 VNB.t2 1154.86
R199 VNB.t11 VNB.t13 1143.31
R200 VNB VNB.t3 1143.31
R201 VNB.t1 VNB.t8 1120.21
R202 VNB.t2 VNB.t1 1027.82
R203 VNB.t13 VNB.t10 1004.72
R204 VNB.t3 VNB.t0 993.177
R205 A2.n4 A2.t4 242.023
R206 A2.n16 A2.t0 232.53
R207 A2.n15 A2.t5 226.809
R208 A2.n1 A2.t1 226.809
R209 A2.n8 A2.t2 226.809
R210 A2.n3 A2.n2 196.013
R211 A2.n9 A2.t3 196.013
R212 A2.n14 A2.n0 196.013
R213 A2.n17 A2.n16 152
R214 A2.n13 A2.n12 152
R215 A2.n11 A2.n10 152
R216 A2.n7 A2.n6 152
R217 A2.n5 A2.n4 152
R218 A2.n15 A2.n14 44.549
R219 A2.n7 A2.n3 43.8187
R220 A2.n9 A2.n8 38.7066
R221 A2.n13 A2.n1 25.5611
R222 A2.n10 A2.n1 24.1005
R223 A2.n10 A2.n9 10.2247
R224 A2.n12 A2.n11 10.1214
R225 A2.n6 A2 9.97259
R226 A2.n5 A2 8.48422
R227 A2 A2.n17 8.18655
R228 A2.n17 A2 6.10283
R229 A2.n4 A2.n3 5.84292
R230 A2 A2.n5 5.80515
R231 A2.n6 A2 4.31678
R232 A2.n12 A2 4.0191
R233 A2.n14 A2.n13 2.92171
R234 A2.n16 A2.n15 2.19141
R235 A2.n8 A2.n7 0.730803
R236 A2.n11 A2 0.149337
R237 VGND.n4 VGND.t7 242.133
R238 VGND.n9 VGND.t6 242.133
R239 VGND.n6 VGND.n5 213.531
R240 VGND.n14 VGND.n2 204.201
R241 VGND.n17 VGND.n16 201.097
R242 VGND.n10 VGND.n1 36.1417
R243 VGND.n16 VGND.t1 35.6762
R244 VGND.n16 VGND.t2 35.6762
R245 VGND.n15 VGND.n14 34.2593
R246 VGND.n5 VGND.t4 34.0546
R247 VGND.n8 VGND.n4 30.1181
R248 VGND.n10 VGND.n9 27.1064
R249 VGND.n2 VGND.t3 23.514
R250 VGND.n5 VGND.t5 22.7032
R251 VGND.n2 VGND.t0 22.7032
R252 VGND.n9 VGND.n8 20.3299
R253 VGND.n17 VGND.n15 16.9417
R254 VGND.n14 VGND.n1 13.177
R255 VGND.n15 VGND.n0 9.3005
R256 VGND.n14 VGND.n13 9.3005
R257 VGND.n12 VGND.n1 9.3005
R258 VGND.n11 VGND.n10 9.3005
R259 VGND.n9 VGND.n3 9.3005
R260 VGND.n8 VGND.n7 9.3005
R261 VGND.n18 VGND.n17 7.45461
R262 VGND.n6 VGND.n4 6.40205
R263 VGND VGND.n18 1.13953
R264 VGND.n7 VGND.n6 0.499311
R265 VGND.n18 VGND.n0 0.152559
R266 VGND.n7 VGND.n3 0.122949
R267 VGND.n11 VGND.n3 0.122949
R268 VGND.n12 VGND.n11 0.122949
R269 VGND.n13 VGND.n12 0.122949
R270 VGND.n13 VGND.n0 0.122949
R271 a_1330_368.n5 a_1330_368.n4 350.399
R272 a_1330_368.n4 a_1330_368.n3 299.95
R273 a_1330_368.n2 a_1330_368.n0 255.934
R274 a_1330_368.n2 a_1330_368.n1 205.487
R275 a_1330_368.n4 a_1330_368.n2 88.8476
R276 a_1330_368.n3 a_1330_368.t7 35.1791
R277 a_1330_368.n0 a_1330_368.t1 26.3844
R278 a_1330_368.n0 a_1330_368.t3 26.3844
R279 a_1330_368.n1 a_1330_368.t0 26.3844
R280 a_1330_368.n1 a_1330_368.t2 26.3844
R281 a_1330_368.n3 a_1330_368.t4 26.3844
R282 a_1330_368.t6 a_1330_368.n5 26.3844
R283 a_1330_368.n5 a_1330_368.t5 26.3844
R284 VPWR.n1 VPWR.n0 618.13
R285 VPWR.n33 VPWR.n3 618.13
R286 VPWR.n15 VPWR.t6 349.789
R287 VPWR.n11 VPWR.n10 315.928
R288 VPWR.n12 VPWR.t1 264.483
R289 VPWR.n16 VPWR.n8 36.1417
R290 VPWR.n20 VPWR.n8 36.1417
R291 VPWR.n21 VPWR.n20 36.1417
R292 VPWR.n22 VPWR.n21 36.1417
R293 VPWR.n22 VPWR.n6 36.1417
R294 VPWR.n26 VPWR.n6 36.1417
R295 VPWR.n27 VPWR.n26 36.1417
R296 VPWR.n28 VPWR.n27 36.1417
R297 VPWR.n28 VPWR.n4 36.1417
R298 VPWR.n32 VPWR.n4 36.1417
R299 VPWR.n35 VPWR.n34 36.1417
R300 VPWR.n37 VPWR.n1 35.5093
R301 VPWR.n10 VPWR.t7 35.1791
R302 VPWR.n10 VPWR.t0 35.1791
R303 VPWR.n15 VPWR.n14 31.2476
R304 VPWR.n3 VPWR.t2 28.1434
R305 VPWR.n0 VPWR.t4 26.3844
R306 VPWR.n0 VPWR.t3 26.3844
R307 VPWR.n3 VPWR.t5 26.3844
R308 VPWR.n34 VPWR.n33 23.3417
R309 VPWR.n16 VPWR.n15 22.2123
R310 VPWR.n14 VPWR.n11 21.4593
R311 VPWR.n33 VPWR.n32 12.8005
R312 VPWR.n14 VPWR.n13 9.3005
R313 VPWR.n15 VPWR.n9 9.3005
R314 VPWR.n17 VPWR.n16 9.3005
R315 VPWR.n18 VPWR.n8 9.3005
R316 VPWR.n20 VPWR.n19 9.3005
R317 VPWR.n21 VPWR.n7 9.3005
R318 VPWR.n23 VPWR.n22 9.3005
R319 VPWR.n24 VPWR.n6 9.3005
R320 VPWR.n26 VPWR.n25 9.3005
R321 VPWR.n27 VPWR.n5 9.3005
R322 VPWR.n29 VPWR.n28 9.3005
R323 VPWR.n30 VPWR.n4 9.3005
R324 VPWR.n32 VPWR.n31 9.3005
R325 VPWR.n34 VPWR.n2 9.3005
R326 VPWR.n36 VPWR.n35 9.3005
R327 VPWR.n35 VPWR.n1 8.28285
R328 VPWR.n12 VPWR.n11 6.8344
R329 VPWR.n13 VPWR.n12 0.569119
R330 VPWR VPWR.n37 0.527539
R331 VPWR.n37 VPWR.n36 0.149442
R332 VPWR.n13 VPWR.n9 0.122949
R333 VPWR.n17 VPWR.n9 0.122949
R334 VPWR.n18 VPWR.n17 0.122949
R335 VPWR.n19 VPWR.n18 0.122949
R336 VPWR.n19 VPWR.n7 0.122949
R337 VPWR.n23 VPWR.n7 0.122949
R338 VPWR.n24 VPWR.n23 0.122949
R339 VPWR.n25 VPWR.n24 0.122949
R340 VPWR.n25 VPWR.n5 0.122949
R341 VPWR.n29 VPWR.n5 0.122949
R342 VPWR.n30 VPWR.n29 0.122949
R343 VPWR.n31 VPWR.n30 0.122949
R344 VPWR.n31 VPWR.n2 0.122949
R345 VPWR.n36 VPWR.n2 0.122949
R346 A1.n1 A1.t1 306.046
R347 A1.n2 A1.t4 226.809
R348 A1.n4 A1.t0 226.809
R349 A1.n8 A1.t3 226.809
R350 A1.n7 A1.t5 216.463
R351 A1.n6 A1.t2 196.013
R352 A1.n13 A1.n3 196.013
R353 A1.n1 A1.n0 196.013
R354 A1.n15 A1.n14 152
R355 A1.n12 A1.n11 152
R356 A1.n10 A1.n9 152
R357 A1.n7 A1.n5 152
R358 A1.n6 A1.n4 35.7853
R359 A1.n14 A1.n13 33.5944
R360 A1.n9 A1.n8 27.0217
R361 A1.n8 A1.n7 22.6399
R362 A1.n2 A1.n1 19.7187
R363 A1.n14 A1.n2 19.7187
R364 A1.n13 A1.n12 16.0672
R365 A1.n12 A1.n4 10.955
R366 A1.n10 A1.n5 10.1214
R367 A1.n11 A1 9.97259
R368 A1 A1.n15 8.48422
R369 A1.n15 A1 5.80515
R370 A1.n11 A1 4.31678
R371 A1.n5 A1 4.0191
R372 A1.n9 A1.n6 2.92171
R373 A1 A1.n10 0.149337
C0 VPWR VGND 0.172712f
C1 A2 Y 0.023084f
C2 B2 VGND 0.026198f
C3 A2 VPB 0.16242f
C4 A1 Y 2.77e-19
C5 A2 VPWR 0.026701f
C6 B1 VGND 0.026842f
C7 A1 VPB 0.167317f
C8 A1 VPWR 0.102796f
C9 A3 VGND 0.051871f
C10 Y VPB 0.019401f
C11 Y VPWR 0.06532f
C12 A2 A3 0.034166f
C13 VPWR VPB 0.266197f
C14 Y B2 0.324812f
C15 VPB B2 0.138144f
C16 VPWR B2 0.025233f
C17 Y B1 0.460299f
C18 VPB B1 0.150882f
C19 VPWR B1 0.049508f
C20 Y A3 0.356339f
C21 B2 B1 0.080598f
C22 VPB A3 0.14985f
C23 VPWR A3 0.02413f
C24 B1 A3 0.059441f
C25 A2 VGND 0.069798f
C26 A1 VGND 0.07276f
C27 Y VGND 0.055692f
C28 A2 A1 0.068007f
C29 VPB VGND 0.012569f
C30 VGND VNB 1.22224f
C31 VPWR VNB 1.01915f
C32 Y VNB 0.054103f
C33 A1 VNB 0.487347f
C34 A2 VNB 0.449071f
C35 A3 VNB 0.434389f
C36 B1 VNB 0.425683f
C37 B2 VNB 0.442296f
C38 VPB VNB 2.54894f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o32ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32ai_2 VNB VPB VPWR VGND B2 B1 A3 A2 A1 Y
X0 Y.t3 B2.t0 a_27_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_499_368.t3 A2.t0 a_768_368.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_27_74.t9 A2.t1 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1221 ps=1.07 w=0.74 l=0.15
X3 a_27_74.t4 A1.t0 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.3367 ps=1.65 w=0.74 l=0.15
X4 a_768_368.t2 A2.t2 a_499_368.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_27_74.t2 B1.t0 Y.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X6 a_499_368.t1 A3.t0 Y.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t1 B2.t1 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VGND.t4 A2.t3 a_27_74.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.12765 ps=1.085 w=0.74 l=0.15
X9 Y.t4 A3.t1 a_499_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X10 Y.t7 B1.t1 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 a_27_74.t5 A3.t2 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12765 pd=1.085 as=0.2993 ps=1.6 w=0.74 l=0.15
X12 a_27_368.t3 B1.t2 VPWR.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VPWR.t0 B1.t3 a_27_368.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_27_368.t0 B2.t2 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_768_368.t1 A1.t1 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.3864 ps=2.93 w=1.12 l=0.15
X16 a_27_74.t0 B2.t3 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t0 A1.t2 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.3367 pd=1.65 as=0.11285 ps=1.045 w=0.74 l=0.15
X18 VPWR.t2 A1.t3 a_768_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1708 ps=1.425 w=1.12 l=0.15
X19 VGND.t3 A3.t3 a_27_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2993 pd=1.6 as=0.1295 ps=1.09 w=0.74 l=0.15
R0 B2.n0 B2.t2 231.19
R1 B2.n3 B2.t0 226.809
R2 B2.n2 B2.t1 196.013
R3 B2.n0 B2.t3 196.013
R4 B2.n5 B2.n4 152
R5 B2.n2 B2.n1 152
R6 B2.n4 B2.n3 48.2005
R7 B2.n4 B2.n0 13.146
R8 B2.n1 B2 10.1214
R9 B2 B2.n5 8.33538
R10 B2.n5 B2 5.95399
R11 B2.n1 B2 4.16794
R12 B2.n3 B2.n2 1.46111
R13 a_27_368.n0 a_27_368.t3 393.846
R14 a_27_368.n0 a_27_368.t1 321.233
R15 a_27_368.n1 a_27_368.n0 285.967
R16 a_27_368.n1 a_27_368.t2 26.3844
R17 a_27_368.t0 a_27_368.n1 26.3844
R18 Y.n2 Y 594.697
R19 Y.n3 Y.n2 585
R20 Y.n1 Y.n0 452.798
R21 Y.n6 Y.n4 251.565
R22 Y.n6 Y.n5 185
R23 Y Y.n6 142.395
R24 Y.n5 Y.t7 34.0546
R25 Y.n2 Y.t6 26.3844
R26 Y.n2 Y.t4 26.3844
R27 Y.n0 Y.t2 26.3844
R28 Y.n0 Y.t3 26.3844
R29 Y.n5 Y.t5 22.7032
R30 Y.n4 Y.t0 22.7032
R31 Y.n4 Y.t1 22.7032
R32 Y Y.n1 11.055
R33 Y.n3 Y.n1 1.93989
R34 Y Y.n3 1.35808
R35 VPB.t0 VPB.t6 541.399
R36 VPB.t9 VPB.t5 515.861
R37 VPB VPB.t3 257.93
R38 VPB.t6 VPB.t4 232.393
R39 VPB.t1 VPB.t0 229.839
R40 VPB.t8 VPB.t1 229.839
R41 VPB.t5 VPB.t8 229.839
R42 VPB.t7 VPB.t9 229.839
R43 VPB.t2 VPB.t7 229.839
R44 VPB.t3 VPB.t2 229.839
R45 A2.n0 A2.t0 226.809
R46 A2.n1 A2.t2 226.809
R47 A2.n1 A2.t3 198.204
R48 A2.n0 A2.t1 198.204
R49 A2.n3 A2.n2 152
R50 A2.n2 A2.n0 54.7732
R51 A2.n2 A2.n1 10.955
R52 A2.n3 A2 9.67492
R53 A2 A2.n3 4.61445
R54 a_768_368.n1 a_768_368.n0 600.081
R55 a_768_368.t0 a_768_368.n1 27.2639
R56 a_768_368.n0 a_768_368.t3 26.3844
R57 a_768_368.n0 a_768_368.t2 26.3844
R58 a_768_368.n1 a_768_368.t1 26.3844
R59 a_499_368.n0 a_499_368.t0 393.745
R60 a_499_368.n0 a_499_368.t3 384.464
R61 a_499_368.n1 a_499_368.n0 215.828
R62 a_499_368.t2 a_499_368.n1 26.3844
R63 a_499_368.n1 a_499_368.t1 26.3844
R64 VGND.n11 VGND.n4 209.631
R65 VGND.n1 VGND.n0 192.925
R66 VGND.n8 VGND.n7 187.329
R67 VGND.n6 VGND.n5 185
R68 VGND.n7 VGND.n6 102.162
R69 VGND.n0 VGND.t2 55.1356
R70 VGND.n0 VGND.t3 55.1356
R71 VGND.n13 VGND.n12 35.8746
R72 VGND.n11 VGND.n3 32.0005
R73 VGND.n4 VGND.t5 30.0005
R74 VGND.n4 VGND.t4 23.514
R75 VGND.n7 VGND.t1 22.7032
R76 VGND.n6 VGND.t0 22.7032
R77 VGND.n5 VGND.n3 19.8139
R78 VGND.n12 VGND.n11 15.4358
R79 VGND.n15 VGND.n1 11.8726
R80 VGND.n14 VGND.n13 9.3005
R81 VGND.n12 VGND.n2 9.3005
R82 VGND.n9 VGND.n3 9.3005
R83 VGND.n11 VGND.n10 9.3005
R84 VGND.n13 VGND.n1 6.127
R85 VGND.n8 VGND.n5 4.71819
R86 VGND.n9 VGND.n8 3.09216
R87 VGND VGND.n15 0.648083
R88 VGND.n15 VGND.n14 0.151892
R89 VGND.n10 VGND.n9 0.122949
R90 VGND.n10 VGND.n2 0.122949
R91 VGND.n14 VGND.n2 0.122949
R92 a_27_74.n1 a_27_74.t4 236.486
R93 a_27_74.t1 a_27_74.n7 209.268
R94 a_27_74.n5 a_27_74.n4 185
R95 a_27_74.n7 a_27_74.n6 185
R96 a_27_74.n1 a_27_74.n0 101.71
R97 a_27_74.n3 a_27_74.n2 92.7788
R98 a_27_74.n5 a_27_74.n3 80.3156
R99 a_27_74.n7 a_27_74.n5 64.0437
R100 a_27_74.n3 a_27_74.n1 59.3797
R101 a_27_74.n6 a_27_74.t0 34.0546
R102 a_27_74.n4 a_27_74.t2 34.0546
R103 a_27_74.n2 a_27_74.t8 33.2437
R104 a_27_74.n0 a_27_74.t9 26.7573
R105 a_27_74.n6 a_27_74.t7 22.7032
R106 a_27_74.n4 a_27_74.t6 22.7032
R107 a_27_74.n2 a_27_74.t5 22.7032
R108 a_27_74.n0 a_27_74.t3 22.7032
R109 VNB.t3 VNB.t4 2448.29
R110 VNB.t6 VNB.t5 1917.06
R111 VNB.t2 VNB.t6 1154.86
R112 VNB.t7 VNB.t2 1154.86
R113 VNB.t0 VNB.t7 1154.86
R114 VNB.t5 VNB.t8 1143.31
R115 VNB VNB.t1 1143.31
R116 VNB.t8 VNB.t9 1108.66
R117 VNB.t9 VNB.t3 1050.92
R118 VNB.t1 VNB.t0 993.177
R119 A1.n1 A1.t3 226.809
R120 A1.n3 A1.t1 226.809
R121 A1.n5 A1.t2 209.16
R122 A1.n1 A1.t0 198.204
R123 A1.n2 A1.n0 152
R124 A1.n7 A1.n6 152
R125 A1.n5 A1.n4 152
R126 A1.n6 A1.n5 49.6611
R127 A1.n2 A1.n1 40.1672
R128 A1.n3 A1.n2 26.2914
R129 A1.n6 A1.n3 23.3702
R130 A1.n0 A1 13.6935
R131 A1 A1.n7 9.52608
R132 A1.n4 A1 8.93073
R133 A1.n4 A1 5.35864
R134 A1.n7 A1 4.76329
R135 A1 A1.n0 0.595849
R136 B1.n1 B1.t3 229.73
R137 B1.n0 B1.t2 226.809
R138 B1.n0 B1.t0 208.677
R139 B1.n1 B1.t1 196.013
R140 B1 B1.n2 154.522
R141 B1.n2 B1.n1 32.8641
R142 B1.n2 B1.n0 29.9429
R143 A3.n0 A3.t0 234.026
R144 A3.n1 A3.t1 226.809
R145 A3.n2 A3.t3 209.16
R146 A3.n0 A3.t2 196.013
R147 A3.n3 A3.n2 152
R148 A3.n1 A3.n0 56.9641
R149 A3.n2 A3.n1 51.1217
R150 A3.n3 A3 13.0982
R151 A3 A3.n3 1.1912
R152 VPWR.n15 VPWR.n1 611.88
R153 VPWR.n4 VPWR.t3 351.106
R154 VPWR.n5 VPWR.t2 264.471
R155 VPWR.n8 VPWR.n7 36.1417
R156 VPWR.n9 VPWR.n8 36.1417
R157 VPWR.n9 VPWR.n2 36.1417
R158 VPWR.n13 VPWR.n2 36.1417
R159 VPWR.n14 VPWR.n13 36.1417
R160 VPWR.n15 VPWR.n14 33.5064
R161 VPWR.n1 VPWR.t1 26.3844
R162 VPWR.n1 VPWR.t0 26.3844
R163 VPWR.n7 VPWR.n4 20.7064
R164 VPWR.n7 VPWR.n6 9.3005
R165 VPWR.n8 VPWR.n3 9.3005
R166 VPWR.n10 VPWR.n9 9.3005
R167 VPWR.n11 VPWR.n2 9.3005
R168 VPWR.n13 VPWR.n12 9.3005
R169 VPWR.n14 VPWR.n0 9.3005
R170 VPWR.n16 VPWR.n15 6.92964
R171 VPWR.n5 VPWR.n4 6.87272
R172 VPWR.n6 VPWR.n5 0.565013
R173 VPWR VPWR.n16 0.393166
R174 VPWR.n16 VPWR.n0 0.160603
R175 VPWR.n6 VPWR.n3 0.122949
R176 VPWR.n10 VPWR.n3 0.122949
R177 VPWR.n11 VPWR.n10 0.122949
R178 VPWR.n12 VPWR.n11 0.122949
R179 VPWR.n12 VPWR.n0 0.122949
C0 Y VPWR 0.036676f
C1 B1 VPWR 0.02832f
C2 A3 Y 0.227813f
C3 B1 A3 0.073439f
C4 Y VGND 0.033642f
C5 A2 Y 0.022736f
C6 B1 VGND 0.011958f
C7 A3 VPWR 0.014152f
C8 Y VPB 0.015868f
C9 B1 VPB 0.066448f
C10 VPWR VGND 0.100126f
C11 A2 VPWR 0.013004f
C12 A1 Y 3.88e-19
C13 A3 VGND 0.02784f
C14 A3 A2 0.057953f
C15 VPWR VPB 0.169135f
C16 Y B2 0.17516f
C17 A3 VPB 0.08805f
C18 B1 B2 0.095431f
C19 A1 VPWR 0.067915f
C20 A2 VGND 0.035703f
C21 VGND VPB 0.009953f
C22 VPWR B2 0.013532f
C23 A2 VPB 0.066241f
C24 A1 VGND 0.041198f
C25 A2 A1 0.075182f
C26 VGND B2 0.014264f
C27 A1 VPB 0.10421f
C28 VPB B2 0.070824f
C29 B1 Y 0.112151f
C30 VGND VNB 0.70994f
C31 VPWR VNB 0.617045f
C32 Y VNB 0.031051f
C33 A1 VNB 0.315827f
C34 A2 VNB 0.19504f
C35 A3 VNB 0.246319f
C36 B1 VNB 0.198119f
C37 B2 VNB 0.251746f
C38 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o32ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32ai_1 VNB VPB VPWR VGND Y B2 B1 A3 A2 A1
X0 a_456_368.t0 A2.t0 a_342_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X1 a_128_368.t1 B1.t0 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3752 ps=2.91 w=1.12 l=0.15
X2 VPWR.t1 A1.t0 a_456_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X3 Y.t3 B1.t1 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.21645 pd=1.325 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 VGND.t2 A3.t0 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1665 pd=1.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 a_27_74.t0 A2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1665 ps=1.19 w=0.74 l=0.15
X6 Y.t0 B2.t0 a_128_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.28 pd=1.62 as=0.1512 ps=1.39 w=1.12 l=0.15
X7 a_27_74.t1 B2.t1 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.21645 ps=1.325 w=0.74 l=0.15
X8 VGND.t1 A1.t1 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_342_368.t0 A3.t1 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.28 ps=1.62 w=1.12 l=0.15
R0 A2.n0 A2.t0 250.909
R1 A2.n0 A2.t1 220.113
R2 A2 A2.n0 154.081
R3 a_342_368.t0 a_342_368.t1 73.8755
R4 a_456_368.t0 a_456_368.t1 73.8755
R5 VPB.t0 VPB.t1 331.99
R6 VPB.t2 VPB.t4 291.13
R7 VPB.t1 VPB.t2 291.13
R8 VPB VPB.t3 288.575
R9 VPB.t3 VPB.t0 214.517
R10 B1.n0 B1.t0 281.305
R11 B1.n0 B1.t1 171.72
R12 B1 B1.n0 158.788
R13 VPWR.n0 VPWR.t0 263.995
R14 VPWR.n0 VPWR.t1 257.271
R15 VPWR VPWR.n0 0.101024
R16 a_128_368.t0 a_128_368.t1 47.4916
R17 A1.n0 A1.t0 276.767
R18 A1.n0 A1.t1 169.389
R19 A1 A1.n0 158.31
R20 a_27_74.n1 a_27_74.t4 219.373
R21 a_27_74.n2 a_27_74.n1 167.793
R22 a_27_74.n1 a_27_74.n0 88.3339
R23 a_27_74.n0 a_27_74.t1 34.0546
R24 a_27_74.n0 a_27_74.t3 22.7032
R25 a_27_74.n2 a_27_74.t2 22.7032
R26 a_27_74.t0 a_27_74.n2 22.7032
R27 Y Y.n0 587.163
R28 Y.n2 Y.n0 290.995
R29 Y.n2 Y.n1 257.971
R30 Y.n0 Y.t1 61.563
R31 Y.n1 Y.t3 52.7032
R32 Y.n1 Y.t2 42.1627
R33 Y.n0 Y.t0 26.3844
R34 Y Y.n2 6.90434
R35 VNB.t4 VNB.t1 1697.64
R36 VNB.t3 VNB.t0 1385.83
R37 VNB.t1 VNB.t3 1154.86
R38 VNB VNB.t4 1143.31
R39 VNB.t0 VNB.t2 993.177
R40 A3.n0 A3.t1 250.909
R41 A3.n0 A3.t0 220.113
R42 A3 A3.n0 154.522
R43 VGND.n1 VGND.n0 215.202
R44 VGND.n1 VGND.t1 150.775
R45 VGND.n0 VGND.t0 38.9194
R46 VGND.n0 VGND.t2 34.0546
R47 VGND VGND.n1 0.844743
R48 B2.n0 B2.t0 246.206
R49 B2.n0 B2.t1 215.411
R50 B2 B2.n0 154.447
C0 B2 VPB 0.037707f
C1 VPWR Y 0.186164f
C2 A1 VGND 0.047144f
C3 B1 VGND 0.008813f
C4 A2 A1 0.075023f
C5 A3 VPWR 0.02109f
C6 B2 Y 0.11268f
C7 B2 A3 0.079365f
C8 A1 VPB 0.044611f
C9 B1 VPB 0.041907f
C10 A1 Y 0.002185f
C11 B1 Y 0.054504f
C12 B2 VPWR 0.005809f
C13 A3 A1 2.79e-19
C14 A2 VGND 0.016975f
C15 VGND VPB 0.00783f
C16 A1 VPWR 0.048639f
C17 A2 VPB 0.039366f
C18 B2 A1 1.49e-19
C19 B1 VPWR 0.049012f
C20 Y VGND 0.013475f
C21 B1 B2 0.049063f
C22 A3 VGND 0.013481f
C23 A2 Y 0.01358f
C24 A3 A2 0.146267f
C25 Y VPB 0.008911f
C26 A3 VPB 0.037949f
C27 VPWR VGND 0.057105f
C28 B2 VGND 0.006955f
C29 A2 VPWR 0.092133f
C30 A3 Y 0.061064f
C31 VPWR VPB 0.116366f
C32 VGND VNB 0.461038f
C33 Y VNB 0.025685f
C34 VPWR VNB 0.434056f
C35 A1 VNB 0.175437f
C36 A2 VNB 0.112639f
C37 A3 VNB 0.105599f
C38 B2 VNB 0.115149f
C39 B1 VNB 0.17491f
C40 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o32a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32a_4 VNB VPB VPWR VGND B2 A3 A2 A1 X B1
X0 VPWR.t7 B1.t0 a_534_388.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.15 ps=1.3 w=1 l=0.15
X1 X.t7 a_83_256.t8 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_534_388.t1 B2.t0 a_83_256.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X3 X.t0 a_83_256.t9 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.14985 pd=1.145 as=0.1554 ps=1.16 w=0.74 l=0.15
X4 a_564_74.t3 A2.t0 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
X5 a_83_256.t0 B2.t1 a_534_388.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.22 ps=1.44 w=1 l=0.15
X6 a_961_392.t1 A2.t1 a_1234_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X7 VGND.t2 A3.t0 a_564_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.01 as=0.1216 ps=1.02 w=0.64 l=0.15
X8 a_1234_392.t3 A1.t0 VPWR.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.16 ps=1.32 w=1 l=0.15
X9 a_564_74.t1 B2.t2 a_83_256.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1216 pd=1.02 as=0.112 ps=0.99 w=0.64 l=0.15
X10 a_534_388.t2 B1.t1 VPWR.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.44 as=0.2262 ps=1.54 w=1 l=0.15
X11 a_83_256.t3 A3.t1 a_961_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.295 ps=2.59 w=1 l=0.15
X12 X.t6 a_83_256.t10 VPWR.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X13 VGND.t1 A2.t2 a_564_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.096 ps=0.94 w=0.64 l=0.15
X14 VPWR.t2 a_83_256.t11 X.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2262 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X15 a_83_256.t2 B2.t3 a_564_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.112 ps=0.99 w=0.64 l=0.15
X16 VPWR.t4 A1.t1 a_1234_392.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.245 ps=1.49 w=1 l=0.15
X17 a_83_256.t7 B1.t2 a_564_74.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X18 X.t3 a_83_256.t12 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2543 ps=2.19 w=0.74 l=0.15
X19 VPWR.t3 a_83_256.t13 X.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_564_74.t6 B1.t3 a_83_256.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X21 a_564_74.t5 A1.t2 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.152 ps=1.115 w=0.64 l=0.15
X22 VGND.t5 a_83_256.t14 X.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_1234_392.t0 A2.t3 a_961_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.245 pd=1.49 as=0.15 ps=1.3 w=1 l=0.15
X24 a_961_392.t3 A3.t2 a_83_256.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.16 ps=1.32 w=1 l=0.15
X25 VGND.t4 a_83_256.t15 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.14985 ps=1.145 w=0.74 l=0.15
R0 B1.n2 B1.t0 1335.89
R1 B1.n0 B1.t3 266.707
R2 B1.n1 B1.t1 230.251
R3 B1.n1 B1.n0 218.737
R4 B1.n2 B1.n1 152
R5 B1.n0 B1.t2 128.534
R6 B1 B1.n2 5.23686
R7 a_534_388.n1 a_534_388.n0 1217.75
R8 a_534_388.t0 a_534_388.n1 43.3405
R9 a_534_388.n1 a_534_388.t2 43.3405
R10 a_534_388.n0 a_534_388.t3 29.5505
R11 a_534_388.n0 a_534_388.t1 29.5505
R12 VPWR.n8 VPWR.t7 805.801
R13 VPWR.n9 VPWR.n7 611.359
R14 VPWR.n19 VPWR.n2 317.527
R15 VPWR.n21 VPWR.t0 259.171
R16 VPWR.n4 VPWR.n3 222.361
R17 VPWR.n3 VPWR.t6 53.1905
R18 VPWR.n12 VPWR.n6 36.1417
R19 VPWR.n13 VPWR.n12 36.1417
R20 VPWR.n14 VPWR.n13 36.1417
R21 VPWR.n2 VPWR.t3 35.1791
R22 VPWR.n7 VPWR.t5 31.5205
R23 VPWR.n7 VPWR.t4 31.5205
R24 VPWR.n18 VPWR.n4 30.4946
R25 VPWR.n21 VPWR.n20 26.7299
R26 VPWR.n2 VPWR.t1 26.3844
R27 VPWR.n20 VPWR.n19 25.977
R28 VPWR.n3 VPWR.t2 25.9148
R29 VPWR.n19 VPWR.n18 21.4593
R30 VPWR.n14 VPWR.n4 16.9417
R31 VPWR.n9 VPWR.n8 10.2842
R32 VPWR.n10 VPWR.n6 9.3005
R33 VPWR.n12 VPWR.n11 9.3005
R34 VPWR.n13 VPWR.n5 9.3005
R35 VPWR.n15 VPWR.n14 9.3005
R36 VPWR.n16 VPWR.n4 9.3005
R37 VPWR.n18 VPWR.n17 9.3005
R38 VPWR.n19 VPWR.n1 9.3005
R39 VPWR.n20 VPWR.n0 9.3005
R40 VPWR.n22 VPWR.n21 9.3005
R41 VPWR.n8 VPWR.n6 8.65932
R42 VPWR.n10 VPWR.n9 0.150996
R43 VPWR.n11 VPWR.n10 0.122949
R44 VPWR.n11 VPWR.n5 0.122949
R45 VPWR.n15 VPWR.n5 0.122949
R46 VPWR.n16 VPWR.n15 0.122949
R47 VPWR.n17 VPWR.n16 0.122949
R48 VPWR.n17 VPWR.n1 0.122949
R49 VPWR.n1 VPWR.n0 0.122949
R50 VPWR.n22 VPWR.n0 0.122949
R51 VPWR VPWR.n22 0.0617245
R52 VPB.t13 VPB.t4 556.721
R53 VPB.t3 VPB.t10 326.882
R54 VPB.t12 VPB.t1 301.344
R55 VPB.t8 VPB.t12 291.13
R56 VPB.t7 VPB.t8 291.13
R57 VPB VPB.t0 257.93
R58 VPB.t9 VPB.t7 255.376
R59 VPB.t10 VPB.t11 240.054
R60 VPB.t4 VPB.t6 240.054
R61 VPB.t11 VPB.t2 229.839
R62 VPB.t6 VPB.t3 229.839
R63 VPB.t5 VPB.t13 229.839
R64 VPB.t1 VPB.t5 229.839
R65 VPB.t0 VPB.t9 229.839
R66 a_83_256.n16 a_83_256.n0 765.078
R67 a_83_256.n17 a_83_256.n16 586.553
R68 a_83_256.n2 a_83_256.t8 335.526
R69 a_83_256.n3 a_83_256.t13 293.752
R70 a_83_256.n9 a_83_256.t11 245.553
R71 a_83_256.n6 a_83_256.t10 245.553
R72 a_83_256.n14 a_83_256.n12 243.399
R73 a_83_256.n14 a_83_256.n13 195.093
R74 a_83_256.n10 a_83_256.t15 186.666
R75 a_83_256.n2 a_83_256.t12 173.52
R76 a_83_256.n4 a_83_256.t14 173.52
R77 a_83_256.n7 a_83_256.t9 173.52
R78 a_83_256.n5 a_83_256.n1 165.189
R79 a_83_256.n8 a_83_256.n1 152
R80 a_83_256.n11 a_83_256.n10 152
R81 a_83_256.n3 a_83_256.n2 102.828
R82 a_83_256.n5 a_83_256.n4 85.1538
R83 a_83_256.n15 a_83_256.n11 78.8768
R84 a_83_256.n12 a_83_256.t2 39.3755
R85 a_83_256.n9 a_83_256.n8 38.7066
R86 a_83_256.n4 a_83_256.n3 35.3472
R87 a_83_256.n0 a_83_256.t5 33.4905
R88 a_83_256.n16 a_83_256.n15 33.3581
R89 a_83_256.n0 a_83_256.t3 29.5505
R90 a_83_256.n17 a_83_256.t4 29.5505
R91 a_83_256.t0 a_83_256.n17 29.5505
R92 a_83_256.n7 a_83_256.n6 26.2914
R93 a_83_256.n13 a_83_256.t6 26.2505
R94 a_83_256.n13 a_83_256.t7 26.2505
R95 a_83_256.n12 a_83_256.t1 26.2505
R96 a_83_256.n8 a_83_256.n7 18.2581
R97 a_83_256.n11 a_83_256.n1 13.1884
R98 a_83_256.n10 a_83_256.n9 10.955
R99 a_83_256.n15 a_83_256.n14 7.97439
R100 a_83_256.n6 a_83_256.n5 5.11262
R101 X.n5 X.n3 258.822
R102 X.n5 X.n4 208.375
R103 X.n2 X.n0 150.042
R104 X.n2 X.n1 98.9958
R105 X.n6 X.n5 46.3704
R106 X.n0 X.t1 42.9735
R107 X.n3 X.t5 38.6969
R108 X.n3 X.t6 35.1791
R109 X.n6 X.n2 32.6051
R110 X.n4 X.t4 26.3844
R111 X.n4 X.t7 26.3844
R112 X.n1 X.t2 22.7032
R113 X.n1 X.t3 22.7032
R114 X.n0 X.t0 22.7032
R115 X X.n6 0.835283
R116 B2.n0 B2.t1 329.368
R117 B2.n1 B2.t2 242.607
R118 B2.n0 B2.t0 184.768
R119 B2 B2.n2 157.625
R120 B2.n2 B2.n0 143.286
R121 B2.n1 B2.t3 139.488
R122 B2.n2 B2.n1 39.4369
R123 VGND.n7 VGND.t3 252.44
R124 VGND.n6 VGND.t2 239.114
R125 VGND.n27 VGND.n2 206.721
R126 VGND.n9 VGND.n8 205.171
R127 VGND.n29 VGND.t6 150.923
R128 VGND.n22 VGND.t4 138.363
R129 VGND.n8 VGND.t1 39.3755
R130 VGND.n15 VGND.n14 36.1417
R131 VGND.n16 VGND.n15 36.1417
R132 VGND.n16 VGND.n4 36.1417
R133 VGND.n20 VGND.n4 36.1417
R134 VGND.n21 VGND.n20 36.1417
R135 VGND.n23 VGND.n1 36.1417
R136 VGND.n28 VGND.n27 35.0123
R137 VGND.n2 VGND.t7 34.0546
R138 VGND.n2 VGND.t5 34.0546
R139 VGND.n10 VGND.n6 33.1299
R140 VGND.n8 VGND.t0 26.2505
R141 VGND.n10 VGND.n9 17.3181
R142 VGND.n29 VGND.n28 15.4358
R143 VGND.n14 VGND.n6 14.3064
R144 VGND.n27 VGND.n1 12.424
R145 VGND.n30 VGND.n29 9.3005
R146 VGND.n11 VGND.n10 9.3005
R147 VGND.n12 VGND.n6 9.3005
R148 VGND.n14 VGND.n13 9.3005
R149 VGND.n15 VGND.n5 9.3005
R150 VGND.n17 VGND.n16 9.3005
R151 VGND.n18 VGND.n4 9.3005
R152 VGND.n20 VGND.n19 9.3005
R153 VGND.n21 VGND.n3 9.3005
R154 VGND.n24 VGND.n23 9.3005
R155 VGND.n25 VGND.n1 9.3005
R156 VGND.n27 VGND.n26 9.3005
R157 VGND.n28 VGND.n0 9.3005
R158 VGND.n9 VGND.n7 6.95646
R159 VGND.n23 VGND.n22 6.02403
R160 VGND.n22 VGND.n21 5.27109
R161 VGND.n11 VGND.n7 0.593202
R162 VGND.n12 VGND.n11 0.122949
R163 VGND.n13 VGND.n12 0.122949
R164 VGND.n13 VGND.n5 0.122949
R165 VGND.n17 VGND.n5 0.122949
R166 VGND.n18 VGND.n17 0.122949
R167 VGND.n19 VGND.n18 0.122949
R168 VGND.n19 VGND.n3 0.122949
R169 VGND.n24 VGND.n3 0.122949
R170 VGND.n25 VGND.n24 0.122949
R171 VGND.n26 VGND.n25 0.122949
R172 VGND.n26 VGND.n0 0.122949
R173 VGND.n30 VGND.n0 0.122949
R174 VGND VGND.n30 0.0617245
R175 VNB.t2 VNB.t5 2436.75
R176 VNB.t6 VNB.t11 2286.61
R177 VNB.t4 VNB.t3 2240.42
R178 VNB VNB.t8 1466.67
R179 VNB.t7 VNB.t9 1316.54
R180 VNB.t9 VNB.t6 1281.89
R181 VNB.t1 VNB.t4 1224.15
R182 VNB.t3 VNB.t2 1154.86
R183 VNB.t0 VNB.t1 1154.86
R184 VNB.t10 VNB.t0 1154.86
R185 VNB.t11 VNB.t10 993.177
R186 VNB.t8 VNB.t7 993.177
R187 A2.n4 A2.t1 388.983
R188 A2.n0 A2.t2 250.596
R189 A2.n2 A2.t3 227.411
R190 A2.n0 A2.t0 192.8
R191 A2.n1 A2 163.055
R192 A2.n3 A2.n2 152
R193 A2.n2 A2.n1 40.9705
R194 A2.n5 A2 30.0805
R195 A2 A2.n4 19.8405
R196 A2.n1 A2.n0 13.858
R197 A2.n4 A2 4.07323
R198 A2.n3 A2 2.13383
R199 A2.n5 A2.n3 1.74595
R200 A2 A2.n5 0.6405
R201 a_564_74.n1 a_564_74.t7 187.696
R202 a_564_74.n2 a_564_74.t5 187.238
R203 a_564_74.n1 a_564_74.n0 185
R204 a_564_74.n2 a_564_74.t3 134.332
R205 a_564_74.n3 a_564_74.t2 131.755
R206 a_564_74.n5 a_564_74.n4 89.2338
R207 a_564_74.n4 a_564_74.n1 68.1392
R208 a_564_74.n4 a_564_74.n3 57.3741
R209 a_564_74.n3 a_564_74.n2 51.3983
R210 a_564_74.n0 a_564_74.t6 39.3755
R211 a_564_74.t1 a_564_74.n5 39.3755
R212 a_564_74.n5 a_564_74.t4 31.8755
R213 a_564_74.n0 a_564_74.t0 26.2505
R214 a_1234_392.n1 a_1234_392.n0 1224.59
R215 a_1234_392.n1 a_1234_392.t2 48.2655
R216 a_1234_392.t0 a_1234_392.n1 48.2655
R217 a_1234_392.n0 a_1234_392.t1 29.5505
R218 a_1234_392.n0 a_1234_392.t3 29.5505
R219 a_961_392.n1 a_961_392.t2 854.109
R220 a_961_392.n1 a_961_392.n0 585
R221 a_961_392.t1 a_961_392.n1 368.7
R222 a_961_392.n0 a_961_392.t0 29.5505
R223 a_961_392.n0 a_961_392.t3 29.5505
R224 A3.n1 A3.t2 301.324
R225 A3.n2 A3.t1 285.183
R226 A3.n2 A3.t0 162.565
R227 A3.n1 A3.n0 157.453
R228 A3 A3.n3 68.5584
R229 A3.n3 A3.n1 34.4317
R230 A3.n3 A3.n2 29.6871
R231 A1.n0 A1.t1 258.673
R232 A1.n2 A1.t2 247.428
R233 A1.n0 A1.t0 195.721
R234 A1 A1.n3 163.256
R235 A1.n2 A1.n1 139.488
R236 A1.n3 A1.n0 76.6823
R237 A1.n3 A1.n2 17.5278
C0 A1 VGND 0.028485f
C1 VPB B1 0.302875f
C2 A3 VPWR 0.011854f
C3 VPB B2 0.097103f
C4 A2 VPWR 0.019904f
C5 A3 B1 0.136509f
C6 A1 VPWR 0.02741f
C7 VGND VPWR 0.131115f
C8 A3 B2 0.025298f
C9 A2 B1 0.020406f
C10 A3 VPB 0.071963f
C11 VGND X 0.329869f
C12 A2 B2 2.03e-19
C13 A1 B1 0.001756f
C14 A2 VPB 0.103538f
C15 A1 B2 2.02e-20
C16 VGND B1 0.018485f
C17 A1 VPB 0.07936f
C18 VGND B2 0.013321f
C19 VPWR X 0.460245f
C20 VGND VPB 0.012886f
C21 A3 A2 0.089502f
C22 VPWR B1 0.169094f
C23 A3 A1 2.39e-20
C24 X B1 0.01004f
C25 VPWR B2 0.013561f
C26 A3 VGND 0.02875f
C27 A2 A1 0.181152f
C28 VPB VPWR 0.222186f
C29 A2 VGND 0.033215f
C30 VPB X 0.015376f
C31 B1 B2 0.175679f
C32 VGND VNB 0.980853f
C33 A1 VNB 0.263042f
C34 A2 VNB 0.286049f
C35 A3 VNB 0.220074f
C36 B2 VNB 0.257054f
C37 B1 VNB 0.326801f
C38 X VNB 0.058008f
C39 VPWR VNB 0.79106f
C40 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o32a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32a_2 VNB VPB VPWR VGND A1 A2 A3 B1 B2 X
X0 X.t3 a_83_264.t4 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t4 a_83_264.t5 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_83_264.t1 B2.t0 a_349_74.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.33855 pd=1.655 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 a_349_74.t4 B1.t0 a_83_264.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.33855 ps=1.655 w=0.74 l=0.15
X4 a_349_74.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 X.t0 a_83_264.t6 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3404 ps=2.4 w=0.74 l=0.15
X6 a_430_368.t1 A2.t0 a_346_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t2 A2.t1 a_349_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_346_368.t0 A1.t0 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2909 ps=1.67 w=1 l=0.15
X9 a_83_264.t2 A3.t1 a_430_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.195 ps=1.39 w=1 l=0.15
X10 VPWR.t1 a_83_264.t7 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2909 pd=1.67 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_652_368.t1 B2.t1 a_83_264.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 a_349_74.t1 A1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X13 VPWR.t3 B1.t1 a_652_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.21 ps=1.42 w=1 l=0.15
R0 a_83_264.n1 a_83_264.t4 327.224
R1 a_83_264.n4 a_83_264.n3 295.279
R2 a_83_264.n3 a_83_264.t7 258.233
R3 a_83_264.n4 a_83_264.n0 223.724
R4 a_83_264.n5 a_83_264.n4 200.472
R5 a_83_264.n2 a_83_264.t5 197.006
R6 a_83_264.n1 a_83_264.t6 186.374
R7 a_83_264.n0 a_83_264.t1 66.0842
R8 a_83_264.n2 a_83_264.n1 62.6605
R9 a_83_264.n0 a_83_264.t3 60.9872
R10 a_83_264.t0 a_83_264.n5 41.3705
R11 a_83_264.n5 a_83_264.t2 41.3705
R12 a_83_264.n3 a_83_264.n2 12.7593
R13 VPWR.n1 VPWR.t3 355.524
R14 VPWR.n3 VPWR.n2 297.404
R15 VPWR.n5 VPWR.t2 259.171
R16 VPWR.n2 VPWR.t0 53.8788
R17 VPWR.n2 VPWR.t1 50.7141
R18 VPWR.n5 VPWR.n4 26.7299
R19 VPWR.n4 VPWR.n3 25.977
R20 VPWR.n4 VPWR.n0 9.3005
R21 VPWR.n6 VPWR.n5 9.3005
R22 VPWR.n3 VPWR.n1 5.49975
R23 VPWR.n1 VPWR.n0 0.184181
R24 VPWR.n6 VPWR.n0 0.122949
R25 VPWR VPWR.n6 0.0617245
R26 X.n2 X 589.444
R27 X.n2 X.n0 585
R28 X.n3 X.n2 585
R29 X X.n1 163.876
R30 X.n2 X.t2 26.3844
R31 X.n2 X.t3 26.3844
R32 X.n1 X.t1 22.7032
R33 X.n1 X.t0 22.7032
R34 X X.n3 11.9116
R35 X X.n0 10.3116
R36 X X.n0 2.84494
R37 X.n3 X 1.24494
R38 VPB.t4 VPB.t3 357.527
R39 VPB.t0 VPB.t6 291.13
R40 VPB.t2 VPB.t0 291.13
R41 VPB.t1 VPB.t2 275.807
R42 VPB VPB.t5 257.93
R43 VPB.t5 VPB.t4 229.839
R44 VPB.t3 VPB.t1 214.517
R45 VGND.n4 VGND.n3 217.058
R46 VGND.n8 VGND.t3 140.049
R47 VGND.n2 VGND.n1 116.644
R48 VGND.n7 VGND.n6 36.1417
R49 VGND.n3 VGND.t0 34.0546
R50 VGND.n3 VGND.t2 34.0546
R51 VGND.n1 VGND.t1 34.0546
R52 VGND.n1 VGND.t4 34.0546
R53 VGND.n4 VGND.n2 16.5413
R54 VGND.n8 VGND.n7 13.5534
R55 VGND.n9 VGND.n8 9.3005
R56 VGND.n6 VGND.n5 9.3005
R57 VGND.n7 VGND.n0 9.3005
R58 VGND.n6 VGND.n2 1.50638
R59 VGND.n5 VGND.n4 1.00231
R60 VGND.n5 VGND.n0 0.122949
R61 VGND.n9 VGND.n0 0.122949
R62 VGND VGND.n9 0.0617245
R63 VNB.t1 VNB.t4 2459.84
R64 VNB VNB.t5 1547.51
R65 VNB.t3 VNB.t0 1316.54
R66 VNB.t6 VNB.t2 1316.54
R67 VNB.t0 VNB.t1 1154.86
R68 VNB.t2 VNB.t3 993.177
R69 VNB.t5 VNB.t6 993.177
R70 B2.n0 B2.t1 231.629
R71 B2.n0 B2.t0 220.113
R72 B2 B2.n0 159.591
R73 a_349_74.n1 a_349_74.t4 231.97
R74 a_349_74.n1 a_349_74.n0 165.535
R75 a_349_74.n2 a_349_74.n1 88.3339
R76 a_349_74.n2 a_349_74.t2 34.0546
R77 a_349_74.n0 a_349_74.t3 22.7032
R78 a_349_74.n0 a_349_74.t1 22.7032
R79 a_349_74.t0 a_349_74.n2 22.7032
R80 B1.n0 B1.t1 374.598
R81 B1.n1 B1.n0 193.627
R82 B1.n0 B1.t0 154.24
R83 B1 B1.n1 7.56414
R84 B1.n1 B1 6.78838
R85 A3.n0 A3.t1 231.629
R86 A3.n0 A3.t0 220.113
R87 A3 A3.n0 156.019
R88 A2.n0 A2.t0 231.629
R89 A2.n0 A2.t1 220.113
R90 A2 A2.n0 154.233
R91 a_346_368.t0 a_346_368.t1 53.1905
R92 a_430_368.t0 a_430_368.t1 76.8305
R93 A1.n0 A1.t0 226.15
R94 A1.n0 A1.t1 220.113
R95 A1 A1.n0 154.19
R96 a_652_368.t0 a_652_368.t1 82.7405
C0 B2 VGND 0.008037f
C1 X VGND 0.170467f
C2 VPB B2 0.036867f
C3 X A2 4.33e-19
C4 VPB X 0.006067f
C5 VPWR A3 0.007311f
C6 B2 B1 0.047479f
C7 X A1 0.001282f
C8 A3 VGND 0.01218f
C9 VPWR VGND 0.089679f
C10 A2 A3 0.083113f
C11 VPB A3 0.035177f
C12 VPWR A2 0.011045f
C13 VPB VPWR 0.163592f
C14 X B2 5.79e-20
C15 A2 VGND 0.013802f
C16 VPWR B1 0.094857f
C17 VPB VGND 0.012098f
C18 VPWR A1 0.016148f
C19 VPB A2 0.032908f
C20 B1 VGND 0.013521f
C21 A1 VGND 0.030399f
C22 A3 B2 0.079408f
C23 VPB B1 0.093383f
C24 VPWR B2 0.010674f
C25 X A3 2.14e-19
C26 A1 A2 0.094752f
C27 VPWR X 0.198204f
C28 VPB A1 0.037132f
C29 VGND VNB 0.627785f
C30 B1 VNB 0.267297f
C31 B2 VNB 0.114302f
C32 A3 VNB 0.104229f
C33 A2 VNB 0.102602f
C34 A1 VNB 0.104883f
C35 X VNB 0.035514f
C36 VPWR VNB 0.519409f
C37 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o211a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211a_1 VNB VPB VPWR VGND X C1 B1 A2 A1
X0 a_83_264.t2 C1.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.44 ps=1.88 w=1 l=0.15
X1 VPWR.t1 a_83_264.t4 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.6459 pd=2.38 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_257_136.t0 A2.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2352 pd=1.375 as=0.1632 ps=1.15 w=0.64 l=0.15
X3 a_83_264.t3 C1.t1 a_662_136.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2112 pd=1.94 as=0.104 ps=0.965 w=0.64 l=0.15
X4 VGND.t1 a_83_264.t5 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_662_136.t1 B1.t0 a_257_136.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.2352 ps=1.375 w=0.64 l=0.15
X6 VPWR.t2 B1.t1 a_83_264.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.44 pd=1.88 as=0.15 ps=1.3 w=1 l=0.15
X7 a_83_264.t1 A2.t1 a_398_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X8 a_398_392.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.6459 ps=2.38 w=1 l=0.15
X9 VGND.t2 A1.t1 a_257_136.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1632 pd=1.15 as=0.2112 ps=1.94 w=0.64 l=0.15
R0 C1.n0 C1.t0 231.629
R1 C1.n0 C1.t1 175.127
R2 C1 C1.n0 160.053
R3 VPWR.n11 VPWR.n10 292.5
R4 VPWR.n3 VPWR.n2 292.5
R5 VPWR.n9 VPWR.n8 292.5
R6 VPWR.n5 VPWR.n4 139.267
R7 VPWR.n9 VPWR.n2 89.6355
R8 VPWR.n10 VPWR.n9 89.6355
R9 VPWR.n4 VPWR.t2 80.1031
R10 VPWR.n4 VPWR.t3 80.1028
R11 VPWR.n10 VPWR.t1 37.541
R12 VPWR.n5 VPWR.n3 32.282
R13 VPWR.n2 VPWR.t0 29.5505
R14 VPWR.n7 VPWR.n6 9.3005
R15 VPWR.n1 VPWR.n0 9.3005
R16 VPWR.n12 VPWR.n11 8.17702
R17 VPWR.n8 VPWR.n7 5.15525
R18 VPWR.n11 VPWR.n1 4.86566
R19 VPWR.n8 VPWR.n1 0.40593
R20 VPWR.n6 VPWR.n5 0.362433
R21 VPWR VPWR.n12 0.160723
R22 VPWR.n12 VPWR.n0 0.147088
R23 VPWR.n6 VPWR.n0 0.122949
R24 VPWR.n7 VPWR.n3 0.116337
R25 a_83_264.n0 a_83_264.t2 318.577
R26 a_83_264.n0 a_83_264.t3 250.386
R27 a_83_264.n2 a_83_264.n1 245.262
R28 a_83_264.n1 a_83_264.t4 234.841
R29 a_83_264.n3 a_83_264.n2 201.906
R30 a_83_264.n1 a_83_264.t5 187.834
R31 a_83_264.t0 a_83_264.n3 29.5505
R32 a_83_264.n3 a_83_264.t1 29.5505
R33 a_83_264.n2 a_83_264.n0 12.1605
R34 VPB.t4 VPB.t0 720.162
R35 VPB.t1 VPB.t3 526.076
R36 VPB VPB.t4 257.93
R37 VPB.t2 VPB.t1 229.839
R38 VPB.t0 VPB.t2 214.517
R39 X.n1 X 589.444
R40 X.n1 X.n0 585
R41 X.n2 X.n1 585
R42 X X.t1 206.201
R43 X.n1 X.t0 26.3844
R44 X X.n2 11.9116
R45 X X.n0 10.3116
R46 X X.n0 2.84494
R47 X.n2 X 1.24494
R48 A2.t0 A2.t1 443.709
R49 A2 A2.t0 313.264
R50 VGND.n1 VGND.n0 217.827
R51 VGND.n1 VGND.t1 160.394
R52 VGND.n0 VGND.t0 59.063
R53 VGND.n0 VGND.t2 36.563
R54 VGND VGND.n1 0.322267
R55 a_257_136.n0 a_257_136.t2 296.688
R56 a_257_136.n0 a_257_136.t1 64.459
R57 a_257_136.t0 a_257_136.n0 58.489
R58 VNB.t2 VNB.t4 2760.1
R59 VNB.t0 VNB.t3 2044.09
R60 VNB.t4 VNB.t0 1524.41
R61 VNB VNB.t2 1143.31
R62 VNB.t3 VNB.t1 1097.11
R63 a_662_136.t0 a_662_136.t1 60.938
R64 B1.n0 B1.t1 263.762
R65 B1.n0 B1.t0 160.522
R66 B1 B1.n0 157.575
R67 a_398_392.t0 a_398_392.t1 53.1905
R68 A1.n0 A1.t0 228.129
R69 A1.n0 A1.t1 161.982
R70 A1 A1.n0 80.7578
C0 VPWR A2 0.014909f
C1 B1 VPB 0.064531f
C2 VGND A1 0.013404f
C3 B1 C1 0.054678f
C4 VGND X 0.105052f
C5 A1 A2 0.051382f
C6 X A2 2.45e-19
C7 VPWR A1 0.025048f
C8 X VPWR 0.10285f
C9 VGND VPB 0.009024f
C10 VGND C1 0.007153f
C11 VPB A2 0.030541f
C12 C1 A2 0.004528f
C13 VPWR VPB 0.114727f
C14 X A1 5.32e-19
C15 C1 VPWR 0.019209f
C16 VGND B1 0.00577f
C17 VPB A1 0.071305f
C18 B1 A2 0.051046f
C19 X VPB 0.014857f
C20 B1 VPWR 0.022147f
C21 C1 VPB 0.053305f
C22 VGND A2 0.209163f
C23 VGND VPWR 0.073719f
C24 VGND VNB 0.563366f
C25 VPWR VNB 0.418079f
C26 X VNB 0.11394f
C27 C1 VNB 0.131012f
C28 B1 VNB 0.119335f
C29 A2 VNB 0.186501f
C30 A1 VNB 0.128532f
C31 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o211a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211a_2 VNB VPB VPWR VGND A2 C1 A1 B1 X
X0 VGND.t2 A2.t0 a_195_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1751 pd=1.33 as=0.1332 ps=1.1 w=0.74 l=0.15
X1 VPWR.t2 a_27_368.t4 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_117_74.t0 C1.t0 a_27_368.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 X.t2 a_27_368.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3759 ps=1.84 w=1.12 l=0.15
X4 VPWR.t0 A1.t0 a_314_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3759 pd=1.84 as=0.16 ps=1.32 w=1 l=0.15
X5 a_195_74.t2 B1.t0 a_117_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X6 a_27_368.t0 B1.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.31 as=0.195 ps=1.39 w=1 l=0.15
X7 X.t1 a_27_368.t6 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1998 ps=2.02 w=0.74 l=0.15
X8 VPWR.t4 C1.t1 a_27_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.285 ps=2.57 w=1 l=0.15
X9 a_314_368.t1 A2.t1 a_27_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X10 VGND.t1 a_27_368.t7 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_195_74.t1 A1.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1751 ps=1.33 w=0.74 l=0.15
R0 A2.n0 A2.t1 231.629
R1 A2.n0 A2.t0 220.113
R2 A2 A2.n0 154.828
R3 a_195_74.n0 a_195_74.t1 493.135
R4 a_195_74.n0 a_195_74.t2 34.8654
R5 a_195_74.t0 a_195_74.n0 23.514
R6 VGND.n2 VGND.t0 279.909
R7 VGND.n5 VGND.n4 218.306
R8 VGND.n1 VGND.t1 173.418
R9 VGND.n4 VGND.t3 33.2437
R10 VGND.n4 VGND.t2 33.2437
R11 VGND.n3 VGND.n2 29.3652
R12 VGND.n5 VGND.n3 28.9887
R13 VGND.n3 VGND.n0 9.3005
R14 VGND.n6 VGND.n5 7.18735
R15 VGND.n2 VGND.n1 6.65317
R16 VGND.n1 VGND.n0 0.645433
R17 VGND VGND.n6 0.397267
R18 VGND.n6 VGND.n0 0.156565
R19 VNB.t3 VNB.t0 2217.32
R20 VNB.t2 VNB.t3 1293.44
R21 VNB.t5 VNB.t2 1177.95
R22 VNB VNB.t4 1177.95
R23 VNB.t0 VNB.t1 993.177
R24 VNB.t4 VNB.t5 900.788
R25 a_27_368.n3 a_27_368.t3 296.077
R26 a_27_368.n4 a_27_368.t2 281.884
R27 a_27_368.n0 a_27_368.t4 254.924
R28 a_27_368.n2 a_27_368.t5 231.972
R29 a_27_368.n5 a_27_368.n4 202.177
R30 a_27_368.n3 a_27_368.n2 157.562
R31 a_27_368.n0 a_27_368.t7 153.28
R32 a_27_368.n1 a_27_368.t6 142.994
R33 a_27_368.n4 a_27_368.n3 117.46
R34 a_27_368.n1 a_27_368.n0 43.8749
R35 a_27_368.t0 a_27_368.n5 31.5205
R36 a_27_368.n5 a_27_368.t1 29.5505
R37 a_27_368.n2 a_27_368.n1 26.5723
R38 X X.n0 245.106
R39 X.n2 X.n1 185
R40 X.n3 X.n2 185
R41 X.n0 X.t3 26.3844
R42 X.n0 X.t2 26.3844
R43 X.n2 X.t0 22.7032
R44 X.n2 X.t1 22.7032
R45 X.n3 X 16.3142
R46 X.n1 X 12.735
R47 X.n1 X 6.27501
R48 X X.n3 2.25932
R49 VPWR.n8 VPWR.n1 319.615
R50 VPWR.n4 VPWR.t2 265.825
R51 VPWR.n3 VPWR.n2 142.832
R52 VPWR.n2 VPWR.t1 69.8091
R53 VPWR.n2 VPWR.t0 61.9592
R54 VPWR.n1 VPWR.t4 39.4005
R55 VPWR.n1 VPWR.t3 37.4305
R56 VPWR.n7 VPWR.n6 36.1417
R57 VPWR.n6 VPWR.n3 25.977
R58 VPWR.n8 VPWR.n7 19.9534
R59 VPWR.n6 VPWR.n5 9.3005
R60 VPWR.n7 VPWR.n0 9.3005
R61 VPWR.n9 VPWR.n8 7.40447
R62 VPWR.n4 VPWR.n3 3.84167
R63 VPWR.n5 VPWR.n4 0.45173
R64 VPWR VPWR.n9 0.159703
R65 VPWR.n9 VPWR.n0 0.148095
R66 VPWR.n5 VPWR.n0 0.122949
R67 VPB.t0 VPB.t1 444.356
R68 VPB.t5 VPB.t3 275.807
R69 VPB VPB.t5 252.823
R70 VPB.t4 VPB.t0 240.054
R71 VPB.t3 VPB.t4 234.946
R72 VPB.t1 VPB.t2 229.839
R73 C1.n0 C1.t1 258.909
R74 C1.n0 C1.t0 170.81
R75 C1 C1.n0 158.788
R76 a_117_74.t0 a_117_74.t1 38.9194
R77 A1.n0 A1.t0 226.464
R78 A1.n0 A1.t1 214.95
R79 A1 A1.n0 154.522
R80 a_314_368.t0 a_314_368.t1 63.0405
R81 B1.n0 B1.t1 231.629
R82 B1.n0 B1.t0 220.113
R83 B1 B1.n0 161.674
C0 VPB X 0.005779f
C1 C1 VPWR 0.015541f
C2 A2 VGND 0.012104f
C3 C1 B1 0.086254f
C4 VPB A2 0.033006f
C5 VPWR VGND 0.077642f
C6 C1 A1 1.7e-19
C7 VPB VPWR 0.127928f
C8 B1 VGND 0.011561f
C9 A2 X 3.44e-19
C10 VPB B1 0.035389f
C11 VPWR X 0.195282f
C12 A1 VGND 0.011177f
C13 VPB A1 0.042449f
C14 A2 VPWR 0.012318f
C15 B1 X 9.71e-20
C16 C1 VGND 0.007751f
C17 VPB C1 0.04095f
C18 B1 A2 0.088537f
C19 A1 X 9.94e-19
C20 A2 A1 0.093918f
C21 B1 VPWR 0.018804f
C22 VPB VGND 0.008696f
C23 C1 A2 3.64e-19
C24 A1 VPWR 0.020251f
C25 X VGND 0.138504f
C26 VGND VNB 0.524466f
C27 X VNB 0.028311f
C28 VPWR VNB 0.429353f
C29 A1 VNB 0.116208f
C30 A2 VNB 0.10466f
C31 B1 VNB 0.109286f
C32 C1 VNB 0.166903f
C33 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o211a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211a_4 VNB VPB VPWR VGND A1 A2 B1 C1 X
X0 VPWR.t2 A1.t0 a_968_391.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.15 ps=1.3 w=1 l=0.15
X1 a_91_48.t5 C1.t0 a_597_125.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 a_510_125.t5 B1.t0 a_597_125.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1152 pd=1 as=0.112 ps=0.99 w=0.64 l=0.15
X3 VGND.t6 A1.t1 a_510_125.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0992 pd=0.95 as=0.1152 ps=1 w=0.64 l=0.15
X4 a_968_391.t3 A2.t0 a_91_48.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X5 X.t7 a_91_48.t8 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6 a_968_391.t1 A1.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2103 ps=1.435 w=1 l=0.15
X7 a_597_125.t2 C1.t1 a_91_48.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X8 a_510_125.t1 A1.t3 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.112 ps=0.99 w=0.64 l=0.15
X9 a_91_48.t0 A2.t1 a_968_391.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X10 VPWR.t8 a_91_48.t9 X.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_510_125.t0 A2.t2 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1072 pd=0.975 as=0.0992 ps=0.95 w=0.64 l=0.15
X12 VGND.t0 a_91_48.t10 X.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 X.t5 a_91_48.t11 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 VPWR.t0 B1.t1 a_91_48.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2103 pd=1.435 as=0.126 ps=1.14 w=0.84 l=0.15
X15 VGND.t7 A2.t3 a_510_125.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1072 ps=0.975 w=0.64 l=0.15
X16 a_91_48.t3 C1.t2 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1743 ps=1.255 w=0.84 l=0.15
X17 VPWR.t7 C1.t3 a_91_48.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1743 pd=1.255 as=0.126 ps=1.14 w=0.84 l=0.15
X18 X.t2 a_91_48.t12 VPWR.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X19 VPWR.t4 a_91_48.t13 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2789 pd=1.68 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_91_48.t6 B1.t2 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2789 ps=1.68 w=0.84 l=0.15
X21 X.t0 a_91_48.t14 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X22 a_597_125.t0 B1.t3 a_510_125.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1817 ps=1.85 w=0.64 l=0.15
X23 VGND.t2 a_91_48.t15 X.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A1.t3 A1.t1 907.768
R1 A1.t1 A1.t2 456.293
R2 A1.n0 A1.t0 235.644
R3 A1.n0 A1.t3 186.374
R4 A1 A1.n0 158.012
R5 a_968_391.n1 a_968_391.n0 569.886
R6 a_968_391.n0 a_968_391.t2 29.5505
R7 a_968_391.n0 a_968_391.t3 29.5505
R8 a_968_391.t0 a_968_391.n1 29.5505
R9 a_968_391.n1 a_968_391.t1 29.5505
R10 VPWR.n13 VPWR.n7 618.939
R11 VPWR.n22 VPWR.t9 352.519
R12 VPWR.n4 VPWR.n3 317.555
R13 VPWR.n20 VPWR.n2 317.341
R14 VPWR.n9 VPWR.n8 317.223
R15 VPWR.n10 VPWR.t2 269.32
R16 VPWR.n3 VPWR.t3 87.94
R17 VPWR.n8 VPWR.t0 58.0483
R18 VPWR.n7 VPWR.t6 50.4231
R19 VPWR.n7 VPWR.t7 46.9053
R20 VPWR.n8 VPWR.t1 36.7809
R21 VPWR.n15 VPWR.n14 36.1417
R22 VPWR.n13 VPWR.n12 35.7652
R23 VPWR.n3 VPWR.t4 35.4904
R24 VPWR.n2 VPWR.t5 35.1791
R25 VPWR.n2 VPWR.t8 35.1791
R26 VPWR.n19 VPWR.n4 32.7534
R27 VPWR.n21 VPWR.n20 29.7417
R28 VPWR.n22 VPWR.n21 20.7064
R29 VPWR.n12 VPWR.n9 18.4476
R30 VPWR.n20 VPWR.n19 17.6946
R31 VPWR.n15 VPWR.n4 14.6829
R32 VPWR.n14 VPWR.n13 11.6711
R33 VPWR.n12 VPWR.n11 9.3005
R34 VPWR.n13 VPWR.n6 9.3005
R35 VPWR.n14 VPWR.n5 9.3005
R36 VPWR.n16 VPWR.n15 9.3005
R37 VPWR.n17 VPWR.n4 9.3005
R38 VPWR.n19 VPWR.n18 9.3005
R39 VPWR.n20 VPWR.n1 9.3005
R40 VPWR.n21 VPWR.n0 9.3005
R41 VPWR.n23 VPWR.n22 9.3005
R42 VPWR.n10 VPWR.n9 7.38057
R43 VPWR.n11 VPWR.n10 0.167197
R44 VPWR.n11 VPWR.n6 0.122949
R45 VPWR.n6 VPWR.n5 0.122949
R46 VPWR.n16 VPWR.n5 0.122949
R47 VPWR.n17 VPWR.n16 0.122949
R48 VPWR.n18 VPWR.n17 0.122949
R49 VPWR.n18 VPWR.n1 0.122949
R50 VPWR.n1 VPWR.n0 0.122949
R51 VPWR.n23 VPWR.n0 0.122949
R52 VPWR VPWR.n23 0.0617245
R53 VPB.t5 VPB.t4 362.635
R54 VPB.t1 VPB.t2 298.791
R55 VPB.t8 VPB.t7 288.575
R56 VPB VPB.t10 283.469
R57 VPB.t9 VPB.t6 280.914
R58 VPB.t0 VPB.t11 255.376
R59 VPB.t11 VPB.t3 229.839
R60 VPB.t2 VPB.t0 229.839
R61 VPB.t7 VPB.t1 229.839
R62 VPB.t4 VPB.t8 229.839
R63 VPB.t6 VPB.t5 229.839
R64 VPB.t10 VPB.t9 229.839
R65 C1.n1 C1.t3 199.601
R66 C1.n0 C1.t1 166.757
R67 C1.n1 C1.t0 162.274
R68 C1.n0 C1.t2 159.06
R69 C1 C1.n2 155.88
R70 C1.n2 C1.n1 30.8261
R71 C1.n2 C1.n0 12.8912
R72 a_597_125.n1 a_597_125.n0 347.75
R73 a_597_125.n0 a_597_125.t2 39.3755
R74 a_597_125.n0 a_597_125.t1 26.2505
R75 a_597_125.n1 a_597_125.t3 26.2505
R76 a_597_125.t0 a_597_125.n1 26.2505
R77 a_91_48.n16 a_91_48.n14 390.68
R78 a_91_48.n13 a_91_48.n12 300.702
R79 a_91_48.n17 a_91_48.n16 300.702
R80 a_91_48.n16 a_91_48.n15 268.584
R81 a_91_48.n1 a_91_48.t13 256.995
R82 a_91_48.n9 a_91_48.t14 240.197
R83 a_91_48.n2 a_91_48.t9 240.197
R84 a_91_48.n4 a_91_48.t12 240.197
R85 a_91_48.n4 a_91_48.t11 183.81
R86 a_91_48.n8 a_91_48.t8 179.947
R87 a_91_48.n3 a_91_48.t10 179.947
R88 a_91_48.n1 a_91_48.t15 179.947
R89 a_91_48.n6 a_91_48.n5 165.189
R90 a_91_48.n7 a_91_48.n6 152
R91 a_91_48.n8 a_91_48.n0 152
R92 a_91_48.n11 a_91_48.n10 152
R93 a_91_48.n13 a_91_48.n11 82.9039
R94 a_91_48.n16 a_91_48.n13 51.577
R95 a_91_48.n8 a_91_48.n7 49.6611
R96 a_91_48.n14 a_91_48.t0 39.4005
R97 a_91_48.n10 a_91_48.n9 35.7853
R98 a_91_48.n12 a_91_48.t2 35.1791
R99 a_91_48.n12 a_91_48.t6 35.1791
R100 a_91_48.n17 a_91_48.t1 35.1791
R101 a_91_48.t3 a_91_48.n17 35.1791
R102 a_91_48.n5 a_91_48.n4 32.8641
R103 a_91_48.n14 a_91_48.t7 29.5505
R104 a_91_48.n5 a_91_48.n3 26.2914
R105 a_91_48.n15 a_91_48.t4 26.2505
R106 a_91_48.n15 a_91_48.t5 26.2505
R107 a_91_48.n7 a_91_48.n2 16.7975
R108 a_91_48.n9 a_91_48.n8 13.8763
R109 a_91_48.n11 a_91_48.n0 13.1884
R110 a_91_48.n6 a_91_48.n0 13.1884
R111 a_91_48.n10 a_91_48.n1 13.146
R112 a_91_48.n3 a_91_48.n2 6.57323
R113 VNB.t0 VNB.t4 2355.91
R114 VNB VNB.t1 1224.15
R115 VNB.t6 VNB.t8 1177.95
R116 VNB.t11 VNB.t7 1154.86
R117 VNB.t9 VNB.t6 1154.86
R118 VNB.t2 VNB.t3 1154.86
R119 VNB.t5 VNB.t11 1120.21
R120 VNB.t8 VNB.t5 1062.47
R121 VNB.t10 VNB.t9 993.177
R122 VNB.t4 VNB.t10 993.177
R123 VNB.t3 VNB.t0 993.177
R124 VNB.t1 VNB.t2 993.177
R125 B1.n1 B1.t0 1201.88
R126 B1.t0 B1.t1 418.774
R127 B1.n0 B1.t2 189.855
R128 B1.n0 B1.t3 164.637
R129 B1 B1.n1 156.268
R130 B1.n1 B1.n0 5.10403
R131 a_510_125.n4 a_510_125.n3 300.627
R132 a_510_125.n1 a_510_125.t1 186.352
R133 a_510_125.n1 a_510_125.n0 100.812
R134 a_510_125.n3 a_510_125.n2 88.228
R135 a_510_125.n3 a_510_125.n1 64.7165
R136 a_510_125.n2 a_510_125.t2 41.2505
R137 a_510_125.n0 a_510_125.t0 36.563
R138 a_510_125.n2 a_510_125.t5 26.2505
R139 a_510_125.n0 a_510_125.t3 26.2505
R140 a_510_125.n5 a_510_125.n4 2.11673
R141 a_510_125.n4 a_510_125.t4 2.06136
R142 VGND.n23 VGND.t1 285.764
R143 VGND.n7 VGND.n6 220.421
R144 VGND.n9 VGND.n8 213.569
R145 VGND.n21 VGND.n2 207.109
R146 VGND.n17 VGND.t2 164.077
R147 VGND.n6 VGND.t5 39.3755
R148 VGND.n11 VGND.n10 36.1417
R149 VGND.n11 VGND.n4 36.1417
R150 VGND.n15 VGND.n4 36.1417
R151 VGND.n16 VGND.n15 36.1417
R152 VGND.n2 VGND.t3 34.0546
R153 VGND.n8 VGND.t4 30.938
R154 VGND.n17 VGND.n16 27.8593
R155 VGND.n8 VGND.t6 27.188
R156 VGND.n6 VGND.t7 26.2505
R157 VGND.n21 VGND.n1 25.6005
R158 VGND.n23 VGND.n22 24.0946
R159 VGND.n2 VGND.t0 22.7032
R160 VGND.n22 VGND.n21 21.8358
R161 VGND.n10 VGND.n9 20.3299
R162 VGND.n17 VGND.n1 19.577
R163 VGND.n24 VGND.n23 9.3005
R164 VGND.n22 VGND.n0 9.3005
R165 VGND.n21 VGND.n20 9.3005
R166 VGND.n19 VGND.n1 9.3005
R167 VGND.n18 VGND.n17 9.3005
R168 VGND.n10 VGND.n5 9.3005
R169 VGND.n12 VGND.n11 9.3005
R170 VGND.n13 VGND.n4 9.3005
R171 VGND.n15 VGND.n14 9.3005
R172 VGND.n16 VGND.n3 9.3005
R173 VGND.n9 VGND.n7 6.79986
R174 VGND.n7 VGND.n5 0.580041
R175 VGND.n12 VGND.n5 0.122949
R176 VGND.n13 VGND.n12 0.122949
R177 VGND.n14 VGND.n13 0.122949
R178 VGND.n14 VGND.n3 0.122949
R179 VGND.n18 VGND.n3 0.122949
R180 VGND.n19 VGND.n18 0.122949
R181 VGND.n20 VGND.n19 0.122949
R182 VGND.n20 VGND.n0 0.122949
R183 VGND.n24 VGND.n0 0.122949
R184 VGND VGND.n24 0.0617245
R185 A2.n2 A2.t1 214.56
R186 A2.n0 A2.t0 211.544
R187 A2.n0 A2.t3 163.734
R188 A2.n2 A2.t2 162.274
R189 A2 A2.n1 161.115
R190 A2.n4 A2.n3 152
R191 A2.n3 A2.n1 49.6611
R192 A2.n4 A2 14.546
R193 A2.n3 A2.n2 13.146
R194 A2.n1 A2.n0 6.57323
R195 A2 A2.n4 4.07323
R196 X.n2 X.n0 258.046
R197 X.n2 X.n1 207.6
R198 X.n5 X.n3 153.22
R199 X.n5 X.n4 102.019
R200 X X.n2 36.5509
R201 X.n0 X.t1 26.3844
R202 X.n0 X.t0 26.3844
R203 X.n1 X.t3 26.3844
R204 X.n1 X.t2 26.3844
R205 X X.n5 26.1243
R206 X.n3 X.t4 22.7032
R207 X.n3 X.t7 22.7032
R208 X.n4 X.t6 22.7032
R209 X.n4 X.t5 22.7032
C0 VGND X 0.311651f
C1 VPB X 0.015799f
C2 VGND A1 0.091405f
C3 VPWR X 0.426209f
C4 VPB A1 0.084696f
C5 VPWR A1 0.070581f
C6 X A1 2.51e-21
C7 A2 B1 0.001148f
C8 B1 C1 0.144486f
C9 A2 VGND 0.024997f
C10 A2 VPB 0.079813f
C11 B1 VGND 0.085304f
C12 A2 VPWR 0.012148f
C13 B1 VPB 0.103991f
C14 C1 VGND 0.00745f
C15 B1 VPWR 0.029492f
C16 C1 VPB 0.083001f
C17 VGND VPB 0.012178f
C18 B1 X 0.005212f
C19 A2 A1 0.157742f
C20 C1 VPWR 0.030159f
C21 C1 X 7.6e-21
C22 B1 A1 0.051883f
C23 VGND VPWR 0.112013f
C24 VPB VPWR 0.20723f
C25 VGND VNB 0.806935f
C26 C1 VNB 0.160888f
C27 B1 VNB 0.540103f
C28 A2 VNB 0.167649f
C29 A1 VNB 0.4207f
C30 X VNB 0.07194f
C31 VPWR VNB 0.685076f
C32 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211ai_1 VNB VPB VPWR VGND B1 Y C1 A2 A1
X0 a_116_368.t0 A1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t0 A1.t1 a_31_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t1 B1.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3192 ps=1.69 w=1.12 l=0.15
X3 Y.t2 C1.t0 a_311_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.4588 pd=2.72 as=0.1554 ps=1.16 w=0.74 l=0.15
X4 Y.t3 A2.t0 a_116_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=1.69 as=0.1512 ps=1.39 w=1.12 l=0.15
X5 a_311_74.t0 B1.t1 a_31_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.11655 ps=1.055 w=0.74 l=0.15
X6 a_31_74.t2 A2.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 Y.t0 C1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
R0 A1.n0 A1.t0 256.428
R1 A1.n0 A1.t1 196.178
R2 A1 A1.n0 155.067
R3 VPWR.n1 VPWR.n0 323.759
R4 VPWR.n1 VPWR.t2 264.69
R5 VPWR.n0 VPWR.t0 35.1791
R6 VPWR.n0 VPWR.t1 26.3844
R7 VPWR VPWR.n1 0.131264
R8 a_116_368.t0 a_116_368.t1 47.4916
R9 VPB.t3 VPB.t1 367.743
R10 VPB VPB.t2 257.93
R11 VPB.t1 VPB.t0 255.376
R12 VPB.t2 VPB.t3 214.517
R13 a_31_74.t0 a_31_74.n0 300.423
R14 a_31_74.n0 a_31_74.t1 28.3789
R15 a_31_74.n0 a_31_74.t2 22.7032
R16 VGND VGND.n0 214.809
R17 VGND.n0 VGND.t0 34.0546
R18 VGND.n0 VGND.t1 22.7032
R19 VNB.t2 VNB.t0 1316.54
R20 VNB VNB.t1 1189.5
R21 VNB.t1 VNB.t3 1154.86
R22 VNB.t3 VNB.t2 1074.02
R23 B1.n0 B1.t0 264.298
R24 B1.n0 B1.t1 204.048
R25 B1.n1 B1.n0 157.416
R26 B1 B1.n1 5.0092
R27 B1.n1 B1 2.95435
R28 Y.n1 Y.n0 264.07
R29 Y.n1 Y.t0 228.797
R30 Y.n2 Y.t2 96.5208
R31 Y Y.n1 62.516
R32 Y.n0 Y.t3 51.0094
R33 Y.n0 Y.t1 49.2505
R34 Y Y.n2 8.08471
R35 Y.n2 Y 2.69524
R36 C1.n0 C1.t1 285.719
R37 C1.n0 C1.t0 178.34
R38 C1 C1.n0 158.788
R39 a_311_74.t0 a_311_74.t1 68.1086
R40 A2.n0 A2.t0 264.298
R41 A2.n0 A2.t1 204.048
R42 A2.n1 A2.n0 187.553
R43 A2.n1 A2 17.8092
R44 A2.n1 A2 13.6005
R45 A2 A2.n1 2.78311
C0 VPB A2 0.03967f
C1 VPWR Y 0.28234f
C2 VGND VPB 0.006311f
C3 A1 VPWR 0.046395f
C4 A2 C1 2.6e-19
C5 VPB Y 0.033323f
C6 VGND C1 0.010283f
C7 VPB A1 0.042712f
C8 C1 Y 0.103266f
C9 A2 B1 0.071475f
C10 VPB VPWR 0.089663f
C11 VGND B1 0.035099f
C12 B1 Y 0.097668f
C13 C1 VPWR 0.015476f
C14 VPB C1 0.035208f
C15 A1 B1 3.24e-19
C16 VGND A2 0.018842f
C17 A2 Y 0.087554f
C18 B1 VPWR 0.018599f
C19 VGND Y 0.07152f
C20 A1 A2 0.111403f
C21 VPB B1 0.034114f
C22 VGND A1 0.016848f
C23 A1 Y 3.56e-19
C24 A2 VPWR 0.103971f
C25 B1 C1 0.084012f
C26 VGND VPWR 0.046737f
C27 VGND VNB 0.379002f
C28 Y VNB 0.118626f
C29 VPWR VNB 0.347109f
C30 C1 VNB 0.138028f
C31 B1 VNB 0.116707f
C32 A2 VNB 0.112196f
C33 A1 VNB 0.170075f
C34 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o211ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211ai_2 VNB VPB VPWR VGND C1 B1 A2 A1 Y
X0 Y.t4 C1.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_303_84.t5 B1.t0 a_30_84.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X2 VPWR.t4 A1.t0 a_505_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_505_368.t3 A2.t0 Y.t7 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_30_84.t1 C1.t1 Y.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 Y.t2 A2.t1 a_505_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 VGND.t1 A1.t1 a_303_84.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2294 pd=2.1 as=0.12025 ps=1.065 w=0.74 l=0.15
X7 a_303_84.t2 A1.t2 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.10545 ps=1.025 w=0.74 l=0.15
X8 VPWR.t1 B1.t1 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_303_84.t0 A2.t2 VGND.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 Y.t0 B1.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t2 C1.t2 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VGND.t2 A2.t3 a_303_84.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_30_84.t2 B1.t3 a_303_84.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2183 pd=2.07 as=0.1295 ps=1.09 w=0.74 l=0.15
X14 Y.t5 C1.t3 a_30_84.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 a_505_368.t1 A1.t3 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
R0 C1.n0 C1.t2 247.944
R1 C1.n2 C1.t0 246.446
R2 C1.n1 C1.t3 196.608
R3 C1.n0 C1.t1 179.947
R4 C1 C1.n2 158.847
R5 C1.n1 C1.n0 54.2255
R6 C1.n2 C1.n1 2.97581
R7 VPWR.n5 VPWR.t1 349.789
R8 VPWR.n2 VPWR.n1 331.5
R9 VPWR.n4 VPWR.n3 323.38
R10 VPWR.n11 VPWR.t3 257.433
R11 VPWR.n10 VPWR.n9 36.1417
R12 VPWR.n6 VPWR.n2 35.3887
R13 VPWR.n3 VPWR.t5 35.1791
R14 VPWR.n1 VPWR.t0 26.3844
R15 VPWR.n1 VPWR.t2 26.3844
R16 VPWR.n3 VPWR.t4 26.3844
R17 VPWR.n6 VPWR.n5 25.977
R18 VPWR.n11 VPWR.n10 24.4711
R19 VPWR.n7 VPWR.n6 9.3005
R20 VPWR.n9 VPWR.n8 9.3005
R21 VPWR.n10 VPWR.n0 9.3005
R22 VPWR.n12 VPWR.n11 9.3005
R23 VPWR.n5 VPWR.n4 7.31736
R24 VPWR.n9 VPWR.n2 0.753441
R25 VPWR.n7 VPWR.n4 0.167001
R26 VPWR.n8 VPWR.n7 0.122949
R27 VPWR.n8 VPWR.n0 0.122949
R28 VPWR.n12 VPWR.n0 0.122949
R29 VPWR VPWR.n12 0.0617245
R30 Y Y.n0 589.85
R31 Y.n7 Y.n0 585
R32 Y.n6 Y.n0 585
R33 Y.n3 Y.n1 385.033
R34 Y.n3 Y.n2 205.487
R35 Y.n5 Y.n4 162.719
R36 Y.n5 Y.n3 42.9181
R37 Y.n0 Y.t3 26.3844
R38 Y.n0 Y.t4 26.3844
R39 Y.n1 Y.t7 26.3844
R40 Y.n1 Y.t2 26.3844
R41 Y.n2 Y.t1 26.3844
R42 Y.n2 Y.t0 26.3844
R43 Y.n4 Y.t6 22.7032
R44 Y.n4 Y.t5 22.7032
R45 Y Y.n7 8.72777
R46 Y Y.n6 7.95202
R47 Y.n7 Y 5.62474
R48 Y.n6 Y.n5 3.10353
R49 VPB.t1 VPB.t2 515.861
R50 VPB VPB.t4 273.253
R51 VPB.t5 VPB.t7 255.376
R52 VPB.t6 VPB.t5 229.839
R53 VPB.t2 VPB.t6 229.839
R54 VPB.t0 VPB.t1 229.839
R55 VPB.t3 VPB.t0 229.839
R56 VPB.t4 VPB.t3 229.839
R57 B1.n2 B1.t2 227.538
R58 B1.n0 B1.t1 226.809
R59 B1.n0 B1.t3 187.981
R60 B1.n2 B1.t0 179.947
R61 B1 B1.n1 159.591
R62 B1.n4 B1.n3 152
R63 B1.n3 B1.n1 49.6611
R64 B1.n4 B1 11.7586
R65 B1.n3 B1.n2 10.2247
R66 B1.n1 B1.n0 5.11262
R67 B1 B1.n4 2.53073
R68 a_30_84.n0 a_30_84.t2 301.721
R69 a_30_84.n0 a_30_84.t0 212.569
R70 a_30_84.n1 a_30_84.n0 95.184
R71 a_30_84.t1 a_30_84.n1 34.0546
R72 a_30_84.n1 a_30_84.t3 22.7032
R73 a_303_84.n3 a_303_84.n2 287.791
R74 a_303_84.n2 a_303_84.n1 162.905
R75 a_303_84.n2 a_303_84.n0 101.391
R76 a_303_84.n3 a_303_84.t5 34.0546
R77 a_303_84.n1 a_303_84.t3 30.0005
R78 a_303_84.n1 a_303_84.t2 22.7032
R79 a_303_84.n0 a_303_84.t1 22.7032
R80 a_303_84.n0 a_303_84.t0 22.7032
R81 a_303_84.t4 a_303_84.n3 22.7032
R82 VNB.t6 VNB.t0 2309.71
R83 VNB VNB.t1 1177.95
R84 VNB.t7 VNB.t6 1154.86
R85 VNB.t2 VNB.t7 1154.86
R86 VNB.t4 VNB.t5 1097.11
R87 VNB.t3 VNB.t4 1004.72
R88 VNB.t0 VNB.t3 993.177
R89 VNB.t1 VNB.t2 993.177
R90 A1.n1 A1.t0 236.219
R91 A1.n2 A1.t3 234.841
R92 A1.n2 A1.n0 185.573
R93 A1.n1 A1.t2 179.947
R94 A1.n3 A1.t1 179.947
R95 A1 A1.n4 80.0331
R96 A1.n4 A1.n3 31.9471
R97 A1.n4 A1.n1 27.4463
R98 A1.n0 A1 4.26717
R99 A1 A1.n0 2.13383
R100 A1.n3 A1.n2 2.06621
R101 a_505_368.n0 a_505_368.t0 430.075
R102 a_505_368.n0 a_505_368.t1 321.748
R103 a_505_368.n1 a_505_368.n0 181.951
R104 a_505_368.t2 a_505_368.n1 26.3844
R105 a_505_368.n1 a_505_368.t3 26.3844
R106 A2.n1 A2.t0 234.841
R107 A2.n4 A2.t1 234.841
R108 A2.n5 A2.n4 195.089
R109 A2.n1 A2.t3 190.025
R110 A2.n3 A2.t2 186.374
R111 A2.n2 A2 159.311
R112 A2.n3 A2.n0 152
R113 A2.n3 A2.n2 49.6611
R114 A2.n2 A2.n1 9.49444
R115 A2.n5 A2.n0 9.46137
R116 A2.n4 A2.n3 6.57323
R117 A2 A2.n0 2.64398
R118 A2 A2.n5 1.25267
R119 VGND.n5 VGND.t3 232.139
R120 VGND.n3 VGND.n2 209.436
R121 VGND.n1 VGND.t1 159.315
R122 VGND.n2 VGND.t0 23.514
R123 VGND.n2 VGND.t2 22.7032
R124 VGND.n4 VGND.n3 22.5887
R125 VGND.n5 VGND.n4 17.3181
R126 VGND.n4 VGND.n0 9.3005
R127 VGND.n6 VGND.n5 7.43989
R128 VGND.n3 VGND.n1 6.65145
R129 VGND.n1 VGND.n0 0.677131
R130 VGND VGND.n6 0.647175
R131 VGND.n6 VGND.n0 0.152785
C0 Y VGND 0.013378f
C1 Y A2 0.097466f
C2 VGND B1 0.011482f
C3 B1 A2 0.043589f
C4 VGND A2 0.037628f
C5 A1 VPB 0.082348f
C6 A1 VPWR 0.043232f
C7 VPWR VPB 0.145309f
C8 A1 C1 2.57e-20
C9 VPB C1 0.075512f
C10 A1 Y 0.001095f
C11 A1 B1 1.01e-19
C12 Y VPB 0.021213f
C13 VPWR C1 0.060955f
C14 VPB B1 0.069106f
C15 VPWR Y 0.396348f
C16 A1 VGND 0.075636f
C17 VPWR B1 0.031461f
C18 A1 A2 0.082607f
C19 VGND VPB 0.009102f
C20 Y C1 0.116138f
C21 C1 B1 0.057926f
C22 VPB A2 0.087168f
C23 VPWR VGND 0.078553f
C24 VGND C1 0.013168f
C25 VPWR A2 0.014049f
C26 Y B1 0.15174f
C27 C1 A2 2.65e-20
C28 VGND VNB 0.60489f
C29 Y VNB 0.021204f
C30 VPWR VNB 0.501806f
C31 A1 VNB 0.283705f
C32 A2 VNB 0.242145f
C33 B1 VNB 0.202999f
C34 C1 VNB 0.252213f
C35 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o211ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211ai_4 VNB VPB VPWR VGND A1 A2 B1 C1 Y
X0 VPWR.t5 C1.t0 Y.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.9688 pd=3.97 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_30_368.t4 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t6 B1.t0 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.2184 ps=1.51 w=1.12 l=0.15
X3 a_27_74.t11 B1.t1 a_834_74.t7 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2016 ps=1.48 w=1.12 l=0.15
X5 a_27_74.t6 A2.t0 VGND.t7 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VPWR.t1 A1.t1 a_30_368.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_30_368.t2 A1.t2 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Y.t8 C1.t1 a_834_74.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_27_74.t5 A1.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 VGND.t6 A2.t1 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VGND.t2 A1.t4 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 a_27_74.t10 B1.t2 a_834_74.t6 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 Y.t7 C1.t2 a_834_74.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 a_30_368.t0 A2.t2 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X15 VGND.t5 A2.t3 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_834_74.t1 C1.t3 Y.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t1 A1.t5 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_834_74.t5 B1.t3 a_27_74.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_834_74.t0 C1.t4 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_834_74.t4 B1.t4 a_27_74.t8 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VPWR.t2 A1.t6 a_30_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X22 Y.t2 A2.t4 a_30_368.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_30_368.t6 A2.t5 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_27_74.t2 A1.t7 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X25 Y.t4 A2.t6 a_30_368.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X26 Y.t0 B1.t5 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.3304 ps=2.83 w=1.12 l=0.15
X27 a_27_74.t1 A2.t7 VGND.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.111 ps=1.04 w=0.74 l=0.15
R0 C1.n0 C1.t3 318.12
R1 C1.n4 C1.n3 249.447
R2 C1.n2 C1.t0 226.809
R3 C1.n7 C1.t2 179.947
R4 C1.n0 C1.t1 179.947
R5 C1.n1 C1.t4 179.947
R6 C1.n9 C1.n8 152
R7 C1.n7 C1.n6 152
R8 C1.n5 C1.n4 152
R9 C1.n1 C1.n0 125.028
R10 C1.n8 C1.n7 49.6611
R11 C1.n4 C1.n2 43.0884
R12 C1.n8 C1.n1 13.146
R13 C1.n6 C1.n5 10.1214
R14 C1.n9 C1 9.52608
R15 C1.n7 C1.n2 6.57323
R16 C1 C1.n9 4.76329
R17 C1.n5 C1 3.57259
R18 C1.n6 C1 0.595849
R19 Y.n2 Y.n0 346.634
R20 Y.n2 Y.n1 299.95
R21 Y.n9 Y.n7 252.766
R22 Y.n5 Y.t5 231.87
R23 Y.n4 Y.n3 205.487
R24 Y.n9 Y.n8 199.934
R25 Y.n4 Y.n2 92.6123
R26 Y.n6 Y.n5 82.4476
R27 Y.n5 Y.n4 50.4476
R28 Y.n1 Y.t2 35.1791
R29 Y.n3 Y.t0 35.1791
R30 Y.n3 Y.t10 33.4201
R31 Y Y.n9 32.9292
R32 Y.n0 Y.t3 26.3844
R33 Y.n0 Y.t4 26.3844
R34 Y.n1 Y.t1 26.3844
R35 Y.n8 Y.t6 22.7032
R36 Y.n8 Y.t8 22.7032
R37 Y.n7 Y.t9 22.7032
R38 Y.n7 Y.t7 22.7032
R39 Y.n6 Y 6.84887
R40 Y Y.n6 1.62438
R41 VPWR.n8 VPWR.t6 344.825
R42 VPWR.n10 VPWR.t3 343.067
R43 VPWR.n21 VPWR.n2 331.5
R44 VPWR.n23 VPWR.n1 331.5
R45 VPWR.n7 VPWR.t5 206.565
R46 VPWR.n14 VPWR.n5 36.1417
R47 VPWR.n15 VPWR.n14 36.1417
R48 VPWR.n16 VPWR.n15 36.1417
R49 VPWR.n16 VPWR.n3 36.1417
R50 VPWR.n20 VPWR.n3 36.1417
R51 VPWR.n23 VPWR.n22 34.2593
R52 VPWR.n22 VPWR.n21 33.5064
R53 VPWR.n9 VPWR.n8 30.1181
R54 VPWR.n10 VPWR.n5 27.1064
R55 VPWR.n1 VPWR.t4 26.3844
R56 VPWR.n1 VPWR.t2 26.3844
R57 VPWR.n2 VPWR.t0 26.3844
R58 VPWR.n2 VPWR.t1 26.3844
R59 VPWR.n10 VPWR.n9 20.3299
R60 VPWR.n24 VPWR.n23 9.58614
R61 VPWR.n9 VPWR.n6 9.3005
R62 VPWR.n11 VPWR.n10 9.3005
R63 VPWR.n12 VPWR.n5 9.3005
R64 VPWR.n14 VPWR.n13 9.3005
R65 VPWR.n15 VPWR.n4 9.3005
R66 VPWR.n17 VPWR.n16 9.3005
R67 VPWR.n18 VPWR.n3 9.3005
R68 VPWR.n20 VPWR.n19 9.3005
R69 VPWR.n22 VPWR.n0 9.3005
R70 VPWR.n8 VPWR.n7 6.52323
R71 VPWR.n21 VPWR.n20 2.63579
R72 VPWR.n7 VPWR.n6 0.370393
R73 VPWR VPWR.n24 0.163644
R74 VPWR.n24 VPWR.n0 0.144205
R75 VPWR.n11 VPWR.n6 0.122949
R76 VPWR.n12 VPWR.n11 0.122949
R77 VPWR.n13 VPWR.n12 0.122949
R78 VPWR.n13 VPWR.n4 0.122949
R79 VPWR.n17 VPWR.n4 0.122949
R80 VPWR.n18 VPWR.n17 0.122949
R81 VPWR.n19 VPWR.n18 0.122949
R82 VPWR.n19 VPWR.n0 0.122949
R83 VPB.t4 VPB.t3 541.399
R84 VPB.t10 VPB.t9 490.324
R85 VPB.t3 VPB.t10 275.807
R86 VPB VPB.t2 265.591
R87 VPB.t6 VPB.t4 255.376
R88 VPB.t0 VPB.t8 255.376
R89 VPB.t7 VPB.t6 229.839
R90 VPB.t8 VPB.t7 229.839
R91 VPB.t1 VPB.t0 229.839
R92 VPB.t5 VPB.t1 229.839
R93 VPB.t2 VPB.t5 229.839
R94 A1.n0 A1.t0 226.809
R95 A1.n3 A1.t1 226.809
R96 A1.n9 A1.t2 226.809
R97 A1.n4 A1.t6 226.809
R98 A1.n0 A1.t3 204.048
R99 A1.n4 A1.t4 199.666
R100 A1.n10 A1.t7 196.013
R101 A1.n2 A1.t5 196.013
R102 A1 A1.n1 152.298
R103 A1.n12 A1.n11 152
R104 A1.n8 A1.n7 152
R105 A1.n6 A1.n5 152
R106 A1.n8 A1.n5 49.6611
R107 A1.n11 A1.n10 39.4369
R108 A1.n1 A1.n0 38.7066
R109 A1.n2 A1.n1 26.2914
R110 A1.n11 A1.n3 22.6399
R111 A1.n6 A1 12.8005
R112 A1 A1.n12 9.82376
R113 A1.n5 A1.n4 9.49444
R114 A1.n7 A1 8.63306
R115 A1.n9 A1.n8 6.57323
R116 A1.n7 A1 5.65631
R117 A1.n12 A1 4.46562
R118 A1.n10 A1.n9 3.65202
R119 A1 A1.n6 1.48887
R120 A1.n3 A1.n2 0.730803
R121 a_30_368.n1 a_30_368.t0 389.12
R122 a_30_368.n1 a_30_368.n0 305.998
R123 a_30_368.n3 a_30_368.t1 274.788
R124 a_30_368.n3 a_30_368.n2 205.487
R125 a_30_368.n5 a_30_368.n4 189.115
R126 a_30_368.n4 a_30_368.n1 72.7633
R127 a_30_368.n4 a_30_368.n3 59.2899
R128 a_30_368.n5 a_30_368.t7 35.1791
R129 a_30_368.n2 a_30_368.t3 26.3844
R130 a_30_368.n2 a_30_368.t2 26.3844
R131 a_30_368.n0 a_30_368.t5 26.3844
R132 a_30_368.n0 a_30_368.t6 26.3844
R133 a_30_368.t4 a_30_368.n5 26.3844
R134 B1.n4 B1.t4 281.168
R135 B1.n2 B1.t0 226.809
R136 B1.n6 B1.t5 226.809
R137 B1.n2 B1.t1 198.204
R138 B1.n7 B1.t3 196.013
R139 B1.n3 B1.n0 152
R140 B1 B1.n7 152
R141 B1.n5 B1.n1 152
R142 B1.n4 B1.t2 142.994
R143 B1.n7 B1.n3 49.6611
R144 B1.n6 B1.n5 31.4035
R145 B1.n7 B1.n6 18.2581
R146 B1.n5 B1.n4 17.966
R147 B1.n3 B1.n2 10.955
R148 B1 B1.n0 10.1214
R149 B1 B1.n1 10.1214
R150 B1.n0 B1 4.16794
R151 B1.n1 B1 4.16794
R152 a_834_74.n2 a_834_74.n0 212.869
R153 a_834_74.n4 a_834_74.t1 196.345
R154 a_834_74.n2 a_834_74.n1 185
R155 a_834_74.n5 a_834_74.n4 185
R156 a_834_74.n3 a_834_74.t2 152.828
R157 a_834_74.n3 a_834_74.n2 58.4726
R158 a_834_74.n4 a_834_74.n3 43.5166
R159 a_834_74.n0 a_834_74.t6 22.7032
R160 a_834_74.n0 a_834_74.t4 22.7032
R161 a_834_74.n1 a_834_74.t7 22.7032
R162 a_834_74.n1 a_834_74.t5 22.7032
R163 a_834_74.t3 a_834_74.n5 22.7032
R164 a_834_74.n5 a_834_74.t0 22.7032
R165 a_27_74.n8 a_27_74.t11 262.591
R166 a_27_74.n4 a_27_74.t4 200.344
R167 a_27_74.n9 a_27_74.n8 185
R168 a_27_74.n4 a_27_74.n3 104.579
R169 a_27_74.n5 a_27_74.n2 103.65
R170 a_27_74.n6 a_27_74.n1 103.65
R171 a_27_74.n7 a_27_74.n0 97.9062
R172 a_27_74.n6 a_27_74.n5 64.7534
R173 a_27_74.n7 a_27_74.n6 62.8815
R174 a_27_74.n5 a_27_74.n4 57.6005
R175 a_27_74.n8 a_27_74.n7 30.5783
R176 a_27_74.n0 a_27_74.t8 22.7032
R177 a_27_74.n0 a_27_74.t1 22.7032
R178 a_27_74.n3 a_27_74.t3 22.7032
R179 a_27_74.n3 a_27_74.t2 22.7032
R180 a_27_74.n2 a_27_74.t7 22.7032
R181 a_27_74.n2 a_27_74.t5 22.7032
R182 a_27_74.n1 a_27_74.t0 22.7032
R183 a_27_74.n1 a_27_74.t6 22.7032
R184 a_27_74.n9 a_27_74.t9 22.7032
R185 a_27_74.t10 a_27_74.n9 22.7032
R186 VNB.t15 VNB.t10 2286.61
R187 VNB.t3 VNB.t5 1154.86
R188 VNB.t4 VNB.t2 1154.86
R189 VNB VNB.t4 1143.31
R190 VNB.t0 VNB.t1 1039.37
R191 VNB.t11 VNB.t9 993.177
R192 VNB.t8 VNB.t11 993.177
R193 VNB.t10 VNB.t8 993.177
R194 VNB.t13 VNB.t15 993.177
R195 VNB.t14 VNB.t13 993.177
R196 VNB.t12 VNB.t14 993.177
R197 VNB.t1 VNB.t12 993.177
R198 VNB.t6 VNB.t0 993.177
R199 VNB.t7 VNB.t6 993.177
R200 VNB.t5 VNB.t7 993.177
R201 VNB.t2 VNB.t3 993.177
R202 A2.n1 A2.t2 226.444
R203 A2.n10 A2.t4 214.758
R204 A2.n7 A2.t5 214.758
R205 A2.n2 A2.t6 214.758
R206 A2.n2 A2.t3 197.941
R207 A2.n6 A2.t0 196.013
R208 A2.n9 A2.t1 196.013
R209 A2.n1 A2.t7 196.013
R210 A2.n12 A2.n11 152
R211 A2.n8 A2.n0 152
R212 A2.n6 A2.n5 152
R213 A2.n4 A2.n3 152
R214 A2.n6 A2.n3 43.7018
R215 A2.n8 A2.n7 39.2032
R216 A2.n11 A2.n1 25.7072
R217 A2.n11 A2.n10 25.0645
R218 A2.n9 A2.n8 11.5685
R219 A2.n4 A2 11.0145
R220 A2.n12 A2.n0 10.1214
R221 A2.n3 A2.n2 9.6405
R222 A2.n5 A2 7.44236
R223 A2.n10 A2.n9 7.06983
R224 A2.n5 A2 6.84701
R225 A2.n7 A2.n6 4.49917
R226 A2 A2.n4 3.27492
R227 A2 A2.n0 2.67957
R228 A2 A2.n12 1.48887
R229 VGND.n6 VGND.n5 214.816
R230 VGND.n4 VGND.n3 209.631
R231 VGND.n9 VGND.n2 209.631
R232 VGND.n12 VGND.n11 208.079
R233 VGND.n2 VGND.t1 34.0546
R234 VGND.n11 VGND.t2 34.0546
R235 VGND.n10 VGND.n9 25.977
R236 VGND.n5 VGND.t4 25.9464
R237 VGND.n5 VGND.t6 22.7032
R238 VGND.n3 VGND.t7 22.7032
R239 VGND.n3 VGND.t5 22.7032
R240 VGND.n2 VGND.t3 22.7032
R241 VGND.n11 VGND.t0 22.7032
R242 VGND.n9 VGND.n1 21.4593
R243 VGND.n12 VGND.n10 19.2005
R244 VGND.n4 VGND.n1 18.4476
R245 VGND.n7 VGND.n1 9.3005
R246 VGND.n9 VGND.n8 9.3005
R247 VGND.n10 VGND.n0 9.3005
R248 VGND.n13 VGND.n12 7.43488
R249 VGND.n6 VGND.n4 6.78149
R250 VGND.n7 VGND.n6 0.706558
R251 VGND VGND.n13 0.160103
R252 VGND.n13 VGND.n0 0.1477
R253 VGND.n8 VGND.n7 0.122949
R254 VGND.n8 VGND.n0 0.122949
C0 Y VGND 0.025309f
C1 A2 VPWR 0.026849f
C2 B1 C1 0.06736f
C3 A1 Y 9.54e-20
C4 VPB VGND 0.011692f
C5 VPB A1 0.141601f
C6 A2 Y 0.207592f
C7 A1 VGND 0.071856f
C8 B1 VPWR 0.045612f
C9 VPB A2 0.143508f
C10 A2 VGND 0.071562f
C11 B1 Y 0.140634f
C12 A1 A2 0.089257f
C13 VPB B1 0.101901f
C14 B1 VGND 0.020692f
C15 A2 B1 0.068435f
C16 C1 VPWR 0.048099f
C17 C1 Y 0.280159f
C18 VPB C1 0.125718f
C19 VPWR Y 0.605729f
C20 C1 VGND 0.023223f
C21 VPB VPWR 0.219634f
C22 VPWR VGND 0.131104f
C23 A1 VPWR 0.064445f
C24 VPB Y 0.068638f
C25 VGND VNB 0.915256f
C26 Y VNB 0.086553f
C27 VPWR VNB 0.740561f
C28 C1 VNB 0.410418f
C29 B1 VNB 0.349892f
C30 A2 VNB 0.406172f
C31 A1 VNB 0.450801f
C32 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o221a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221a_1 VNB VPB VPWR VGND C1 A1 A2 B1 B2 X
X0 a_83_264.t1 C1.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.43 ps=1.86 w=1 l=0.15
X1 VPWR.t0 a_83_264.t4 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3109 pd=1.71 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_264_392.t1 A1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.3109 ps=1.71 w=1 l=0.15
X3 a_462_392.t1 B2.t0 a_83_264.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X4 a_456_74.t2 B1.t0 a_245_94.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 VPWR.t1 B1.t1 a_462_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.43 pd=1.86 as=0.21 ps=1.42 w=1 l=0.15
X6 VGND.t0 a_83_264.t5 X.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 VGND.t1 A2.t0 a_245_94.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.112 ps=0.99 w=0.64 l=0.15
X8 a_245_94.t0 B2.t1 a_456_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2336 ps=2.01 w=0.64 l=0.15
X9 a_245_94.t3 A1.t1 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.15535 ps=1.17 w=0.64 l=0.15
X10 a_83_264.t0 C1.t1 a_456_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2944 pd=2.2 as=0.112 ps=0.99 w=0.64 l=0.15
X11 a_83_264.t3 A2.t1 a_264_392.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
R0 C1.n0 C1.t0 229.603
R1 C1.n1 C1.t1 157.571
R2 C1 C1.n0 153.695
R3 C1.n2 C1.n1 152
R4 C1.n1 C1.n0 39.9712
R5 C1 C1.n2 11.1064
R6 C1.n2 C1 2.82403
R7 VPWR.n2 VPWR.n1 318.507
R8 VPWR.n2 VPWR.n0 138.398
R9 VPWR.n0 VPWR.t3 82.2737
R10 VPWR.n0 VPWR.t1 72.4241
R11 VPWR.n1 VPWR.t2 59.1005
R12 VPWR.n1 VPWR.t0 55.271
R13 VPWR VPWR.n2 0.214998
R14 a_83_264.n2 a_83_264.n1 258.553
R15 a_83_264.n1 a_83_264.t4 256.337
R16 a_83_264.t1 a_83_264.n3 234.934
R17 a_83_264.n3 a_83_264.t0 216.156
R18 a_83_264.n1 a_83_264.t5 207.869
R19 a_83_264.n2 a_83_264.n0 205.1
R20 a_83_264.n3 a_83_264.n2 137.036
R21 a_83_264.n0 a_83_264.t2 53.1905
R22 a_83_264.n0 a_83_264.t3 29.5505
R23 VPB.t1 VPB.t3 515.861
R24 VPB.t0 VPB.t2 377.957
R25 VPB.t4 VPB.t1 291.13
R26 VPB.t5 VPB.t4 291.13
R27 VPB VPB.t0 257.93
R28 VPB.t2 VPB.t5 214.517
R29 X.n0 X.t0 293.673
R30 X.t1 X.n0 279.738
R31 X.n1 X.t1 279.738
R32 X.n1 X 10.2721
R33 X.n0 X 3.95112
R34 X X.n1 1.42272
R35 A1.n0 A1.t0 236.983
R36 A1.n0 A1.t1 236.18
R37 A1 A1.n0 154.133
R38 a_264_392.t0 a_264_392.t1 53.1905
R39 B2.n0 B2.t1 274.74
R40 B2.n0 B2.t0 236.983
R41 B2 B2.n0 161.504
R42 a_462_392.t0 a_462_392.t1 82.7405
R43 B1.n0 B1.t0 271.527
R44 B1.n0 B1.t1 253.075
R45 B1 B1.n0 154.133
R46 a_245_94.n1 a_245_94.n0 397.993
R47 a_245_94.n0 a_245_94.t2 39.3755
R48 a_245_94.n0 a_245_94.t3 26.2505
R49 a_245_94.n1 a_245_94.t1 26.2505
R50 a_245_94.t0 a_245_94.n1 26.2505
R51 a_456_74.n0 a_456_74.t1 284.541
R52 a_456_74.n0 a_456_74.t2 39.3755
R53 a_456_74.t0 a_456_74.n0 26.2505
R54 VNB.t4 VNB.t2 2471.39
R55 VNB.t0 VNB.t5 1339.63
R56 VNB VNB.t0 1316.54
R57 VNB.t3 VNB.t1 1154.86
R58 VNB.t5 VNB.t4 1154.86
R59 VNB.t2 VNB.t3 993.177
R60 VGND.n1 VGND.t1 245.688
R61 VGND.n1 VGND.n0 121.951
R62 VGND.n0 VGND.t2 41.2505
R63 VGND.n0 VGND.t0 30.6984
R64 VGND VGND.n1 0.479817
R65 A2.n0 A2.t1 236.983
R66 A2.n0 A2.t0 236.18
R67 A2 A2.n0 157.625
C0 A1 VPWR 0.015747f
C1 VPB VGND 0.010233f
C2 B1 C1 0.083783f
C3 B2 X 1.17e-19
C4 VPB A2 0.040583f
C5 A2 VGND 0.015037f
C6 B2 VPWR 0.012608f
C7 A1 C1 7.8e-20
C8 VPB X 0.012817f
C9 X VGND 0.109491f
C10 VPB VPWR 0.117243f
C11 VPWR VGND 0.070901f
C12 B2 C1 8.92e-19
C13 A2 X 2.79e-19
C14 A2 VPWR 0.009489f
C15 VPB C1 0.055532f
C16 A1 B1 1.02e-20
C17 C1 VGND 0.013325f
C18 X VPWR 0.089093f
C19 B2 B1 0.088978f
C20 A2 C1 1.23e-19
C21 C1 X 3.05e-19
C22 VPB B1 0.059314f
C23 B1 VGND 0.006383f
C24 C1 VPWR 0.020842f
C25 A2 B1 1.69e-20
C26 VPB A1 0.044887f
C27 A1 VGND 0.019637f
C28 B1 X 1.24e-20
C29 VPB B2 0.049727f
C30 A1 A2 0.08546f
C31 B1 VPWR 0.023096f
C32 B2 VGND 0.008546f
C33 A1 X 0.00165f
C34 A2 B2 0.069736f
C35 VGND VNB 0.542718f
C36 VPWR VNB 0.427728f
C37 X VNB 0.114149f
C38 C1 VNB 0.165609f
C39 B1 VNB 0.121254f
C40 B2 VNB 0.160211f
C41 A2 VNB 0.107807f
C42 A1 VNB 0.10856f
C43 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o221a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221a_2 VNB VPB VPWR VGND A1 A2 B2 C1 X B1
X0 X.t1 a_27_368.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2957 ps=1.67 w=1.12 l=0.15
X1 VPWR.t4 C1.t0 a_27_368.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.465 pd=1.93 as=0.295 ps=2.59 w=1 l=0.15
X2 VGND.t2 A1.t0 a_264_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_332_368.t1 B1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.465 ps=1.93 w=1 l=0.15
X4 a_530_368.t1 A2.t0 a_27_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X5 VPWR.t3 A1.t1 a_530_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2957 pd=1.67 as=0.21 ps=1.42 w=1 l=0.15
X6 a_165_74.t0 B2.t0 a_264_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.13135 ps=1.095 w=0.74 l=0.15
X7 X.t3 a_27_368.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8 VGND.t0 a_27_368.t6 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.3108 pd=2.32 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_264_74.t0 B1.t1 a_165_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.13135 pd=1.095 as=0.12765 ps=1.085 w=0.74 l=0.15
X10 a_27_368.t1 B2.t1 a_332_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X11 a_165_74.t2 C1.t1 a_27_368.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.12765 pd=1.085 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 a_264_74.t3 A2.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 VPWR.t0 a_27_368.t7 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 a_27_368.n0 a_27_368.t7 323.209
R1 a_27_368.n4 a_27_368.n2 274.95
R2 a_27_368.n2 a_27_368.t4 258.233
R3 a_27_368.n3 a_27_368.t3 243.072
R4 a_27_368.n5 a_27_368.n4 202.177
R5 a_27_368.n3 a_27_368.t2 202.173
R6 a_27_368.n1 a_27_368.t5 197.006
R7 a_27_368.n0 a_27_368.t6 186.374
R8 a_27_368.n4 a_27_368.n3 100.757
R9 a_27_368.n1 a_27_368.n0 75.5138
R10 a_27_368.t0 a_27_368.n5 53.1905
R11 a_27_368.n5 a_27_368.t1 29.5505
R12 a_27_368.n2 a_27_368.n1 12.7593
R13 VPWR.n3 VPWR.n1 585
R14 VPWR.n2 VPWR.n1 585
R15 VPWR.n9 VPWR.n8 315.926
R16 VPWR.n5 VPWR.n4 266.478
R17 VPWR.n7 VPWR.t0 266.221
R18 VPWR.n8 VPWR.t3 68.9505
R19 VPWR.n4 VPWR.n3 52.0482
R20 VPWR.n4 VPWR.n2 52.0482
R21 VPWR.n3 VPWR.t4 39.4005
R22 VPWR.n10 VPWR.n6 36.1417
R23 VPWR.n14 VPWR.n6 36.1417
R24 VPWR.n15 VPWR.n14 36.1417
R25 VPWR.n8 VPWR.t1 35.2408
R26 VPWR.n2 VPWR.t2 29.5505
R27 VPWR.n10 VPWR.n9 21.4593
R28 VPWR.n16 VPWR.n15 11.6711
R29 VPWR.n11 VPWR.n10 9.3005
R30 VPWR.n12 VPWR.n6 9.3005
R31 VPWR.n14 VPWR.n13 9.3005
R32 VPWR.n15 VPWR.n0 9.3005
R33 VPWR.n16 VPWR.n5 8.65105
R34 VPWR.n9 VPWR.n7 6.8344
R35 VPWR.n5 VPWR.n1 4.78292
R36 VPWR.n17 VPWR.n16 4.09689
R37 VPWR.n11 VPWR.n7 0.569119
R38 VPWR VPWR.n17 0.225146
R39 VPWR.n17 VPWR.n0 0.204827
R40 VPWR.n12 VPWR.n11 0.122949
R41 VPWR.n13 VPWR.n12 0.122949
R42 VPWR.n13 VPWR.n0 0.122949
R43 X.n1 X.n0 265.277
R44 X.n2 X.n1 185
R45 X.n3 X.n2 185
R46 X.n0 X.t0 26.3844
R47 X.n0 X.t1 26.3844
R48 X.n2 X.t2 22.7032
R49 X.n2 X.t3 22.7032
R50 X.n3 X 8.75839
R51 X.n1 X 3.36892
R52 X X.n3 1.21313
R53 VPB.t6 VPB.t3 551.614
R54 VPB.t5 VPB.t1 357.527
R55 VPB.t2 VPB.t5 291.13
R56 VPB.t4 VPB.t2 291.13
R57 VPB VPB.t6 257.93
R58 VPB.t1 VPB.t0 229.839
R59 VPB.t3 VPB.t4 214.517
R60 C1.n0 C1.t0 242.339
R61 C1 C1.n0 193.113
R62 C1.n0 C1.t1 190.025
R63 A1.n0 A1.t1 231.629
R64 A1.n0 A1.t0 220.113
R65 A1 A1.n0 157.507
R66 a_264_74.n1 a_264_74.n0 388.817
R67 a_264_74.n1 a_264_74.t2 29.1897
R68 a_264_74.t0 a_264_74.n1 28.3789
R69 a_264_74.n0 a_264_74.t1 22.7032
R70 a_264_74.n0 a_264_74.t3 22.7032
R71 VGND.n5 VGND.t3 233.498
R72 VGND.n1 VGND.t0 176.026
R73 VGND.n3 VGND.n2 116.644
R74 VGND.n2 VGND.t1 34.0546
R75 VGND.n2 VGND.t2 34.0546
R76 VGND.n5 VGND.n4 32.377
R77 VGND.n4 VGND.n3 12.8005
R78 VGND.n4 VGND.n0 9.3005
R79 VGND.n3 VGND.n1 7.24947
R80 VGND.n6 VGND.n5 6.56837
R81 VGND VGND.n6 0.633217
R82 VGND.n1 VGND.n0 0.494123
R83 VGND.n6 VGND.n0 0.166523
R84 VNB.t4 VNB.t5 2286.61
R85 VNB VNB.t6 1732.28
R86 VNB.t3 VNB.t2 1316.54
R87 VNB.t0 VNB.t4 1166.4
R88 VNB.t6 VNB.t0 1143.31
R89 VNB.t2 VNB.t1 993.177
R90 VNB.t5 VNB.t3 993.177
R91 B1.n0 B1.t0 267.413
R92 B1.n0 B1.t1 220.113
R93 B1 B1.n0 155.423
R94 a_332_368.t0 a_332_368.t1 53.1905
R95 A2.n0 A2.t0 231.629
R96 A2.n0 A2.t1 220.113
R97 A2 A2.n0 154.828
R98 a_530_368.t0 a_530_368.t1 82.7405
R99 B2.n0 B2.t0 233.26
R100 B2.n0 B2.t1 231.629
R101 B2 B2.n0 152.149
R102 a_165_74.t0 a_165_74.n0 374.781
R103 a_165_74.n0 a_165_74.t2 33.2437
R104 a_165_74.n0 a_165_74.t1 22.7032
C0 VPB B1 0.052636f
C1 A1 VPWR 0.013223f
C2 VGND VPWR 0.091515f
C3 C1 B1 0.041413f
C4 B2 VPB 0.040906f
C5 A2 VPB 0.035482f
C6 X VPB 0.006067f
C7 B2 B1 0.092135f
C8 A1 VPB 0.039121f
C9 X C1 1.1e-20
C10 VGND VPB 0.010701f
C11 VPWR VPB 0.156073f
C12 VGND C1 0.013733f
C13 X B1 4.38e-20
C14 VPWR C1 0.017889f
C15 VGND B1 0.007324f
C16 VPWR B1 0.02078f
C17 B2 A2 0.075487f
C18 X B2 2.85e-19
C19 VGND B2 0.010016f
C20 X A2 3.93e-19
C21 B2 VPWR 0.013701f
C22 A2 A1 0.088538f
C23 VGND A2 0.017323f
C24 X A1 0.001309f
C25 X VGND 0.185683f
C26 VPB C1 0.054633f
C27 A2 VPWR 0.009084f
C28 X VPWR 0.198422f
C29 VGND A1 0.028404f
C30 VGND VNB 0.636457f
C31 X VNB 0.035517f
C32 VPWR VNB 0.515437f
C33 A1 VNB 0.104758f
C34 A2 VNB 0.105559f
C35 B2 VNB 0.140726f
C36 B1 VNB 0.128132f
C37 C1 VNB 0.197353f
C38 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o221a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221a_4 VNB VPB VPWR VGND X A1 A2 B1 B2 C1
X0 a_763_387.t3 A2.t0 a_114_125.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.1625 ps=1.325 w=1 l=0.15
X1 VPWR.t3 a_114_125.t8 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.475 w=1.12 l=0.15
X2 a_300_125.t4 A2.t1 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 a_114_125.t4 C1.t0 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X4 X.t4 a_114_125.t9 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.475 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_300_125.t7 B1.t0 a_27_125.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1008 pd=0.955 as=0.112 ps=0.99 w=0.64 l=0.15
X6 a_300_125.t1 B2.t0 a_27_125.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0912 pd=0.925 as=0.1008 ps=0.955 w=0.64 l=0.15
X7 a_114_125.t6 A2.t2 a_763_387.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.1625 ps=1.325 w=1 l=0.15
X8 VPWR.t5 B1.t1 a_297_387.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3925 pd=1.785 as=0.15 ps=1.3 w=1 l=0.15
X9 a_297_387.t3 B2.t1 a_114_125.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X10 a_114_125.t0 B2.t2 a_297_387.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1725 ps=1.345 w=1 l=0.15
X11 VGND.t2 a_114_125.t10 X.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.10545 ps=1.025 w=0.74 l=0.15
X12 a_763_387.t1 A1.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.3925 ps=1.785 w=1 l=0.15
X13 a_300_125.t5 A1.t1 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0912 pd=0.925 as=0.1824 ps=1.85 w=0.64 l=0.15
X14 VGND.t6 A1.t2 a_300_125.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1535 pd=1.165 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 a_27_125.t4 C1.t1 a_114_125.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 a_27_125.t0 B1.t2 a_300_125.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0912 ps=0.925 w=0.64 l=0.15
X17 a_114_125.t2 C1.t2 a_27_125.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X18 X.t3 a_114_125.t11 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.495 as=0.1934 ps=1.475 w=1.12 l=0.15
X19 X.t1 a_114_125.t12 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X20 VPWR.t6 C1.t3 a_114_125.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1525 pd=1.305 as=0.15 ps=1.3 w=1 l=0.15
X21 a_27_125.t2 B2.t3 a_300_125.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1008 pd=0.955 as=0.1008 ps=0.955 w=0.64 l=0.15
X22 a_297_387.t0 B1.t3 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.1525 ps=1.305 w=1 l=0.15
X23 VPWR.t0 A1.t3 a_763_387.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.175 ps=1.35 w=1 l=0.15
X24 VGND.t3 A2.t3 a_300_125.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0912 ps=0.925 w=0.64 l=0.15
X25 VGND.t0 a_114_125.t13 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A2.n1 A2.t2 211.911
R1 A2.n0 A2.t0 209.19
R2 A2.n0 A2.t1 170.308
R3 A2.n1 A2.t3 170.308
R4 A2 A2.n2 154.102
R5 A2.n2 A2.n1 41.6278
R6 A2.n2 A2.n0 21.1793
R7 a_114_125.n18 a_114_125.n17 300.733
R8 a_114_125.n13 a_114_125.n12 300.514
R9 a_114_125.n3 a_114_125.t8 252.053
R10 a_114_125.n5 a_114_125.t9 226.809
R11 a_114_125.n7 a_114_125.n2 226.809
R12 a_114_125.n9 a_114_125.t11 226.809
R13 a_114_125.n16 a_114_125.n15 223.911
R14 a_114_125.n16 a_114_125.n14 177.93
R15 a_114_125.n6 a_114_125.n0 165.189
R16 a_114_125.n17 a_114_125.n13 163.388
R17 a_114_125.n9 a_114_125.n8 158.038
R18 a_114_125.n3 a_114_125.t13 155.847
R19 a_114_125.n1 a_114_125.t10 155.847
R20 a_114_125.n4 a_114_125.t12 155.847
R21 a_114_125.n11 a_114_125.n10 152
R22 a_114_125.n1 a_114_125.n0 152
R23 a_114_125.n13 a_114_125.n11 99.0465
R24 a_114_125.n17 a_114_125.n16 74.1652
R25 a_114_125.n4 a_114_125.n3 73.1769
R26 a_114_125.n10 a_114_125.n1 49.6611
R27 a_114_125.n12 a_114_125.t6 34.4755
R28 a_114_125.n7 a_114_125.n6 33.5944
R29 a_114_125.n6 a_114_125.n5 32.1338
R30 a_114_125.n15 a_114_125.t3 29.5505
R31 a_114_125.n15 a_114_125.t4 29.5505
R32 a_114_125.n12 a_114_125.t7 29.5505
R33 a_114_125.n18 a_114_125.t1 29.5505
R34 a_114_125.t0 a_114_125.n18 29.5505
R35 a_114_125.n14 a_114_125.t5 26.2505
R36 a_114_125.n14 a_114_125.t2 26.2505
R37 a_114_125.n1 a_114_125.n7 16.0672
R38 a_114_125.n11 a_114_125.n0 13.1884
R39 a_114_125.n10 a_114_125.n9 10.955
R40 a_114_125.n5 a_114_125.n4 2.19141
R41 a_763_387.n1 a_763_387.n0 658.148
R42 a_763_387.n0 a_763_387.t3 39.4005
R43 a_763_387.t2 a_763_387.n1 34.4755
R44 a_763_387.n0 a_763_387.t0 29.5505
R45 a_763_387.n1 a_763_387.t1 29.5505
R46 VPB.t1 VPB.t2 497.985
R47 VPB.t7 VPB.t5 477.555
R48 VPB.t2 VPB.t3 257.93
R49 VPB.t0 VPB.t1 257.93
R50 VPB VPB.t9 257.93
R51 VPB.t11 VPB.t0 255.376
R52 VPB.t12 VPB.t4 252.823
R53 VPB.t10 VPB.t11 242.608
R54 VPB.t5 VPB.t10 242.608
R55 VPB.t8 VPB.t12 232.393
R56 VPB.t6 VPB.t7 229.839
R57 VPB.t4 VPB.t6 229.839
R58 VPB.t9 VPB.t8 229.839
R59 X.n1 X.t3 293.151
R60 X.n1 X.n0 205.66
R61 X.n3 X.t2 196.163
R62 X.n3 X.n2 99.1033
R63 X.n0 X.t4 36.0585
R64 X.n0 X.t5 26.3844
R65 X.n4 X.n3 24.6724
R66 X.n2 X.t0 22.7032
R67 X.n2 X.t1 22.7032
R68 X X.n4 13.357
R69 X.n4 X.n1 10.4732
R70 VPWR.n9 VPWR.t2 351.026
R71 VPWR.n25 VPWR.n2 324.182
R72 VPWR.n13 VPWR.n8 317.038
R73 VPWR.n10 VPWR.t3 264.486
R74 VPWR.n27 VPWR.t7 261.353
R75 VPWR.n19 VPWR.n5 136.803
R76 VPWR.n5 VPWR.t5 70.6176
R77 VPWR.n5 VPWR.t4 70.6172
R78 VPWR.n8 VPWR.t0 39.4005
R79 VPWR.n20 VPWR.n3 36.1417
R80 VPWR.n24 VPWR.n3 36.1417
R81 VPWR.n14 VPWR.n6 36.1417
R82 VPWR.n18 VPWR.n6 36.1417
R83 VPWR.n19 VPWR.n18 33.8829
R84 VPWR.n2 VPWR.t8 30.5355
R85 VPWR.n2 VPWR.t6 29.5505
R86 VPWR.n26 VPWR.n25 28.2358
R87 VPWR.n13 VPWR.n12 27.8593
R88 VPWR.n8 VPWR.t1 27.1918
R89 VPWR.n12 VPWR.n9 27.1064
R90 VPWR.n27 VPWR.n26 26.7299
R91 VPWR.n25 VPWR.n24 25.224
R92 VPWR.n20 VPWR.n19 20.7064
R93 VPWR.n14 VPWR.n13 19.577
R94 VPWR.n12 VPWR.n11 9.3005
R95 VPWR.n13 VPWR.n7 9.3005
R96 VPWR.n15 VPWR.n14 9.3005
R97 VPWR.n16 VPWR.n6 9.3005
R98 VPWR.n18 VPWR.n17 9.3005
R99 VPWR.n21 VPWR.n20 9.3005
R100 VPWR.n22 VPWR.n3 9.3005
R101 VPWR.n24 VPWR.n23 9.3005
R102 VPWR.n25 VPWR.n1 9.3005
R103 VPWR.n26 VPWR.n0 9.3005
R104 VPWR.n28 VPWR.n27 9.3005
R105 VPWR.n10 VPWR.n9 6.8559
R106 VPWR.n19 VPWR.n4 4.62059
R107 VPWR.n11 VPWR.n10 0.565232
R108 VPWR.n17 VPWR.n4 0.184273
R109 VPWR.n21 VPWR.n4 0.184273
R110 VPWR.n11 VPWR.n7 0.122949
R111 VPWR.n15 VPWR.n7 0.122949
R112 VPWR.n16 VPWR.n15 0.122949
R113 VPWR.n17 VPWR.n16 0.122949
R114 VPWR.n22 VPWR.n21 0.122949
R115 VPWR.n23 VPWR.n22 0.122949
R116 VPWR.n23 VPWR.n1 0.122949
R117 VPWR.n1 VPWR.n0 0.122949
R118 VPWR.n28 VPWR.n0 0.122949
R119 VPWR VPWR.n28 0.0617245
R120 VGND.n14 VGND.t5 281.654
R121 VGND.n12 VGND.n2 213.898
R122 VGND.n6 VGND.n5 205.481
R123 VGND.n4 VGND.t0 166.28
R124 VGND.n8 VGND.t6 162.431
R125 VGND.n5 VGND.t1 39.7302
R126 VGND.n8 VGND.n7 32.7534
R127 VGND.n12 VGND.n1 31.2476
R128 VGND.n5 VGND.t2 28.3789
R129 VGND.n2 VGND.t4 26.2505
R130 VGND.n2 VGND.t3 26.2505
R131 VGND.n14 VGND.n13 24.0946
R132 VGND.n13 VGND.n12 16.1887
R133 VGND.n8 VGND.n1 14.6829
R134 VGND.n7 VGND.n6 12.424
R135 VGND.n13 VGND.n0 9.3005
R136 VGND.n12 VGND.n11 9.3005
R137 VGND.n10 VGND.n1 9.3005
R138 VGND.n7 VGND.n3 9.3005
R139 VGND.n9 VGND.n8 9.3005
R140 VGND.n15 VGND.n14 7.12802
R141 VGND.n6 VGND.n4 6.96039
R142 VGND VGND.n15 0.888238
R143 VGND.n4 VGND.n3 0.594857
R144 VGND.n15 VGND.n0 0.157708
R145 VGND.n9 VGND.n3 0.122949
R146 VGND.n10 VGND.n9 0.122949
R147 VGND.n11 VGND.n10 0.122949
R148 VGND.n11 VGND.n0 0.122949
R149 a_300_125.n5 a_300_125.n4 148.611
R150 a_300_125.n2 a_300_125.n1 136.106
R151 a_300_125.n4 a_300_125.n2 106.007
R152 a_300_125.n4 a_300_125.n3 98.6928
R153 a_300_125.n2 a_300_125.n0 96.0511
R154 a_300_125.n1 a_300_125.t0 32.813
R155 a_300_125.n3 a_300_125.t3 27.188
R156 a_300_125.n0 a_300_125.t2 27.188
R157 a_300_125.n3 a_300_125.t5 26.2505
R158 a_300_125.n0 a_300_125.t1 26.2505
R159 a_300_125.n1 a_300_125.t7 26.2505
R160 a_300_125.n5 a_300_125.t6 26.2505
R161 a_300_125.t4 a_300_125.n5 26.2505
R162 VNB.t5 VNB.t10 2355.91
R163 VNB.t11 VNB.t2 2332.81
R164 VNB.t2 VNB.t1 1316.54
R165 VNB.t7 VNB.t12 1154.86
R166 VNB VNB.t6 1143.31
R167 VNB.t3 VNB.t4 1074.02
R168 VNB.t12 VNB.t3 1074.02
R169 VNB.t10 VNB.t8 1004.72
R170 VNB.t4 VNB.t5 1004.72
R171 VNB.t1 VNB.t0 993.177
R172 VNB.t9 VNB.t11 993.177
R173 VNB.t8 VNB.t9 993.177
R174 VNB.t6 VNB.t7 993.177
R175 C1.n0 C1.t3 211.911
R176 C1.n2 C1.t0 207.529
R177 C1.n4 C1.n3 168.067
R178 C1.n3 C1.t2 160.667
R179 C1.n0 C1.t1 160.667
R180 C1 C1.n1 155.44
R181 C1.n2 C1.n1 32.1338
R182 C1.n1 C1.n0 29.2126
R183 C1 C1.n4 9.55274
R184 C1.n4 C1 8.78856
R185 C1.n3 C1.n2 1.46111
R186 B1.n1 B1.t0 1210.99
R187 B1.t0 B1.t3 450.938
R188 B1.n0 B1.t1 275.812
R189 B1.n0 B1.t2 180.75
R190 B1.n2 B1.n1 152
R191 B1.n1 B1.n0 91.5805
R192 B1 B1.n2 9.36169
R193 B1.n2 B1 8.9796
R194 a_27_125.n1 a_27_125.t0 314.483
R195 a_27_125.n3 a_27_125.n2 201.292
R196 a_27_125.n1 a_27_125.n0 200.516
R197 a_27_125.n2 a_27_125.t3 199.994
R198 a_27_125.n2 a_27_125.n1 51.2233
R199 a_27_125.t1 a_27_125.n3 39.3755
R200 a_27_125.n0 a_27_125.t2 32.813
R201 a_27_125.n0 a_27_125.t5 26.2505
R202 a_27_125.n3 a_27_125.t4 26.2505
R203 B2.n0 B2.t1 207.529
R204 B2.n1 B2.t2 207.529
R205 B2.n1 B2.t3 162.858
R206 B2.n0 B2.t0 160.667
R207 B2.n3 B2.n2 152
R208 B2.n2 B2.n1 54.7732
R209 B2.n2 B2.n0 10.955
R210 B2 B2.n3 10.508
R211 B2.n3 B2 7.83334
R212 a_297_387.n1 a_297_387.n0 650.617
R213 a_297_387.n0 a_297_387.t0 38.4155
R214 a_297_387.n0 a_297_387.t2 29.5505
R215 a_297_387.t1 a_297_387.n1 29.5505
R216 a_297_387.n1 a_297_387.t3 29.5505
R217 A1.t2 A1.t1 840.288
R218 A1.t1 A1.t0 449.57
R219 A1.n0 A1.t3 257.067
R220 A1.n0 A1.t2 163.881
R221 A1 A1.n0 157.953
C0 VPB B1 0.102519f
C1 VPWR B2 0.011409f
C2 X B1 4.86e-19
C3 B1 A1 0.078938f
C4 VPWR VPB 0.212669f
C5 VPB B2 0.0723f
C6 C1 B1 0.049521f
C7 VPWR X 0.402023f
C8 VGND B1 0.07846f
C9 X B2 1.8e-20
C10 VPWR A1 0.034074f
C11 B2 A1 6.26e-20
C12 B1 A2 0.03689f
C13 X VPB 0.014351f
C14 VPWR C1 0.058556f
C15 VPB A1 0.080486f
C16 VPWR VGND 0.127101f
C17 VPWR A2 0.01098f
C18 X A1 0.001963f
C19 VGND B2 0.008343f
C20 VPB C1 0.086888f
C21 VGND VPB 0.011559f
C22 VPB A2 0.072302f
C23 X VGND 0.306354f
C24 X A2 4.19e-19
C25 VGND A1 0.105345f
C26 A1 A2 0.161113f
C27 VGND C1 0.011501f
C28 VGND A2 0.02402f
C29 VPWR B1 0.043351f
C30 B1 B2 0.155795f
C31 VGND VNB 0.92318f
C32 X VNB 0.04126f
C33 VPWR VNB 0.771402f
C34 A2 VNB 0.157572f
C35 A1 VNB 0.364859f
C36 B2 VNB 0.160025f
C37 B1 VNB 0.55289f
C38 C1 VNB 0.231484f
C39 VPB VNB 1.79899f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o41ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o41ai_4 VNB VPB VPWR VGND A1 A2 A3 A4 B1 Y
X0 Y.t4 B1.t0 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_1191_368.t7 A1.t0 VPWR.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_788_368.t4 A3.t0 a_339_368.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VPWR.t0 B1.t1 Y.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4 a_27_74.t4 A4.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.2146 ps=1.32 w=0.74 l=0.15
X5 a_339_368.t1 A3.t1 a_788_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X6 a_339_368.t0 A3.t2 a_788_368.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_27_74.t16 A1.t1 VGND.t10 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.13505 ps=1.105 w=0.74 l=0.15
X8 Y.t5 B1.t2 a_27_74.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 VGND.t5 A2.t0 a_27_74.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_27_74.t13 A3.t3 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 VPWR.t3 A1.t2 a_1191_368.t6 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_1191_368.t5 A1.t3 VPWR.t4 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X13 VGND.t3 A4.t1 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=1.32 as=0.1295 ps=1.09 w=0.74 l=0.15
X14 VGND.t8 A3.t4 a_27_74.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_27_74.t7 B1.t3 Y.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 a_27_74.t11 A3.t5 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 a_788_368.t1 A3.t6 a_339_368.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VPWR.t5 A1.t4 a_1191_368.t4 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VGND.t2 A4.t2 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11285 ps=1.045 w=0.74 l=0.15
X20 a_27_74.t15 A1.t5 VGND.t12 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X21 a_1191_368.t3 A2.t1 a_788_368.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_27_74.t6 B1.t4 Y.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_339_368.t4 A4.t3 Y.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_27_74.t0 A2.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12395 pd=1.075 as=0.11655 ps=1.055 w=0.74 l=0.15
X25 Y.t7 A4.t4 a_339_368.t5 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 a_788_368.t5 A2.t3 a_1191_368.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 a_1191_368.t0 A2.t4 a_788_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 a_339_368.t6 A4.t5 Y.t8 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 Y.t9 A4.t6 a_339_368.t7 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X30 a_788_368.t6 A2.t5 a_1191_368.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X31 a_27_74.t1 A4.t7 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 Y.t0 B1.t5 a_27_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 VGND.t6 A3.t7 a_27_74.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X34 VGND.t11 A1.t6 a_27_74.t14 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 B1.n1 B1.t3 303.661
R1 B1.n2 B1.t1 261.62
R2 B1.n6 B1.t0 261.62
R3 B1.n8 B1.n7 177.751
R4 B1.n4 B1.n3 163.762
R5 B1.n5 B1.n4 152
R6 B1.n1 B1.t5 142.994
R7 B1.n7 B1.t2 142.994
R8 B1.n0 B1.t4 142.994
R9 B1.n2 B1.n1 79.3654
R10 B1.n5 B1.n0 37.6361
R11 B1.n6 B1.n5 17.8279
R12 B1.n8 B1 11.5897
R13 B1.n3 B1.n2 9.90461
R14 B1.n3 B1.n0 7.26351
R15 B1 B1.n8 5.01672
R16 B1.n7 B1.n6 1.32105
R17 B1.n4 B1 0.173473
R18 VPWR.n34 VPWR.t0 413.724
R19 VPWR.n12 VPWR.n9 323.921
R20 VPWR.n11 VPWR.n10 318.236
R21 VPWR.n36 VPWR.t1 250.081
R22 VPWR.n15 VPWR.n8 36.1417
R23 VPWR.n16 VPWR.n15 36.1417
R24 VPWR.n17 VPWR.n16 36.1417
R25 VPWR.n17 VPWR.n6 36.1417
R26 VPWR.n21 VPWR.n6 36.1417
R27 VPWR.n22 VPWR.n21 36.1417
R28 VPWR.n23 VPWR.n22 36.1417
R29 VPWR.n23 VPWR.n4 36.1417
R30 VPWR.n27 VPWR.n4 36.1417
R31 VPWR.n28 VPWR.n27 36.1417
R32 VPWR.n29 VPWR.n28 36.1417
R33 VPWR.n29 VPWR.n2 36.1417
R34 VPWR.n33 VPWR.n2 36.1417
R35 VPWR.n10 VPWR.t4 35.1791
R36 VPWR.n9 VPWR.t3 35.1791
R37 VPWR.n35 VPWR.n34 29.7417
R38 VPWR.n10 VPWR.t5 26.3844
R39 VPWR.n9 VPWR.t2 26.3844
R40 VPWR.n36 VPWR.n35 20.7064
R41 VPWR.n11 VPWR.n8 19.9534
R42 VPWR.n34 VPWR.n33 17.6946
R43 VPWR.n13 VPWR.n8 9.3005
R44 VPWR.n15 VPWR.n14 9.3005
R45 VPWR.n16 VPWR.n7 9.3005
R46 VPWR.n18 VPWR.n17 9.3005
R47 VPWR.n19 VPWR.n6 9.3005
R48 VPWR.n21 VPWR.n20 9.3005
R49 VPWR.n22 VPWR.n5 9.3005
R50 VPWR.n24 VPWR.n23 9.3005
R51 VPWR.n25 VPWR.n4 9.3005
R52 VPWR.n27 VPWR.n26 9.3005
R53 VPWR.n28 VPWR.n3 9.3005
R54 VPWR.n30 VPWR.n29 9.3005
R55 VPWR.n31 VPWR.n2 9.3005
R56 VPWR.n33 VPWR.n32 9.3005
R57 VPWR.n34 VPWR.n1 9.3005
R58 VPWR.n35 VPWR.n0 9.3005
R59 VPWR.n37 VPWR.n36 9.3005
R60 VPWR.n12 VPWR.n11 6.94321
R61 VPWR.n13 VPWR.n12 0.516733
R62 VPWR.n14 VPWR.n13 0.122949
R63 VPWR.n14 VPWR.n7 0.122949
R64 VPWR.n18 VPWR.n7 0.122949
R65 VPWR.n19 VPWR.n18 0.122949
R66 VPWR.n20 VPWR.n19 0.122949
R67 VPWR.n20 VPWR.n5 0.122949
R68 VPWR.n24 VPWR.n5 0.122949
R69 VPWR.n25 VPWR.n24 0.122949
R70 VPWR.n26 VPWR.n25 0.122949
R71 VPWR.n26 VPWR.n3 0.122949
R72 VPWR.n30 VPWR.n3 0.122949
R73 VPWR.n31 VPWR.n30 0.122949
R74 VPWR.n32 VPWR.n31 0.122949
R75 VPWR.n32 VPWR.n1 0.122949
R76 VPWR.n1 VPWR.n0 0.122949
R77 VPWR.n37 VPWR.n0 0.122949
R78 VPWR VPWR.n37 0.0617245
R79 Y Y.n0 301.837
R80 Y.n7 Y.n1 297.224
R81 Y.n6 Y.n2 250.608
R82 Y.n5 Y.n3 245.613
R83 Y.n5 Y.n4 187.522
R84 Y.n2 Y.t3 35.1791
R85 Y.n2 Y.t4 35.1791
R86 Y.n6 Y.n5 34.1338
R87 Y.n4 Y.t0 34.0546
R88 Y.n7 Y.n6 30.1444
R89 Y.n1 Y.t8 26.3844
R90 Y.n1 Y.t9 26.3844
R91 Y.n0 Y.t6 26.3844
R92 Y.n0 Y.t7 26.3844
R93 Y.n4 Y.t2 22.7032
R94 Y.n3 Y.t1 22.7032
R95 Y.n3 Y.t5 22.7032
R96 Y Y.n7 7.88887
R97 VPB.t0 VPB.t10 515.861
R98 VPB.t5 VPB.t14 515.861
R99 VPB.t1 VPB.t3 280.914
R100 VPB.t6 VPB.t5 280.914
R101 VPB VPB.t6 257.93
R102 VPB.t15 VPB.t7 255.376
R103 VPB.t17 VPB.t16 255.376
R104 VPB.t16 VPB.t15 229.839
R105 VPB.t11 VPB.t17 229.839
R106 VPB.t8 VPB.t11 229.839
R107 VPB.t4 VPB.t8 229.839
R108 VPB.t10 VPB.t4 229.839
R109 VPB.t2 VPB.t0 229.839
R110 VPB.t3 VPB.t2 229.839
R111 VPB.t9 VPB.t1 229.839
R112 VPB.t12 VPB.t9 229.839
R113 VPB.t13 VPB.t12 229.839
R114 VPB.t14 VPB.t13 229.839
R115 A1.n1 A1.t0 261.62
R116 A1.n7 A1.t2 261.62
R117 A1.n10 A1.t3 261.62
R118 A1.n12 A1.t4 261.62
R119 A1.n1 A1.t5 155.702
R120 A1.n12 A1.n11 154.24
R121 A1.n9 A1.t1 154.24
R122 A1.n6 A1.t6 154.24
R123 A1.n3 A1.n2 152
R124 A1.n5 A1.n4 152
R125 A1.n8 A1.n0 152
R126 A1.n14 A1.n13 152
R127 A1.n5 A1.n2 49.6611
R128 A1.n13 A1.n12 45.2793
R129 A1.n8 A1.n7 41.6278
R130 A1.n13 A1.n10 25.5611
R131 A1.n9 A1.n8 19.7187
R132 A1.n2 A1.n1 15.3369
R133 A1.n14 A1.n0 11.7627
R134 A1.n4 A1 11.5897
R135 A1.n3 A1 9.85996
R136 A1 A1.n3 6.74645
R137 A1.n6 A1.n5 6.57323
R138 A1.n4 A1 5.01672
R139 A1 A1.n14 4.67077
R140 A1.n10 A1.n9 4.38232
R141 A1.n7 A1.n6 1.46111
R142 A1 A1.n0 0.173473
R143 a_1191_368.n2 a_1191_368.t2 458.132
R144 a_1191_368.n2 a_1191_368.n1 304.668
R145 a_1191_368.n4 a_1191_368.t7 289.856
R146 a_1191_368.n5 a_1191_368.n4 210.334
R147 a_1191_368.n3 a_1191_368.n0 186.477
R148 a_1191_368.n4 a_1191_368.n3 76.995
R149 a_1191_368.n3 a_1191_368.n2 69.6245
R150 a_1191_368.n0 a_1191_368.t4 26.3844
R151 a_1191_368.n0 a_1191_368.t3 26.3844
R152 a_1191_368.n1 a_1191_368.t1 26.3844
R153 a_1191_368.n1 a_1191_368.t0 26.3844
R154 a_1191_368.t6 a_1191_368.n5 26.3844
R155 a_1191_368.n5 a_1191_368.t5 26.3844
R156 A3.n9 A3.t6 360.894
R157 A3.n1 A3.t2 214.758
R158 A3.n8 A3.t0 214.758
R159 A3.n10 A3.t1 214.758
R160 A3.n3 A3.t5 203.171
R161 A3.n7 A3.t3 154.24
R162 A3.n9 A3.t4 154.24
R163 A3.n2 A3.t7 154.24
R164 A3.n4 A3.n3 152
R165 A3.n6 A3.n5 152
R166 A3.n7 A3.n0 152
R167 A3.n12 A3.n11 152
R168 A3.n3 A3.n2 32.7195
R169 A3.n7 A3.n6 32.452
R170 A3.n11 A3.n8 29.1114
R171 A3.n11 A3.n10 13.8401
R172 A3.n12 A3.n0 11.7627
R173 A3.n4 A3 11.5897
R174 A3.n5 A3 9.85996
R175 A3.n6 A3.n1 7.15892
R176 A3.n5 A3 6.74645
R177 A3 A3.n4 5.01672
R178 A3.n8 A3.n7 3.34109
R179 A3 A3.n12 2.94104
R180 A3 A3.n0 1.9032
R181 A3.n2 A3.n1 1.43218
R182 A3.n10 A3.n9 1.43218
R183 a_339_368.t0 a_339_368.n5 462
R184 a_339_368.n1 a_339_368.t7 450.51
R185 a_339_368.n5 a_339_368.n4 305.055
R186 a_339_368.n1 a_339_368.n0 303.534
R187 a_339_368.n3 a_339_368.n2 211.363
R188 a_339_368.n5 a_339_368.n3 50.4476
R189 a_339_368.n3 a_339_368.n1 46.6829
R190 a_339_368.n0 a_339_368.t5 26.3844
R191 a_339_368.n0 a_339_368.t6 26.3844
R192 a_339_368.n2 a_339_368.t2 26.3844
R193 a_339_368.n2 a_339_368.t4 26.3844
R194 a_339_368.n4 a_339_368.t3 26.3844
R195 a_339_368.n4 a_339_368.t1 26.3844
R196 a_788_368.n3 a_788_368.n1 363.43
R197 a_788_368.n4 a_788_368.n0 357.262
R198 a_788_368.n5 a_788_368.n4 309.587
R199 a_788_368.n3 a_788_368.n2 309.389
R200 a_788_368.n4 a_788_368.n3 92.6123
R201 a_788_368.n0 a_788_368.t3 35.1791
R202 a_788_368.n0 a_788_368.t1 35.1791
R203 a_788_368.n1 a_788_368.t7 26.3844
R204 a_788_368.n1 a_788_368.t5 26.3844
R205 a_788_368.n2 a_788_368.t0 26.3844
R206 a_788_368.n2 a_788_368.t6 26.3844
R207 a_788_368.n5 a_788_368.t2 26.3844
R208 a_788_368.t4 a_788_368.n5 26.3844
R209 A4.n1 A4.t7 278.745
R210 A4.n9 A4.t6 247.322
R211 A4.n2 A4.t3 214.758
R212 A4.n0 A4.t4 214.758
R213 A4.n7 A4.t5 214.758
R214 A4.n5 A4.n4 163.762
R215 A4.n6 A4.n5 152
R216 A4.n10 A4.n9 152
R217 A4.n8 A4.t1 142.994
R218 A4.n3 A4.t0 142.994
R219 A4.n1 A4.t2 140.059
R220 A4.n3 A4.n2 29.4561
R221 A4.n6 A4.n0 27.6709
R222 A4.n2 A4.n1 17.2592
R223 A4.n8 A4.n7 14.282
R224 A4.n7 A4.n6 12.4968
R225 A4.n10 A4 8.3032
R226 A4 A4.n10 8.3032
R227 A4.n4 A4.n3 8.03383
R228 A4.n9 A4.n8 3.57087
R229 A4.n5 A4 3.45996
R230 A4.n4 A4.n0 2.67828
R231 VGND.n9 VGND.t10 240.387
R232 VGND.n11 VGND.n10 212.028
R233 VGND.n15 VGND.n14 206.333
R234 VGND.n22 VGND.n21 206.333
R235 VGND.n5 VGND.n4 206.333
R236 VGND.n1 VGND.n0 185
R237 VGND.n28 VGND.n3 132.637
R238 VGND.n0 VGND.t3 48.6491
R239 VGND.n0 VGND.t4 45.4059
R240 VGND.n30 VGND.n29 36.1417
R241 VGND.n10 VGND.t11 34.0546
R242 VGND.n21 VGND.t6 34.0546
R243 VGND.n4 VGND.t8 34.0546
R244 VGND.n27 VGND.n5 33.1299
R245 VGND.n23 VGND.n22 30.8711
R246 VGND.n20 VGND.n7 28.6123
R247 VGND.n14 VGND.t0 28.3789
R248 VGND.n15 VGND.n13 26.3534
R249 VGND.n28 VGND.n27 24.4711
R250 VGND.n10 VGND.t12 22.7032
R251 VGND.n14 VGND.t5 22.7032
R252 VGND.n21 VGND.t7 22.7032
R253 VGND.n4 VGND.t9 22.7032
R254 VGND.n3 VGND.t1 22.7032
R255 VGND.n3 VGND.t2 22.7032
R256 VGND.n13 VGND.n9 21.4593
R257 VGND.n16 VGND.n15 21.0829
R258 VGND.n16 VGND.n7 18.824
R259 VGND.n22 VGND.n20 16.5652
R260 VGND.n30 VGND.n1 14.6471
R261 VGND.n23 VGND.n5 14.3064
R262 VGND.n29 VGND.n28 11.6711
R263 VGND.n31 VGND.n30 9.3005
R264 VGND.n29 VGND.n2 9.3005
R265 VGND.n27 VGND.n26 9.3005
R266 VGND.n25 VGND.n5 9.3005
R267 VGND.n13 VGND.n12 9.3005
R268 VGND.n15 VGND.n8 9.3005
R269 VGND.n17 VGND.n16 9.3005
R270 VGND.n18 VGND.n7 9.3005
R271 VGND.n20 VGND.n19 9.3005
R272 VGND.n22 VGND.n6 9.3005
R273 VGND.n24 VGND.n23 9.3005
R274 VGND.n32 VGND.n1 8.98103
R275 VGND.n11 VGND.n9 6.88087
R276 VGND VGND.n32 0.644923
R277 VGND.n12 VGND.n11 0.513127
R278 VGND.n32 VGND.n31 0.155002
R279 VGND.n12 VGND.n8 0.122949
R280 VGND.n17 VGND.n8 0.122949
R281 VGND.n18 VGND.n17 0.122949
R282 VGND.n19 VGND.n18 0.122949
R283 VGND.n19 VGND.n6 0.122949
R284 VGND.n24 VGND.n6 0.122949
R285 VGND.n25 VGND.n24 0.122949
R286 VGND.n26 VGND.n25 0.122949
R287 VGND.n26 VGND.n2 0.122949
R288 VGND.n31 VGND.n2 0.122949
R289 a_27_74.n5 a_27_74.t15 191.471
R290 a_27_74.n1 a_27_74.t8 191.417
R291 a_27_74.n1 a_27_74.n0 185
R292 a_27_74.n7 a_27_74.t9 141.788
R293 a_27_74.n8 a_27_74.t11 141.036
R294 a_27_74.n6 a_27_74.t0 133.886
R295 a_27_74.n13 a_27_74.n12 102.121
R296 a_27_74.n10 a_27_74.n9 97.4677
R297 a_27_74.n5 a_27_74.n4 96.3134
R298 a_27_74.n12 a_27_74.n11 96.3134
R299 a_27_74.n14 a_27_74.n13 96.2058
R300 a_27_74.n3 a_27_74.n2 88.6891
R301 a_27_74.n13 a_27_74.n3 72.0013
R302 a_27_74.n3 a_27_74.n1 69.9489
R303 a_27_74.n7 a_27_74.n6 60.9887
R304 a_27_74.n8 a_27_74.n7 57.6005
R305 a_27_74.n10 a_27_74.n8 51.2005
R306 a_27_74.n12 a_27_74.n10 51.2005
R307 a_27_74.n6 a_27_74.n5 50.4476
R308 a_27_74.n2 a_27_74.t7 34.0546
R309 a_27_74.t4 a_27_74.n14 26.7573
R310 a_27_74.n2 a_27_74.t3 22.7032
R311 a_27_74.n0 a_27_74.t5 22.7032
R312 a_27_74.n0 a_27_74.t6 22.7032
R313 a_27_74.n11 a_27_74.t12 22.7032
R314 a_27_74.n11 a_27_74.t1 22.7032
R315 a_27_74.n4 a_27_74.t14 22.7032
R316 a_27_74.n4 a_27_74.t16 22.7032
R317 a_27_74.n9 a_27_74.t10 22.7032
R318 a_27_74.n9 a_27_74.t13 22.7032
R319 a_27_74.n14 a_27_74.t2 22.7032
R320 VNB.t11 VNB.t9 3141.21
R321 VNB.t0 VNB.t16 2309.71
R322 VNB.t3 VNB.t4 1686.09
R323 VNB.t14 VNB.t15 1154.86
R324 VNB.t10 VNB.t11 1154.86
R325 VNB.t12 VNB.t13 1154.86
R326 VNB.t7 VNB.t3 1154.86
R327 VNB.t5 VNB.t7 1154.86
R328 VNB VNB.t8 1143.31
R329 VNB.t9 VNB.t0 1074.02
R330 VNB.t4 VNB.t2 1050.92
R331 VNB.t16 VNB.t14 993.177
R332 VNB.t13 VNB.t10 993.177
R333 VNB.t1 VNB.t12 993.177
R334 VNB.t2 VNB.t1 993.177
R335 VNB.t6 VNB.t5 993.177
R336 VNB.t8 VNB.t6 993.177
R337 A2.n3 A2.t1 264.541
R338 A2.n2 A2.t3 261.62
R339 A2.n10 A2.t4 261.62
R340 A2.n13 A2.t5 261.62
R341 A2.n13 A2.n12 163.734
R342 A2.n11 A2.n1 154.24
R343 A2.n8 A2.t0 154.24
R344 A2.n3 A2.t2 154.24
R345 A2.n5 A2.n4 152
R346 A2.n7 A2.n6 152
R347 A2.n9 A2.n0 152
R348 A2.n15 A2.n14 152
R349 A2.n4 A2.n2 47.4702
R350 A2.n9 A2.n8 46.7399
R351 A2.n14 A2.n11 33.5944
R352 A2.n14 A2.n13 29.9429
R353 A2.n4 A2.n3 15.3369
R354 A2.n10 A2.n9 13.8763
R355 A2.n15 A2.n0 11.7627
R356 A2.n6 A2 11.5897
R357 A2.n5 A2 9.85996
R358 A2 A2.n5 6.74645
R359 A2.n6 A2 5.01672
R360 A2 A2.n15 4.67077
R361 A2.n8 A2.n7 2.92171
R362 A2.n7 A2.n2 2.19141
R363 A2.n11 A2.n10 2.19141
R364 A2 A2.n0 0.173473
C0 VPB A2 0.1307f
C1 VPB B1 0.105569f
C2 A4 A3 0.06705f
C3 VPB A1 0.134231f
C4 A3 VPWR 0.026588f
C5 A2 A1 0.084206f
C6 VPB A4 0.138986f
C7 VPB VPWR 0.24259f
C8 A2 VPWR 0.02455f
C9 A3 Y 0.001026f
C10 B1 A4 0.033281f
C11 B1 VPWR 0.078258f
C12 VPB Y 0.023204f
C13 A2 Y 8.09e-20
C14 A1 VPWR 0.089684f
C15 VGND A3 0.068348f
C16 A4 VPWR 0.026296f
C17 B1 Y 0.209363f
C18 A1 Y 4.37e-20
C19 VPB VGND 0.010672f
C20 VGND A2 0.068371f
C21 A4 Y 0.221484f
C22 VPWR Y 0.273263f
C23 B1 VGND 0.023806f
C24 VGND A1 0.067172f
C25 A4 VGND 0.064861f
C26 VGND VPWR 0.159687f
C27 VGND Y 0.024968f
C28 VPB A3 0.158208f
C29 A3 A2 0.067648f
C30 VGND VNB 1.1295f
C31 Y VNB 0.032045f
C32 VPWR VNB 0.937005f
C33 A1 VNB 0.46345f
C34 A2 VNB 0.413264f
C35 A3 VNB 0.436522f
C36 A4 VNB 0.447385f
C37 B1 VNB 0.423301f
C38 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4_2 VNB VPB VPWR VGND Y C D B A
X0 Y.t5 B.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3696 ps=1.78 w=1.12 l=0.15
X1 a_27_74.t1 C.t0 a_304_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.23225 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_515_74.t1 A.t0 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.22325 pd=2.15 as=0.111 ps=1.04 w=0.74 l=0.15
X3 VPWR.t0 D.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.1904 ps=1.46 w=1.12 l=0.15
X4 Y.t9 D.t1 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.336 ps=2.84 w=1.12 l=0.15
X5 VPWR.t5 C.t1 Y.t6 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3696 pd=1.78 as=0.1792 ps=1.44 w=1.12 l=0.15
X6 VGND.t1 D.t2 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1369 pd=1.11 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 a_304_74.t1 C.t2 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 Y.t8 A.t1 a_515_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 Y.t7 C.t3 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.1904 ps=1.46 w=1.12 l=0.15
X10 a_27_74.t2 D.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1369 ps=1.11 w=0.74 l=0.15
X11 a_304_74.t2 B.t1 a_515_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1983 ps=2.05 w=0.74 l=0.15
X12 VPWR.t2 A.t2 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X13 Y.t1 A.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2296 ps=1.53 w=1.12 l=0.15
X14 a_515_74.t2 B.t2 a_304_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VPWR.t3 B.t3 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2296 pd=1.53 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B.n0 B.t0 237.762
R1 B.n2 B.t3 226.809
R2 B.n3 B.t2 209.16
R3 B.n1 B.t1 196.013
R4 B.n0 B 157.656
R5 B.n4 B.n3 152
R6 B.n2 B.n1 41.6278
R7 B.n1 B.n0 13.146
R8 B.n3 B.n2 8.03383
R9 B B.n4 7.14469
R10 B.n4 B 7.14469
R11 VPWR.n5 VPWR.t2 349.962
R12 VPWR.n13 VPWR.n2 316.353
R13 VPWR.n7 VPWR.n6 316.353
R14 VPWR.n15 VPWR.t7 249.968
R15 VPWR.n4 VPWR.n3 145.525
R16 VPWR.n3 VPWR.t5 54.9544
R17 VPWR.n3 VPWR.t4 54.9541
R18 VPWR.n6 VPWR.t1 36.938
R19 VPWR.n8 VPWR.n4 35.3887
R20 VPWR.n6 VPWR.t3 35.1791
R21 VPWR.n2 VPWR.t6 31.6612
R22 VPWR.n12 VPWR.n4 30.1181
R23 VPWR.n2 VPWR.t0 28.1434
R24 VPWR.n14 VPWR.n13 26.3534
R25 VPWR.n13 VPWR.n12 21.0829
R26 VPWR.n15 VPWR.n14 20.3299
R27 VPWR.n8 VPWR.n7 15.8123
R28 VPWR.n9 VPWR.n8 9.3005
R29 VPWR.n12 VPWR.n11 9.3005
R30 VPWR.n13 VPWR.n1 9.3005
R31 VPWR.n14 VPWR.n0 9.3005
R32 VPWR.n16 VPWR.n15 9.3005
R33 VPWR.n7 VPWR.n5 6.98267
R34 VPWR.n10 VPWR.n4 4.62059
R35 VPWR.n9 VPWR.n5 0.63499
R36 VPWR.n10 VPWR.n9 0.184273
R37 VPWR.n11 VPWR.n10 0.184273
R38 VPWR.n11 VPWR.n1 0.122949
R39 VPWR.n1 VPWR.n0 0.122949
R40 VPWR.n16 VPWR.n0 0.122949
R41 VPWR VPWR.n16 0.0617245
R42 Y.n2 Y.n0 258.303
R43 Y Y.n7 222.785
R44 Y.n6 Y.n5 204.101
R45 Y.n2 Y.n1 203.27
R46 Y.n4 Y.n3 203.27
R47 Y.n4 Y.n2 70.024
R48 Y.n6 Y.n4 51.6391
R49 Y.n0 Y.t0 33.4201
R50 Y.n1 Y.t7 29.9023
R51 Y.n0 Y.t9 26.3844
R52 Y.n1 Y.t6 26.3844
R53 Y.n3 Y.t4 26.3844
R54 Y.n3 Y.t5 26.3844
R55 Y.n5 Y.t2 26.3844
R56 Y.n5 Y.t1 26.3844
R57 Y Y.n6 26.2813
R58 Y.n7 Y.t3 25.9464
R59 Y.n7 Y.t8 22.7032
R60 VPB.t5 VPB.t4 413.711
R61 VPB.t3 VPB.t1 286.022
R62 VPB VPB.t7 260.485
R63 VPB.t0 VPB.t6 250.269
R64 VPB.t7 VPB.t0 250.269
R65 VPB.t6 VPB.t5 240.054
R66 VPB.t1 VPB.t2 229.839
R67 VPB.t4 VPB.t3 229.839
R68 C.n0 C.t1 226.809
R69 C.n1 C.t3 226.809
R70 C C.n0 203.964
R71 C.n1 C.t2 203.762
R72 C.n3 C.t0 196.013
R73 C.n5 C.n4 152
R74 C.n2 C 152
R75 C.n3 C.n2 40.8975
R76 C.n2 C.n1 15.3369
R77 C.n5 C 10.1214
R78 C.n4 C.n3 8.76414
R79 C C.n5 4.16794
R80 C.n4 C.n0 3.65202
R81 a_304_74.n1 a_304_74.n0 477.512
R82 a_304_74.n0 a_304_74.t3 22.7032
R83 a_304_74.n0 a_304_74.t2 22.7032
R84 a_304_74.t0 a_304_74.n1 22.7032
R85 a_304_74.n1 a_304_74.t1 22.7032
R86 a_27_74.n2 a_27_74.n1 297.454
R87 a_27_74.n1 a_27_74.t3 227.159
R88 a_27_74.n1 a_27_74.n0 84.741
R89 a_27_74.n3 a_27_74.n2 69.6005
R90 a_27_74.n0 a_27_74.t0 22.7032
R91 a_27_74.n0 a_27_74.t2 22.7032
R92 a_27_74.n2 a_27_74.t1 17.8444
R93 VNB.t1 VNB.t6 2448.29
R94 VNB.t3 VNB.t2 1201.05
R95 VNB VNB.t3 1143.31
R96 VNB.t7 VNB.t4 1039.37
R97 VNB.t5 VNB.t7 993.177
R98 VNB.t6 VNB.t5 993.177
R99 VNB.t0 VNB.t1 993.177
R100 VNB.t2 VNB.t0 993.177
R101 A.n1 A.t3 228.877
R102 A.n0 A.t2 226.809
R103 A.n0 A.t0 198.204
R104 A.n1 A.t1 196.013
R105 A A.n2 154.522
R106 A.n2 A.n1 37.246
R107 A.n2 A.n0 26.2914
R108 a_515_74.n1 a_515_74.t3 274.486
R109 a_515_74.n2 a_515_74.n1 262.671
R110 a_515_74.n1 a_515_74.n0 111.294
R111 a_515_74.n3 a_515_74.n2 69.6005
R112 a_515_74.n0 a_515_74.t0 22.7032
R113 a_515_74.n0 a_515_74.t2 22.7032
R114 a_515_74.n2 a_515_74.t1 17.8444
R115 D.n0 D.t0 226.809
R116 D.n2 D.t1 226.809
R117 D.n2 D.t2 198.204
R118 D.n0 D.t3 198.204
R119 D D.n1 160.633
R120 D.n4 D.n3 152
R121 D.n3 D.n1 49.6611
R122 D.n4 D 12.8005
R123 D.n1 D.n0 10.955
R124 D.n3 D.n2 10.955
R125 D D.n4 1.48887
R126 VGND VGND.n0 215.621
R127 VGND.n0 VGND.t1 34.0546
R128 VGND.n0 VGND.t0 25.9464
C0 VPB VGND 0.0072f
C1 C B 0.065205f
C2 D VPWR 0.07506f
C3 C VPWR 0.043359f
C4 D Y 0.068759f
C5 B A 0.094837f
C6 D VGND 0.035529f
C7 C Y 0.126621f
C8 B VPWR 0.037909f
C9 B Y 0.126813f
C10 C VGND 0.014615f
C11 A VPWR 0.037135f
C12 A Y 0.164599f
C13 B VGND 0.013808f
C14 D VPB 0.070397f
C15 VPWR Y 0.825586f
C16 A VGND 0.012282f
C17 C VPB 0.088365f
C18 VPWR VGND 0.080192f
C19 B VPB 0.073539f
C20 Y VGND 0.017642f
C21 A VPB 0.064387f
C22 VPB VPWR 0.141782f
C23 VPB Y 0.022849f
C24 D C 0.076674f
C25 VGND VNB 0.566902f
C26 Y VNB 0.076642f
C27 VPWR VNB 0.514414f
C28 A VNB 0.216854f
C29 B VNB 0.211396f
C30 C VNB 0.23989f
C31 D VNB 0.248389f
C32 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4_4 VNB VPB VPWR VGND C D A Y B
X0 VPWR.t3 C.t0 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.4872 pd=1.99 as=0.3808 ps=1.8 w=1.12 l=0.15
X1 Y.t0 B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.4872 ps=1.99 w=1.12 l=0.15
X2 Y.t8 D.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=1.736 ps=5.34 w=1.12 l=0.15
X3 a_923_74.t7 A.t0 Y.t2 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t3 D.t1 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_27_74.t4 C.t1 a_554_74.t7 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.19515 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_27_74.t6 C.t2 a_554_74.t6 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 Y.t5 A.t1 a_923_74.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VGND.t2 D.t2 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=1.29 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 Y.t6 A.t2 a_923_74.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_923_74.t4 A.t3 Y.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1962 pd=2.05 as=0.1628 ps=1.18 w=0.74 l=0.15
X11 a_554_74.t5 C.t3 a_27_74.t7 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_554_74.t3 B.t1 a_923_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_554_74.t4 C.t4 a_27_74.t5 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X14 VPWR.t1 B.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.9296 pd=2.78 as=0.3808 ps=1.8 w=1.12 l=0.15
X15 a_27_74.t1 D.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 a_923_74.t3 B.t3 a_554_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_554_74.t1 B.t4 a_923_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1969 ps=2.05 w=0.74 l=0.15
X18 Y.t3 C.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VPWR.t6 A.t4 Y.t10 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.4368 ps=1.9 w=1.12 l=0.15
X20 a_27_74.t0 D.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2035 ps=1.29 w=0.74 l=0.15
X21 VPWR.t5 D.t5 Y.t9 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.4368 pd=1.9 as=0.9296 ps=2.78 w=1.12 l=0.15
X23 a_923_74.t0 B.t5 a_554_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 C.n7 C.t0 226.809
R1 C.n1 C.t5 226.809
R2 C.n9 C.t1 222.304
R3 C.n1 C.t4 198.204
R4 C.n0 C.t2 196.013
R5 C.n8 C.t3 196.013
R6 C.n10 C.n9 152
R7 C.n6 C.n5 152
R8 C.n4 C.n0 152
R9 C.n3 C.n2 152
R10 C.n6 C.n0 49.6611
R11 C.n2 C.n0 49.6611
R12 C.n9 C.n8 36.5157
R13 C.n7 C.n6 10.955
R14 C.n2 C.n1 10.955
R15 C.n5 C.n4 10.1214
R16 C.n10 C 8.63306
R17 C C.n3 7.44236
R18 C.n3 C 6.84701
R19 C C.n10 5.65631
R20 C.n4 C 2.67957
R21 C.n8 C.n7 2.19141
R22 C.n5 C 1.48887
R23 Y.n15 Y.n14 585
R24 Y.n14 Y.n12 585
R25 Y.n16 Y.n15 585
R26 Y.n16 Y.n12 585
R27 Y.n3 Y.n1 292.502
R28 Y.n8 Y.n6 292.502
R29 Y.n2 Y.n1 292.5
R30 Y.n7 Y.n6 292.5
R31 Y.n5 Y.n4 276.695
R32 Y.n10 Y.n9 276.695
R33 Y.n13 Y.n11 272.815
R34 Y.n5 Y.n0 253.53
R35 Y.n19 Y.n17 233.129
R36 Y.n19 Y.n18 185
R37 Y.n16 Y.n10 153.601
R38 Y.n10 Y.n5 93.3652
R39 Y Y.n16 46.0281
R40 Y.n15 Y.n13 39.3741
R41 Y.n13 Y.n12 39.3741
R42 Y.n18 Y.t7 35.6762
R43 Y.n18 Y.t5 35.6762
R44 Y.n0 Y.t9 35.1791
R45 Y Y.n19 32.6127
R46 Y.n4 Y.n3 31.6146
R47 Y.n4 Y.n2 31.6146
R48 Y.n9 Y.n8 31.6146
R49 Y.n9 Y.n7 31.6146
R50 Y.n0 Y.t8 26.3844
R51 Y.n2 Y.t4 26.3844
R52 Y.n3 Y.t3 26.3844
R53 Y.n7 Y.t1 26.3844
R54 Y.n8 Y.t0 26.3844
R55 Y.n12 Y.t10 26.3844
R56 Y.n17 Y.t2 22.7032
R57 Y.n17 Y.t6 22.7032
R58 Y.n5 Y.n1 10.0437
R59 Y.n10 Y.n6 10.0437
R60 Y.n14 Y.n11 7.42079
R61 Y.n16 Y.n11 7.04978
R62 VPWR.n20 VPWR.n14 352.305
R63 VPWR.n15 VPWR.t6 349.438
R64 VPWR.n35 VPWR.n7 315.928
R65 VPWR.n22 VPWR.n11 292.5
R66 VPWR.n24 VPWR.n23 292.5
R67 VPWR.n21 VPWR.n13 292.5
R68 VPWR.n20 VPWR.n19 292.5
R69 VPWR.n44 VPWR.n43 265.358
R70 VPWR.n4 VPWR.n3 195
R71 VPWR.n41 VPWR.n2 195
R72 VPWR.n43 VPWR.n42 195
R73 VPWR.n9 VPWR.n8 133.587
R74 VPWR.n43 VPWR.n2 71.2371
R75 VPWR.n3 VPWR.n2 70.3576
R76 VPWR.n8 VPWR.t3 69.1811
R77 VPWR.n8 VPWR.t0 69.1808
R78 VPWR.n21 VPWR.n20 59.8041
R79 VPWR.n23 VPWR.n21 59.8041
R80 VPWR.n23 VPWR.n22 59.8041
R81 VPWR.n37 VPWR.n36 36.1417
R82 VPWR.n34 VPWR.n9 36.1417
R83 VPWR.n30 VPWR.n29 36.1417
R84 VPWR.n35 VPWR.n34 35.3887
R85 VPWR.n15 VPWR.n14 31.7058
R86 VPWR.n29 VPWR.n28 31.6675
R87 VPWR.n3 VPWR.t4 27.2639
R88 VPWR.n22 VPWR.t1 26.3844
R89 VPWR.n7 VPWR.t2 26.3844
R90 VPWR.n7 VPWR.t5 26.3844
R91 VPWR.n36 VPWR.n35 12.0476
R92 VPWR.n45 VPWR.n44 10.0432
R93 VPWR.n17 VPWR.n16 9.3005
R94 VPWR.n18 VPWR.n12 9.3005
R95 VPWR.n26 VPWR.n25 9.3005
R96 VPWR.n28 VPWR.n27 9.3005
R97 VPWR.n29 VPWR.n10 9.3005
R98 VPWR.n31 VPWR.n30 9.3005
R99 VPWR.n34 VPWR.n33 9.3005
R100 VPWR.n35 VPWR.n6 9.3005
R101 VPWR.n36 VPWR.n5 9.3005
R102 VPWR.n38 VPWR.n37 9.3005
R103 VPWR.n40 VPWR.n39 9.3005
R104 VPWR.n1 VPWR.n0 9.3005
R105 VPWR.n32 VPWR.n9 4.62059
R106 VPWR.n30 VPWR.n9 4.51815
R107 VPWR.n24 VPWR.n11 3.86894
R108 VPWR.n19 VPWR.n17 3.69828
R109 VPWR.n42 VPWR.n41 3.53907
R110 VPWR.n44 VPWR.n1 3.45169
R111 VPWR.n25 VPWR.n13 3.35694
R112 VPWR.n37 VPWR.n4 3.30779
R113 VPWR.n40 VPWR.n4 2.88378
R114 VPWR.n18 VPWR.n13 2.10539
R115 VPWR.n19 VPWR.n18 1.76406
R116 VPWR.n28 VPWR.n11 1.08139
R117 VPWR.n41 VPWR.n40 0.612104
R118 VPWR.n16 VPWR.n15 0.541527
R119 VPWR.n25 VPWR.n24 0.5125
R120 VPWR.n32 VPWR.n31 0.184273
R121 VPWR.n33 VPWR.n32 0.184273
R122 VPWR.n17 VPWR.n14 0.171167
R123 VPWR.n16 VPWR.n12 0.122949
R124 VPWR.n26 VPWR.n12 0.122949
R125 VPWR.n27 VPWR.n26 0.122949
R126 VPWR.n27 VPWR.n10 0.122949
R127 VPWR.n31 VPWR.n10 0.122949
R128 VPWR.n33 VPWR.n6 0.122949
R129 VPWR.n6 VPWR.n5 0.122949
R130 VPWR.n38 VPWR.n5 0.122949
R131 VPWR.n39 VPWR.n38 0.122949
R132 VPWR.n39 VPWR.n0 0.122949
R133 VPWR.n45 VPWR.n0 0.122949
R134 VPWR VPWR.n45 0.0617245
R135 VPWR.n42 VPWR.n1 0.044186
R136 VPB.t1 VPB.t6 1399.46
R137 VPB VPB.t4 898.926
R138 VPB.t3 VPB.t0 520.968
R139 VPB.t0 VPB.t1 423.925
R140 VPB.t2 VPB.t3 423.925
R141 VPB.t4 VPB.t5 255.376
R142 VPB.t5 VPB.t2 229.839
R143 B.n3 B.t0 237.762
R144 B.n0 B.t3 235.451
R145 B.n8 B.t2 226.809
R146 B.n2 B.t4 196.013
R147 B.n9 B.t5 196.013
R148 B.n1 B.t1 196.013
R149 B B.n0 154.381
R150 B.n11 B.n10 152
R151 B.n7 B.n6 152
R152 B.n5 B.n2 152
R153 B.n4 B.n3 152
R154 B.n7 B.n2 49.6611
R155 B.n3 B.n2 49.6611
R156 B.n10 B.n9 36.5157
R157 B.n10 B.n1 26.2914
R158 B.n1 B.n0 23.3702
R159 B.n8 B.n7 10.955
R160 B.n6 B.n5 10.1214
R161 B B.n4 9.52608
R162 B B.n11 7.74003
R163 B.n11 B 6.54934
R164 B.n4 B 4.76329
R165 B.n6 B 3.57259
R166 B.n9 B.n8 2.19141
R167 B.n5 B 0.595849
R168 D.n0 D.t5 236.303
R169 D.n4 D.t1 232.53
R170 D.n10 D.t0 226.809
R171 D.n3 D.t3 196.013
R172 D.n9 D.t2 196.013
R173 D.n0 D.t4 196.013
R174 D D.n1 152.893
R175 D.n12 D.n11 152
R176 D.n8 D.n7 152
R177 D.n6 D.n2 152
R178 D.n5 D.n4 152
R179 D.n11 D.n1 49.6611
R180 D.n8 D.n2 49.6611
R181 D.n10 D.n9 38.7066
R182 D.n4 D.n3 36.5157
R183 D.n1 D.n0 13.146
R184 D.n3 D.n2 13.146
R185 D.n9 D.n8 10.2247
R186 D.n6 D.n5 10.1214
R187 D D.n12 9.22841
R188 D.n7 D 9.22841
R189 D.n12 D 5.06097
R190 D.n7 D 5.06097
R191 D.n5 D 3.27492
R192 D D.n6 0.893523
R193 D.n11 D.n10 0.730803
R194 A.n0 A.t4 226.809
R195 A.n3 A.n2 226.809
R196 A.n5 A.t2 225.957
R197 A.n0 A.t3 198.204
R198 A.n4 A.t0 196.013
R199 A.n9 A.t1 196.013
R200 A A.n1 154.53
R201 A.n11 A.n10 152
R202 A.n8 A.n7 152
R203 A.n6 A.n5 152
R204 A.n10 A.n1 49.6611
R205 A.n9 A.n8 46.0096
R206 A.n5 A.n4 32.8641
R207 A.n1 A.n0 30.6732
R208 A.n4 A.n3 10.955
R209 A.n7 A.n6 10.1214
R210 A A.n11 7.5912
R211 A.n11 A 6.69817
R212 A.n8 A.n3 5.84292
R213 A.n10 A.n9 3.65202
R214 A.n7 A 3.42376
R215 A.n6 A 0.744686
R216 a_923_74.n4 a_923_74.t4 274.582
R217 a_923_74.n1 a_923_74.t2 262.204
R218 a_923_74.n1 a_923_74.n0 185
R219 a_923_74.n3 a_923_74.n2 185
R220 a_923_74.n5 a_923_74.n4 185
R221 a_923_74.n3 a_923_74.n1 51.6397
R222 a_923_74.n4 a_923_74.n3 51.6397
R223 a_923_74.n2 a_923_74.t5 22.7032
R224 a_923_74.n2 a_923_74.t3 22.7032
R225 a_923_74.n0 a_923_74.t1 22.7032
R226 a_923_74.n0 a_923_74.t0 22.7032
R227 a_923_74.t6 a_923_74.n5 22.7032
R228 a_923_74.n5 a_923_74.t7 22.7032
R229 VNB.t15 VNB.t5 2286.61
R230 VNB.t2 VNB.t0 1616.8
R231 VNB.t10 VNB.t8 1362.73
R232 VNB.t0 VNB.t12 1154.86
R233 VNB.t1 VNB.t2 1154.86
R234 VNB.t3 VNB.t1 1154.86
R235 VNB VNB.t3 1143.31
R236 VNB.t11 VNB.t10 993.177
R237 VNB.t9 VNB.t11 993.177
R238 VNB.t6 VNB.t9 993.177
R239 VNB.t7 VNB.t6 993.177
R240 VNB.t4 VNB.t7 993.177
R241 VNB.t5 VNB.t4 993.177
R242 VNB.t13 VNB.t15 993.177
R243 VNB.t14 VNB.t13 993.177
R244 VNB.t12 VNB.t14 993.177
R245 a_27_74.n3 a_27_74.t4 244.835
R246 a_27_74.n1 a_27_74.t3 199.591
R247 a_27_74.n3 a_27_74.n2 185
R248 a_27_74.n1 a_27_74.n0 101.71
R249 a_27_74.n5 a_27_74.n4 89.8175
R250 a_27_74.n4 a_27_74.n1 70.6456
R251 a_27_74.n4 a_27_74.n3 41.4406
R252 a_27_74.n0 a_27_74.t1 34.0546
R253 a_27_74.n5 a_27_74.t5 34.0546
R254 a_27_74.n0 a_27_74.t2 22.7032
R255 a_27_74.n2 a_27_74.t7 22.7032
R256 a_27_74.n2 a_27_74.t6 22.7032
R257 a_27_74.t0 a_27_74.n5 22.7032
R258 VGND.n2 VGND.n0 216.785
R259 VGND.n2 VGND.n1 216.68
R260 VGND.n0 VGND.t0 55.1356
R261 VGND.n0 VGND.t2 34.0546
R262 VGND.n1 VGND.t3 34.0546
R263 VGND.n1 VGND.t1 22.7032
R264 VGND VGND.n2 0.483401
R265 a_554_74.n5 a_554_74.n4 229.032
R266 a_554_74.n2 a_554_74.n0 224.315
R267 a_554_74.n2 a_554_74.n1 185
R268 a_554_74.n4 a_554_74.n3 185
R269 a_554_74.n4 a_554_74.n2 71.7994
R270 a_554_74.n3 a_554_74.t0 22.7032
R271 a_554_74.n3 a_554_74.t1 22.7032
R272 a_554_74.n0 a_554_74.t6 22.7032
R273 a_554_74.n0 a_554_74.t4 22.7032
R274 a_554_74.n1 a_554_74.t7 22.7032
R275 a_554_74.n1 a_554_74.t5 22.7032
R276 a_554_74.n5 a_554_74.t2 22.7032
R277 a_554_74.t3 a_554_74.n5 22.7032
C0 VPWR Y 1.11826f
C1 VPB Y 0.030245f
C2 D VPWR 0.194778f
C3 VPB D 0.141083f
C4 VPWR VGND 0.148095f
C5 D Y 0.070983f
C6 VPB VGND 0.009539f
C7 C VPWR 0.044611f
C8 VPB C 0.118164f
C9 Y VGND 0.031344f
C10 B VPWR 0.050725f
C11 C Y 0.182074f
C12 D VGND 0.066321f
C13 D C 0.083321f
C14 VPB B 0.147411f
C15 C VGND 0.02244f
C16 B Y 0.192252f
C17 A VPWR 0.049474f
C18 VPB A 0.132643f
C19 A Y 0.342747f
C20 B VGND 0.02736f
C21 C B 0.055408f
C22 A VGND 0.02637f
C23 B A 0.061828f
C24 VPB VPWR 0.230836f
C25 VGND VNB 0.974056f
C26 Y VNB 0.083651f
C27 VPWR VNB 0.809734f
C28 A VNB 0.395533f
C29 B VNB 0.395508f
C30 C VNB 0.355934f
C31 D VNB 0.452898f
C32 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4b_1 VNB VPB VPWR VGND A_N D Y C B
X0 a_341_74.t0 C.t0 a_263_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 VPWR.t2 C.t1 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t0 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.231 ps=1.555 w=1.12 l=0.15
X3 VPWR.t3 a_27_112.t2 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t3 B.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2352 ps=1.54 w=1.12 l=0.15
X5 VPWR.t0 A_N.t0 a_27_112.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 a_263_74.t0 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1348 ps=1.13 w=0.74 l=0.15
X7 a_443_74.t0 B.t1 a_341_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1332 ps=1.1 w=0.74 l=0.15
X8 Y.t4 a_27_112.t3 a_443_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.3404 pd=2.4 as=0.1443 ps=1.13 w=0.74 l=0.15
X9 VGND.t1 A_N.t1 a_27_112.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1348 pd=1.13 as=0.2695 ps=2.08 w=0.55 l=0.15
R0 C.n0 C.t1 285.719
R1 C.n0 C.t0 178.34
R2 C C.n0 158.788
R3 a_263_74.t0 a_263_74.t1 38.9194
R4 a_341_74.t0 a_341_74.t1 58.3789
R5 VNB VNB.t3 1616.8
R6 VNB.t2 VNB.t4 1247.24
R7 VNB.t3 VNB.t0 1247.24
R8 VNB.t1 VNB.t2 1177.95
R9 VNB.t0 VNB.t1 900.788
R10 Y.n1 Y.t4 236.754
R11 Y Y.n2 217.413
R12 Y.n1 Y.n0 200.579
R13 Y.n2 Y.t1 26.3844
R14 Y.n2 Y.t0 26.3844
R15 Y.n0 Y.t2 26.3844
R16 Y.n0 Y.t3 26.3844
R17 Y Y.n1 11.5635
R18 VPWR.n3 VPWR.n2 316.399
R19 VPWR.n4 VPWR.t3 262.95
R20 VPWR.n8 VPWR.n1 231.036
R21 VPWR.n1 VPWR.t0 56.9831
R22 VPWR.n2 VPWR.t4 38.6969
R23 VPWR.n1 VPWR.t1 36.6184
R24 VPWR.n7 VPWR.n6 36.1417
R25 VPWR.n2 VPWR.t2 35.1791
R26 VPWR.n9 VPWR.n8 12.5979
R27 VPWR.n4 VPWR.n3 10.5045
R28 VPWR.n6 VPWR.n5 9.3005
R29 VPWR.n7 VPWR.n0 9.3005
R30 VPWR.n6 VPWR.n3 7.90638
R31 VPWR.n8 VPWR.n7 6.4005
R32 VPWR.n5 VPWR.n4 0.647735
R33 VPWR VPWR.n9 0.163644
R34 VPWR.n9 VPWR.n0 0.144205
R35 VPWR.n5 VPWR.n0 0.122949
R36 VPB VPB.t0 326.882
R37 VPB.t0 VPB.t1 298.791
R38 VPB.t2 VPB.t4 291.13
R39 VPB.t4 VPB.t3 229.839
R40 VPB.t1 VPB.t2 229.839
R41 D.n0 D.t0 285.719
R42 D.n0 D.t1 178.34
R43 D D.n0 158.788
R44 a_27_112.t0 a_27_112.n1 464.87
R45 a_27_112.n1 a_27_112.n0 330.509
R46 a_27_112.n0 a_27_112.t2 285.719
R47 a_27_112.n1 a_27_112.t1 215.546
R48 a_27_112.n0 a_27_112.t3 178.34
R49 B.n0 B.t0 285.719
R50 B.n0 B.t1 178.34
R51 B B.n0 158.4
R52 A_N.n0 A_N.t0 240.732
R53 A_N A_N.n0 158.054
R54 A_N.n0 A_N.t1 147.814
R55 VGND VGND.n0 216.599
R56 VGND.n0 VGND.t1 53.455
R57 VGND.n0 VGND.t0 22.2054
R58 a_443_74.t0 a_443_74.t1 63.2437
C0 VPWR Y 0.45044f
C1 VPWR C 0.01392f
C2 Y VPB 0.021146f
C3 A_N D 0.071893f
C4 VPB C 0.030512f
C5 A_N Y 0.001016f
C6 Y D 0.015163f
C7 D C 0.091805f
C8 Y C 0.050945f
C9 B VGND 0.007695f
C10 VPWR VGND 0.055912f
C11 B VPWR 0.013944f
C12 VGND VPB 0.007501f
C13 B VPB 0.030408f
C14 A_N VGND 0.009283f
C15 VGND D 0.014412f
C16 VPWR VPB 0.112499f
C17 Y VGND 0.053592f
C18 VPWR A_N 0.021568f
C19 B Y 0.05601f
C20 VGND C 0.009785f
C21 VPWR D 0.031473f
C22 B C 0.081362f
C23 A_N VPB 0.041234f
C24 VPB D 0.033379f
C25 VGND VNB 0.448087f
C26 Y VNB 0.092909f
C27 A_N VNB 0.140541f
C28 VPWR VNB 0.391945f
C29 B VNB 0.105474f
C30 C VNB 0.103549f
C31 D VNB 0.10938f
C32 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4b_2 VNB VPB VPWR VGND Y A_N D C B
X0 a_719_123.t3 D.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.111 ps=1.04 w=0.74 l=0.15
X1 a_225_74.t1 a_27_74.t2 Y.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1147 ps=1.05 w=0.74 l=0.15
X2 VGND.t2 A_N.t0 a_27_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1726 pd=1.85 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 a_719_123.t1 C.t0 a_490_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_225_74.t2 B.t0 a_490_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.197775 pd=2.05 as=0.1773 ps=1.28 w=0.74 l=0.15
X5 VPWR.t8 B.t1 Y.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t6 A_N.t1 a_27_74.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.213 pd=1.51 as=0.295 ps=2.59 w=1 l=0.15
X7 Y.t8 B.t2 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3724 ps=1.785 w=1.12 l=0.15
X8 VGND.t0 D.t1 a_719_123.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t3 a_27_74.t3 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3724 pd=1.785 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t1 a_27_74.t4 a_225_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.1962 ps=2.05 w=0.74 l=0.15
X11 Y.t2 a_27_74.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.213 ps=1.51 w=1.12 l=0.15
X12 a_490_74.t0 C.t1 a_719_123.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.204075 ps=2.05 w=0.74 l=0.15
X13 a_490_74.t3 B.t3 a_225_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1773 pd=1.28 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 Y.t6 D.t2 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.28 ps=1.62 w=1.12 l=0.15
X15 VPWR.t1 C.t2 Y.t9 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.28 pd=1.62 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VPWR.t4 D.t3 Y.t5 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.168 ps=1.42 w=1.12 l=0.15
X17 Y.t0 C.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
R0 D.n1 D.t2 228.877
R1 D.n0 D.t3 226.809
R2 D.n0 D.t0 182.138
R3 D.n1 D.t1 179.947
R4 D.n3 D.n2 152
R5 D.n2 D.n0 50.3914
R6 D.n2 D.n1 13.146
R7 D.n3 D 12.8005
R8 D D.n3 1.48887
R9 VGND.n1 VGND.t2 240.626
R10 VGND.n1 VGND.n0 214.44
R11 VGND.n0 VGND.t1 25.9464
R12 VGND.n0 VGND.t0 22.7032
R13 VGND VGND.n1 0.189719
R14 a_719_123.n0 a_719_123.t0 257.418
R15 a_719_123.n0 a_719_123.t3 189.924
R16 a_719_123.n1 a_719_123.n0 98.2658
R17 a_719_123.t2 a_719_123.n1 22.7032
R18 a_719_123.n1 a_719_123.t1 22.7032
R19 VNB.t4 VNB.t0 2286.61
R20 VNB.t8 VNB.t7 2286.61
R21 VNB.t5 VNB.t4 1362.73
R22 VNB VNB.t8 1143.31
R23 VNB.t7 VNB.t6 1062.47
R24 VNB.t2 VNB.t3 1039.37
R25 VNB.t1 VNB.t2 993.177
R26 VNB.t0 VNB.t1 993.177
R27 VNB.t6 VNB.t5 993.177
R28 a_27_74.n3 a_27_74.t0 319.014
R29 a_27_74.t1 a_27_74.n3 274.803
R30 a_27_74.n1 a_27_74.t5 234.112
R31 a_27_74.n0 a_27_74.t3 226.809
R32 a_27_74.n0 a_27_74.t2 204.778
R33 a_27_74.n1 a_27_74.t4 196.013
R34 a_27_74.n3 a_27_74.n2 152
R35 a_27_74.n2 a_27_74.n0 48.2005
R36 a_27_74.n2 a_27_74.n1 10.2247
R37 Y.n5 Y.n4 282.209
R38 Y Y.n7 281.041
R39 Y.n2 Y.n0 261.06
R40 Y.n2 Y.n1 203.083
R41 Y.n5 Y.n3 201.483
R42 Y.n6 Y.n2 44.4366
R43 Y.n3 Y.t7 26.3844
R44 Y.n3 Y.t8 26.3844
R45 Y.n4 Y.t4 26.3844
R46 Y.n4 Y.t2 26.3844
R47 Y.n0 Y.t5 26.3844
R48 Y.n0 Y.t6 26.3844
R49 Y.n1 Y.t9 26.3844
R50 Y.n1 Y.t0 26.3844
R51 Y.n7 Y.t3 25.1356
R52 Y.n7 Y.t1 25.1356
R53 Y Y.n6 13.357
R54 Y.n6 Y.n5 8.3205
R55 a_225_74.n0 a_225_74.t2 280.998
R56 a_225_74.n0 a_225_74.t0 251.582
R57 a_225_74.n1 a_225_74.n0 185
R58 a_225_74.n1 a_225_74.t3 22.7032
R59 a_225_74.t1 a_225_74.n1 22.7032
R60 A_N.n0 A_N.t1 264.005
R61 A_N.n0 A_N 159.177
R62 A_N.n1 A_N.t0 157.453
R63 A_N.n2 A_N.n1 154.191
R64 A_N.n1 A_N.n0 47.4702
R65 A_N A_N.n2 12.6066
R66 A_N.n2 A_N 6.01262
R67 C.n0 C.t0 239.685
R68 C.n0 C.t2 226.809
R69 C.n3 C.t3 226.809
R70 C.n2 C.t1 179.947
R71 C.n4 C.n3 153.462
R72 C C.n1 153.042
R73 C.n3 C.n2 37.246
R74 C.n1 C.n0 17.5278
R75 C.n2 C.n1 10.955
R76 C C.n4 9.07957
R77 C.n4 C 5.2098
R78 a_490_74.n1 a_490_74.n0 476.024
R79 a_490_74.n0 a_490_74.t2 35.6762
R80 a_490_74.n0 a_490_74.t3 35.6762
R81 a_490_74.t1 a_490_74.n1 22.7032
R82 a_490_74.n1 a_490_74.t0 22.7032
R83 B.n0 B.t1 253.829
R84 B.n1 B.t2 226.809
R85 B.n2 B.t3 203.316
R86 B.n0 B.t0 196.013
R87 B B.n2 162.419
R88 B.n2 B.n1 40.1672
R89 B.n1 B.n0 38.7066
R90 VPWR.n8 VPWR.n7 316.353
R91 VPWR.n11 VPWR.n10 316.305
R92 VPWR.n6 VPWR.t4 260.113
R93 VPWR.n1 VPWR.n0 223.316
R94 VPWR.n17 VPWR.n3 144.778
R95 VPWR.n3 VPWR.t3 55.312
R96 VPWR.n3 VPWR.t7 55.3117
R97 VPWR.n0 VPWR.t6 46.2955
R98 VPWR.n7 VPWR.t1 45.7326
R99 VPWR.n7 VPWR.t5 42.2148
R100 VPWR.n16 VPWR.n4 36.1417
R101 VPWR.n12 VPWR.n9 36.1417
R102 VPWR.n10 VPWR.t0 35.1791
R103 VPWR.n10 VPWR.t8 35.1791
R104 VPWR.n0 VPWR.t2 27.7937
R105 VPWR.n18 VPWR.n17 23.7181
R106 VPWR.n18 VPWR.n1 23.3417
R107 VPWR.n9 VPWR.n8 18.0711
R108 VPWR.n11 VPWR.n4 10.5417
R109 VPWR.n9 VPWR.n5 9.3005
R110 VPWR.n13 VPWR.n12 9.3005
R111 VPWR.n14 VPWR.n4 9.3005
R112 VPWR.n16 VPWR.n15 9.3005
R113 VPWR.n17 VPWR.n2 9.3005
R114 VPWR.n19 VPWR.n18 9.3005
R115 VPWR.n20 VPWR.n1 7.17142
R116 VPWR.n8 VPWR.n6 6.98558
R117 VPWR.n17 VPWR.n16 3.76521
R118 VPWR.n12 VPWR.n11 0.753441
R119 VPWR.n6 VPWR.n5 0.561428
R120 VPWR VPWR.n20 0.274942
R121 VPWR.n20 VPWR.n19 0.155855
R122 VPWR.n13 VPWR.n5 0.122949
R123 VPWR.n14 VPWR.n13 0.122949
R124 VPWR.n15 VPWR.n14 0.122949
R125 VPWR.n15 VPWR.n2 0.122949
R126 VPWR.n19 VPWR.n2 0.122949
R127 VPB VPB.t6 457.125
R128 VPB.t3 VPB.t7 416.264
R129 VPB.t1 VPB.t5 331.99
R130 VPB.t8 VPB.t0 280.914
R131 VPB.t6 VPB.t2 275.807
R132 VPB.t5 VPB.t4 229.839
R133 VPB.t0 VPB.t1 229.839
R134 VPB.t7 VPB.t8 229.839
R135 VPB.t2 VPB.t3 229.839
C0 VGND Y 0.017772f
C1 Y B 0.207461f
C2 C D 0.076279f
C3 C VPWR 0.034217f
C4 C Y 0.132463f
C5 D VPWR 0.068926f
C6 VPB A_N 0.060039f
C7 VGND VPB 0.011008f
C8 D Y 0.094406f
C9 VPB B 0.083879f
C10 VGND A_N 0.019272f
C11 VPWR Y 0.821575f
C12 VGND B 0.015662f
C13 C VPB 0.076843f
C14 D VPB 0.069648f
C15 VGND C 0.015695f
C16 C B 0.036255f
C17 VPWR VPB 0.172033f
C18 VGND D 0.032718f
C19 Y VPB 0.019404f
C20 VPWR A_N 0.024551f
C21 VGND VPWR 0.095722f
C22 VPWR B 0.035493f
C23 Y A_N 0.00164f
C24 VGND VNB 0.691321f
C25 Y VNB 0.028402f
C26 VPWR VNB 0.578956f
C27 D VNB 0.236856f
C28 C VNB 0.221719f
C29 B VNB 0.236409f
C30 A_N VNB 0.20845f
C31 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4b_4 VNB VPB VPWR VGND A_N C B Y D
X0 a_225_74.t7 B.t0 a_656_74.t5 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VPWR.t2 D.t0 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.1792 ps=1.44 w=1.12 l=0.15
X2 VGND D a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t2 a_27_158.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3976 pd=1.83 as=0.203 ps=1.505 w=1.12 l=0.15
X4 a_225_74.t0 a_27_158.t4 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VPWR.t3 A_N.t0 a_27_158.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.126 ps=1.14 w=0.84 l=0.15
X6 a_656_74.t4 B.t1 a_225_74.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_27_158.t0 A_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2898 ps=2.37 w=0.84 l=0.15
X8 VGND.t0 A_N.t2 a_27_158.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.19515 pd=2.05 as=0.1962 ps=2.05 w=0.74 l=0.15
X9 a_656_74.t1 C.t0 a_1025_158# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VPWR.t9 B.t2 Y.t11 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.6132 pd=2.215 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_656_74.t3 B.t3 a_225_74.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 Y.t10 B.t4 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.7336 ps=2.43 w=1.12 l=0.15
X13 Y.t8 C.t1 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.6132 ps=2.215 w=1.12 l=0.15
X14 a_656_74.t6 C.t2 a_1025_158# VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1962 ps=2.05 w=0.74 l=0.15
X15 Y.t4 a_27_158.t5 a_225_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_1025_158# D.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.14615 ps=1.135 w=0.74 l=0.15
X17 VGND D a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.14615 pd=1.135 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 Y.t5 a_27_158.t6 a_225_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1962 ps=2.05 w=0.74 l=0.15
X19 a_1025_158# C.t3 a_656_74.t7 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t5 a_27_158.t7 Y.t6 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.7336 pd=2.43 as=0.3976 ps=1.83 w=1.12 l=0.15
X21 Y.t0 D.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.6552 ps=2.29 w=1.12 l=0.15
X22 a_225_74.t3 a_27_158.t8 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_1025_158# D.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VPWR.t6 C.t4 Y.t7 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.6552 pd=2.29 as=0.3808 ps=1.8 w=1.12 l=0.15
X25 a_1025_158# C.t5 a_656_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.10915 ps=1.035 w=0.74 l=0.15
X26 a_225_74.t4 B.t5 a_656_74.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.19515 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 B.n0 B.t2 265.899
R1 B.n1 B.t4 226.809
R2 B.n5 B.t3 209.16
R3 B.n4 B.t0 196.013
R4 B.n0 B.t5 196.013
R5 B.n2 B.t1 196.013
R6 B B.n5 160.047
R7 B B.n3 72.6615
R8 B.n5 B.n4 49.6611
R9 B.n1 B.n0 37.641
R10 B.n3 B.n2 35.4519
R11 B.n2 B.n1 27.0217
R12 B.n4 B.n3 20.6197
R13 a_656_74.n2 a_656_74.n0 229.032
R14 a_656_74.n5 a_656_74.n4 222.089
R15 a_656_74.n2 a_656_74.n1 185
R16 a_656_74.n4 a_656_74.n3 185
R17 a_656_74.n4 a_656_74.n2 72.0787
R18 a_656_74.t0 a_656_74.n5 25.1356
R19 a_656_74.n3 a_656_74.t7 22.7032
R20 a_656_74.n3 a_656_74.t6 22.7032
R21 a_656_74.n0 a_656_74.t5 22.7032
R22 a_656_74.n0 a_656_74.t3 22.7032
R23 a_656_74.n1 a_656_74.t2 22.7032
R24 a_656_74.n1 a_656_74.t4 22.7032
R25 a_656_74.n5 a_656_74.t1 22.7032
R26 a_225_74.n4 a_225_74.t4 276.224
R27 a_225_74.n1 a_225_74.t2 262.813
R28 a_225_74.n1 a_225_74.n0 185
R29 a_225_74.n3 a_225_74.n2 185
R30 a_225_74.n5 a_225_74.n4 185
R31 a_225_74.n3 a_225_74.n1 76.5564
R32 a_225_74.n4 a_225_74.n3 73.4123
R33 a_225_74.n2 a_225_74.t5 22.7032
R34 a_225_74.n2 a_225_74.t0 22.7032
R35 a_225_74.n0 a_225_74.t1 22.7032
R36 a_225_74.n0 a_225_74.t3 22.7032
R37 a_225_74.t6 a_225_74.n5 22.7032
R38 a_225_74.n5 a_225_74.t7 22.7032
R39 VNB.t9 VNB.t13 2286.61
R40 VNB.t0 VNB.t5 2286.61
R41 VNB.t1 VNB.t2 2251.97
R42 VNB.t6 VNB.t1 1986.35
R43 VNB VNB.t0 1143.31
R44 VNB.t7 VNB.t6 1027.82
R45 VNB.t14 VNB.t7 993.177
R46 VNB.t13 VNB.t14 993.177
R47 VNB.t11 VNB.t9 993.177
R48 VNB.t12 VNB.t11 993.177
R49 VNB.t10 VNB.t12 993.177
R50 VNB.t3 VNB.t10 993.177
R51 VNB.t4 VNB.t3 993.177
R52 VNB.t8 VNB.t4 993.177
R53 VNB.t5 VNB.t8 993.177
R54 D.n6 D.n5 318.12
R55 D.n0 D.t0 240.197
R56 D.n8 D.t2 240.197
R57 D D.n1 186.331
R58 D.n6 D.t3 179.947
R59 D.n7 D.n4 179.947
R60 D.n1 D.t1 179.947
R61 D.n3 D.n2 152
R62 D.n10 D.n9 152
R63 D.n7 D.n6 125.028
R64 D.n9 D.n3 49.6611
R65 D.n9 D.n8 10.955
R66 D D.n10 8.93383
R67 D.n1 D.n0 8.76414
R68 D.n3 D.n0 8.03383
R69 D.n2 D 7.6005
R70 D.n2 D 5.2005
R71 D.n10 D 3.86717
R72 D.n8 D.n7 2.19141
R73 Y.n5 Y.n0 321.462
R74 Y.n3 Y.n1 292.502
R75 Y.n2 Y.n1 292.5
R76 Y.n8 Y.n6 281.284
R77 Y.n5 Y.n4 276.695
R78 Y.n12 Y.n10 223.761
R79 Y.n8 Y.n7 204.577
R80 Y.n12 Y.n11 185
R81 Y Y.n12 134.631
R82 Y.n9 Y.n5 109.566
R83 Y.n6 Y.t2 56.8172
R84 Y.n6 Y.t6 56.8171
R85 Y Y.n9 33.9483
R86 Y.n4 Y.n3 31.6146
R87 Y.n4 Y.n2 31.6146
R88 Y.n0 Y.t0 29.9023
R89 Y.n0 Y.t1 26.3844
R90 Y.n2 Y.t7 26.3844
R91 Y.n3 Y.t8 26.3844
R92 Y.n7 Y.t11 26.3844
R93 Y.n7 Y.t10 26.3844
R94 Y.n11 Y.t3 22.7032
R95 Y.n11 Y.t4 22.7032
R96 Y.n10 Y.t9 22.7032
R97 Y.n10 Y.t5 22.7032
R98 Y.n5 Y.n1 10.5404
R99 Y.n9 Y.n8 3.48894
R100 VPWR.n48 VPWR.t0 374.26
R101 VPWR.n40 VPWR.n39 292.5
R102 VPWR.n38 VPWR.n5 292.5
R103 VPWR.n37 VPWR.n36 292.5
R104 VPWR.n29 VPWR.n28 292.5
R105 VPWR.n27 VPWR.n8 292.5
R106 VPWR.n26 VPWR.n25 292.5
R107 VPWR.n18 VPWR.n17 292.5
R108 VPWR.n16 VPWR.n11 292.5
R109 VPWR.n15 VPWR.n14 292.5
R110 VPWR.n12 VPWR.t2 260.288
R111 VPWR.n46 VPWR.n2 233.293
R112 VPWR.n38 VPWR.n37 90.5853
R113 VPWR.n39 VPWR.n38 87.0675
R114 VPWR.n16 VPWR.n15 79.1523
R115 VPWR.n17 VPWR.n16 73.8755
R116 VPWR.n28 VPWR.n27 73.8755
R117 VPWR.n27 VPWR.n26 65.9603
R118 VPWR.n2 VPWR.t3 55.1136
R119 VPWR.n45 VPWR.n3 36.1417
R120 VPWR.n23 VPWR.n9 36.1417
R121 VPWR.n2 VPWR.t4 29.6087
R122 VPWR.n34 VPWR.n6 29.1109
R123 VPWR.n19 VPWR.n9 28.1521
R124 VPWR.n48 VPWR.n47 27.4829
R125 VPWR.n15 VPWR.t1 26.3844
R126 VPWR.n17 VPWR.t6 26.3844
R127 VPWR.n26 VPWR.t7 26.3844
R128 VPWR.n28 VPWR.t9 26.3844
R129 VPWR.n37 VPWR.t8 26.3844
R130 VPWR.n39 VPWR.t5 26.3844
R131 VPWR.n47 VPWR.n46 25.6005
R132 VPWR.n46 VPWR.n45 21.8358
R133 VPWR.n40 VPWR.n3 17.6896
R134 VPWR.n29 VPWR.n6 16.9367
R135 VPWR.n25 VPWR.n23 10.5367
R136 VPWR.n13 VPWR.n10 9.3005
R137 VPWR.n20 VPWR.n19 9.3005
R138 VPWR.n21 VPWR.n9 9.3005
R139 VPWR.n23 VPWR.n22 9.3005
R140 VPWR.n24 VPWR.n7 9.3005
R141 VPWR.n31 VPWR.n30 9.3005
R142 VPWR.n32 VPWR.n6 9.3005
R143 VPWR.n34 VPWR.n33 9.3005
R144 VPWR.n35 VPWR.n4 9.3005
R145 VPWR.n42 VPWR.n41 9.3005
R146 VPWR.n43 VPWR.n3 9.3005
R147 VPWR.n45 VPWR.n44 9.3005
R148 VPWR.n46 VPWR.n1 9.3005
R149 VPWR.n47 VPWR.n0 9.3005
R150 VPWR.n14 VPWR.n12 7.48019
R151 VPWR.n49 VPWR.n48 7.03525
R152 VPWR.n14 VPWR.n13 4.89294
R153 VPWR.n36 VPWR.n35 4.83606
R154 VPWR.n18 VPWR.n11 4.77917
R155 VPWR.n41 VPWR.n5 4.43783
R156 VPWR.n30 VPWR.n8 3.47072
R157 VPWR.n25 VPWR.n24 2.27606
R158 VPWR.n24 VPWR.n8 1.99161
R159 VPWR.n30 VPWR.n29 1.30894
R160 VPWR.n41 VPWR.n40 1.19517
R161 VPWR.n35 VPWR.n5 1.0245
R162 VPWR.n36 VPWR.n34 0.626278
R163 VPWR.n12 VPWR.n10 0.604742
R164 VPWR.n19 VPWR.n18 0.455611
R165 VPWR.n13 VPWR.n11 0.228056
R166 VPWR VPWR.n49 0.154841
R167 VPWR.n49 VPWR.n0 0.152893
R168 VPWR.n20 VPWR.n10 0.122949
R169 VPWR.n21 VPWR.n20 0.122949
R170 VPWR.n22 VPWR.n21 0.122949
R171 VPWR.n22 VPWR.n7 0.122949
R172 VPWR.n31 VPWR.n7 0.122949
R173 VPWR.n32 VPWR.n31 0.122949
R174 VPWR.n33 VPWR.n32 0.122949
R175 VPWR.n33 VPWR.n4 0.122949
R176 VPWR.n42 VPWR.n4 0.122949
R177 VPWR.n43 VPWR.n42 0.122949
R178 VPWR.n44 VPWR.n43 0.122949
R179 VPWR.n44 VPWR.n1 0.122949
R180 VPWR.n1 VPWR.n0 0.122949
R181 VPB.t5 VPB.t8 745.699
R182 VPB.t6 VPB.t1 674.194
R183 VPB.t9 VPB.t7 635.888
R184 VPB VPB.t0 482.661
R185 VPB.t4 VPB.t5 439.248
R186 VPB.t7 VPB.t6 423.925
R187 VPB.t3 VPB.t4 273.253
R188 VPB.t1 VPB.t2 240.054
R189 VPB.t8 VPB.t9 229.839
R190 VPB.t0 VPB.t3 229.839
R191 VGND.n7 VGND.t2 249.391
R192 VGND.n8 VGND.t1 231.558
R193 VGND.n28 VGND.t0 231.453
R194 VGND.n10 VGND.n9 36.1417
R195 VGND.n10 VGND.n5 36.1417
R196 VGND.n14 VGND.n5 36.1417
R197 VGND.n15 VGND.n14 36.1417
R198 VGND.n16 VGND.n15 36.1417
R199 VGND.n16 VGND.n3 36.1417
R200 VGND.n20 VGND.n3 36.1417
R201 VGND.n21 VGND.n20 36.1417
R202 VGND.n22 VGND.n21 36.1417
R203 VGND.n22 VGND.n1 36.1417
R204 VGND.n26 VGND.n1 36.1417
R205 VGND.n27 VGND.n26 36.1417
R206 VGND.n28 VGND.n27 24.4711
R207 VGND.n9 VGND.n8 23.3417
R208 VGND.n27 VGND.n0 9.3005
R209 VGND.n26 VGND.n25 9.3005
R210 VGND.n24 VGND.n1 9.3005
R211 VGND.n23 VGND.n22 9.3005
R212 VGND.n21 VGND.n2 9.3005
R213 VGND.n20 VGND.n19 9.3005
R214 VGND.n18 VGND.n3 9.3005
R215 VGND.n17 VGND.n16 9.3005
R216 VGND.n15 VGND.n4 9.3005
R217 VGND.n14 VGND.n13 9.3005
R218 VGND.n12 VGND.n5 9.3005
R219 VGND.n11 VGND.n10 9.3005
R220 VGND.n9 VGND.n6 9.3005
R221 VGND.n29 VGND.n28 7.19894
R222 VGND.n8 VGND.n7 6.62032
R223 VGND.n7 VGND.n6 0.65114
R224 VGND VGND.n29 0.156997
R225 VGND.n29 VGND.n0 0.150766
R226 VGND.n11 VGND.n6 0.122949
R227 VGND.n12 VGND.n11 0.122949
R228 VGND.n13 VGND.n12 0.122949
R229 VGND.n13 VGND.n4 0.122949
R230 VGND.n17 VGND.n4 0.122949
R231 VGND.n18 VGND.n17 0.122949
R232 VGND.n19 VGND.n18 0.122949
R233 VGND.n19 VGND.n2 0.122949
R234 VGND.n23 VGND.n2 0.122949
R235 VGND.n24 VGND.n23 0.122949
R236 VGND.n25 VGND.n24 0.122949
R237 VGND.n25 VGND.n0 0.122949
R238 a_27_158.n7 a_27_158.n6 314.418
R239 a_27_158.n6 a_27_158.t1 278.709
R240 a_27_158.n0 a_27_158.t6 264.37
R241 a_27_158.n1 a_27_158.t7 228.877
R242 a_27_158.n0 a_27_158.t3 226.809
R243 a_27_158.n5 a_27_158.n4 152
R244 a_27_158.n3 a_27_158.t5 142.994
R245 a_27_158.n1 a_27_158.t4 142.994
R246 a_27_158.n0 a_27_158.t8 142.994
R247 a_27_158.n5 a_27_158.n2 90.0435
R248 a_27_158.n7 a_27_158.t2 35.1791
R249 a_27_158.t0 a_27_158.n7 35.1791
R250 a_27_158.n6 a_27_158.n5 34.3045
R251 a_27_158.n4 a_27_158.n3 33.1076
R252 a_27_158.n2 a_27_158.n1 24.5851
R253 a_27_158.n3 a_27_158.n2 14.1958
R254 a_27_158.n4 a_27_158.n0 8.76414
R255 A_N.n0 A_N.t0 286.822
R256 A_N.n2 A_N.t2 179.947
R257 A_N.n3 A_N.n2 170.714
R258 A_N.n0 A_N.t1 169.772
R259 A_N.n1 A_N 152.934
R260 A_N.n1 A_N.n0 31.1887
R261 A_N.n2 A_N.n1 19.8476
R262 A_N.n3 A_N 8.13383
R263 A_N A_N.n3 4.66717
R264 C.n0 C.t4 226.809
R265 C.n5 C.t1 226.809
R266 C.n3 C.t2 224.495
R267 C.n0 C.t5 198.204
R268 C.n4 C.t3 196.013
R269 C.n1 C.t0 196.013
R270 C.n11 C.n10 152
R271 C.n9 C.n8 152
R272 C.n7 C.n6 152
R273 C.n3 C.n2 152
R274 C.n10 C.n9 49.6611
R275 C.n6 C.n1 47.4702
R276 C.n4 C.n3 34.3247
R277 C.n10 C.n0 10.955
R278 C.n6 C.n5 10.955
R279 C.n8 C.n7 10.1214
R280 C.n11 C 9.07957
R281 C.n2 C 7.29352
R282 C.n2 C 6.99585
R283 C C.n11 5.2098
R284 C.n5 C.n4 4.38232
R285 C.n7 C 3.12608
R286 C.n9 C.n1 2.19141
R287 C.n8 C 1.04236
C0 VPB VGND 0.013876f
C1 B Y 0.303975f
C2 D VPWR 0.083815f
C3 C Y 0.289971f
C4 B VGND 0.022711f
C5 a_1025_158# VPB 7.12e-19
C6 C VGND 0.032129f
C7 a_1025_158# B 0.001383f
C8 VPWR A_N 0.074304f
C9 D Y 0.092614f
C10 a_1025_158# C 0.234644f
C11 VPWR Y 1.14333f
C12 D VGND 0.06808f
C13 VPB B 0.128097f
C14 A_N Y 9.88e-19
C15 VPWR VGND 0.154796f
C16 a_1025_158# D 0.1695f
C17 VPB C 0.132143f
C18 A_N VGND 0.020864f
C19 a_1025_158# VPWR 0.005844f
C20 B C 0.027147f
C21 Y VGND 0.033987f
C22 VPB D 0.121155f
C23 a_1025_158# Y 0.011042f
C24 VPB VPWR 0.276401f
C25 VPB A_N 0.117689f
C26 B VPWR 0.054876f
C27 C D 0.077523f
C28 a_1025_158# VGND 0.331107f
C29 B A_N 8e-20
C30 VPB Y 0.02716f
C31 C VPWR 0.054151f
C32 VGND VNB 1.04119f
C33 Y VNB 0.034382f
C34 A_N VNB 0.265843f
C35 VPWR VNB 0.858049f
C36 D VNB 0.438091f
C37 C VNB 0.37645f
C38 B VNB 0.372331f
C39 VPB VNB 2.1204f
C40 a_1025_158# VNB 0.061403f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4bb_1 VNB VPB VPWR VGND B_N A_N D Y C
X0 a_513_74.t1 a_226_398.t2 a_435_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 VGND.t1 D.t0 a_627_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.266 pd=2.34 as=0.1554 ps=1.16 w=0.74 l=0.15
X2 VPWR.t3 A_N.t0 a_27_398.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X3 Y.t3 D.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4 a_226_398.t1 B_N.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.168 ps=1.24 w=0.84 l=0.15
X5 a_435_74.t1 a_27_398.t2 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.19585 ps=2.05 w=0.74 l=0.15
X6 VGND.t2 A_N.t1 a_27_398.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.122175 pd=1.025 as=0.150975 ps=1.67 w=0.55 l=0.15
X7 VPWR.t5 C.t0 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.196 ps=1.47 w=1.12 l=0.15
X8 a_627_74.t0 C.t1 a_513_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 VPWR.t1 a_27_398.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2464 pd=1.56 as=0.3304 ps=2.83 w=1.12 l=0.15
X10 a_226_398.t0 B_N.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15055 pd=1.69 as=0.122175 ps=1.025 w=0.55 l=0.15
X11 Y.t0 a_226_398.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2464 ps=1.56 w=1.12 l=0.15
R0 a_226_398.t1 a_226_398.n1 490.2
R1 a_226_398.n1 a_226_398.t0 309.221
R2 a_226_398.n0 a_226_398.t3 285.719
R3 a_226_398.n0 a_226_398.t2 178.34
R4 a_226_398.n1 a_226_398.n0 152
R5 a_435_74.t0 a_435_74.t1 38.9194
R6 a_513_74.t0 a_513_74.t1 68.1086
R7 VNB.t1 VNB.t4 2309.71
R8 VNB.t5 VNB.t1 1339.63
R9 VNB.t0 VNB.t3 1316.54
R10 VNB.t2 VNB.t0 1316.54
R11 VNB VNB.t5 1201.05
R12 VNB.t4 VNB.t2 900.788
R13 D.n0 D.t1 250.909
R14 D.n0 D.t0 220.113
R15 D D.n0 158.102
R16 a_627_74.t0 a_627_74.t1 68.1086
R17 VGND.n1 VGND.t1 278.536
R18 VGND.n1 VGND.n0 221.553
R19 VGND.n0 VGND.t2 45.9805
R20 VGND.n0 VGND.t0 34.7215
R21 VGND VGND.n1 0.202699
R22 A_N.t1 A_N.t0 433.8
R23 A_N A_N.t1 310.591
R24 a_27_398.t1 a_27_398.n1 449.353
R25 a_27_398.n0 a_27_398.t3 277.849
R26 a_27_398.n1 a_27_398.n0 254.668
R27 a_27_398.n1 a_27_398.t0 216.948
R28 a_27_398.n0 a_27_398.t2 170.471
R29 VPWR.n5 VPWR.n4 600.696
R30 VPWR.n11 VPWR.n1 322.757
R31 VPWR.n6 VPWR.n3 321.24
R32 VPWR.n1 VPWR.t4 46.9053
R33 VPWR.n1 VPWR.t3 46.9053
R34 VPWR.n4 VPWR.t1 43.0943
R35 VPWR.n9 VPWR.n2 36.1417
R36 VPWR.n10 VPWR.n9 36.1417
R37 VPWR.n3 VPWR.t2 35.1791
R38 VPWR.n3 VPWR.t5 35.1791
R39 VPWR.n4 VPWR.t0 34.2996
R40 VPWR.n11 VPWR.n10 19.2005
R41 VPWR.n6 VPWR.n5 10.5157
R42 VPWR.n7 VPWR.n2 9.3005
R43 VPWR.n9 VPWR.n8 9.3005
R44 VPWR.n10 VPWR.n0 9.3005
R45 VPWR.n12 VPWR.n11 7.43488
R46 VPWR.n5 VPWR.n2 1.12991
R47 VPWR.n7 VPWR.n6 0.628027
R48 VPWR VPWR.n12 0.160103
R49 VPWR.n12 VPWR.n0 0.1477
R50 VPWR.n8 VPWR.n7 0.122949
R51 VPWR.n8 VPWR.n0 0.122949
R52 VPB.t4 VPB.t1 515.861
R53 VPB.t1 VPB.t0 301.344
R54 VPB.t5 VPB.t2 280.914
R55 VPB.t3 VPB.t4 280.914
R56 VPB VPB.t3 257.93
R57 VPB.t0 VPB.t5 255.376
R58 Y.n0 Y.t2 423.582
R59 Y Y.t1 364.983
R60 Y.n0 Y.t3 228.94
R61 Y.n2 Y.n1 196.423
R62 Y.n2 Y.n0 53.6476
R63 Y.n1 Y.t0 35.1791
R64 Y.n1 Y.t4 26.3844
R65 Y Y.n2 7.27323
R66 B_N.n0 B_N.t0 213.954
R67 B_N.n0 B_N.t1 199.227
R68 B_N.n1 B_N.n0 152
R69 B_N.n1 B_N 14.546
R70 B_N B_N.n1 4.07323
R71 C.n0 C.t0 285.719
R72 C.n0 C.t1 178.34
R73 C C.n0 158.788
C0 VPWR B_N 0.051994f
C1 VGND A_N 0.095608f
C2 VPB C 0.031199f
C3 VGND B_N 0.012655f
C4 VPWR Y 0.416057f
C5 VGND Y 0.271608f
C6 A_N B_N 0.053264f
C7 D Y 0.142469f
C8 A_N Y 6.81e-19
C9 VPWR VPB 0.132491f
C10 B_N Y 0.002697f
C11 VPWR C 0.015574f
C12 VGND VPB 0.010198f
C13 VPB D 0.039168f
C14 VGND C 0.008765f
C15 VPB A_N 0.041432f
C16 C D 0.070502f
C17 VPB B_N 0.060499f
C18 VPB Y 0.033891f
C19 VPWR VGND 0.070589f
C20 C Y 0.109813f
C21 VPWR D 0.016849f
C22 VPWR A_N 0.019051f
C23 VGND D 0.009611f
C24 VGND VNB 0.577313f
C25 VPWR VNB 0.430495f
C26 Y VNB 0.115268f
C27 B_N VNB 0.114589f
C28 A_N VNB 0.20742f
C29 D VNB 0.136538f
C30 C VNB 0.109926f
C31 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4bb_2 VNB VPB VPWR VGND A_N Y C D B_N
X0 VPWR.t0 A_N.t0 a_27_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.24225 pd=1.52 as=0.295 ps=2.59 w=1 l=0.15
X1 a_678_74.t3 C.t0 a_886_74# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t6 a_231_74.t2 Y.t7 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.4648 pd=1.95 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t6 a_231_74.t3 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X4 VGND.t1 A_N.t1 a_27_368.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.1824 ps=1.85 w=0.64 l=0.15
X5 a_231_74.t0 B_N.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1344 ps=1.06 w=0.64 l=0.15
X6 a_373_74.t3 a_231_74.t4 a_678_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2516 pd=2.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 Y.t4 D.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.224 ps=1.52 w=1.12 l=0.15
X8 a_886_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 a_678_74.t1 a_231_74.t5 a_373_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1773 ps=1.28 w=0.74 l=0.15
X10 VPWR.t8 D.t1 Y.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3416 pd=2.85 as=0.1904 ps=1.46 w=1.12 l=0.15
X11 a_886_74# C.t1 a_678_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X12 VPWR.t2 a_27_368.t2 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_231_74.t1 B_N.t1 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.395 pd=2.79 as=0.24225 ps=1.52 w=1 l=0.15
X14 Y.t1 a_27_368.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X15 VGND D a_886_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 Y.t9 C.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4648 ps=1.95 w=1.12 l=0.15
X17 VPWR.t9 C.t3 Y.t8 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X18 Y.t3 a_27_368.t4 a_373_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.2442 ps=2.14 w=0.74 l=0.15
X19 a_373_74.t0 a_27_368.t5 Y.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1773 pd=1.28 as=0.11285 ps=1.045 w=0.74 l=0.15
R0 A_N.n0 A_N.t0 243.641
R1 A_N.n0 A_N.t1 218.737
R2 A_N A_N.n0 155.68
R3 a_27_368.n2 a_27_368.n1 319.385
R4 a_27_368.n1 a_27_368.t3 270.991
R5 a_27_368.n0 a_27_368.t2 266.44
R6 a_27_368.t0 a_27_368.n2 224.377
R7 a_27_368.n2 a_27_368.t1 217.454
R8 a_27_368.n0 a_27_368.t4 200.566
R9 a_27_368.n0 a_27_368.t5 166.023
R10 a_27_368.n1 a_27_368.n0 30.7949
R11 VPWR.n2 VPWR.t1 823.319
R12 VPWR.n22 VPWR.n1 607.692
R13 VPWR.n15 VPWR.n4 316.87
R14 VPWR.n9 VPWR.n8 315.928
R15 VPWR.n7 VPWR.t8 257.207
R16 VPWR.n6 VPWR.n5 136.322
R17 VPWR.n5 VPWR.t6 66.5907
R18 VPWR.n5 VPWR.t3 66.5904
R19 VPWR.n1 VPWR.t4 46.2955
R20 VPWR.n1 VPWR.t0 46.2955
R21 VPWR.n21 VPWR.n20 36.1417
R22 VPWR.n4 VPWR.t7 35.1791
R23 VPWR.n4 VPWR.t2 35.1791
R24 VPWR.n8 VPWR.t5 35.1791
R25 VPWR.n8 VPWR.t9 35.1791
R26 VPWR.n16 VPWR.n2 35.0123
R27 VPWR.n10 VPWR.n6 32.7534
R28 VPWR.n15 VPWR.n14 32.0005
R29 VPWR.n14 VPWR.n6 18.4476
R30 VPWR.n10 VPWR.n9 17.6946
R31 VPWR.n22 VPWR.n21 16.5652
R32 VPWR.n16 VPWR.n15 15.4358
R33 VPWR.n20 VPWR.n2 12.424
R34 VPWR.n11 VPWR.n10 9.3005
R35 VPWR.n14 VPWR.n13 9.3005
R36 VPWR.n15 VPWR.n3 9.3005
R37 VPWR.n17 VPWR.n16 9.3005
R38 VPWR.n18 VPWR.n2 9.3005
R39 VPWR.n20 VPWR.n19 9.3005
R40 VPWR.n21 VPWR.n0 9.3005
R41 VPWR.n23 VPWR.n22 7.53404
R42 VPWR.n9 VPWR.n7 6.96039
R43 VPWR.n12 VPWR.n6 4.62059
R44 VPWR.n11 VPWR.n7 0.594857
R45 VPWR.n12 VPWR.n11 0.184273
R46 VPWR.n13 VPWR.n12 0.184273
R47 VPWR VPWR.n23 0.161409
R48 VPWR.n23 VPWR.n0 0.146411
R49 VPWR.n13 VPWR.n3 0.122949
R50 VPWR.n17 VPWR.n3 0.122949
R51 VPWR.n18 VPWR.n17 0.122949
R52 VPWR.n19 VPWR.n18 0.122949
R53 VPWR.n19 VPWR.n0 0.122949
R54 VPB.t4 VPB.t1 592.473
R55 VPB.t6 VPB.t3 500.538
R56 VPB.t0 VPB.t4 316.668
R57 VPB.t9 VPB.t5 280.914
R58 VPB.t2 VPB.t7 280.914
R59 VPB VPB.t0 257.93
R60 VPB.t5 VPB.t8 250.269
R61 VPB.t3 VPB.t9 229.839
R62 VPB.t7 VPB.t6 229.839
R63 VPB.t1 VPB.t2 229.839
R64 C.n2 C.t2 237.762
R65 C.n1 C.t3 226.809
R66 C.n0 C.t1 206.238
R67 C.n2 C.t0 196.013
R68 C C.n0 159.888
R69 C.n4 C.n3 152
R70 C.n3 C.n1 41.6278
R71 C.n3 C.n2 13.146
R72 C.n4 C 12.0563
R73 C.n1 C.n0 8.03383
R74 C C.n4 2.23306
R75 a_678_74.n1 a_678_74.n0 480.005
R76 a_678_74.n1 a_678_74.t3 34.0546
R77 a_678_74.n0 a_678_74.t0 22.7032
R78 a_678_74.n0 a_678_74.t1 22.7032
R79 a_678_74.t2 a_678_74.n1 22.7032
R80 VNB.t0 VNB.t3 2748.56
R81 VNB.t4 VNB.t7 2413.65
R82 VNB.t2 VNB.t5 1362.73
R83 VNB.t1 VNB.t0 1316.54
R84 VNB VNB.t1 1177.95
R85 VNB.t7 VNB.t6 1154.86
R86 VNB.t3 VNB.t2 1050.92
R87 VNB.t5 VNB.t4 993.177
R88 a_231_74.t1 a_231_74.n5 819.967
R89 a_231_74.n3 a_231_74.t3 227.538
R90 a_231_74.n0 a_231_74.t2 226.809
R91 a_231_74.n0 a_231_74.t4 197.475
R92 a_231_74.n2 a_231_74.t5 196.013
R93 a_231_74.n4 a_231_74.n1 169.409
R94 a_231_74.n4 a_231_74.n3 152
R95 a_231_74.n5 a_231_74.n4 142.849
R96 a_231_74.n5 a_231_74.t0 134.773
R97 a_231_74.n2 a_231_74.n1 46.0096
R98 a_231_74.n1 a_231_74.n0 15.3369
R99 a_231_74.n3 a_231_74.n2 3.65202
R100 Y Y.n7 315.325
R101 Y.n5 Y.n4 258.046
R102 Y.n2 Y.n0 253.624
R103 Y.n2 Y.n1 205.487
R104 Y.n5 Y.n3 204.577
R105 Y.n6 Y.n2 49.1229
R106 Y Y.n6 35.6179
R107 Y.n0 Y.t5 33.4201
R108 Y.n7 Y.t3 26.7573
R109 Y.n3 Y.t7 26.3844
R110 Y.n3 Y.t6 26.3844
R111 Y.n4 Y.t2 26.3844
R112 Y.n4 Y.t1 26.3844
R113 Y.n0 Y.t4 26.3844
R114 Y.n1 Y.t8 26.3844
R115 Y.n1 Y.t9 26.3844
R116 Y.n7 Y.t0 22.7032
R117 Y.n6 Y.n5 19.2005
R118 VGND VGND.n0 121.715
R119 VGND.n0 VGND.t0 39.3755
R120 VGND.n0 VGND.t1 39.3755
R121 B_N.n0 B_N.t1 277.151
R122 B_N.n0 B_N.t0 181.554
R123 B_N B_N.n0 157.237
R124 a_373_74.n1 a_373_74.t3 303.24
R125 a_373_74.t1 a_373_74.n1 285.606
R126 a_373_74.n1 a_373_74.n0 185
R127 a_373_74.n0 a_373_74.t2 35.6762
R128 a_373_74.n0 a_373_74.t0 35.6762
R129 D.n1 D.t0 227.538
R130 D.n3 D.t1 226.809
R131 D.n3 D.n2 198.204
R132 D.n1 D.n0 196.013
R133 D D.n4 78.7237
R134 D.n4 D.n1 32.5869
R135 D.n4 D.n3 31.5319
C0 D VGND 0.034537f
C1 a_886_74# D 0.110929f
C2 Y VGND 0.019515f
C3 D VPWR 0.07092f
C4 Y A_N 1.11e-19
C5 a_886_74# Y 0.016728f
C6 VGND A_N 0.035447f
C7 Y VPWR 0.823857f
C8 a_886_74# VGND 0.187529f
C9 VPB D 0.07084f
C10 Y B_N 6.14e-19
C11 D C 0.080849f
C12 VGND VPWR 0.111828f
C13 A_N VPWR 0.015849f
C14 VPB Y 0.024517f
C15 a_886_74# VPWR 0.004167f
C16 VGND B_N 0.019743f
C17 Y C 0.151253f
C18 A_N B_N 0.070573f
C19 VPB VGND 0.011745f
C20 VPB A_N 0.039948f
C21 a_886_74# B_N 1.03e-19
C22 a_886_74# VPB 8.28e-19
C23 VGND C 0.017106f
C24 VPWR B_N 0.01359f
C25 a_886_74# C 0.105944f
C26 VPB VPWR 0.20072f
C27 VPWR C 0.039039f
C28 VPB B_N 0.039264f
C29 VPB C 0.075444f
C30 D Y 0.071792f
C31 VGND VNB 0.785127f
C32 Y VNB 0.035908f
C33 D VNB 0.246438f
C34 C VNB 0.219213f
C35 B_N VNB 0.128822f
C36 VPWR VNB 0.653778f
C37 A_N VNB 0.151217f
C38 VPB VNB 1.58472f
C39 a_886_74# VNB 0.056742f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4bb_4 VNB VPB VPWR VGND C D A_N B_N Y
X0 VPWR.t12 D.t0 Y.t16 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_374_74.t6 a_27_114.t3 Y.t5 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t19 C.t0 Y.t19 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VGND.t4 D.t1 a_1229_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VPWR.t13 B_N.t0 a_232_114.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2765 pd=1.69 as=0.126 ps=1.14 w=0.84 l=0.15
X5 Y.t15 D.t2 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t0 C.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VPWR.t10 D.t3 Y.t14 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_232_114.t1 B_N.t1 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X9 Y.t6 a_27_114.t4 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2765 ps=1.69 w=1.12 l=0.15
X10 VPWR.t1 a_232_114.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t15 A_N.t0 a_27_114.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X12 Y.t13 D.t4 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X13 Y.t7 a_27_114.t5 a_374_74.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.14245 pd=1.125 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 Y.t2 a_232_114.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X15 a_374_74.t0 a_232_114.t5 a_828_74.t7 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1657 ps=1.2 w=0.74 l=0.15
X16 a_828_74.t6 a_232_114.t6 a_374_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_1229_74.t6 D.t5 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_232_114.t0 B_N.t2 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2368 pd=2.12 as=0.21935 ps=1.57 w=0.74 l=0.15
X19 Y.t8 a_27_114.t6 a_374_74.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1073 ps=1.03 w=0.74 l=0.15
X20 a_1229_74.t2 C.t2 a_828_74.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VPWR.t3 a_232_114.t7 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X22 Y.t4 a_232_114.t8 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 VPWR.t16 C.t3 Y.t17 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_1229_74.t0 C.t4 a_828_74.t2 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 VPWR.t6 a_27_114.t7 Y.t9 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 Y.t18 C.t5 VPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X27 Y.t10 a_27_114.t8 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 a_27_114.t2 A_N.t1 VPWR.t18 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2478 ps=2.27 w=0.84 l=0.15
X29 VGND.t0 A_N.t2 a_27_114.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.21935 pd=1.57 as=0.2109 ps=2.05 w=0.74 l=0.15
X30 a_828_74.t1 C.t6 a_1229_74.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 a_374_74.t3 a_27_114.t9 Y.t11 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.14245 ps=1.125 w=0.74 l=0.15
X32 a_828_74.t5 a_232_114.t9 a_374_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1657 pd=1.2 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 a_1229_74.t5 D.t6 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X34 a_828_74.t0 C.t7 a_1229_74.t3 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X35 VPWR.t8 a_27_114.t10 Y.t12 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X36 VGND.t1 D.t7 a_1229_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X37 a_374_74.t7 a_232_114.t10 a_828_74.t4 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 D.n11 D.t4 242.704
R1 D.n3 D.t0 240.197
R2 D.n1 D.t2 240.197
R3 D.n9 D.t3 240.197
R4 D.n11 D.t1 180.649
R5 D.n7 D.t7 179.947
R6 D.n10 D.t5 179.947
R7 D.n2 D.t6 179.947
R8 D.n2 D 178.559
R9 D.n5 D.n4 152
R10 D.n7 D.n6 152
R11 D.n8 D.n0 152
R12 D.n13 D.n12 152
R13 D.n8 D.n7 49.6611
R14 D.n4 D.n1 43.8187
R15 D.n12 D.n10 36.5157
R16 D.n12 D.n11 25.5905
R17 D.n4 D.n3 21.9096
R18 D.n9 D.n8 10.2247
R19 D.n13 D.n0 9.06717
R20 D.n5 D 8.8005
R21 D.n6 D 7.73383
R22 D.n7 D.n1 5.84292
R23 D.n6 D 5.06717
R24 D D.n5 4.0005
R25 D.n10 D.n9 2.92171
R26 D D.n13 2.4005
R27 D.n3 D.n2 1.46111
R28 D D.n0 1.33383
R29 Y Y.n0 588.928
R30 Y.n19 Y.n0 585
R31 Y.n18 Y.n0 585
R32 Y.n4 Y.n2 248.405
R33 Y.n11 Y.n10 247.724
R34 Y.n12 Y.n11 216.471
R35 Y.n13 Y.n1 215.304
R36 Y.n4 Y.n3 205.487
R37 Y.n17 Y.n16 205.206
R38 Y.n6 Y.n5 203.127
R39 Y.n8 Y.n7 202.457
R40 Y.n15 Y.n14 200.487
R41 Y.n11 Y.n9 185.754
R42 Y.n15 Y.n13 57.7113
R43 Y.n12 Y.n8 53.3092
R44 Y.n17 Y.n15 52.794
R45 Y.n8 Y.n6 51.1192
R46 Y.n18 Y.n17 50.4476
R47 Y.n6 Y.n4 46.6829
R48 Y.n0 Y.t12 35.1791
R49 Y.n10 Y.t11 33.2437
R50 Y.n10 Y.t7 29.1897
R51 Y.n1 Y.t1 26.3844
R52 Y.n1 Y.t2 26.3844
R53 Y.n7 Y.t19 26.3844
R54 Y.n7 Y.t0 26.3844
R55 Y.n2 Y.t16 26.3844
R56 Y.n2 Y.t15 26.3844
R57 Y.n3 Y.t14 26.3844
R58 Y.n3 Y.t13 26.3844
R59 Y.n5 Y.t17 26.3844
R60 Y.n5 Y.t18 26.3844
R61 Y.n14 Y.t3 26.3844
R62 Y.n14 Y.t4 26.3844
R63 Y.n16 Y.t9 26.3844
R64 Y.n16 Y.t10 26.3844
R65 Y.n0 Y.t6 26.3844
R66 Y.n9 Y.t5 22.7032
R67 Y.n9 Y.t8 22.7032
R68 Y Y.n19 5.96414
R69 Y Y.n18 5.09141
R70 Y.n19 Y 4.8005
R71 Y.n13 Y.n12 2.25932
R72 VPWR.n48 VPWR.t18 351.104
R73 VPWR.n20 VPWR.n18 331.5
R74 VPWR.n12 VPWR.n11 325.01
R75 VPWR.n16 VPWR.n15 323.406
R76 VPWR.n33 VPWR.n10 316.87
R77 VPWR.n27 VPWR.n14 315.928
R78 VPWR.n46 VPWR.n2 314.962
R79 VPWR.n4 VPWR.n3 314.962
R80 VPWR.n39 VPWR.n6 314.962
R81 VPWR.n8 VPWR.n7 314.962
R82 VPWR.n19 VPWR.t12 262.974
R83 VPWR.n3 VPWR.t5 73.2134
R84 VPWR.n3 VPWR.t13 56.2862
R85 VPWR.n20 VPWR.n19 40.1055
R86 VPWR.n41 VPWR.n40 36.1417
R87 VPWR.n22 VPWR.n21 36.1417
R88 VPWR.n2 VPWR.t14 35.1791
R89 VPWR.n2 VPWR.t15 35.1791
R90 VPWR.n10 VPWR.t3 35.1791
R91 VPWR.n14 VPWR.t17 35.1791
R92 VPWR.n14 VPWR.t19 35.1791
R93 VPWR.n15 VPWR.t9 35.1791
R94 VPWR.n38 VPWR.n8 32.7534
R95 VPWR.n34 VPWR.n33 32.0005
R96 VPWR.n26 VPWR.n16 32.0005
R97 VPWR.n32 VPWR.n12 27.4829
R98 VPWR.n28 VPWR.n27 26.7299
R99 VPWR.n6 VPWR.t7 26.3844
R100 VPWR.n6 VPWR.t8 26.3844
R101 VPWR.n7 VPWR.t4 26.3844
R102 VPWR.n7 VPWR.t6 26.3844
R103 VPWR.n10 VPWR.t2 26.3844
R104 VPWR.n11 VPWR.t0 26.3844
R105 VPWR.n11 VPWR.t1 26.3844
R106 VPWR.n15 VPWR.t16 26.3844
R107 VPWR.n18 VPWR.t11 26.3844
R108 VPWR.n18 VPWR.t10 26.3844
R109 VPWR.n28 VPWR.n12 25.977
R110 VPWR.n46 VPWR.n45 25.224
R111 VPWR.n45 VPWR.n4 24.4711
R112 VPWR.n41 VPWR.n4 22.9652
R113 VPWR.n47 VPWR.n46 22.2123
R114 VPWR.n22 VPWR.n16 21.4593
R115 VPWR.n48 VPWR.n47 20.7064
R116 VPWR.n27 VPWR.n26 20.7064
R117 VPWR.n33 VPWR.n32 15.4358
R118 VPWR.n34 VPWR.n8 14.6829
R119 VPWR.n39 VPWR.n38 10.1652
R120 VPWR.n21 VPWR.n17 9.3005
R121 VPWR.n23 VPWR.n22 9.3005
R122 VPWR.n24 VPWR.n16 9.3005
R123 VPWR.n26 VPWR.n25 9.3005
R124 VPWR.n27 VPWR.n13 9.3005
R125 VPWR.n29 VPWR.n28 9.3005
R126 VPWR.n30 VPWR.n12 9.3005
R127 VPWR.n32 VPWR.n31 9.3005
R128 VPWR.n33 VPWR.n9 9.3005
R129 VPWR.n35 VPWR.n34 9.3005
R130 VPWR.n36 VPWR.n8 9.3005
R131 VPWR.n38 VPWR.n37 9.3005
R132 VPWR.n40 VPWR.n5 9.3005
R133 VPWR.n42 VPWR.n41 9.3005
R134 VPWR.n43 VPWR.n4 9.3005
R135 VPWR.n45 VPWR.n44 9.3005
R136 VPWR.n46 VPWR.n1 9.3005
R137 VPWR.n47 VPWR.n0 9.3005
R138 VPWR.n49 VPWR.n48 9.3005
R139 VPWR.n19 VPWR.n17 2.0514
R140 VPWR.n21 VPWR.n20 1.50638
R141 VPWR.n40 VPWR.n39 1.12991
R142 VPWR.n23 VPWR.n17 0.122949
R143 VPWR.n24 VPWR.n23 0.122949
R144 VPWR.n25 VPWR.n24 0.122949
R145 VPWR.n25 VPWR.n13 0.122949
R146 VPWR.n29 VPWR.n13 0.122949
R147 VPWR.n30 VPWR.n29 0.122949
R148 VPWR.n31 VPWR.n30 0.122949
R149 VPWR.n31 VPWR.n9 0.122949
R150 VPWR.n35 VPWR.n9 0.122949
R151 VPWR.n36 VPWR.n35 0.122949
R152 VPWR.n37 VPWR.n36 0.122949
R153 VPWR.n37 VPWR.n5 0.122949
R154 VPWR.n42 VPWR.n5 0.122949
R155 VPWR.n43 VPWR.n42 0.122949
R156 VPWR.n44 VPWR.n43 0.122949
R157 VPWR.n44 VPWR.n1 0.122949
R158 VPWR.n1 VPWR.n0 0.122949
R159 VPWR.n49 VPWR.n0 0.122949
R160 VPWR VPWR.n49 0.0617245
R161 VPB.t13 VPB.t5 367.743
R162 VPB.t19 VPB.t17 280.914
R163 VPB VPB.t18 257.93
R164 VPB.t16 VPB.t9 255.376
R165 VPB.t3 VPB.t2 255.376
R166 VPB.t5 VPB.t8 255.376
R167 VPB.t11 VPB.t12 229.839
R168 VPB.t10 VPB.t11 229.839
R169 VPB.t9 VPB.t10 229.839
R170 VPB.t17 VPB.t16 229.839
R171 VPB.t0 VPB.t19 229.839
R172 VPB.t1 VPB.t0 229.839
R173 VPB.t2 VPB.t1 229.839
R174 VPB.t4 VPB.t3 229.839
R175 VPB.t6 VPB.t4 229.839
R176 VPB.t7 VPB.t6 229.839
R177 VPB.t8 VPB.t7 229.839
R178 VPB.t14 VPB.t13 229.839
R179 VPB.t15 VPB.t14 229.839
R180 VPB.t18 VPB.t15 229.839
R181 a_27_114.n12 a_27_114.n11 417.442
R182 a_27_114.n1 a_27_114.t7 300.113
R183 a_27_114.n2 a_27_114.t8 214.758
R184 a_27_114.n4 a_27_114.t10 214.758
R185 a_27_114.n8 a_27_114.t4 214.758
R186 a_27_114.n1 a_27_114.t3 187.981
R187 a_27_114.n11 a_27_114.n10 170.546
R188 a_27_114.n5 a_27_114.n0 164.8
R189 a_27_114.n9 a_27_114.t5 162.831
R190 a_27_114.n6 a_27_114.t9 154.24
R191 a_27_114.n3 a_27_114.t6 154.24
R192 a_27_114.n10 a_27_114.n9 152
R193 a_27_114.n7 a_27_114.n0 152
R194 a_27_114.n11 a_27_114.t0 131.315
R195 a_27_114.n3 a_27_114.n2 36.6814
R196 a_27_114.t1 a_27_114.n12 35.1791
R197 a_27_114.n12 a_27_114.t2 35.1791
R198 a_27_114.n9 a_27_114.n8 24.3391
R199 a_27_114.n6 a_27_114.n5 22.4302
R200 a_27_114.n2 a_27_114.n1 13.2555
R201 a_27_114.n10 a_27_114.n0 12.8005
R202 a_27_114.n4 a_27_114.n3 12.4084
R203 a_27_114.n7 a_27_114.n6 10.0223
R204 a_27_114.n8 a_27_114.n7 8.11337
R205 a_27_114.n5 a_27_114.n4 7.15892
R206 a_374_74.n1 a_374_74.t0 278.579
R207 a_374_74.n3 a_374_74.t5 193.653
R208 a_374_74.n3 a_374_74.n2 185
R209 a_374_74.n1 a_374_74.n0 185
R210 a_374_74.n5 a_374_74.n4 185
R211 a_374_74.n4 a_374_74.n1 68.5934
R212 a_374_74.n4 a_374_74.n3 60.1329
R213 a_374_74.n2 a_374_74.t4 23.514
R214 a_374_74.n2 a_374_74.t3 23.514
R215 a_374_74.n0 a_374_74.t2 22.7032
R216 a_374_74.n0 a_374_74.t7 22.7032
R217 a_374_74.n5 a_374_74.t1 22.7032
R218 a_374_74.t6 a_374_74.n5 22.7032
R219 VNB.t8 VNB.t11 2644.62
R220 VNB.t0 VNB.t16 2286.61
R221 VNB.t2 VNB.t0 1362.73
R222 VNB.t3 VNB.t8 1362.73
R223 VNB.t11 VNB.t9 1235.7
R224 VNB.t4 VNB.t5 1154.86
R225 VNB VNB.t3 1143.31
R226 VNB.t9 VNB.t10 1016.27
R227 VNB.t6 VNB.t4 993.177
R228 VNB.t7 VNB.t6 993.177
R229 VNB.t13 VNB.t7 993.177
R230 VNB.t15 VNB.t13 993.177
R231 VNB.t14 VNB.t15 993.177
R232 VNB.t16 VNB.t14 993.177
R233 VNB.t17 VNB.t2 993.177
R234 VNB.t1 VNB.t17 993.177
R235 VNB.t12 VNB.t1 993.177
R236 VNB.t10 VNB.t12 993.177
R237 C.n1 C.t1 256.75
R238 C.n2 C.t3 234.841
R239 C.n5 C.t5 234.841
R240 C.n9 C.t0 234.841
R241 C.n2 C.t2 198.751
R242 C.n8 C.t7 186.374
R243 C.n7 C.t4 186.374
R244 C.n4 C.t6 186.374
R245 C.n3 C.n0 165.189
R246 C.n11 C.n1 165.189
R247 C.n6 C.n0 152
R248 C.n11 C.n10 152
R249 C.n3 C.n2 40.8975
R250 C.n9 C.n8 32.1338
R251 C.n6 C.n5 24.8308
R252 C.n7 C.n6 24.8308
R253 C.n10 C.n7 24.8308
R254 C.n5 C.n4 13.146
R255 C.n4 C.n3 11.6853
R256 C.n8 C.n1 11.6853
R257 C C.n12 8.36973
R258 C.n10 C.n9 5.84292
R259 C.n12 C.n0 5.62474
R260 C C.n11 4.26717
R261 C.n12 C 3.29747
R262 a_1229_74.n4 a_1229_74.t3 276.553
R263 a_1229_74.n1 a_1229_74.t5 204.804
R264 a_1229_74.n5 a_1229_74.n4 194.036
R265 a_1229_74.n3 a_1229_74.n2 106.285
R266 a_1229_74.n1 a_1229_74.n0 100.181
R267 a_1229_74.n4 a_1229_74.n3 59.8593
R268 a_1229_74.n3 a_1229_74.n1 58.3534
R269 a_1229_74.n2 a_1229_74.t7 22.7032
R270 a_1229_74.n2 a_1229_74.t2 22.7032
R271 a_1229_74.n0 a_1229_74.t4 22.7032
R272 a_1229_74.n0 a_1229_74.t6 22.7032
R273 a_1229_74.n5 a_1229_74.t1 22.7032
R274 a_1229_74.t0 a_1229_74.n5 22.7032
R275 VGND.n1 VGND.n0 286.38
R276 VGND.n12 VGND.n11 212.583
R277 VGND.n10 VGND.n9 207.109
R278 VGND.n15 VGND.n14 36.1417
R279 VGND.n16 VGND.n15 36.1417
R280 VGND.n16 VGND.n7 36.1417
R281 VGND.n20 VGND.n7 36.1417
R282 VGND.n21 VGND.n20 36.1417
R283 VGND.n22 VGND.n21 36.1417
R284 VGND.n22 VGND.n5 36.1417
R285 VGND.n26 VGND.n5 36.1417
R286 VGND.n27 VGND.n26 36.1417
R287 VGND.n28 VGND.n27 36.1417
R288 VGND.n28 VGND.n3 36.1417
R289 VGND.n32 VGND.n3 36.1417
R290 VGND.n33 VGND.n32 36.1417
R291 VGND.n34 VGND.n33 36.1417
R292 VGND.n0 VGND.t5 35.6762
R293 VGND.n0 VGND.t0 35.6762
R294 VGND.n11 VGND.t2 34.0546
R295 VGND.n14 VGND.n10 26.7299
R296 VGND.n11 VGND.t1 22.7032
R297 VGND.n9 VGND.t3 22.7032
R298 VGND.n9 VGND.t4 22.7032
R299 VGND.n34 VGND.n1 22.1206
R300 VGND.n35 VGND.n34 9.3005
R301 VGND.n33 VGND.n2 9.3005
R302 VGND.n32 VGND.n31 9.3005
R303 VGND.n30 VGND.n3 9.3005
R304 VGND.n29 VGND.n28 9.3005
R305 VGND.n27 VGND.n4 9.3005
R306 VGND.n26 VGND.n25 9.3005
R307 VGND.n24 VGND.n5 9.3005
R308 VGND.n23 VGND.n22 9.3005
R309 VGND.n21 VGND.n6 9.3005
R310 VGND.n20 VGND.n19 9.3005
R311 VGND.n18 VGND.n7 9.3005
R312 VGND.n17 VGND.n16 9.3005
R313 VGND.n15 VGND.n8 9.3005
R314 VGND.n14 VGND.n13 9.3005
R315 VGND.n36 VGND.n1 9.10055
R316 VGND.n12 VGND.n10 6.44389
R317 VGND.n13 VGND.n12 0.645025
R318 VGND VGND.n36 0.161517
R319 VGND.n36 VGND.n35 0.146304
R320 VGND.n13 VGND.n8 0.122949
R321 VGND.n17 VGND.n8 0.122949
R322 VGND.n18 VGND.n17 0.122949
R323 VGND.n19 VGND.n18 0.122949
R324 VGND.n19 VGND.n6 0.122949
R325 VGND.n23 VGND.n6 0.122949
R326 VGND.n24 VGND.n23 0.122949
R327 VGND.n25 VGND.n24 0.122949
R328 VGND.n25 VGND.n4 0.122949
R329 VGND.n29 VGND.n4 0.122949
R330 VGND.n30 VGND.n29 0.122949
R331 VGND.n31 VGND.n30 0.122949
R332 VGND.n31 VGND.n2 0.122949
R333 VGND.n35 VGND.n2 0.122949
R334 B_N.n0 B_N.t2 264.89
R335 B_N.n1 B_N.t0 213.589
R336 B_N.n0 B_N.t1 180.482
R337 B_N B_N.n1 157.237
R338 B_N.n1 B_N.n0 23.5766
R339 a_232_114.n10 a_232_114.t0 353.712
R340 a_232_114.n11 a_232_114.n10 304.598
R341 a_232_114.n2 a_232_114.t3 300.788
R342 a_232_114.n8 a_232_114.t6 238.518
R343 a_232_114.n3 a_232_114.t4 226.809
R344 a_232_114.n6 a_232_114.t7 226.809
R345 a_232_114.n8 a_232_114.t8 226.809
R346 a_232_114.n10 a_232_114.n9 212.225
R347 a_232_114.n4 a_232_114.n1 169.409
R348 a_232_114.n9 a_232_114.n0 152
R349 a_232_114.n7 a_232_114.n1 152
R350 a_232_114.n0 a_232_114.t10 142.994
R351 a_232_114.n5 a_232_114.t9 142.994
R352 a_232_114.n2 a_232_114.t5 142.994
R353 a_232_114.t2 a_232_114.n11 35.1791
R354 a_232_114.n11 a_232_114.t1 35.1791
R355 a_232_114.n0 a_232_114.n7 33.1076
R356 a_232_114.n5 a_232_114.n4 24.8308
R357 a_232_114.n4 a_232_114.n3 18.9884
R358 a_232_114.n9 a_232_114.n1 17.4085
R359 a_232_114.n3 a_232_114.n2 13.6328
R360 a_232_114.n0 a_232_114.n8 7.30353
R361 a_232_114.n6 a_232_114.n5 4.86919
R362 a_232_114.n7 a_232_114.n6 3.40858
R363 A_N.n0 A_N.t0 218.507
R364 A_N.n1 A_N.t2 186.603
R365 A_N.n0 A_N.t1 169.389
R366 A_N A_N.n1 153.135
R367 A_N.n1 A_N.n0 48.8891
R368 a_828_74.n5 a_828_74.n4 238.02
R369 a_828_74.n2 a_828_74.n0 222.023
R370 a_828_74.n2 a_828_74.n1 185
R371 a_828_74.n4 a_828_74.n3 185
R372 a_828_74.n4 a_828_74.n2 98.3985
R373 a_828_74.n1 a_828_74.t7 35.6762
R374 a_828_74.n1 a_828_74.t5 35.6762
R375 a_828_74.n3 a_828_74.t2 22.7032
R376 a_828_74.n3 a_828_74.t0 22.7032
R377 a_828_74.n0 a_828_74.t4 22.7032
R378 a_828_74.n0 a_828_74.t6 22.7032
R379 a_828_74.t3 a_828_74.n5 22.7032
R380 a_828_74.n5 a_828_74.t1 22.7032
C0 C D 0.070053f
C1 Y VGND 0.036562f
C2 Y VPB 0.034303f
C3 VGND VPB 0.011033f
C4 VPWR Y 1.48907f
C5 VGND A_N 0.012558f
C6 Y B_N 0.001494f
C7 VPWR VGND 0.165681f
C8 VPB A_N 0.094919f
C9 VPWR VPB 0.275417f
C10 Y C 0.220349f
C11 VGND B_N 0.009511f
C12 VPB B_N 0.114175f
C13 VPWR A_N 0.038646f
C14 VGND C 0.028448f
C15 Y D 0.180892f
C16 A_N B_N 0.05439f
C17 VPB C 0.143718f
C18 VPWR B_N 0.037508f
C19 VGND D 0.071406f
C20 VPB D 0.151651f
C21 VPWR C 0.071823f
C22 VPWR D 0.096924f
C23 VGND VNB 1.13546f
C24 Y VNB 0.041175f
C25 VPWR VNB 0.956425f
C26 D VNB 0.47377f
C27 C VNB 0.417098f
C28 B_N VNB 0.163826f
C29 A_N VNB 0.15647f
C30 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2_1 VNB VPB VPWR VGND B Y A
X0 a_116_368.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t1 A.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 Y.t2 B.t0 a_116_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X3 VGND.t0 B.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t0 257.118
R1 A.n0 A.t1 196.869
R2 A A.n0 155.601
R3 VPWR VPWR.t0 255.82
R4 a_116_368.t0 a_116_368.t1 47.4916
R5 VPB VPB.t0 257.93
R6 VPB.t0 VPB.t1 214.517
R7 VGND.n0 VGND.t1 178.476
R8 VGND.n0 VGND.t0 170.718
R9 VGND VGND.n0 0.584638
R10 Y Y.n0 587.389
R11 Y.n3 Y.n0 585
R12 Y.n2 Y.n0 585
R13 Y.n2 Y.n1 171.266
R14 Y.n0 Y.t2 26.3844
R15 Y.n1 Y.t0 22.7032
R16 Y.n1 Y.t1 22.7032
R17 Y Y.n3 4.29901
R18 Y Y.n2 3.91692
R19 Y.n3 Y 2.77065
R20 VNB VNB.t1 1189.5
R21 VNB.t1 VNB.t0 993.177
R22 B.n0 B.t0 256.765
R23 B.n0 B.t1 196.516
R24 B B.n0 156.462
C0 B Y 0.107242f
C1 VPWR Y 0.142492f
C2 VGND B 0.052706f
C3 VGND VPWR 0.026685f
C4 VGND Y 0.16016f
C5 VPB A 0.041449f
C6 VPB B 0.041972f
C7 VPB VPWR 0.052201f
C8 A B 0.061434f
C9 A VPWR 0.055467f
C10 VPB Y 0.014849f
C11 A Y 0.064507f
C12 VPB VGND 0.004969f
C13 B VPWR 0.007487f
C14 A VGND 0.044652f
C15 VGND VNB 0.299108f
C16 Y VNB 0.065308f
C17 VPWR VNB 0.222166f
C18 B VNB 0.166986f
C19 A VNB 0.166689f
C20 VPB VNB 0.406224f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2b_2 VNB VPB VPWR VGND A B_N Y
X0 a_228_368.t2 A.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t1 A.t1 a_228_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t3 A.t2 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=2.09 as=0.1221 ps=1.07 w=0.74 l=0.15
X3 a_228_368.t0 a_27_392.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t5 a_27_392.t3 a_228_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 Y.t2 A.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.111 ps=1.04 w=0.74 l=0.15
X6 Y.t4 a_27_392.t4 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.16335 ps=1.195 w=0.74 l=0.15
X7 VGND.t1 B_N.t0 a_27_392.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.16335 pd=1.195 as=0.1824 ps=1.85 w=0.64 l=0.15
X8 VGND.t0 a_27_392.t5 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1221 ps=1.07 w=0.74 l=0.15
X9 VPWR.t0 B_N.t1 a_27_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.29 ps=2.58 w=1 l=0.15
R0 A.n0 A.t0 228.47
R1 A.n1 A.t1 226.809
R2 A.n1 A.t3 202.587
R3 A.n0 A.t2 196.013
R4 A.n3 A.n2 152
R5 A.n2 A.n0 56.9641
R6 A.n3 A 11.3121
R7 A.n2 A.n1 6.57323
R8 A A.n3 2.97724
R9 VPWR.n1 VPWR.n0 329.921
R10 VPWR.n1 VPWR.t0 257.546
R11 VPWR.n0 VPWR.t2 26.3844
R12 VPWR.n0 VPWR.t1 26.3844
R13 VPWR VPWR.n1 0.199785
R14 a_228_368.n1 a_228_368.t3 301.219
R15 a_228_368.t2 a_228_368.n1 295.856
R16 a_228_368.n1 a_228_368.n0 188.462
R17 a_228_368.n0 a_228_368.t1 26.3844
R18 a_228_368.n0 a_228_368.t0 26.3844
R19 VPB.t1 VPB.t4 515.861
R20 VPB VPB.t1 255.376
R21 VPB.t2 VPB.t3 229.839
R22 VPB.t0 VPB.t2 229.839
R23 VPB.t4 VPB.t0 229.839
R24 Y.n2 Y.n0 361.702
R25 Y.n4 Y.n3 103.299
R26 Y.n2 Y.n1 99.1624
R27 Y.n4 Y.n2 44.5096
R28 Y.n3 Y.t3 30.8113
R29 Y.n1 Y.t1 30.8113
R30 Y Y.n4 27.257
R31 Y.n0 Y.t0 26.3844
R32 Y.n0 Y.t5 26.3844
R33 Y.n3 Y.t2 22.7032
R34 Y.n1 Y.t4 22.7032
R35 VGND.n1 VGND.t3 243.756
R36 VGND.n3 VGND.n2 209.243
R37 VGND.n6 VGND.n5 116.436
R38 VGND.n5 VGND.t1 45.938
R39 VGND.n5 VGND.t4 30.2643
R40 VGND.n6 VGND.n4 27.4829
R41 VGND.n2 VGND.t0 25.9464
R42 VGND.n4 VGND.n3 22.9652
R43 VGND.n2 VGND.t2 22.7032
R44 VGND.n4 VGND.n0 9.3005
R45 VGND.n7 VGND.n6 6.93371
R46 VGND.n3 VGND.n1 6.6595
R47 VGND.n1 VGND.n0 0.655456
R48 VGND VGND.n7 0.271269
R49 VGND.n7 VGND.n0 0.159472
R50 VNB VNB.t1 1917.06
R51 VNB.t1 VNB.t4 1397.38
R52 VNB.t2 VNB.t3 1108.66
R53 VNB.t4 VNB.t0 1108.66
R54 VNB.t0 VNB.t2 1039.37
R55 a_27_392.t0 a_27_392.n3 277.205
R56 a_27_392.n0 a_27_392.t2 251.114
R57 a_27_392.n1 a_27_392.t3 235.512
R58 a_27_392.n3 a_27_392.n2 202.649
R59 a_27_392.n2 a_27_392.t4 154.24
R60 a_27_392.n0 a_27_392.t5 154.24
R61 a_27_392.n3 a_27_392.t1 135.77
R62 a_27_392.n1 a_27_392.n0 53.762
R63 a_27_392.n2 a_27_392.n1 5.56204
R64 B_N.n0 B_N.t0 238.226
R65 B_N.n0 B_N.t1 236.011
R66 B_N B_N.n0 154.327
C0 VPB VPWR 0.101949f
C1 B_N VPWR 0.054145f
C2 VPWR Y 0.010294f
C3 A VPWR 0.036289f
C4 VPB B_N 0.064313f
C5 VPWR VGND 0.055171f
C6 VPB Y 0.004819f
C7 VPB A 0.067058f
C8 B_N Y 0.008082f
C9 VPB VGND 0.007844f
C10 A Y 0.134979f
C11 B_N VGND 0.014654f
C12 Y VGND 0.313761f
C13 A VGND 0.035199f
C14 VGND VNB 0.457483f
C15 Y VNB 0.047099f
C16 VPWR VNB 0.344854f
C17 A VNB 0.237768f
C18 B_N VNB 0.154154f
C19 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2b_1 VNB VPB VPWR VGND B_N Y A
X0 Y.t0 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.13135 pd=1.095 as=0.153575 ps=1.2 w=0.74 l=0.15
X1 Y.t1 a_27_112.t2 a_278_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.42 pd=2.99 as=0.1512 ps=1.39 w=1.12 l=0.15
X2 a_278_368.t1 A.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.2345 ps=1.58 w=1.12 l=0.15
X3 VGND.t0 B_N.t0 a_27_112.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.153575 pd=1.2 as=0.2805 ps=2.12 w=0.55 l=0.15
X4 VGND.t2 a_27_112.t3 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.13135 ps=1.095 w=0.74 l=0.15
X5 VPWR.t1 B_N.t1 a_27_112.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2345 pd=1.58 as=0.2478 ps=2.27 w=0.84 l=0.15
R0 A.n0 A.t1 283.113
R1 A.n0 A.t0 175.736
R2 A A.n0 158.788
R3 VGND.n1 VGND.t2 244.565
R4 VGND.n1 VGND.n0 126.425
R5 VGND.n0 VGND.t0 69.1152
R6 VGND.n0 VGND.t1 21.9332
R7 VGND VGND.n1 0.633775
R8 Y.n2 Y 588.636
R9 Y.n2 Y.n0 585
R10 Y.n3 Y.n2 585
R11 Y Y.n1 190.779
R12 Y.n1 Y.t0 34.8654
R13 Y.n2 Y.t1 27.2639
R14 Y.n1 Y.t2 22.7032
R15 Y Y.n3 9.74595
R16 Y Y.n0 8.43686
R17 Y Y.n0 2.32777
R18 Y.n3 Y 1.01868
R19 VNB VNB.t0 1662.99
R20 VNB.t0 VNB.t1 1408.92
R21 VNB.t1 VNB.t2 1166.4
R22 a_27_112.t1 a_27_112.n1 409.457
R23 a_27_112.n1 a_27_112.t0 276.375
R24 a_27_112.n0 a_27_112.t2 258.942
R25 a_27_112.n1 a_27_112.n0 234.287
R26 a_27_112.n0 a_27_112.t3 210.474
R27 a_278_368.t0 a_278_368.t1 47.4916
R28 VPB VPB.t2 360.082
R29 VPB.t2 VPB.t1 311.56
R30 VPB.t1 VPB.t0 214.517
R31 VPWR VPWR.n0 238.133
R32 VPWR.n0 VPWR.t1 72.7029
R33 VPWR.n0 VPWR.t0 29.6087
R34 B_N.n0 B_N.t1 219.846
R35 B_N B_N.n0 219.404
R36 B_N.n0 B_N.t0 128.288
C0 Y VPB 0.018501f
C1 Y VGND 0.155163f
C2 VGND VPB 0.007567f
C3 Y A 0.01216f
C4 VPB A 0.034167f
C5 Y VPWR 0.085391f
C6 VGND A 0.045283f
C7 VPB VPWR 0.079209f
C8 Y B_N 7.99e-19
C9 VGND VPWR 0.04023f
C10 VPB B_N 0.058201f
C11 A VPWR 0.022418f
C12 VGND B_N 0.012616f
C13 A B_N 0.035287f
C14 VPWR B_N 0.014609f
C15 VGND VNB 0.37126f
C16 Y VNB 0.096599f
C17 B_N VNB 0.194145f
C18 VPWR VNB 0.278425f
C19 A VNB 0.118889f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2_8 VNB VPB VPWR VGND A B Y
X0 a_27_368.t7 B.t0 Y.t11 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X1 VPWR.t7 A.t0 a_27_368.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VGND.t3 A.t1 Y.t12 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 VGND.t2 A.t2 Y.t13 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2775 pd=1.49 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 VPWR.t6 A.t3 a_27_368.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_27_368.t10 A.t4 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t4 A.t5 a_27_368.t11 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t10 B.t1 a_27_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_27_368.t5 B.t2 Y.t9 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t14 A.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2775 ps=1.49 w=0.74 l=0.15
X10 a_27_368.t12 A.t7 VPWR.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X11 Y.t8 B.t3 a_27_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X12 a_27_368.t13 A.t8 VPWR.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X13 Y.t15 A.t9 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.7881 ps=3.61 w=0.74 l=0.15
X14 VGND.t7 B.t4 Y.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_27_368.t3 B.t5 Y.t7 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X16 Y.t6 B.t6 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_27_368.t1 B.t7 Y.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 Y.t3 B.t8 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X19 Y.t4 B.t9 a_27_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X20 Y.t2 B.t10 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.35705 pd=1.705 as=0.1295 ps=1.09 w=0.74 l=0.15
X21 VPWR.t1 A.t10 a_27_368.t14 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_27_368.t15 A.t11 VPWR.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X23 VGND.t4 B.t11 Y.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.35705 ps=1.705 w=0.74 l=0.15
R0 B.n1 B.t0 339.274
R1 B.n8 B.t5 339.274
R2 B.n0 B.t1 319.192
R3 B.n2 B.t9 319.192
R4 B.n4 B.t7 319.192
R5 B.n6 B.t6 319.192
R6 B.n9 B.t3 319.192
R7 B.n9 B.t2 319.192
R8 B.n0 B.t10 173.52
R9 B.n3 B.t11 142.994
R10 B.n5 B.t8 142.994
R11 B.n7 B.t4 142.994
R12 B.n4 B.n3 138.173
R13 B.n1 B.n0 131.748
R14 B.n2 B.n1 131.748
R15 B.n10 B.n8 102.828
R16 B.n6 B.n5 99.6138
R17 B.n8 B.n7 77.1205
R18 B.n11 B.n10 71.1166
R19 B.n5 B.n4 44.9872
R20 B.n7 B.n6 38.5605
R21 B.n11 B 9.45419
R22 B.n3 B.n2 6.42717
R23 B.n10 B.n9 5.7386
R24 B B.n11 4.22497
R25 Y.n5 Y.n3 264.574
R26 Y.n5 Y.n4 217.921
R27 Y Y.n0 212.524
R28 Y.n7 Y.n1 209.547
R29 Y.n17 Y.n16 185
R30 Y.n14 Y.n13 185
R31 Y.n11 Y.n9 182.275
R32 Y.n6 Y.n2 103.457
R33 Y.n11 Y.n10 101.71
R34 Y.n15 Y.n14 80.5048
R35 Y.n17 Y.n8 80.3516
R36 Y.n12 Y.n11 72.3314
R37 Y.n15 Y.n8 48.2927
R38 Y.n0 Y.t10 35.1791
R39 Y.n9 Y.t13 34.0546
R40 Y.n10 Y.t12 34.0546
R41 Y.n3 Y.t9 26.3844
R42 Y.n3 Y.t8 26.3844
R43 Y.n4 Y.t7 26.3844
R44 Y.n4 Y.t6 26.3844
R45 Y.n1 Y.t5 26.3844
R46 Y.n1 Y.t4 26.3844
R47 Y.n0 Y.t11 26.3844
R48 Y.n13 Y.n8 24.2999
R49 Y.n16 Y.n15 23.9934
R50 Y.n13 Y.t1 22.7032
R51 Y.n16 Y.t2 22.7032
R52 Y.n9 Y.t15 22.7032
R53 Y.n10 Y.t14 22.7032
R54 Y.n2 Y.t0 22.7032
R55 Y.n2 Y.t3 22.7032
R56 Y.n7 Y.n6 13.7162
R57 Y.n18 Y.n17 7.36794
R58 Y.n18 Y.n7 5.1005
R59 Y.n14 Y.n12 4.68887
R60 Y.n6 Y.n5 4.13831
R61 Y.n17 Y.n12 2.0098
R62 Y Y.n18 1.78655
R63 a_27_368.n9 a_27_368.t5 296.887
R64 a_27_368.n1 a_27_368.t8 293.865
R65 a_27_368.n11 a_27_368.n10 219.754
R66 a_27_368.n9 a_27_368.n8 214.609
R67 a_27_368.n13 a_27_368.n12 212.934
R68 a_27_368.n1 a_27_368.n0 208.185
R69 a_27_368.n3 a_27_368.n2 205.916
R70 a_27_368.n5 a_27_368.n4 205.916
R71 a_27_368.n7 a_27_368.n6 188.462
R72 a_27_368.n12 a_27_368.n7 72.6101
R73 a_27_368.n7 a_27_368.n5 65.3196
R74 a_27_368.n3 a_27_368.n1 61.3652
R75 a_27_368.n5 a_27_368.n3 52.7064
R76 a_27_368.n11 a_27_368.n9 52.3299
R77 a_27_368.n12 a_27_368.n11 51.9534
R78 a_27_368.n8 a_27_368.t3 35.1791
R79 a_27_368.t7 a_27_368.n13 35.1791
R80 a_27_368.n8 a_27_368.t4 26.3844
R81 a_27_368.n10 a_27_368.t2 26.3844
R82 a_27_368.n10 a_27_368.t1 26.3844
R83 a_27_368.n0 a_27_368.t11 26.3844
R84 a_27_368.n0 a_27_368.t13 26.3844
R85 a_27_368.n2 a_27_368.t9 26.3844
R86 a_27_368.n2 a_27_368.t10 26.3844
R87 a_27_368.n4 a_27_368.t14 26.3844
R88 a_27_368.n4 a_27_368.t15 26.3844
R89 a_27_368.n6 a_27_368.t6 26.3844
R90 a_27_368.n6 a_27_368.t12 26.3844
R91 a_27_368.n13 a_27_368.t0 26.3844
R92 VPB.t14 VPB.t12 280.914
R93 VPB VPB.t8 257.93
R94 VPB.t3 VPB.t4 255.376
R95 VPB.t7 VPB.t0 255.376
R96 VPB.t6 VPB.t7 255.376
R97 VPB.t9 VPB.t15 255.376
R98 VPB.t8 VPB.t13 255.376
R99 VPB.t4 VPB.t5 229.839
R100 VPB.t2 VPB.t3 229.839
R101 VPB.t1 VPB.t2 229.839
R102 VPB.t0 VPB.t1 229.839
R103 VPB.t12 VPB.t6 229.839
R104 VPB.t15 VPB.t14 229.839
R105 VPB.t10 VPB.t9 229.839
R106 VPB.t11 VPB.t10 229.839
R107 VPB.t13 VPB.t11 229.839
R108 A.n5 A.t0 360.5
R109 A.n1 A.t7 236.496
R110 A.n17 A.t10 214.758
R111 A.n14 A.t11 214.758
R112 A.n3 A.t3 214.758
R113 A.n8 A.t4 214.758
R114 A.n5 A.t8 204.048
R115 A.n6 A.t5 204.048
R116 A.n7 A.t9 196.013
R117 A.n4 A.t2 196.013
R118 A.n16 A.t6 196.013
R119 A.n1 A.t1 196.013
R120 A.n19 A.n18 152
R121 A.n15 A.n0 152
R122 A.n13 A.n12 152
R123 A.n11 A.n2 152
R124 A.n10 A.n9 152
R125 A.n6 A.n5 132.423
R126 A.n7 A.n6 93.5254
R127 A.n13 A.n2 43.7018
R128 A.n18 A.n1 37.2752
R129 A.n9 A.n4 32.1338
R130 A.n15 A.n14 28.9205
R131 A.n9 A.n8 19.9232
R132 A.n16 A.n15 16.7098
R133 A.n18 A.n17 14.7818
R134 A.n14 A.n13 14.7818
R135 A.n10 A 13.8424
R136 A.n17 A.n16 12.2112
R137 A.n8 A.n7 12.2112
R138 A.n19 A.n0 10.1214
R139 A.n11 A 9.67492
R140 A.n12 A 8.7819
R141 A.n3 A.n2 5.7845
R142 A.n4 A.n3 5.7845
R143 A.n12 A 5.50748
R144 A A.n11 4.61445
R145 A A.n19 2.82841
R146 A A.n0 1.34003
R147 A A.n10 0.447012
R148 VPWR.n7 VPWR.n6 321.514
R149 VPWR.n12 VPWR.n1 317.526
R150 VPWR.n10 VPWR.n3 315.928
R151 VPWR.n5 VPWR.n4 315.928
R152 VPWR.n1 VPWR.t7 35.1791
R153 VPWR.n4 VPWR.t6 35.1791
R154 VPWR.n6 VPWR.t3 35.1791
R155 VPWR.n6 VPWR.t1 35.1791
R156 VPWR.n1 VPWR.t2 26.3844
R157 VPWR.n3 VPWR.t5 26.3844
R158 VPWR.n3 VPWR.t4 26.3844
R159 VPWR.n4 VPWR.t0 26.3844
R160 VPWR.n11 VPWR.n10 23.7181
R161 VPWR.n10 VPWR.n9 23.7181
R162 VPWR.n9 VPWR.n5 22.9652
R163 VPWR.n12 VPWR.n11 19.2005
R164 VPWR.n9 VPWR.n8 9.3005
R165 VPWR.n10 VPWR.n2 9.3005
R166 VPWR.n11 VPWR.n0 9.3005
R167 VPWR.n13 VPWR.n12 7.43488
R168 VPWR.n7 VPWR.n5 6.7615
R169 VPWR.n8 VPWR.n7 0.551893
R170 VPWR VPWR.n13 0.160103
R171 VPWR.n13 VPWR.n0 0.1477
R172 VPWR.n8 VPWR.n2 0.122949
R173 VPWR.n2 VPWR.n0 0.122949
R174 VGND.n7 VGND.n6 211.183
R175 VGND.n19 VGND.n4 185
R176 VGND.n21 VGND.n20 185
R177 VGND.n3 VGND.n0 185
R178 VGND.n28 VGND.n27 185
R179 VGND.n29 VGND.n28 185
R180 VGND.n28 VGND.n0 185
R181 VGND.n9 VGND.t7 160.166
R182 VGND.n11 VGND.n10 115.841
R183 VGND.n3 VGND.n2 91.5754
R184 VGND.n20 VGND.n19 76.2167
R185 VGND.n13 VGND.n12 36.1417
R186 VGND.n18 VGND.n17 36.1417
R187 VGND.n26 VGND.n25 35.4941
R188 VGND.n13 VGND.n7 35.3887
R189 VGND.n10 VGND.t6 34.0546
R190 VGND.n10 VGND.t4 34.0546
R191 VGND.n6 VGND.t5 34.0546
R192 VGND.n12 VGND.n11 30.4946
R193 VGND.n28 VGND.t0 25.3526
R194 VGND.t0 VGND.n3 25.3526
R195 VGND.n20 VGND.t1 22.7032
R196 VGND.n19 VGND.t2 22.7032
R197 VGND.n6 VGND.t3 22.7032
R198 VGND.n25 VGND.n4 17.3426
R199 VGND.n17 VGND.n7 12.0476
R200 VGND.n31 VGND.n30 9.3005
R201 VGND.n12 VGND.n8 9.3005
R202 VGND.n14 VGND.n13 9.3005
R203 VGND.n15 VGND.n7 9.3005
R204 VGND.n17 VGND.n16 9.3005
R205 VGND.n18 VGND.n5 9.3005
R206 VGND.n23 VGND.n22 9.3005
R207 VGND.n25 VGND.n24 9.3005
R208 VGND.n26 VGND.n1 9.3005
R209 VGND.n32 VGND.n0 9.2982
R210 VGND.n11 VGND.n9 6.37487
R211 VGND.n22 VGND.n21 4.91293
R212 VGND.n21 VGND.n18 3.57392
R213 VGND.n30 VGND.n0 3.31902
R214 VGND.n27 VGND.n2 1.85225
R215 VGND.n29 VGND.n2 1.85225
R216 VGND.n22 VGND.n4 1.59185
R217 VGND.n27 VGND.n26 0.895973
R218 VGND.n9 VGND.n8 0.499401
R219 VGND.n30 VGND.n29 0.421899
R220 VGND VGND.n32 0.16175
R221 VGND.n32 VGND.n31 0.146075
R222 VGND.n14 VGND.n8 0.122949
R223 VGND.n15 VGND.n14 0.122949
R224 VGND.n16 VGND.n15 0.122949
R225 VGND.n16 VGND.n5 0.122949
R226 VGND.n23 VGND.n5 0.122949
R227 VGND.n24 VGND.n23 0.122949
R228 VGND.n24 VGND.n1 0.122949
R229 VGND.n31 VGND.n1 0.122949
R230 VNB VNB.t0 4180.58
R231 VNB.t5 VNB.t4 2575.33
R232 VNB.t2 VNB.t1 2078.74
R233 VNB.t4 VNB.t6 1316.54
R234 VNB.t3 VNB.t5 1154.86
R235 VNB.t1 VNB.t3 1154.86
R236 VNB.t0 VNB.t2 1154.86
R237 VNB.t6 VNB.t7 993.177
C0 VPB VGND 0.008989f
C1 B Y 0.397665f
C2 A VGND 0.112181f
C3 VPWR Y 0.0493f
C4 B VGND 0.193066f
C5 VPWR VGND 0.132435f
C6 Y VGND 0.829006f
C7 VPB A 0.290559f
C8 VPB B 0.246123f
C9 A B 0.049503f
C10 VPB VPWR 0.182009f
C11 VPB Y 0.020532f
C12 A VPWR 0.164771f
C13 B VPWR 0.044843f
C14 A Y 0.241778f
C15 VGND VNB 1.00792f
C16 Y VNB 0.087975f
C17 VPWR VNB 0.73751f
C18 B VNB 0.992507f
C19 A VNB 0.697252f
C20 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2_4 VNB VPB VPWR VGND Y A B
X0 VPWR.t3 A.t0 a_27_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t4 A.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.4218 pd=1.88 as=0.2294 ps=2.1 w=0.74 l=0.15
X2 Y.t5 B.t0 a_27_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X3 Y.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1221 ps=1.07 w=0.74 l=0.15
X4 a_27_368.t0 B.t2 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VGND.t1 A.t2 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.4218 ps=1.88 w=0.74 l=0.15
X6 Y.t2 B.t3 a_27_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_27_368.t2 A.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t1 A.t4 a_27_368.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_27_368.t4 A.t5 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_27_368.t7 B.t4 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3976 pd=2.95 as=0.196 ps=1.47 w=1.12 l=0.15
X11 VGND.t3 B.t5 Y.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.0138 pd=4.22 as=0.111 ps=1.04 w=0.74 l=0.15
R0 A.n1 A.t3 268.815
R1 A.n8 A.t0 263.81
R2 A.n3 A.t4 261.62
R3 A.n0 A.t5 261.62
R4 A.n8 A.t1 154.24
R5 A.n1 A.t2 154.24
R6 A.n2 A 153.212
R7 A.n5 A.n4 152
R8 A.n7 A.n6 152
R9 A.n10 A.n9 152
R10 A.n9 A.n7 49.6611
R11 A.n4 A.n0 48.9308
R12 A.n3 A.n2 32.8641
R13 A.n2 A.n1 26.2914
R14 A.n4 A.n3 16.7975
R15 A A.n10 15.741
R16 A.n9 A.n8 13.146
R17 A.n6 A 10.8978
R18 A.n5 A 10.5519
R19 A A.n5 6.05455
R20 A.n6 A 5.70861
R21 A.n10 A 0.865365
R22 A.n7 A.n0 0.730803
R23 a_27_368.n4 a_27_368.t7 290.063
R24 a_27_368.n1 a_27_368.t3 280.005
R25 a_27_368.n1 a_27_368.n0 210.702
R26 a_27_368.n5 a_27_368.n4 208.577
R27 a_27_368.n3 a_27_368.n2 186.857
R28 a_27_368.n4 a_27_368.n3 76.8239
R29 a_27_368.n3 a_27_368.n1 69.5234
R30 a_27_368.t0 a_27_368.n5 35.1791
R31 a_27_368.n2 a_27_368.t1 26.3844
R32 a_27_368.n2 a_27_368.t2 26.3844
R33 a_27_368.n0 a_27_368.t5 26.3844
R34 a_27_368.n0 a_27_368.t4 26.3844
R35 a_27_368.n5 a_27_368.t6 26.3844
R36 VPWR.n2 VPWR.n1 344.329
R37 VPWR.n2 VPWR.n0 342.296
R38 VPWR.n0 VPWR.t0 26.3844
R39 VPWR.n0 VPWR.t3 26.3844
R40 VPWR.n1 VPWR.t2 26.3844
R41 VPWR.n1 VPWR.t1 26.3844
R42 VPWR VPWR.n2 0.518338
R43 VPB VPB.t5 257.93
R44 VPB.t6 VPB.t7 255.376
R45 VPB.t0 VPB.t6 255.376
R46 VPB.t1 VPB.t0 229.839
R47 VPB.t4 VPB.t1 229.839
R48 VPB.t3 VPB.t4 229.839
R49 VPB.t2 VPB.t3 229.839
R50 VPB.t5 VPB.t2 229.839
R51 VGND.n3 VGND.n2 206.333
R52 VGND.n9 VGND.t2 136.739
R53 VGND.n4 VGND.t3 83.95
R54 VGND.n7 VGND.n1 36.1417
R55 VGND.n8 VGND.n7 36.1417
R56 VGND.n2 VGND.t0 30.8113
R57 VGND.n2 VGND.t1 22.7032
R58 VGND.n9 VGND.n8 18.824
R59 VGND.n3 VGND.n1 13.5534
R60 VGND.n10 VGND.n9 9.3005
R61 VGND.n5 VGND.n1 9.3005
R62 VGND.n7 VGND.n6 9.3005
R63 VGND.n8 VGND.n0 9.3005
R64 VGND.n4 VGND.n3 7.27433
R65 VGND.n5 VGND.n4 0.422662
R66 VGND.n6 VGND.n5 0.122949
R67 VGND.n6 VGND.n0 0.122949
R68 VGND.n10 VGND.n0 0.122949
R69 VGND VGND.n10 0.0617245
R70 Y.n2 Y.n0 259.024
R71 Y.n2 Y.n1 208.577
R72 Y.n5 Y.n3 95.9272
R73 Y.n5 Y.n4 70.6316
R74 Y.n4 Y.t4 66.9203
R75 Y.n4 Y.t3 60.884
R76 Y.n0 Y.t5 35.1791
R77 Y.n1 Y.t1 26.3844
R78 Y.n1 Y.t2 26.3844
R79 Y.n0 Y.t7 26.3844
R80 Y.n3 Y.t0 25.9464
R81 Y.n3 Y.t6 22.7032
R82 Y.n6 Y.n2 19.7823
R83 Y Y.n5 10.2747
R84 Y Y.n6 7.7918
R85 Y.n6 Y 3.29747
R86 VNB.t2 VNB.t1 2979.53
R87 VNB VNB.t2 1201.05
R88 VNB.t1 VNB.t0 1108.66
R89 VNB.t0 VNB.t3 1039.37
R90 B.n0 B.t4 261.62
R91 B.n6 B.t0 261.62
R92 B.n5 B.t2 261.62
R93 B.n3 B.t3 261.62
R94 B B.n0 189.764
R95 B.n3 B.t1 156.431
R96 B.n4 B.t5 154.24
R97 B.n2 B.n1 152
R98 B.n8 B.n7 152
R99 B.n6 B.n5 73.0308
R100 B.n4 B.n3 63.5369
R101 B.n7 B.n2 49.6611
R102 B.n2 B.n0 12.4157
R103 B.n1 B 11.2437
R104 B.n7 B.n6 10.955
R105 B B.n8 10.2059
R106 B.n8 B 6.4005
R107 B.n1 B 5.36266
R108 B.n5 B.n4 2.19141
C0 VPB B 0.148195f
C1 VGND VPWR 0.072331f
C2 A B 0.054778f
C3 VPB VPWR 0.103466f
C4 VGND Y 0.378655f
C5 VPB Y 0.009132f
C6 A VPWR 0.06943f
C7 B VPWR 0.024856f
C8 A Y 0.148654f
C9 B Y 0.224289f
C10 VPWR Y 0.023409f
C11 VGND VPB 0.006374f
C12 VGND A 0.076873f
C13 VPB A 0.127101f
C14 VGND B 0.160967f
C15 VGND VNB 0.585935f
C16 Y VNB 0.04079f
C17 VPWR VNB 0.425675f
C18 B VNB 0.432842f
C19 A VNB 0.402447f
C20 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2_2 VNB VPB VPWR VGND B Y A
X0 a_35_368.t3 B.t0 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t3 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X2 Y.t1 B.t2 a_35_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 VGND.t0 A.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_35_368.t0 A.t1 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t0 A.t2 a_35_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B.n0 B.t0 318.12
R1 B.n0 B.t2 223.588
R2 B.n1 B.t1 169.389
R3 B B.n1 158.788
R4 B.n1 B.n0 51.6247
R5 Y.n0 Y 594.413
R6 Y.n1 Y.n0 585
R7 Y Y.n2 134.726
R8 Y.n0 Y.t2 26.3844
R9 Y.n0 Y.t1 26.3844
R10 Y.n2 Y.t0 22.7032
R11 Y.n2 Y.t3 22.7032
R12 Y.n1 Y 12.6123
R13 Y Y.n1 1.31815
R14 a_35_368.t2 a_35_368.n1 339.568
R15 a_35_368.n1 a_35_368.t0 322.969
R16 a_35_368.n1 a_35_368.n0 181.875
R17 a_35_368.n0 a_35_368.t1 26.3844
R18 a_35_368.n0 a_35_368.t3 26.3844
R19 VPB VPB.t2 278.361
R20 VPB.t1 VPB.t0 229.839
R21 VPB.t3 VPB.t1 229.839
R22 VPB.t2 VPB.t3 229.839
R23 VGND.n0 VGND.t0 160.304
R24 VGND.n0 VGND.t1 156.738
R25 VGND VGND.n0 0.440377
R26 VNB VNB.t1 1304.99
R27 VNB.t1 VNB.t0 993.177
R28 A.n1 A.t1 487.892
R29 A.n0 A.t0 269.385
R30 A.n0 A.t2 250.909
R31 A A.n1 158.611
R32 A.n4 A.n3 152
R33 A.n3 A.n2 134.736
R34 A.n1 A.n0 62.482
R35 A.n3 A.n1 12.4157
R36 A.n4 A 7.08135
R37 A.n2 A 5.48544
R38 A.n2 A 4.42139
R39 A A.n4 2.99624
R40 VPWR VPWR.n0 331.99
R41 VPWR.n0 VPWR.t1 26.3844
R42 VPWR.n0 VPWR.t0 26.3844
C0 A VPWR 0.041155f
C1 VPB VGND 0.006362f
C2 B VPWR 0.012175f
C3 A VGND 0.143282f
C4 Y VPWR 0.010345f
C5 B VGND 0.05451f
C6 Y VGND 0.159285f
C7 VPWR VGND 0.039532f
C8 VPB A 0.074595f
C9 VPB B 0.076044f
C10 B A 0.055802f
C11 VPB Y 0.004411f
C12 A Y 0.035491f
C13 VPB VPWR 0.063783f
C14 B Y 0.0875f
C15 VGND VNB 0.37006f
C16 VPWR VNB 0.264268f
C17 Y VNB 0.028308f
C18 A VNB 0.452763f
C19 B VNB 0.219612f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3b_1 VNB VPB VPWR VGND Y C_N A B
X0 VGND.t0 B.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1184 ps=1.06 w=0.74 l=0.15
X1 VPWR.t0 C_N.t0 a_27_112.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2177 pd=1.54 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 a_344_368.t0 B.t1 a_260_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X3 a_260_368.t1 A.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.2177 ps=1.54 w=1.12 l=0.15
X4 Y.t1 a_27_112.t2 a_344_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X5 Y.t2 a_27_112.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X6 Y.t3 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.137175 ps=1.13 w=0.74 l=0.15
X7 VGND.t2 C_N.t1 a_27_112.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.137175 pd=1.13 as=0.2695 ps=2.08 w=0.55 l=0.15
R0 B.n0 B.t1 250.909
R1 B.n0 B.t0 220.113
R2 B B.n0 155.721
R3 Y.n1 Y.t1 411.062
R4 Y.t2 Y.n2 279.738
R5 Y.n3 Y.t2 279.738
R6 Y.n1 Y.n0 152.159
R7 Y.n0 Y.t3 29.1897
R8 Y.n0 Y.t0 22.7032
R9 Y.n3 Y 8.94674
R10 Y.n2 Y.n1 3.57899
R11 Y.n2 Y 3.44136
R12 Y Y.n3 1.23921
R13 VGND.n2 VGND.n0 216.605
R14 VGND.n2 VGND.n1 126.115
R15 VGND.n1 VGND.t2 49.0811
R16 VGND.n0 VGND.t1 34.0546
R17 VGND.n0 VGND.t0 34.0546
R18 VGND.n1 VGND.t3 24.2235
R19 VGND VGND.n2 0.538326
R20 VNB VNB.t2 1616.8
R21 VNB.t0 VNB.t1 1316.54
R22 VNB.t2 VNB.t3 1247.24
R23 VNB.t3 VNB.t0 1085.56
R24 C_N.n0 C_N.t0 240.732
R25 C_N C_N.n0 158.054
R26 C_N.n0 C_N.t1 147.814
R27 a_27_112.t0 a_27_112.n0 387.56
R28 a_27_112.n0 a_27_112.n1 300.329
R29 a_27_112.n0 a_27_112.t1 293.592
R30 a_27_112.n1 a_27_112.t2 250.909
R31 a_27_112.n1 a_27_112.t3 220.113
R32 VPWR VPWR.n0 343.911
R33 VPWR.n0 VPWR.t0 63.3219
R34 VPWR.n0 VPWR.t1 29.6087
R35 VPB VPB.t1 334.543
R36 VPB.t0 VPB.t2 291.13
R37 VPB.t1 VPB.t3 291.13
R38 VPB.t3 VPB.t0 214.517
R39 a_260_368.t0 a_260_368.t1 47.4916
R40 a_344_368.t0 a_344_368.t1 73.8755
R41 A.n0 A.t0 250.909
R42 A.n0 A.t1 220.113
R43 A A.n0 154.522
C0 VPB C_N 0.040031f
C1 C_N Y 0.00376f
C2 A C_N 0.060042f
C3 C_N VGND 0.016423f
C4 B C_N 4.14e-19
C5 VPB Y 0.023944f
C6 VPWR C_N 0.010853f
C7 VPB A 0.035741f
C8 VPB VGND 0.007716f
C9 A Y 0.00982f
C10 Y VGND 0.27144f
C11 VPB B 0.032857f
C12 B Y 0.048752f
C13 A VGND 0.030969f
C14 A B 0.087181f
C15 VPB VPWR 0.086098f
C16 VPWR Y 0.07323f
C17 B VGND 0.013361f
C18 A VPWR 0.017387f
C19 VPWR VGND 0.046859f
C20 B VPWR 0.011289f
C21 VGND VNB 0.402345f
C22 Y VNB 0.128622f
C23 C_N VNB 0.144277f
C24 VPWR VNB 0.318352f
C25 B VNB 0.105065f
C26 A VNB 0.110554f
C27 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3_4 VNB VPB VPWR VGND A B C Y
X0 Y.t9 C.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1 a_295_368.t7 C.t1 Y.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2744 pd=1.7 as=0.26145 ps=1.64 w=1.12 l=0.15
X2 VGND.t3 B.t0 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 a_27_368.t7 A.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_295_368.t2 B.t1 a_27_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2713 pd=1.695 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_295_368.t3 B.t2 a_27_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VPWR.t1 A.t2 a_27_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_27_368.t5 A.t3 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_27_368.t1 B.t3 a_295_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2744 ps=1.7 w=1.12 l=0.15
X10 a_27_368.t0 B.t4 a_295_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t1 B.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1517 ps=1.15 w=0.74 l=0.15
X12 VGND.t2 A.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1517 pd=1.15 as=0.1073 ps=1.03 w=0.74 l=0.15
X13 VGND.t4 C.t2 Y.t8 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.40425 pd=2.58 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 Y.t6 C.t3 a_295_368.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.26145 pd=1.64 as=0.2713 ps=1.695 w=1.12 l=0.15
X15 Y.t5 C.t4 a_295_368.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.26145 pd=1.64 as=0.2744 ps=1.7 w=1.12 l=0.15
X16 VPWR.t3 A.t5 a_27_368.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
X17 a_295_368.t4 C.t5 Y.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2744 pd=1.7 as=0.26145 ps=1.64 w=1.12 l=0.15
R0 C.n1 C.t3 371.409
R1 C.n6 C.n5 318.777
R2 C.n1 C.t0 258.673
R3 C.n3 C.t2 258.673
R4 C.n5 C.t5 242.875
R5 C.n2 C.t1 222.792
R6 C.n4 C.t4 204.048
R7 C.n5 C.n4 154.679
R8 C.n6 C 153.745
R9 C.n9 C.n0 152
R10 C.n8 C.n7 152
R11 C.n10 C.n0 133.218
R12 C.n3 C.n2 102.828
R13 C.n4 C.n3 83.9853
R14 C.n7 C.n0 49.6611
R15 C.n7 C.n6 49.6611
R16 C.n2 C.n1 35.3472
R17 C C.n9 12.6066
R18 C C.n10 12.099
R19 C.n8 C 11.4429
R20 C C.n8 7.17626
R21 C.n10 C 6.04708
R22 C.n9 C 6.01262
R23 VGND.n5 VGND.t4 263.688
R24 VGND.n8 VGND.n2 211.183
R25 VGND.n4 VGND.n3 206.333
R26 VGND.n10 VGND.t0 171.77
R27 VGND.n3 VGND.t5 34.0546
R28 VGND.n3 VGND.t3 34.0546
R29 VGND.n2 VGND.t1 34.0546
R30 VGND.n2 VGND.t2 32.4329
R31 VGND.n4 VGND.n1 27.4829
R32 VGND.n10 VGND.n9 26.7299
R33 VGND.n9 VGND.n8 24.4711
R34 VGND.n8 VGND.n1 22.9652
R35 VGND.n11 VGND.n10 9.3005
R36 VGND.n6 VGND.n1 9.3005
R37 VGND.n8 VGND.n7 9.3005
R38 VGND.n9 VGND.n0 9.3005
R39 VGND.n5 VGND.n4 6.58038
R40 VGND.n6 VGND.n5 0.497297
R41 VGND.n7 VGND.n6 0.122949
R42 VGND.n7 VGND.n0 0.122949
R43 VGND.n11 VGND.n0 0.122949
R44 VGND VGND.n11 0.0617245
R45 Y.n3 Y.n1 645.105
R46 Y.n3 Y.n2 585
R47 Y.n5 Y.n3 349.565
R48 Y.n5 Y.n4 96.3134
R49 Y.n6 Y.n0 95.9272
R50 Y.n8 Y.n7 88.3339
R51 Y.n8 Y.n6 69.6083
R52 Y.n6 Y.n5 51.2526
R53 Y.n2 Y.t4 39.5764
R54 Y.n2 Y.t5 39.5764
R55 Y.n1 Y.t7 39.5764
R56 Y.n1 Y.t6 39.5764
R57 Y.n7 Y.t2 24.3248
R58 Y.n7 Y.t0 22.7032
R59 Y.n0 Y.t3 22.7032
R60 Y.n0 Y.t1 22.7032
R61 Y.n4 Y.t8 22.7032
R62 Y.n4 Y.t9 22.7032
R63 Y Y.n8 10.0806
R64 VNB.t4 VNB 11016.2
R65 VNB VNB.n0 4268.12
R66 VNB.t3 VNB.t5 1366.76
R67 VNB.t1 VNB.t2 1293.44
R68 VNB.t0 VNB 1143.31
R69 VNB.t5 VNB.t4 1031.06
R70 VNB.t2 VNB.t0 1016.27
R71 VNB.n0 VNB.t1 658.269
R72 VNB.n0 VNB.t3 347.685
R73 a_295_368.n5 a_295_368.n4 653.552
R74 a_295_368.n2 a_295_368.n0 650.698
R75 a_295_368.n2 a_295_368.n1 585
R76 a_295_368.n4 a_295_368.n3 585
R77 a_295_368.n4 a_295_368.n2 68.8361
R78 a_295_368.n5 a_295_368.t2 40.4559
R79 a_295_368.n3 a_295_368.t5 40.4559
R80 a_295_368.n3 a_295_368.t7 40.4559
R81 a_295_368.n1 a_295_368.t0 40.4559
R82 a_295_368.n1 a_295_368.t4 40.4559
R83 a_295_368.t6 a_295_368.n5 39.5764
R84 a_295_368.n0 a_295_368.t1 26.3844
R85 a_295_368.n0 a_295_368.t3 26.3844
R86 VPB.t8 VPB 1948.52
R87 VPB VPB.n0 876.167
R88 VPB.t8 VPB.t0 307.659
R89 VPB.t11 VPB.t9 300.26
R90 VPB.t9 VPB.t8 295.337
R91 VPB.t10 VPB.t11 295.337
R92 VPB.t2 VPB 255.376
R93 VPB.t6 VPB.t4 229.839
R94 VPB.t1 VPB.t6 229.839
R95 VPB.t5 VPB.t1 229.839
R96 VPB.t0 VPB.t5 229.839
R97 VPB.t3 VPB.t7 229.839
R98 VPB.t7 VPB.t2 229.839
R99 VPB.n0 VPB.t3 194.087
R100 VPB.n0 VPB.t10 110.751
R101 B.n0 B.t4 338.058
R102 B.n1 B.t3 298.019
R103 B.n0 B.t2 272.33
R104 B.n3 B.t1 250.909
R105 B.n2 B.t0 234.573
R106 B B.n3 190.024
R107 B.n2 B.t5 153.948
R108 B B.n1 142.107
R109 B.n3 B.n2 37.246
R110 B.n1 B.n0 33.3172
R111 A A.n0 409.267
R112 A.n1 A.t3 229
R113 A.n0 A.t2 228.877
R114 A.n0 A.t1 228.877
R115 A.n2 A.t5 206.865
R116 A.n2 A.t0 197.465
R117 A.n1 A.t4 196.013
R118 A A.n3 168.874
R119 A.n3 A.n2 38.7131
R120 A.n3 A.n1 24.1005
R121 VPWR.n2 VPWR.n0 612.751
R122 VPWR.n2 VPWR.n1 611.798
R123 VPWR.n1 VPWR.t0 26.3844
R124 VPWR.n1 VPWR.t3 26.3844
R125 VPWR.n0 VPWR.t2 26.3844
R126 VPWR.n0 VPWR.t1 26.3844
R127 VPWR VPWR.n2 0.19128
R128 a_27_368.n3 a_27_368.n2 585
R129 a_27_368.n1 a_27_368.n0 298.132
R130 a_27_368.n5 a_27_368.n4 293.13
R131 a_27_368.n1 a_27_368.t7 288.197
R132 a_27_368.n4 a_27_368.t4 285.731
R133 a_27_368.n4 a_27_368.n3 246.794
R134 a_27_368.n3 a_27_368.n1 64.2665
R135 a_27_368.n2 a_27_368.t2 26.3844
R136 a_27_368.n2 a_27_368.t1 26.3844
R137 a_27_368.n0 a_27_368.t6 26.3844
R138 a_27_368.n0 a_27_368.t0 26.3844
R139 a_27_368.t3 a_27_368.n5 26.3844
R140 a_27_368.n5 a_27_368.t5 26.3844
C0 VPB A 0.134955f
C1 VPB C 0.18606f
C2 VPB B 0.134923f
C3 A C 0.09844f
C4 VPB Y 0.015339f
C5 VPB VPWR 0.149567f
C6 A B 0.193763f
C7 VPB VGND 0.008381f
C8 A Y 0.407894f
C9 B C 0.191763f
C10 A VPWR 0.091626f
C11 C Y 0.23509f
C12 VPWR C 0.020247f
C13 A VGND 0.097975f
C14 B Y 0.634772f
C15 B VPWR 0.031624f
C16 C VGND 0.234007f
C17 B VGND 0.048569f
C18 VPWR Y 0.01923f
C19 Y VGND 0.505644f
C20 VPWR VGND 0.103916f
C21 VGND VNB 0.838362f
C22 Y VNB 0.064409f
C23 C VNB 0.65987f
C24 VPWR VNB 0.631469f
C25 B VNB 0.40104f
C26 A VNB 0.589002f
C27 VPB VNB 1.60194f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3_2 VNB VPB VPWR VGND Y A B C
X0 a_306_368.t2 A.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X1 Y.t3 C.t0 a_27_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VGND.t2 C.t1 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.32745 pd=1.625 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_306_368.t3 B.t0 a_27_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t0 A.t1 a_306_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.1848 ps=1.45 w=1.12 l=0.15
X5 a_27_368.t2 C.t2 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6 VGND.t1 A.t2 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 Y.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.32745 ps=1.625 w=0.74 l=0.15
X8 a_27_368.t0 B.t2 a_306_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n0 A.t1 349.719
R1 A.n1 A.t0 339.274
R2 A A.n1 207.256
R3 A.n0 A.t2 142.994
R4 A.n1 A.n0 91.5805
R5 VPWR VPWR.n0 321.695
R6 VPWR.n0 VPWR.t0 29.9023
R7 VPWR.n0 VPWR.t1 26.3844
R8 a_306_368.n1 a_306_368.n0 456.05
R9 a_306_368.n0 a_306_368.t1 31.6612
R10 a_306_368.n0 a_306_368.t3 26.3844
R11 a_306_368.n1 a_306_368.t0 26.3844
R12 a_306_368.t2 a_306_368.n1 26.3844
R13 VPB VPB.t5 257.93
R14 VPB.t5 VPB.t4 255.376
R15 VPB.t3 VPB.t1 245.161
R16 VPB.t1 VPB.t2 240.054
R17 VPB.t2 VPB.t0 229.839
R18 VPB.t4 VPB.t3 229.839
R19 C.n0 C.t0 248.101
R20 C.n0 C.t2 213.419
R21 C.n1 C.t1 212.081
R22 C C.n1 158.054
R23 C.n1 C.n0 32.1338
R24 a_27_368.t0 a_27_368.n1 407.296
R25 a_27_368.n1 a_27_368.t3 330.507
R26 a_27_368.n1 a_27_368.n0 181.875
R27 a_27_368.n0 a_27_368.t1 26.3844
R28 a_27_368.n0 a_27_368.t2 26.3844
R29 Y.n3 Y.t4 279.738
R30 Y.t4 Y.n2 262.896
R31 Y Y.n1 240.155
R32 Y.n2 Y.n0 188.237
R33 Y.n1 Y.t3 35.1791
R34 Y.n0 Y.t0 34.0546
R35 Y.n1 Y.t2 26.3844
R36 Y.n0 Y.t1 22.7032
R37 Y.n2 Y 13.9641
R38 Y Y.n3 12.6066
R39 Y Y.n2 3.29747
R40 Y.n3 Y 1.74595
R41 VGND.n4 VGND.n3 185
R42 VGND.n2 VGND.n0 185
R43 VGND.n1 VGND.t1 159.198
R44 VGND.n3 VGND.n2 86.7573
R45 VGND.n2 VGND.t2 34.0546
R46 VGND.n4 VGND.n1 24.3676
R47 VGND.n3 VGND.t0 22.7032
R48 VGND.n6 VGND.n5 9.3005
R49 VGND.n7 VGND.n0 8.54972
R50 VGND.n5 VGND.n0 7.31479
R51 VGND.n5 VGND.n4 2.00322
R52 VGND.n6 VGND.n1 1.29816
R53 VGND VGND.n7 0.161024
R54 VGND.n7 VGND.n6 0.146791
R55 VNB.t2 VNB.t0 2390.55
R56 VNB.t0 VNB.t1 1154.86
R57 VNB VNB.t2 1143.31
R58 B.n1 B.t2 422.214
R59 B.n0 B.t0 285.719
R60 B.n1 B.n0 258.632
R61 B.n0 B.t1 178.34
R62 B B.n1 6.78838
C0 VPB VGND 0.005038f
C1 C VPWR 0.011702f
C2 B VPWR 0.02294f
C3 C VGND 0.021436f
C4 A VPWR 0.036837f
C5 B VGND 0.052001f
C6 VPB C 0.064689f
C7 A VGND 0.168714f
C8 Y VPWR 0.012795f
C9 VPB B 0.070574f
C10 Y VGND 0.291425f
C11 C B 0.073859f
C12 VPB A 0.060242f
C13 VPB Y 0.006526f
C14 C A 2.99e-19
C15 B A 0.184267f
C16 C Y 0.154447f
C17 B Y 0.057607f
C18 A Y 0.014269f
C19 VPWR VGND 0.054353f
C20 VPB VPWR 0.080762f
C21 VGND VNB 0.436777f
C22 VPWR VNB 0.341607f
C23 Y VNB 0.090648f
C24 A VNB 0.38522f
C25 B VNB 0.242641f
C26 C VNB 0.20177f
C27 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3_1 VNB VPB VPWR VGND Y C B A
X0 a_198_368.t1 B.t0 a_114_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.1512 ps=1.39 w=1.12 l=0.15
X1 Y.t1 C.t0 a_198_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.2016 ps=1.48 w=1.12 l=0.15
X2 Y.t0 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 Y.t2 C.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 a_114_368.t0 A.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3192 ps=2.81 w=1.12 l=0.15
X5 VGND.t2 B.t1 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 B.n0 B.t0 264.298
R1 B.n0 B.t1 204.048
R2 B B.n0 156.133
R3 a_114_368.t0 a_114_368.t1 47.4916
R4 a_198_368.t0 a_198_368.t1 63.3219
R5 VPB.t2 VPB.t0 260.485
R6 VPB VPB.t1 252.823
R7 VPB.t1 VPB.t2 214.517
R8 C.n0 C.t0 256.765
R9 C.n0 C.t1 196.516
R10 C C.n0 156.462
R11 Y.n0 Y.t1 224.066
R12 Y.n2 Y.t2 184.821
R13 Y.n3 Y.n2 111.406
R14 Y.n2 Y.n1 98.0421
R15 Y.n1 Y.t3 22.7032
R16 Y.n1 Y.t0 22.7032
R17 Y.n3 Y.n0 3.86287
R18 Y.n0 Y 1.83356
R19 Y Y.n3 1.41445
R20 A.n0 A.t1 278.188
R21 A.n0 A.t0 170.81
R22 A.n1 A.n0 152
R23 A A.n1 9.78874
R24 A.n1 A 8.78481
R25 VGND.n1 VGND.n0 211.031
R26 VGND.n1 VGND.t1 145.026
R27 VGND.n0 VGND.t0 34.0546
R28 VGND.n0 VGND.t2 22.7032
R29 VGND VGND.n1 0.5838
R30 VNB.t2 VNB.t0 1154.86
R31 VNB VNB.t1 1143.31
R32 VNB.t1 VNB.t2 993.177
R33 VPWR VPWR.t0 256.259
C0 VPB B 0.031776f
C1 VGND C 0.014622f
C2 VPB C 0.043247f
C3 A B 0.064836f
C4 B C 0.102248f
C5 VPWR Y 0.216649f
C6 VPWR VGND 0.034583f
C7 VPWR VPB 0.06115f
C8 Y VGND 0.225201f
C9 VPWR A 0.047188f
C10 Y VPB 0.018696f
C11 Y A 0.081317f
C12 VPWR B 0.00579f
C13 VGND VPB 0.004899f
C14 VPWR C 0.005673f
C15 VGND A 0.045184f
C16 Y B 0.156766f
C17 VPB A 0.03991f
C18 VGND B 0.016548f
C19 Y C 0.102193f
C20 VGND VNB 0.30715f
C21 Y VNB 0.101234f
C22 VPWR VNB 0.261552f
C23 C VNB 0.168108f
C24 B VNB 0.103448f
C25 A VNB 0.173976f
C26 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor2b_4 VNB VPB VPWR VGND A B_N Y
X0 a_116_368.t7 A.t0 VPWR.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t3 A.t1 Y.t7 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t4 A.t2 a_116_368.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.196 ps=1.47 w=1.12 l=0.15
X3 Y.t0 a_353_323.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3223 ps=2.57 w=0.74 l=0.15
X4 a_353_323.t1 B_N.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.518 pd=2.88 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 Y.t6 A.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.4097 ps=1.84 w=0.74 l=0.15
X6 a_116_368.t0 a_353_323.t4 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t2 a_353_323.t5 a_116_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_116_368.t2 a_353_323.t6 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t4 a_353_323.t7 a_116_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VPWR.t5 B_N.t1 a_353_323.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X11 a_116_368.t5 A.t4 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_353_323.t0 B_N.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.231 ps=1.555 w=0.84 l=0.15
X13 VPWR.t2 A.t5 a_116_368.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VGND.t1 a_353_323.t8 Y.t5 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.4097 pd=1.84 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n2 A.t0 384.574
R1 A.n3 A.t4 333.92
R2 A.n2 A.t5 317.853
R3 A A.n1 308.943
R4 A.n1 A.t2 281.502
R5 A.n0 A.t3 187.981
R6 A.n0 A.t1 163.278
R7 A.n2 A 158.002
R8 A.n4 A.n3 152
R9 A.n3 A.n2 49.6611
R10 A.n1 A.n0 10.8455
R11 A A.n4 9.6005
R12 A.n4 A 5.7605
R13 VPWR.n7 VPWR.t5 429.935
R14 VPWR.n17 VPWR.n1 332.039
R15 VPWR.n19 VPWR.t1 258.772
R16 VPWR.n6 VPWR.n5 221.766
R17 VPWR.n5 VPWR.t0 55.1136
R18 VPWR.n5 VPWR.t4 36.905
R19 VPWR.n10 VPWR.n4 36.1417
R20 VPWR.n11 VPWR.n10 36.1417
R21 VPWR.n12 VPWR.n11 36.1417
R22 VPWR.n12 VPWR.n2 36.1417
R23 VPWR.n16 VPWR.n2 36.1417
R24 VPWR.n18 VPWR.n17 34.6358
R25 VPWR.n19 VPWR.n18 26.7299
R26 VPWR.n1 VPWR.t3 26.3844
R27 VPWR.n1 VPWR.t2 26.3844
R28 VPWR.n6 VPWR.n4 16.1887
R29 VPWR.n8 VPWR.n4 9.3005
R30 VPWR.n10 VPWR.n9 9.3005
R31 VPWR.n11 VPWR.n3 9.3005
R32 VPWR.n13 VPWR.n12 9.3005
R33 VPWR.n14 VPWR.n2 9.3005
R34 VPWR.n16 VPWR.n15 9.3005
R35 VPWR.n18 VPWR.n0 9.3005
R36 VPWR.n20 VPWR.n19 9.3005
R37 VPWR.n7 VPWR.n6 7.07648
R38 VPWR.n17 VPWR.n16 1.50638
R39 VPWR.n8 VPWR.n7 0.544235
R40 VPWR.n9 VPWR.n8 0.122949
R41 VPWR.n9 VPWR.n3 0.122949
R42 VPWR.n13 VPWR.n3 0.122949
R43 VPWR.n14 VPWR.n13 0.122949
R44 VPWR.n15 VPWR.n14 0.122949
R45 VPWR.n15 VPWR.n0 0.122949
R46 VPWR.n20 VPWR.n0 0.122949
R47 VPWR VPWR.n20 0.0617245
R48 a_116_368.n4 a_116_368.n3 302.161
R49 a_116_368.n2 a_116_368.n0 270.921
R50 a_116_368.n5 a_116_368.n4 255.26
R51 a_116_368.n2 a_116_368.n1 186.974
R52 a_116_368.n4 a_116_368.n2 76.012
R53 a_116_368.n5 a_116_368.t0 35.1791
R54 a_116_368.n1 a_116_368.t3 26.3844
R55 a_116_368.n1 a_116_368.t5 26.3844
R56 a_116_368.n0 a_116_368.t4 26.3844
R57 a_116_368.n0 a_116_368.t7 26.3844
R58 a_116_368.n3 a_116_368.t1 26.3844
R59 a_116_368.n3 a_116_368.t2 26.3844
R60 a_116_368.t6 a_116_368.n5 26.3844
R61 VPB.t7 VPB.t0 298.791
R62 VPB VPB.t8 257.93
R63 VPB.t1 VPB.t7 255.376
R64 VPB.t0 VPB.t9 229.839
R65 VPB.t2 VPB.t1 229.839
R66 VPB.t3 VPB.t2 229.839
R67 VPB.t4 VPB.t3 229.839
R68 VPB.t6 VPB.t4 229.839
R69 VPB.t5 VPB.t6 229.839
R70 VPB.t8 VPB.t5 229.839
R71 Y.n2 Y.n1 355.812
R72 Y.n2 Y.n0 295.8
R73 Y.n5 Y.n3 286.308
R74 Y.n5 Y.n4 185
R75 Y Y.n2 160.909
R76 Y Y.n5 139.921
R77 Y.n0 Y.t3 26.3844
R78 Y.n0 Y.t4 26.3844
R79 Y.n1 Y.t1 26.3844
R80 Y.n1 Y.t2 26.3844
R81 Y.n4 Y.t5 22.7032
R82 Y.n4 Y.t0 22.7032
R83 Y.n3 Y.t7 22.7032
R84 Y.n3 Y.t6 22.7032
R85 VGND.n12 VGND.t0 334.122
R86 VGND.n3 VGND.n2 224.238
R87 VGND.n4 VGND.n1 185
R88 VGND.n6 VGND.n5 185
R89 VGND.n5 VGND.n4 62.6092
R90 VGND.n11 VGND.n10 32.4027
R91 VGND.n4 VGND.t1 31.0757
R92 VGND.n5 VGND.t2 31.0757
R93 VGND.n6 VGND.n3 26.1139
R94 VGND.n2 VGND.t4 22.7032
R95 VGND.n2 VGND.t3 22.7032
R96 VGND.n12 VGND.n11 21.0829
R97 VGND.n11 VGND.n0 9.3005
R98 VGND.n10 VGND.n9 9.3005
R99 VGND.n8 VGND.n7 9.3005
R100 VGND.n7 VGND.n1 8.42443
R101 VGND.n13 VGND.n12 7.27891
R102 VGND.n7 VGND.n6 2.07913
R103 VGND.n10 VGND.n1 2.07913
R104 VGND.n8 VGND.n3 1.60491
R105 VGND VGND.n13 0.398725
R106 VGND.n13 VGND.n0 0.155131
R107 VGND.n9 VGND.n8 0.122949
R108 VGND.n9 VGND.n0 0.122949
R109 VNB VNB.t0 4642.52
R110 VNB.t1 VNB.t2 2471.39
R111 VNB.t3 VNB.t4 993.177
R112 VNB.t2 VNB.t3 993.177
R113 VNB.t0 VNB.t1 993.177
R114 a_353_323.n10 a_353_323.n9 314.714
R115 a_353_323.n1 a_353_323.t7 236.448
R116 a_353_323.n7 a_353_323.t4 217.808
R117 a_353_323.n6 a_353_323.t5 204.048
R118 a_353_323.n2 a_353_323.t6 204.048
R119 a_353_323.n3 a_353_323.n0 165.189
R120 a_353_323.n1 a_353_323.t3 155.847
R121 a_353_323.n4 a_353_323.t8 155.847
R122 a_353_323.n5 a_353_323.n0 152
R123 a_353_323.n8 a_353_323.n7 152
R124 a_353_323.n9 a_353_323.t1 142.254
R125 a_353_323.n9 a_353_323.n8 97.2212
R126 a_353_323.n10 a_353_323.t2 35.1791
R127 a_353_323.t0 a_353_323.n10 35.1791
R128 a_353_323.n7 a_353_323.n6 27.2246
R129 a_353_323.n2 a_353_323.n1 26.332
R130 a_353_323.n5 a_353_323.n4 24.9931
R131 a_353_323.n8 a_353_323.n0 13.1884
R132 a_353_323.n3 a_353_323.n2 6.69494
R133 a_353_323.n4 a_353_323.n3 5.35606
R134 a_353_323.n6 a_353_323.n5 3.12457
R135 B_N.n0 B_N.t0 242.607
R136 B_N B_N.n1 171.317
R137 B_N.n0 B_N.t2 169.573
R138 B_N.n1 B_N.t1 159.06
R139 B_N.n1 B_N.n0 40.0769
C0 VPWR VPB 0.155812f
C1 Y VPB 0.010117f
C2 B_N VPB 0.11107f
C3 A VPB 0.128422f
C4 VGND VPB 0.00748f
C5 VPWR Y 0.047096f
C6 VPWR B_N 0.064062f
C7 A VPWR 0.070201f
C8 VPWR VGND 0.087424f
C9 Y B_N 1.24e-19
C10 A Y 0.443435f
C11 Y VGND 0.305616f
C12 A B_N 0.045619f
C13 B_N VGND 0.018733f
C14 A VGND 0.070353f
C15 VGND VNB 0.645661f
C16 B_N VNB 0.228919f
C17 Y VNB 0.112039f
C18 VPWR VNB 0.586574f
C19 A VNB 0.47117f
C20 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4bb_4 VNB VPB VPWR VGND A B Y C_N D_N
X0 a_897_349.t1 a_1162_48.t3 Y.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3668 pd=1.775 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t16 a_864_48.t3 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1295 ps=1.09 w=0.74 l=0.15
X2 a_116_368.t3 B.t0 a_27_368# VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 VPWR.t7 A.t0 a_116_368.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_116_368.t5 A.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5 a_116_368.t7 A.t2 VPWR.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.2071 pd=1.57 as=0.2184 ps=1.51 w=1.12 l=0.15
X6 VPWR.t2 D_N.t0 a_1162_48.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X7 Y.t17 B.t1 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1221 ps=1.07 w=0.74 l=0.15
X8 a_864_48.t2 C_N.t0 VGND.t16 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.34965 ps=1.685 w=0.74 l=0.15
X9 VGND.t3 a_1162_48.t4 Y.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2516 pd=1.42 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_1162_48.t0 D_N.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X11 VGND.t11 A.t3 Y.t9 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.12025 ps=1.065 w=0.74 l=0.15
X12 Y.t6 A.t4 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1443 ps=1.13 w=0.74 l=0.15
X13 VGND.t7 a_864_48.t4 Y.t8 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.34965 pd=1.685 as=0.11285 ps=1.045 w=0.74 l=0.15
X14 Y.t12 B.t2 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X15 Y.t7 A.t5 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.13875 ps=1.115 w=0.74 l=0.15
X16 VGND.t6 a_864_48.t5 Y.t15 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 VPWR.t4 A.t6 a_116_368.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X18 a_1162_48.t1 D_N.t2 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X19 Y.t3 a_1162_48.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1332 ps=1.1 w=0.74 l=0.15
X20 a_27_368# B.t3 a_116_368.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.196 ps=1.47 w=1.12 l=0.15
X21 Y.t10 a_864_48.t6 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_27_368# a_864_48.t7 a_897_349.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.364 pd=2.89 as=0.3668 ps=1.775 w=1.12 l=0.15
X23 VPWR.t0 C_N.t1 a_864_48.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X24 a_864_48.t1 C_N.t2 VPWR.t3 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2898 ps=2.37 w=0.84 l=0.15
X25 VGND.t12 A.t7 Y.t11 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.13875 pd=1.115 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 Y.t2 a_1162_48.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.2516 ps=1.42 w=0.74 l=0.15
X27 Y.t4 a_1162_48.t7 a_897_349.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 VGND.t14 B.t4 Y.t13 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.111 ps=1.04 w=0.74 l=0.15
X29 VGND.t0 a_1162_48.t8 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.1258 ps=1.08 w=0.74 l=0.15
X30 a_27_368# a_864_48.t8 a_897_349.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.30235 pd=1.86 as=0.168 ps=1.42 w=1.12 l=0.15
X31 a_116_368.t1 B.t5 a_27_368# VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X32 a_897_349.t4 a_864_48.t9 a_27_368# VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X33 VGND.t15 B.t6 Y.t14 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X34 a_27_368# B.t7 a_116_368.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2071 ps=1.57 w=1.12 l=0.15
R0 a_1162_48.n11 a_1162_48.n10 399.289
R1 a_1162_48.n10 a_1162_48.n9 303.435
R2 a_1162_48.n3 a_1162_48.n2 295.091
R3 a_1162_48.n1 a_1162_48.t7 292.223
R4 a_1162_48.n7 a_1162_48.t3 234.841
R5 a_1162_48.n5 a_1162_48.n0 234.841
R6 a_1162_48.n3 a_1162_48.t5 185.571
R7 a_1162_48.n1 a_1162_48.t8 182.702
R8 a_1162_48.n8 a_1162_48.t6 159.499
R9 a_1162_48.n10 a_1162_48.t0 156.52
R10 a_1162_48.n4 a_1162_48.t4 155.847
R11 a_1162_48.n9 a_1162_48.n8 152
R12 a_1162_48.n4 a_1162_48.n3 100.928
R13 a_1162_48.n3 a_1162_48.n1 86.7605
R14 a_1162_48.n9 a_1162_48.n6 81.6328
R15 a_1162_48.n8 a_1162_48.n7 49.6611
R16 a_1162_48.n6 a_1162_48.n5 38.4293
R17 a_1162_48.n11 a_1162_48.t2 35.1791
R18 a_1162_48.t1 a_1162_48.n11 35.1791
R19 a_1162_48.n7 a_1162_48.n6 20.5774
R20 a_1162_48.n5 a_1162_48.n4 2.19141
R21 Y.n11 Y.t5 866.548
R22 Y.n11 Y.t4 857.518
R23 Y.n16 Y.n15 185
R24 Y.n17 Y.n16 185
R25 Y.n2 Y.n0 147.179
R26 Y.n6 Y.n5 101.507
R27 Y.n10 Y.n9 99.7158
R28 Y.n8 Y.n7 99.3719
R29 Y.n14 Y.n13 99.1033
R30 Y.n4 Y.n3 97.6664
R31 Y.n2 Y.n1 96.3134
R32 Y.n15 Y.n14 73.1271
R33 Y.n6 Y.n4 55.0405
R34 Y.n4 Y.n2 54.2123
R35 Y.n10 Y.n8 51.2005
R36 Y.n8 Y.n6 50.4476
R37 Y.n14 Y.n12 37.5563
R38 Y.n12 Y.n10 35.9007
R39 Y.n5 Y.t14 34.0546
R40 Y.n7 Y.t10 34.0546
R41 Y.n9 Y.t1 32.4329
R42 Y.n1 Y.t7 30.0005
R43 Y.n16 Y.t8 26.7573
R44 Y.n3 Y.t13 25.9464
R45 Y.n16 Y.t2 22.7032
R46 Y.n13 Y.t0 22.7032
R47 Y.n13 Y.t3 22.7032
R48 Y.n9 Y.t16 22.7032
R49 Y.n3 Y.t6 22.7032
R50 Y.n0 Y.t11 22.7032
R51 Y.n0 Y.t12 22.7032
R52 Y.n1 Y.t9 22.7032
R53 Y.n5 Y.t17 22.7032
R54 Y.n7 Y.t15 22.7032
R55 Y.n12 Y.n11 13.1884
R56 Y Y.n17 12.6066
R57 Y Y.n15 1.93989
R58 Y.n17 Y 1.74595
R59 a_897_349.n1 a_897_349.t0 811.551
R60 a_897_349.n2 a_897_349.n1 328.058
R61 a_897_349.n1 a_897_349.n0 273.421
R62 a_897_349.t1 a_897_349.n2 64.3092
R63 a_897_349.n2 a_897_349.t2 46.8546
R64 a_897_349.n0 a_897_349.t3 26.3844
R65 a_897_349.n0 a_897_349.t4 26.3844
R66 VPB.n0 VPB 4430.78
R67 VPB VPB.n1 1205.12
R68 VPB.t0 VPB.t1 660.87
R69 VPB.t8 VPB.t0 519.949
R70 VPB.t1 VPB.t4 391.176
R71 VPB.t4 VPB.n0 281.841
R72 VPB.n1 VPB.t5 268.146
R73 VPB.n0 VPB.t14 260.485
R74 VPB.t16 VPB 257.93
R75 VPB.t6 VPB.t10 255.376
R76 VPB.t10 VPB.t16 255.376
R77 VPB.t15 VPB.t13 245.397
R78 VPB.t12 VPB.t11 242.968
R79 VPB.t3 VPB.t7 229.839
R80 VPB.t2 VPB.t3 229.839
R81 VPB.t14 VPB.t2 229.839
R82 VPB.t5 VPB.t6 229.839
R83 VPB.t11 VPB.t9 223.53
R84 VPB.t9 VPB.t8 218.671
R85 VPB.t13 VPB.t12 218.671
R86 VPB.n1 VPB.t15 3.73576
R87 a_864_48.n11 a_864_48.n10 357.608
R88 a_864_48.n10 a_864_48.n7 322.728
R89 a_864_48.n9 a_864_48.t2 258.288
R90 a_864_48.n9 a_864_48.n8 242.662
R91 a_864_48.n8 a_864_48.t7 242.493
R92 a_864_48.n3 a_864_48.n2 239.224
R93 a_864_48.n4 a_864_48.t8 226.809
R94 a_864_48.n0 a_864_48.t9 226.809
R95 a_864_48.n0 a_864_48.t6 167.679
R96 a_864_48.n5 a_864_48.t5 165.488
R97 a_864_48.n3 a_864_48.t3 165.488
R98 a_864_48.n8 a_864_48.t4 154.24
R99 a_864_48.n7 a_864_48.n6 152
R100 a_864_48.n7 a_864_48.n1 81.6328
R101 a_864_48.n6 a_864_48.n5 43.0884
R102 a_864_48.n1 a_864_48.n0 36.9687
R103 a_864_48.t0 a_864_48.n11 35.1791
R104 a_864_48.n11 a_864_48.t1 35.1791
R105 a_864_48.n6 a_864_48.n3 29.9429
R106 a_864_48.n4 a_864_48.n1 22.038
R107 a_864_48.n10 a_864_48.n9 16.4853
R108 a_864_48.n5 a_864_48.n4 5.11262
R109 VGND.n32 VGND.n8 207.498
R110 VGND.n35 VGND.n34 207.498
R111 VGND.n39 VGND.n5 207.498
R112 VGND.n42 VGND.n41 206.333
R113 VGND.n46 VGND.n2 206.333
R114 VGND.n18 VGND.n17 185
R115 VGND.n16 VGND.n15 185
R116 VGND.n20 VGND.n10 185
R117 VGND.n22 VGND.n21 185
R118 VGND.n48 VGND.t13 154.727
R119 VGND.n14 VGND.t4 140.248
R120 VGND.n28 VGND.n27 116.644
R121 VGND.n16 VGND.t16 75.4059
R122 VGND.n21 VGND.n20 64.8654
R123 VGND.n17 VGND.n16 55.1356
R124 VGND.n26 VGND.n25 35.2632
R125 VGND.n33 VGND.n32 34.2593
R126 VGND.n27 VGND.t2 34.0546
R127 VGND.n8 VGND.t6 34.0546
R128 VGND.n41 VGND.t11 34.0546
R129 VGND.n2 VGND.t12 34.0546
R130 VGND.n40 VGND.n39 33.5064
R131 VGND.n42 VGND.n1 32.7534
R132 VGND.n28 VGND.n7 32.0005
R133 VGND.n35 VGND.n4 31.2476
R134 VGND.n5 VGND.t14 30.8113
R135 VGND.n22 VGND.n19 30.5783
R136 VGND.n47 VGND.n46 29.7417
R137 VGND.n41 VGND.t9 29.1897
R138 VGND.n2 VGND.t10 26.7573
R139 VGND.n27 VGND.t0 24.3248
R140 VGND.n19 VGND.n18 23.4672
R141 VGND.n21 VGND.t1 22.7032
R142 VGND.n20 VGND.t3 22.7032
R143 VGND.n17 VGND.t7 22.7032
R144 VGND.n8 VGND.t8 22.7032
R145 VGND.n34 VGND.t5 22.7032
R146 VGND.n34 VGND.t15 22.7032
R147 VGND.n5 VGND.t17 22.7032
R148 VGND.n48 VGND.n47 20.7064
R149 VGND.n15 VGND.n14 18.8018
R150 VGND.n46 VGND.n1 17.6946
R151 VGND.n35 VGND.n33 16.1887
R152 VGND.n28 VGND.n26 15.4358
R153 VGND.n42 VGND.n40 14.6829
R154 VGND.n39 VGND.n4 13.9299
R155 VGND.n32 VGND.n7 13.177
R156 VGND.n49 VGND.n48 9.3005
R157 VGND.n13 VGND.n12 9.3005
R158 VGND.n19 VGND.n11 9.3005
R159 VGND.n23 VGND.n22 9.3005
R160 VGND.n25 VGND.n24 9.3005
R161 VGND.n26 VGND.n9 9.3005
R162 VGND.n29 VGND.n28 9.3005
R163 VGND.n30 VGND.n7 9.3005
R164 VGND.n32 VGND.n31 9.3005
R165 VGND.n33 VGND.n6 9.3005
R166 VGND.n36 VGND.n35 9.3005
R167 VGND.n37 VGND.n4 9.3005
R168 VGND.n39 VGND.n38 9.3005
R169 VGND.n40 VGND.n3 9.3005
R170 VGND.n43 VGND.n42 9.3005
R171 VGND.n44 VGND.n1 9.3005
R172 VGND.n46 VGND.n45 9.3005
R173 VGND.n47 VGND.n0 9.3005
R174 VGND.n22 VGND.n10 6.69331
R175 VGND.n15 VGND.n12 4.43449
R176 VGND.n25 VGND.n10 1.33906
R177 VGND.n18 VGND.n12 1.2554
R178 VGND.n14 VGND.n13 0.207811
R179 VGND.n13 VGND.n11 0.122949
R180 VGND.n23 VGND.n11 0.122949
R181 VGND.n24 VGND.n23 0.122949
R182 VGND.n24 VGND.n9 0.122949
R183 VGND.n29 VGND.n9 0.122949
R184 VGND.n30 VGND.n29 0.122949
R185 VGND.n31 VGND.n30 0.122949
R186 VGND.n31 VGND.n6 0.122949
R187 VGND.n36 VGND.n6 0.122949
R188 VGND.n37 VGND.n36 0.122949
R189 VGND.n38 VGND.n37 0.122949
R190 VGND.n38 VGND.n3 0.122949
R191 VGND.n43 VGND.n3 0.122949
R192 VGND.n44 VGND.n43 0.122949
R193 VGND.n45 VGND.n44 0.122949
R194 VGND.n45 VGND.n0 0.122949
R195 VGND.n49 VGND.n0 0.122949
R196 VGND VGND.n49 0.0617245
R197 VNB.n0 VNB 20036.7
R198 VNB VNB.n1 6028.73
R199 VNB.t16 VNB.t4 3095.01
R200 VNB.t3 VNB.t1 2017.68
R201 VNB.t7 VNB.n0 1373.48
R202 VNB.t13 VNB 1304.99
R203 VNB.t0 VNB.t2 1239.78
R204 VNB.n0 VNB.t16 1224.15
R205 VNB.t6 VNB.t8 1215.47
R206 VNB.t5 VNB.t6 1215.47
R207 VNB.t17 VNB.t15 1215.47
R208 VNB.t10 VNB.t12 1212.6
R209 VNB.t8 VNB.t0 1191.16
R210 VNB.t14 VNB.t17 1166.85
R211 VNB.n1 VNB.t11 1120.21
R212 VNB.t1 VNB.t7 1106.08
R213 VNB.t11 VNB.t10 1097.11
R214 VNB.t9 VNB.t14 1093.92
R215 VNB.t2 VNB.t3 1045.3
R216 VNB.t15 VNB.t5 1045.3
R217 VNB.t12 VNB.t13 993.177
R218 VNB.n1 VNB.t9 65.1418
R219 B.n9 B.t0 258.942
R220 B.n1 B.t3 226.809
R221 B.n4 B.t5 226.809
R222 B.n6 B.t7 226.809
R223 B.n9 B.t2 207.845
R224 B B.n9 178.571
R225 B.n6 B.t4 167.679
R226 B.n1 B.t6 167.679
R227 B.n3 B.t1 165.488
R228 B.n2 B.n0 165.189
R229 B.n8 B.n7 152
R230 B.n5 B.n0 152
R231 B.n10 B.n8 140.143
R232 B.n7 B.n5 49.6611
R233 B.n3 B.n2 42.3581
R234 B.n2 B.n1 28.4823
R235 B.n8 B.n0 13.1884
R236 B.n7 B.n6 10.955
R237 B.n5 B.n4 5.11262
R238 B B.n10 3.89615
R239 B.n10 B 3.29747
R240 B.n4 B.n3 2.19141
R241 a_116_368.n2 a_116_368.n1 585
R242 a_116_368.n2 a_116_368.n0 380.464
R243 a_116_368.n5 a_116_368.n4 348.467
R244 a_116_368.n4 a_116_368.n3 296.788
R245 a_116_368.n4 a_116_368.n2 59.8141
R246 a_116_368.n1 a_116_368.t0 37.589
R247 a_116_368.n0 a_116_368.t1 35.1791
R248 a_116_368.t3 a_116_368.n5 35.1791
R249 a_116_368.n1 a_116_368.t7 27.1456
R250 a_116_368.n0 a_116_368.t2 26.3844
R251 a_116_368.n3 a_116_368.t4 26.3844
R252 a_116_368.n3 a_116_368.t5 26.3844
R253 a_116_368.n5 a_116_368.t6 26.3844
R254 A.n6 A.t6 262.771
R255 A.n1 A.t2 261.62
R256 A.n5 A.t0 261.62
R257 A.n7 A.t1 261.62
R258 A.n2 A 161.067
R259 A.n1 A.t4 160.083
R260 A.n6 A.t7 155.677
R261 A.n8 A.t5 154.24
R262 A.n3 A.t3 154.24
R263 A.n4 A.n0 152
R264 A.n10 A.n9 152
R265 A.n7 A.n6 73.0551
R266 A.n3 A.n2 48.9308
R267 A.n9 A.n5 44.549
R268 A.n2 A.n1 24.1005
R269 A.n9 A.n8 18.9884
R270 A.n10 A.n0 12.0894
R271 A.n5 A.n4 5.11262
R272 A A.n0 3.02272
R273 A.n8 A.n7 2.19141
R274 A A.n10 1.95606
R275 A.n4 A.n3 0.730803
R276 VPWR.n1 VPWR.n0 604.976
R277 VPWR.n39 VPWR.n3 602.817
R278 VPWR.n13 VPWR.t2 356.622
R279 VPWR.n10 VPWR.t3 352.279
R280 VPWR.n14 VPWR.n12 334.877
R281 VPWR.n14 VPWR.n13 39.5202
R282 VPWR.n3 VPWR.t7 38.6969
R283 VPWR.n21 VPWR.n20 36.1417
R284 VPWR.n22 VPWR.n21 36.1417
R285 VPWR.n22 VPWR.n8 36.1417
R286 VPWR.n26 VPWR.n8 36.1417
R287 VPWR.n27 VPWR.n26 36.1417
R288 VPWR.n28 VPWR.n27 36.1417
R289 VPWR.n28 VPWR.n6 36.1417
R290 VPWR.n32 VPWR.n6 36.1417
R291 VPWR.n33 VPWR.n32 36.1417
R292 VPWR.n34 VPWR.n33 36.1417
R293 VPWR.n34 VPWR.n4 36.1417
R294 VPWR.n38 VPWR.n4 36.1417
R295 VPWR.n16 VPWR.n15 36.1417
R296 VPWR.n0 VPWR.t4 35.1791
R297 VPWR.n12 VPWR.t1 35.1791
R298 VPWR.n12 VPWR.t0 35.1791
R299 VPWR.n3 VPWR.t5 29.9023
R300 VPWR.n20 VPWR.n10 29.3652
R301 VPWR.n40 VPWR.n39 28.9887
R302 VPWR.n0 VPWR.t6 26.3844
R303 VPWR.n16 VPWR.n10 18.0711
R304 VPWR.n40 VPWR.n1 17.6946
R305 VPWR.n39 VPWR.n38 15.4358
R306 VPWR.n15 VPWR.n11 9.3005
R307 VPWR.n17 VPWR.n16 9.3005
R308 VPWR.n18 VPWR.n10 9.3005
R309 VPWR.n20 VPWR.n19 9.3005
R310 VPWR.n21 VPWR.n9 9.3005
R311 VPWR.n23 VPWR.n22 9.3005
R312 VPWR.n24 VPWR.n8 9.3005
R313 VPWR.n26 VPWR.n25 9.3005
R314 VPWR.n27 VPWR.n7 9.3005
R315 VPWR.n29 VPWR.n28 9.3005
R316 VPWR.n30 VPWR.n6 9.3005
R317 VPWR.n32 VPWR.n31 9.3005
R318 VPWR.n33 VPWR.n5 9.3005
R319 VPWR.n35 VPWR.n34 9.3005
R320 VPWR.n36 VPWR.n4 9.3005
R321 VPWR.n38 VPWR.n37 9.3005
R322 VPWR.n39 VPWR.n2 9.3005
R323 VPWR.n41 VPWR.n40 9.3005
R324 VPWR.n42 VPWR.n1 7.42789
R325 VPWR.n13 VPWR.n11 2.34593
R326 VPWR.n15 VPWR.n14 1.50638
R327 VPWR VPWR.n42 0.278906
R328 VPWR.n42 VPWR.n41 0.151952
R329 VPWR.n17 VPWR.n11 0.122949
R330 VPWR.n18 VPWR.n17 0.122949
R331 VPWR.n19 VPWR.n18 0.122949
R332 VPWR.n19 VPWR.n9 0.122949
R333 VPWR.n23 VPWR.n9 0.122949
R334 VPWR.n24 VPWR.n23 0.122949
R335 VPWR.n25 VPWR.n24 0.122949
R336 VPWR.n25 VPWR.n7 0.122949
R337 VPWR.n29 VPWR.n7 0.122949
R338 VPWR.n30 VPWR.n29 0.122949
R339 VPWR.n31 VPWR.n30 0.122949
R340 VPWR.n31 VPWR.n5 0.122949
R341 VPWR.n35 VPWR.n5 0.122949
R342 VPWR.n36 VPWR.n35 0.122949
R343 VPWR.n37 VPWR.n36 0.122949
R344 VPWR.n37 VPWR.n2 0.122949
R345 VPWR.n41 VPWR.n2 0.122949
R346 D_N.n1 D_N.t2 259.964
R347 D_N.n0 D_N.t0 231.377
R348 D_N.n0 D_N.t1 230.298
R349 D_N D_N.n1 154.133
R350 D_N.n1 D_N.n0 35.0943
R351 C_N.n1 C_N.t0 277.954
R352 C_N.n0 C_N.t1 267.243
R353 C_N.n0 C_N.t2 219.554
R354 C_N C_N.n1 152.583
R355 C_N.n1 C_N.n0 13.146
C0 a_27_368# A 0.032926f
C1 a_27_368# VPWR 0.601294f
C2 VPB D_N 0.097459f
C3 D_N VGND 0.023105f
C4 VPB Y 0.011086f
C5 C_N D_N 0.070981f
C6 Y VGND 1.19923f
C7 B Y 0.2124f
C8 VPB VGND 0.01616f
C9 C_N Y 5.36e-19
C10 VPB B 0.15588f
C11 VPB C_N 0.112952f
C12 VPWR D_N 0.036868f
C13 C_N VGND 0.009808f
C14 A Y 0.153054f
C15 B VGND 0.094512f
C16 VPB A 0.14397f
C17 B C_N 1.85e-20
C18 VPWR Y 0.019703f
C19 A VGND 0.063378f
C20 B A 0.289027f
C21 VPB VPWR 0.267049f
C22 A C_N 4.65e-19
C23 VPWR VGND 0.176779f
C24 B VPWR 0.040597f
C25 VPWR C_N 0.052008f
C26 A VPWR 0.053773f
C27 a_27_368# Y 0.016786f
C28 a_27_368# VPB 0.061062f
C29 a_27_368# VGND 0.017295f
C30 a_27_368# B 0.365694f
C31 a_27_368# C_N 0.001733f
C32 VGND VNB 1.28218f
C33 Y VNB 0.055447f
C34 D_N VNB 0.198595f
C35 C_N VNB 0.162286f
C36 VPWR VNB 1.00886f
C37 A VNB 0.424137f
C38 B VNB 0.450196f
C39 VPB VNB 2.61957f
C40 a_27_368# VNB 0.051363f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4bb_2 VNB VPB VPWR VGND C_N D_N A B Y
X0 a_985_368.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t3 C_N.t0 a_27_392.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.585 pd=2.17 as=0.295 ps=2.59 w=1 l=0.15
X2 VGND.t3 C_N.t1 a_27_392.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.180725 pd=1.42 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 Y.t3 A.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.30155 ps=1.555 w=0.74 l=0.15
X4 VPWR.t0 A.t2 a_985_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5 a_493_368.t3 a_311_124.t2 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t5 a_311_124.t3 a_493_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 Y.t7 a_311_124.t4 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.4735 ps=2.86 w=0.74 l=0.15
X8 Y.t6 B.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 VGND.t9 B.t1 Y.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.30155 pd=1.555 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_985_368.t3 B.t2 a_772_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VGND.t8 a_311_124.t5 Y.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2096 pd=1.405 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_772_368.t2 B.t3 a_985_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X13 VGND.t5 A.t3 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.12025 ps=1.065 w=0.74 l=0.15
X14 a_311_124.t1 D_N.t0 VPWR.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.585 ps=2.17 w=1 l=0.15
X15 VGND.t2 a_27_392.t2 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_493_368.t0 a_27_392.t3 a_772_368.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X17 a_311_124.t0 D_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2496 pd=2.06 as=0.180725 ps=1.42 w=0.64 l=0.15
X18 Y.t0 a_27_392.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2096 ps=1.405 w=0.74 l=0.15
X19 a_772_368.t0 a_27_392.t5 a_493_368.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
R0 A.n3 A.t0 226.809
R1 A.n1 A.t2 226.809
R2 A.n1 A.t1 198.204
R3 A.n4 A.t3 196.013
R4 A.n5 A.n4 168.067
R5 A.n2 A.n0 152
R6 A.n2 A.n1 33.5944
R7 A.n3 A.n2 32.1338
R8 A.n5 A.n0 10.1214
R9 A.n0 A 2.3819
R10 A A.n5 1.78655
R11 A.n4 A.n3 1.46111
R12 VPWR.n5 VPWR.n2 585
R13 VPWR.n10 VPWR.n0 339.889
R14 VPWR.n3 VPWR.n1 291.515
R15 VPWR.n7 VPWR.n6 291.515
R16 VPWR.n6 VPWR.n4 274.512
R17 VPWR.n9 VPWR.n8 272.539
R18 VPWR.n4 VPWR.n2 39.9244
R19 VPWR.n8 VPWR.n7 39.9244
R20 VPWR.n4 VPWR.n3 39.9244
R21 VPWR.n8 VPWR.n2 39.9244
R22 VPWR.n3 VPWR.t2 29.5505
R23 VPWR.n7 VPWR.t3 29.5505
R24 VPWR.n0 VPWR.t1 26.3844
R25 VPWR.n0 VPWR.t0 26.3844
R26 VPWR.n10 VPWR.n9 8.59944
R27 VPWR.n5 VPWR.n1 1.97252
R28 VPWR.n6 VPWR.n5 1.97252
R29 VPWR.n9 VPWR.n1 1.97252
R30 VPWR VPWR.n10 0.30541
R31 a_985_368.n1 a_985_368.t2 447.334
R32 a_985_368.t1 a_985_368.n1 272.572
R33 a_985_368.n1 a_985_368.n0 203.27
R34 a_985_368.n0 a_985_368.t3 35.1791
R35 a_985_368.n0 a_985_368.t0 26.3844
R36 VPB.t8 VPB.t7 674.194
R37 VPB.t9 VPB.t4 515.861
R38 VPB.t7 VPB.t3 515.861
R39 VPB VPB.t8 257.93
R40 VPB.t5 VPB.t0 255.376
R41 VPB.t6 VPB.t9 255.376
R42 VPB.t2 VPB.t6 255.376
R43 VPB.t0 VPB.t1 229.839
R44 VPB.t4 VPB.t5 229.839
R45 VPB.t3 VPB.t2 229.839
R46 C_N.n2 C_N.t1 250.641
R47 C_N.n1 C_N.t0 234.549
R48 C_N.n3 C_N.n2 176.101
R49 C_N.n1 C_N.n0 152
R50 C_N.n2 C_N.n1 25.5611
R51 C_N.n3 C_N.n0 13.1884
R52 C_N C_N.n3 3.29747
R53 C_N.n0 C_N 2.13383
R54 a_27_392.n3 a_27_392.n2 400.31
R55 a_27_392.t0 a_27_392.n3 324.945
R56 a_27_392.n0 a_27_392.t3 226.809
R57 a_27_392.n2 a_27_392.t5 226.809
R58 a_27_392.n0 a_27_392.t2 204.411
R59 a_27_392.n1 a_27_392.t4 196.013
R60 a_27_392.n3 a_27_392.t1 130.214
R61 a_27_392.n1 a_27_392.n0 55.5035
R62 a_27_392.n2 a_27_392.n1 17.5278
R63 VGND.n3 VGND.t7 264.637
R64 VGND.n18 VGND.n17 211.183
R65 VGND.n1 VGND.n0 204.201
R66 VGND.n24 VGND.n23 197.537
R67 VGND.n15 VGND.n14 185
R68 VGND.n13 VGND.n12 185
R69 VGND.n8 VGND.t5 169.025
R70 VGND.n14 VGND.n13 86.7573
R71 VGND.n0 VGND.t0 70.8659
R72 VGND.n23 VGND.t1 39.7302
R73 VGND.n23 VGND.t8 38.9194
R74 VGND.n30 VGND.n29 36.1417
R75 VGND.n17 VGND.t2 34.0546
R76 VGND.n0 VGND.t3 33.7505
R77 VGND.n26 VGND.n25 32.3047
R78 VGND.n33 VGND.n1 31.5148
R79 VGND.n12 VGND.n8 31.2928
R80 VGND.n18 VGND.n5 28.2358
R81 VGND.n16 VGND.n15 27.2916
R82 VGND.n22 VGND.n5 26.7943
R83 VGND.n25 VGND.n24 25.1307
R84 VGND.n13 VGND.t4 22.7032
R85 VGND.n14 VGND.t9 22.7032
R86 VGND.n17 VGND.t6 22.7032
R87 VGND.n18 VGND.n16 19.2005
R88 VGND.n31 VGND.n30 18.8752
R89 VGND.n32 VGND.n31 9.3005
R90 VGND.n30 VGND.n2 9.3005
R91 VGND.n29 VGND.n28 9.3005
R92 VGND.n27 VGND.n26 9.3005
R93 VGND.n25 VGND.n4 9.3005
R94 VGND.n22 VGND.n21 9.3005
R95 VGND.n20 VGND.n5 9.3005
R96 VGND.n19 VGND.n18 9.3005
R97 VGND.n16 VGND.n6 9.3005
R98 VGND.n9 VGND.n7 9.3005
R99 VGND.n11 VGND.n10 9.3005
R100 VGND.n29 VGND.n3 7.85819
R101 VGND.n11 VGND.n7 6.64266
R102 VGND.n26 VGND.n3 3.8917
R103 VGND.n10 VGND.n8 2.34593
R104 VGND.n31 VGND.n1 0.8197
R105 VGND.n15 VGND.n7 0.554013
R106 VGND.n24 VGND.n22 0.328705
R107 VGND.n12 VGND.n11 0.208068
R108 VGND VGND.n33 0.163644
R109 VGND.n33 VGND.n32 0.144205
R110 VGND.n10 VGND.n9 0.122949
R111 VGND.n9 VGND.n6 0.122949
R112 VGND.n19 VGND.n6 0.122949
R113 VGND.n20 VGND.n19 0.122949
R114 VGND.n21 VGND.n20 0.122949
R115 VGND.n21 VGND.n4 0.122949
R116 VGND.n27 VGND.n4 0.122949
R117 VGND.n28 VGND.n27 0.122949
R118 VGND.n28 VGND.n2 0.122949
R119 VGND.n32 VGND.n2 0.122949
R120 VNB.t0 VNB.t7 3141.21
R121 VNB.t9 VNB.t5 2228.87
R122 VNB VNB.t3 1997.9
R123 VNB.t8 VNB.t1 1466.67
R124 VNB.t3 VNB.t0 1420.47
R125 VNB.t2 VNB.t6 1154.86
R126 VNB.t5 VNB.t4 1097.11
R127 VNB.t6 VNB.t9 993.177
R128 VNB.t1 VNB.t2 993.177
R129 VNB.t7 VNB.t8 993.177
R130 Y.n8 Y.n0 382.216
R131 Y.n6 Y.n5 248.738
R132 Y.n3 Y.n1 188.156
R133 Y.n3 Y.n2 104.579
R134 Y.n6 Y.n4 92.7788
R135 Y.n7 Y.n3 51.2005
R136 Y.n8 Y.n7 31.1563
R137 Y.n1 Y.t3 30.0005
R138 Y.n0 Y.t4 26.3844
R139 Y.n0 Y.t5 26.3844
R140 Y.n4 Y.t1 22.7032
R141 Y.n4 Y.t0 22.7032
R142 Y.n5 Y.t8 22.7032
R143 Y.n5 Y.t7 22.7032
R144 Y.n1 Y.t2 22.7032
R145 Y.n2 Y.t9 22.7032
R146 Y.n2 Y.t6 22.7032
R147 Y Y.n8 15.3048
R148 Y.n7 Y.n6 8.93268
R149 a_311_124.t1 a_311_124.n3 267.786
R150 a_311_124.n3 a_311_124.t0 255.868
R151 a_311_124.n2 a_311_124.t2 228.47
R152 a_311_124.n0 a_311_124.t3 226.809
R153 a_311_124.n2 a_311_124.t5 196.013
R154 a_311_124.n0 a_311_124.t4 196.013
R155 a_311_124.n1 a_311_124.n0 8.65511
R156 a_311_124.n1 a_311_124.n2 52.9719
R157 a_311_124.n3 a_311_124.n1 71.634
R158 a_493_368.n1 a_493_368.t0 380.717
R159 a_493_368.t2 a_493_368.n1 301.808
R160 a_493_368.n1 a_493_368.n0 288.108
R161 a_493_368.n0 a_493_368.t3 35.1791
R162 a_493_368.n0 a_493_368.t1 26.3844
R163 B.n3 B.t2 242.023
R164 B.n2 B.t3 226.809
R165 B.n0 B.t0 223.766
R166 B.n1 B.t1 196.013
R167 B.n0 B 169.96
R168 B.n4 B.n3 152
R169 B.n3 B.n2 50.3914
R170 B.n1 B.n0 35.055
R171 B B.n4 8.18655
R172 B.n4 B 6.10283
R173 B.n2 B.n1 4.38232
R174 a_772_368.n1 a_772_368.n0 990.072
R175 a_772_368.n1 a_772_368.t0 35.1791
R176 a_772_368.n0 a_772_368.t3 26.3844
R177 a_772_368.n0 a_772_368.t2 26.3844
R178 a_772_368.t1 a_772_368.n1 26.3844
R179 D_N.n0 D_N.t0 231.629
R180 D_N.n0 D_N.t1 196.599
R181 D_N D_N.n0 154.522
C0 A VGND 0.069519f
C1 B VPWR 0.018564f
C2 VPWR Y 0.015298f
C3 A VPWR 0.032098f
C4 VPWR VGND 0.118854f
C5 VPB C_N 0.080866f
C6 VPB D_N 0.066307f
C7 VPB B 0.090252f
C8 C_N D_N 0.069968f
C9 VPB Y 0.014165f
C10 VPB A 0.075451f
C11 C_N Y 2.15e-19
C12 VPB VGND 0.013645f
C13 D_N Y 0.00107f
C14 C_N VGND 0.017435f
C15 VPB VPWR 0.180291f
C16 B Y 0.162782f
C17 D_N VGND 0.017668f
C18 B A 0.075885f
C19 C_N VPWR 0.092611f
C20 B VGND 0.039556f
C21 A Y 0.050465f
C22 Y VGND 0.597022f
C23 D_N VPWR 0.050121f
C24 VGND VNB 0.879403f
C25 Y VNB 0.04476f
C26 VPWR VNB 0.66195f
C27 A VNB 0.266285f
C28 B VNB 0.245342f
C29 D_N VNB 0.147287f
C30 C_N VNB 0.194187f
C31 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4bb_1 VNB VPB VPWR VGND D_N C_N B A Y
X0 VPWR.t2 C_N.t0 a_27_112.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.510675 pd=2.125 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VGND.t1 C_N.t1 a_27_112.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1671 pd=1.225 as=0.3025 ps=2.2 w=0.55 l=0.15
X2 a_530_368.t1 a_27_112.t2 a_397_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2884 ps=1.635 w=1.12 l=0.15
X3 Y.t2 A.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1671 ps=1.225 w=0.74 l=0.15
X4 Y.t1 a_611_244.t2 a_530_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X5 a_397_368.t0 B.t0 a_313_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2884 pd=1.635 as=0.1512 ps=1.39 w=1.12 l=0.15
X6 a_611_244.t1 D_N.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.231 ps=2.23 w=0.84 l=0.15
X7 a_313_368.t1 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.510675 ps=2.125 w=1.12 l=0.15
X8 a_611_244.t0 D_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.331425 ps=1.655 w=0.55 l=0.15
X9 VGND.t3 a_611_244.t3 Y.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.331425 pd=1.655 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 VGND.t4 B.t1 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.25715 pd=1.435 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 Y.t4 a_27_112.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.25715 ps=1.435 w=0.74 l=0.15
R0 C_N.n0 C_N.t0 226.387
R1 C_N C_N.n0 179.968
R2 C_N.n0 C_N.t1 142.649
R3 a_27_112.t0 a_27_112.n1 768.644
R4 a_27_112.t0 a_27_112.n2 768.644
R5 a_27_112.n1 a_27_112.n0 504.205
R6 a_27_112.n2 a_27_112.t1 282.935
R7 a_27_112.n0 a_27_112.t2 250.909
R8 a_27_112.n0 a_27_112.t3 220.113
R9 a_27_112.n2 a_27_112.n1 10.6672
R10 VPWR.n1 VPWR.t1 435.699
R11 VPWR.n1 VPWR.n0 434.277
R12 VPWR.n0 VPWR.t2 107.882
R13 VPWR.n0 VPWR.t0 65.9603
R14 VPWR VPWR.n1 0.256809
R15 VPB.t4 VPB.t1 587.366
R16 VPB.t2 VPB.t0 503.091
R17 VPB.t3 VPB.t5 339.651
R18 VPB.t5 VPB.t4 291.13
R19 VPB VPB.t2 257.93
R20 VPB.t0 VPB.t3 214.517
R21 VGND.n5 VGND.n3 185
R22 VGND.n4 VGND.n3 185
R23 VGND.n12 VGND.n11 185
R24 VGND.n10 VGND.n9 185
R25 VGND.n15 VGND.n14 119.966
R26 VGND.n7 VGND.n6 77.5469
R27 VGND.n11 VGND.n10 67.2978
R28 VGND.n14 VGND.t1 63.21
R29 VGND.n5 VGND.t3 41.3519
R30 VGND.n4 VGND.t0 39.8776
R31 VGND.n14 VGND.t2 32.4229
R32 VGND.n15 VGND.n13 30.4946
R33 VGND.n6 VGND.n5 29.9091
R34 VGND.n6 VGND.n4 29.9091
R35 VGND.n13 VGND.n12 22.7142
R36 VGND.n10 VGND.t5 22.7032
R37 VGND.n11 VGND.t4 22.7032
R38 VGND.n8 VGND.n7 11.8626
R39 VGND.n2 VGND.n1 9.3005
R40 VGND.n13 VGND.n0 9.3005
R41 VGND.n9 VGND.n8 9.23889
R42 VGND.n16 VGND.n15 6.72455
R43 VGND.n9 VGND.n1 6.10769
R44 VGND.n7 VGND.n3 5.65245
R45 VGND.n12 VGND.n1 0.837101
R46 VGND.n8 VGND.n2 0.361413
R47 VGND VGND.n16 0.268037
R48 VGND.n16 VGND.n0 0.162655
R49 VGND.n2 VGND.n0 0.122949
R50 VNB.t3 VNB.t0 2459.84
R51 VNB.t4 VNB.t5 1951.71
R52 VNB VNB.t1 1755.38
R53 VNB.t1 VNB.t2 1466.67
R54 VNB.t5 VNB.t3 1154.86
R55 VNB.t2 VNB.t4 1154.86
R56 a_397_368.t0 a_397_368.t1 90.5853
R57 a_530_368.t0 a_530_368.t1 73.8755
R58 A.n0 A.t1 242.556
R59 A.n0 A.t0 211.762
R60 A A.n0 154.522
R61 Y.n1 Y.t1 844.615
R62 Y.n1 Y.n0 96.6686
R63 Y.n3 Y.n1 90.532
R64 Y.n3 Y.n2 89.4479
R65 Y.n2 Y.t4 34.0546
R66 Y.n0 Y.t3 34.0546
R67 Y.n2 Y.t0 22.7032
R68 Y.n0 Y.t2 22.7032
R69 Y Y.n3 7.64324
R70 a_611_244.n0 a_611_244.t2 205.534
R71 a_611_244.t1 a_611_244.n1 462.527
R72 a_611_244.n0 a_611_244.t3 159.448
R73 a_611_244.n1 a_611_244.t0 228.733
R74 a_611_244.n1 a_611_244.n0 147.236
R75 B.n0 B.t0 245.522
R76 B.n0 B.t1 214.726
R77 B B.n0 154.311
R78 a_313_368.t0 a_313_368.t1 47.4916
R79 D_N.n0 D_N.t0 251.81
R80 D_N.n0 D_N.t1 219.41
R81 D_N D_N.n0 159.177
C0 VGND A 0.0409f
C1 B VPB 0.038694f
C2 B Y 0.11705f
C3 C_N VPB 0.058317f
C4 B VPWR 0.009528f
C5 C_N Y 7.66e-19
C6 Y VPB 0.004552f
C7 B A 0.056729f
C8 C_N VPWR 0.00468f
C9 B VGND 0.018322f
C10 C_N D_N 6.13e-19
C11 VPB VPWR 0.134131f
C12 C_N A 0.032123f
C13 Y VPWR 0.025044f
C14 D_N VPB 0.064446f
C15 C_N VGND 0.012812f
C16 Y D_N 5.19e-19
C17 VPB A 0.047161f
C18 D_N VPWR 0.037291f
C19 VGND VPB 0.010901f
C20 Y A 0.094441f
C21 Y VGND 0.340804f
C22 VPWR A 0.027409f
C23 VGND VPWR 0.081924f
C24 D_N VGND 0.014815f
C25 VGND VNB 0.610253f
C26 D_N VNB 0.15184f
C27 Y VNB 0.025982f
C28 C_N VNB 0.198598f
C29 B VNB 0.118051f
C30 A VNB 0.128315f
C31 VPWR VNB 0.472517f
C32 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4b_4 VNB VPB VPWR VGND D_N C B A Y
X0 a_319_368.t4 a_47_88.t3 Y.t11 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t10 a_47_88.t4 a_319_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_1191_368.t3 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VGND.t10 a_47_88.t5 Y.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1332 ps=1.1 w=0.74 l=0.15
X4 Y.t1 A.t1 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.16465 ps=1.185 w=0.74 l=0.15
X5 VPWR.t3 A.t2 a_1191_368.t2 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t0 C.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.30525 ps=1.565 w=0.74 l=0.15
X7 a_1191_368.t1 A.t3 VPWR.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_319_368.t6 C.t1 a_778_368.t3 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.182 ps=1.445 w=1.12 l=0.15
X9 VGND.t5 A.t4 Y.t12 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VPWR.t4 D_N.t0 a_47_88.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X11 VPWR.t0 A.t5 a_1191_368.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_778_368.t2 C.t2 a_319_368.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.182 pd=1.445 as=0.21 ps=1.495 w=1.12 l=0.15
X13 a_1191_368.t4 B.t0 a_778_368.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X15 a_778_368.t5 B.t1 a_1191_368.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X16 Y.t2 C.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X17 VGND.t4 A.t6 Y.t14 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_319_368.t2 a_47_88.t6 Y.t9 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t7 a_47_88.t7 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.10915 ps=1.035 w=0.74 l=0.15
X20 Y.t8 a_47_88.t8 a_319_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X21 VGND.t8 a_47_88.t9 Y.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X23 a_1191_368.t6 B.t2 a_778_368.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X24 a_47_88.t1 D_N.t1 VPWR.t5 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2478 ps=2.27 w=0.84 l=0.15
X25 a_319_368.t0 C.t4 a_778_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.495 as=0.196 ps=1.47 w=1.12 l=0.15
X26 VGND.t2 C.t5 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.28305 pd=1.505 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.28305 ps=1.505 w=0.74 l=0.15
X28 VGND.t12 D_N.t2 a_47_88.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.31115 ps=2.85 w=0.74 l=0.15
X29 Y.t5 a_47_88.t10 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X30 a_778_368.t7 B.t3 a_1191_368.t7 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X31 VGND.t11 B.t4 Y.t13 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.16465 pd=1.185 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 Y.t15 A.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 a_778_368.t0 C.t6 a_319_368.t7 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X34 VGND.t13 C.t7 Y.t16 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.30525 pd=1.565 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_47_88.n11 a_47_88.n10 338.022
R1 a_47_88.n2 a_47_88.t3 328.228
R2 a_47_88.n5 a_47_88.t6 214.758
R3 a_47_88.n0 a_47_88.t8 214.758
R4 a_47_88.n2 a_47_88.t4 210.254
R5 a_47_88.n8 a_47_88.t7 191.73
R6 a_47_88.n10 a_47_88.t2 189.141
R7 a_47_88.n0 a_47_88.t5 186.374
R8 a_47_88.n4 a_47_88.t10 186.374
R9 a_47_88.n3 a_47_88.t9 186.374
R10 a_47_88.n6 a_47_88.n1 165.189
R11 a_47_88.n9 a_47_88.n8 152
R12 a_47_88.n7 a_47_88.n1 152
R13 a_47_88.n4 a_47_88.n3 51.1758
R14 a_47_88.n8 a_47_88.n7 40.4647
R15 a_47_88.t0 a_47_88.n11 35.1791
R16 a_47_88.n11 a_47_88.t1 35.1791
R17 a_47_88.n6 a_47_88.n5 29.7536
R18 a_47_88.n10 a_47_88.n9 26.3763
R19 a_47_88.n0 a_47_88.n6 23.803
R20 a_47_88.n7 a_47_88.n0 16.6622
R21 a_47_88.n9 a_47_88.n1 13.1884
R22 a_47_88.n5 a_47_88.n4 4.16593
R23 a_47_88.n3 a_47_88.n2 1.8847
R24 Y.n2 Y.n0 255.553
R25 Y.n2 Y.n1 200.526
R26 Y Y.n2 184.304
R27 Y.n12 Y.n10 156.532
R28 Y.n5 Y.n3 154.244
R29 Y.n13 Y.t13 149.99
R30 Y.n12 Y.n11 104.579
R31 Y.n7 Y.n6 104.579
R32 Y.n9 Y.n8 101.71
R33 Y.n5 Y.n4 100.547
R34 Y.n14 Y.n13 96.7534
R35 Y.n9 Y.n7 86.9652
R36 Y.n7 Y.n5 77.7077
R37 Y.n13 Y.n12 52.3299
R38 Y.n3 Y.t7 35.6762
R39 Y.n1 Y.t11 26.3844
R40 Y.n1 Y.t10 26.3844
R41 Y.n0 Y.t9 26.3844
R42 Y.n0 Y.t8 26.3844
R43 Y.n10 Y.t12 22.7032
R44 Y.n10 Y.t15 22.7032
R45 Y.n11 Y.t14 22.7032
R46 Y.n11 Y.t1 22.7032
R47 Y.n6 Y.t16 22.7032
R48 Y.n6 Y.t2 22.7032
R49 Y.n4 Y.t6 22.7032
R50 Y.n4 Y.t5 22.7032
R51 Y.n3 Y.t4 22.7032
R52 Y.n8 Y.t3 22.7032
R53 Y.n8 Y.t0 22.7032
R54 Y.n14 Y.n9 12.8005
R55 Y Y.n14 6.4005
R56 a_319_368.n1 a_319_368.t6 672.992
R57 a_319_368.n1 a_319_368.n0 585
R58 a_319_368.n3 a_319_368.n2 305.301
R59 a_319_368.n3 a_319_368.t1 294.469
R60 a_319_368.n5 a_319_368.n4 288.555
R61 a_319_368.n4 a_319_368.n1 66.9089
R62 a_319_368.n4 a_319_368.n3 65.4258
R63 a_319_368.n0 a_319_368.t0 35.1791
R64 a_319_368.n2 a_319_368.t3 31.6612
R65 a_319_368.n0 a_319_368.t5 30.7817
R66 a_319_368.n2 a_319_368.t2 29.9023
R67 a_319_368.n5 a_319_368.t7 26.3844
R68 a_319_368.t4 a_319_368.n5 26.3844
R69 VPB.t15 VPB.t12 515.861
R70 VPB.t2 VPB.t3 515.861
R71 VPB.t1 VPB.t7 268.146
R72 VPB VPB.t16 257.93
R73 VPB.t10 VPB.t9 255.376
R74 VPB.t12 VPB.t10 255.376
R75 VPB.t17 VPB.t1 255.376
R76 VPB.t4 VPB.t5 255.376
R77 VPB.t7 VPB.t15 242.608
R78 VPB.t14 VPB.t0 229.839
R79 VPB.t11 VPB.t14 229.839
R80 VPB.t13 VPB.t11 229.839
R81 VPB.t8 VPB.t13 229.839
R82 VPB.t9 VPB.t8 229.839
R83 VPB.t6 VPB.t17 229.839
R84 VPB.t5 VPB.t6 229.839
R85 VPB.t3 VPB.t4 229.839
R86 VPB.t16 VPB.t2 229.839
R87 A.n2 A.t0 235.571
R88 A.n9 A.t5 228.549
R89 A.n3 A.t2 226.809
R90 A.n7 A.t3 226.809
R91 A.n9 A.t1 196.725
R92 A.n8 A.t6 196.013
R93 A.n1 A.t7 196.013
R94 A.n2 A.t4 196.013
R95 A A.n4 153.786
R96 A.n6 A.n5 152
R97 A.n8 A.n0 152
R98 A A.n10 152
R99 A.n10 A.n8 49.6611
R100 A.n7 A.n6 46.7399
R101 A.n4 A.n3 30.6732
R102 A.n4 A.n2 26.2914
R103 A.n6 A.n1 13.146
R104 A.n10 A.n9 12.4355
R105 A A.n0 10.1214
R106 A.n5 A 8.33538
R107 A.n5 A 5.95399
R108 A.n3 A.n1 5.84292
R109 A A.n0 4.16794
R110 A.n8 A.n7 2.92171
R111 VPWR.n36 VPWR.t5 417.604
R112 VPWR.n34 VPWR.t4 411.692
R113 VPWR.n12 VPWR.n9 329.329
R114 VPWR.n11 VPWR.n10 323.406
R115 VPWR.n15 VPWR.n8 36.1417
R116 VPWR.n16 VPWR.n15 36.1417
R117 VPWR.n17 VPWR.n16 36.1417
R118 VPWR.n17 VPWR.n6 36.1417
R119 VPWR.n21 VPWR.n6 36.1417
R120 VPWR.n22 VPWR.n21 36.1417
R121 VPWR.n23 VPWR.n22 36.1417
R122 VPWR.n23 VPWR.n4 36.1417
R123 VPWR.n27 VPWR.n4 36.1417
R124 VPWR.n28 VPWR.n27 36.1417
R125 VPWR.n29 VPWR.n28 36.1417
R126 VPWR.n29 VPWR.n2 36.1417
R127 VPWR.n33 VPWR.n2 36.1417
R128 VPWR.n11 VPWR.n8 27.4829
R129 VPWR.n35 VPWR.n34 26.7299
R130 VPWR.n36 VPWR.n35 26.7299
R131 VPWR.n10 VPWR.t2 26.3844
R132 VPWR.n10 VPWR.t0 26.3844
R133 VPWR.n9 VPWR.t1 26.3844
R134 VPWR.n9 VPWR.t3 26.3844
R135 VPWR.n34 VPWR.n33 25.224
R136 VPWR.n13 VPWR.n8 9.3005
R137 VPWR.n15 VPWR.n14 9.3005
R138 VPWR.n16 VPWR.n7 9.3005
R139 VPWR.n18 VPWR.n17 9.3005
R140 VPWR.n19 VPWR.n6 9.3005
R141 VPWR.n21 VPWR.n20 9.3005
R142 VPWR.n22 VPWR.n5 9.3005
R143 VPWR.n24 VPWR.n23 9.3005
R144 VPWR.n25 VPWR.n4 9.3005
R145 VPWR.n27 VPWR.n26 9.3005
R146 VPWR.n28 VPWR.n3 9.3005
R147 VPWR.n30 VPWR.n29 9.3005
R148 VPWR.n31 VPWR.n2 9.3005
R149 VPWR.n33 VPWR.n32 9.3005
R150 VPWR.n34 VPWR.n1 9.3005
R151 VPWR.n35 VPWR.n0 9.3005
R152 VPWR.n37 VPWR.n36 9.3005
R153 VPWR.n12 VPWR.n11 6.92587
R154 VPWR.n13 VPWR.n12 0.478146
R155 VPWR.n14 VPWR.n13 0.122949
R156 VPWR.n14 VPWR.n7 0.122949
R157 VPWR.n18 VPWR.n7 0.122949
R158 VPWR.n19 VPWR.n18 0.122949
R159 VPWR.n20 VPWR.n19 0.122949
R160 VPWR.n20 VPWR.n5 0.122949
R161 VPWR.n24 VPWR.n5 0.122949
R162 VPWR.n25 VPWR.n24 0.122949
R163 VPWR.n26 VPWR.n25 0.122949
R164 VPWR.n26 VPWR.n3 0.122949
R165 VPWR.n30 VPWR.n3 0.122949
R166 VPWR.n31 VPWR.n30 0.122949
R167 VPWR.n32 VPWR.n31 0.122949
R168 VPWR.n32 VPWR.n1 0.122949
R169 VPWR.n1 VPWR.n0 0.122949
R170 VPWR.n37 VPWR.n0 0.122949
R171 VPWR VPWR.n37 0.0617245
R172 a_1191_368.n1 a_1191_368.t7 435.517
R173 a_1191_368.n1 a_1191_368.n0 297.598
R174 a_1191_368.t3 a_1191_368.n5 280.983
R175 a_1191_368.n3 a_1191_368.n2 206.922
R176 a_1191_368.n5 a_1191_368.n4 203.394
R177 a_1191_368.n3 a_1191_368.n1 46.6829
R178 a_1191_368.n5 a_1191_368.n3 46.6829
R179 a_1191_368.n0 a_1191_368.t6 35.1791
R180 a_1191_368.n0 a_1191_368.t5 26.3844
R181 a_1191_368.n2 a_1191_368.t0 26.3844
R182 a_1191_368.n2 a_1191_368.t4 26.3844
R183 a_1191_368.n4 a_1191_368.t2 26.3844
R184 a_1191_368.n4 a_1191_368.t1 26.3844
R185 VGND.n25 VGND.n24 263.649
R186 VGND.n12 VGND.n11 209.825
R187 VGND.n41 VGND.n2 209.243
R188 VGND.n16 VGND.n10 208.077
R189 VGND.n26 VGND.n25 185
R190 VGND.n28 VGND.n4 185
R191 VGND.n30 VGND.n29 185
R192 VGND.n13 VGND.t5 161.357
R193 VGND.n44 VGND.n43 116.644
R194 VGND.n37 VGND.n36 116.644
R195 VGND.n29 VGND.n28 88.3789
R196 VGND.n10 VGND.t6 36.487
R197 VGND.n10 VGND.t11 35.6762
R198 VGND.n36 VGND.t1 34.0546
R199 VGND.n36 VGND.t8 34.0546
R200 VGND.n2 VGND.t7 34.0546
R201 VGND.n23 VGND.n7 31.2252
R202 VGND.n27 VGND.n26 28.7974
R203 VGND.n18 VGND.n17 27.1064
R204 VGND.n37 VGND.n1 27.1064
R205 VGND.n35 VGND.n34 26.9232
R206 VGND.n43 VGND.t12 25.1356
R207 VGND.n30 VGND.n27 24.2798
R208 VGND.n42 VGND.n41 24.0946
R209 VGND.n17 VGND.n16 23.3417
R210 VGND.n41 VGND.n1 23.3417
R211 VGND.n12 VGND.n9 22.9652
R212 VGND.n29 VGND.t0 22.7032
R213 VGND.n28 VGND.t13 22.7032
R214 VGND.n25 VGND.t2 22.7032
R215 VGND.n11 VGND.t3 22.7032
R216 VGND.n11 VGND.t4 22.7032
R217 VGND.n2 VGND.t10 22.7032
R218 VGND.n43 VGND.t9 22.7032
R219 VGND.n16 VGND.n9 22.2123
R220 VGND.n44 VGND.n42 21.8358
R221 VGND.n18 VGND.n7 20.3299
R222 VGND.n37 VGND.n35 20.3299
R223 VGND.n14 VGND.n9 9.3005
R224 VGND.n16 VGND.n15 9.3005
R225 VGND.n17 VGND.n8 9.3005
R226 VGND.n19 VGND.n18 9.3005
R227 VGND.n20 VGND.n7 9.3005
R228 VGND.n23 VGND.n22 9.3005
R229 VGND.n21 VGND.n6 9.3005
R230 VGND.n27 VGND.n5 9.3005
R231 VGND.n32 VGND.n31 9.3005
R232 VGND.n34 VGND.n33 9.3005
R233 VGND.n35 VGND.n3 9.3005
R234 VGND.n38 VGND.n37 9.3005
R235 VGND.n39 VGND.n1 9.3005
R236 VGND.n41 VGND.n40 9.3005
R237 VGND.n42 VGND.n0 9.3005
R238 VGND.n45 VGND.n44 7.24643
R239 VGND.n13 VGND.n12 6.6595
R240 VGND.n24 VGND.n6 6.43509
R241 VGND.n31 VGND.n4 6.43509
R242 VGND.n31 VGND.n30 1.10753
R243 VGND.n14 VGND.n13 0.655456
R244 VGND.n26 VGND.n6 0.277257
R245 VGND VGND.n45 0.276102
R246 VGND.n24 VGND.n23 0.208068
R247 VGND.n34 VGND.n4 0.208068
R248 VGND.n45 VGND.n0 0.154713
R249 VGND.n15 VGND.n14 0.122949
R250 VGND.n15 VGND.n8 0.122949
R251 VGND.n19 VGND.n8 0.122949
R252 VGND.n20 VGND.n19 0.122949
R253 VGND.n22 VGND.n20 0.122949
R254 VGND.n22 VGND.n21 0.122949
R255 VGND.n21 VGND.n5 0.122949
R256 VGND.n32 VGND.n5 0.122949
R257 VGND.n33 VGND.n32 0.122949
R258 VGND.n33 VGND.n3 0.122949
R259 VGND.n38 VGND.n3 0.122949
R260 VGND.n39 VGND.n38 0.122949
R261 VGND.n40 VGND.n39 0.122949
R262 VGND.n40 VGND.n0 0.122949
R263 VNB.t2 VNB.t11 5416.27
R264 VNB VNB.t12 2298.16
R265 VNB.t13 VNB.t0 2251.97
R266 VNB.t11 VNB.t6 1374.28
R267 VNB.t8 VNB.t1 1316.54
R268 VNB.t9 VNB.t10 1177.95
R269 VNB.t10 VNB.t7 1154.86
R270 VNB.t12 VNB.t9 1027.82
R271 VNB.t3 VNB.t5 993.177
R272 VNB.t4 VNB.t3 993.177
R273 VNB.t6 VNB.t4 993.177
R274 VNB.t0 VNB.t2 993.177
R275 VNB.t1 VNB.t13 993.177
R276 VNB.t7 VNB.t8 993.177
R277 C.n0 C.t1 328.832
R278 C.n4 C.t3 240.125
R279 C.n2 C.t2 226.809
R280 C.n3 C.t4 226.809
R281 C.n4 C.t6 226.809
R282 C.n11 C.n10 152
R283 C.n9 C.n8 152
R284 C.n7 C.n6 152
R285 C.n0 C.t5 142.994
R286 C.n5 C.t7 142.994
R287 C.n1 C.t0 142.994
R288 C.n1 C.n0 121.376
R289 C.n10 C.n9 33.1076
R290 C.n6 C.n3 22.3965
R291 C.n6 C.n5 19.9621
R292 C.n9 C.n3 10.7116
R293 C.n8 C.n7 10.1214
R294 C.n11 C 8.63306
R295 C.n10 C.n2 7.30353
R296 C.n5 C.n4 6.32979
R297 C C.n11 5.65631
R298 C.n7 C 2.67957
R299 C.n8 C 1.48887
R300 C.n2 C.n1 1.46111
R301 a_778_368.n4 a_778_368.n3 648.34
R302 a_778_368.n5 a_778_368.n4 585
R303 a_778_368.n2 a_778_368.n0 359.479
R304 a_778_368.n2 a_778_368.n1 302.74
R305 a_778_368.n4 a_778_368.n2 93.5936
R306 a_778_368.n3 a_778_368.t0 35.1791
R307 a_778_368.n1 a_778_368.t7 35.1791
R308 a_778_368.n5 a_778_368.t2 30.7817
R309 a_778_368.n3 a_778_368.t1 26.3844
R310 a_778_368.n0 a_778_368.t4 26.3844
R311 a_778_368.n0 a_778_368.t5 26.3844
R312 a_778_368.n1 a_778_368.t6 26.3844
R313 a_778_368.t3 a_778_368.n5 26.3844
R314 D_N.n0 D_N.t1 296.966
R315 D_N.n0 D_N.t0 201.905
R316 D_N.n2 D_N 168.899
R317 D_N D_N.n1 157.572
R318 D_N.n4 D_N.n3 152
R319 D_N.n2 D_N.t2 144.3
R320 D_N.n3 D_N.n1 19.8647
R321 D_N.n3 D_N.n2 13.6635
R322 D_N.n1 D_N.n0 7.01141
R323 D_N.n4 D_N 6.47579
R324 D_N D_N.n4 4.66874
R325 B.n1 B.t0 247.988
R326 B.n2 B.t1 226.809
R327 B.n12 B.t2 226.809
R328 B.n5 B.t3 226.809
R329 B.n7 B.n6 209.16
R330 B.n11 B.n4 196.013
R331 B.n14 B.n3 196.013
R332 B.n1 B.t4 196.013
R333 B.n16 B.n15 152
R334 B.n13 B.n0 152
R335 B.n10 B.n9 152
R336 B.n8 B.n7 152
R337 B.n2 B.n1 44.549
R338 B.n10 B.n5 44.549
R339 B.n14 B.n13 33.5944
R340 B.n13 B.n12 21.1793
R341 B.n12 B.n11 18.2581
R342 B.n15 B.n14 16.0672
R343 B.n8 B 11.1633
R344 B.n11 B.n10 10.2247
R345 B.n16 B.n0 10.1214
R346 B.n9 B 7.29352
R347 B.n9 B 6.99585
R348 B.n7 B.n5 5.11262
R349 B B.n8 3.12608
R350 B B.n0 2.82841
R351 B.n15 B.n2 2.19141
R352 B B.n16 1.34003
C0 VPB B 0.153721f
C1 D_N C 3.93e-20
C2 A VPWR 0.074373f
C3 Y VGND 1.36656f
C4 A Y 0.19538f
C5 C B 0.022225f
C6 A VGND 0.074246f
C7 VPB VPWR 0.247032f
C8 VPB Y 0.017275f
C9 D_N VPWR 0.066162f
C10 VPB VGND 0.014915f
C11 C VPWR 0.028363f
C12 D_N Y 0.002469f
C13 VPB A 0.138517f
C14 C Y 0.406623f
C15 D_N VGND 0.034261f
C16 B VPWR 0.029798f
C17 C VGND 0.0816f
C18 B Y 0.250075f
C19 B VGND 0.069584f
C20 B A 0.088166f
C21 VPB D_N 0.125949f
C22 VPWR Y 0.035247f
C23 VPB C 0.152308f
C24 VPWR VGND 0.161488f
C25 VGND VNB 1.1706f
C26 Y VNB 0.086503f
C27 VPWR VNB 0.935178f
C28 A VNB 0.440687f
C29 B VNB 0.432256f
C30 C VNB 0.471577f
C31 D_N VNB 0.303524f
C32 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4b_2 VNB VPB VPWR VGND A B C D_N Y
X0 a_498_368.t3 B.t0 a_701_368.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t2 D_N.t0 a_27_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.295 ps=2.59 w=1 l=0.15
X2 VGND.t8 a_27_392.t2 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=1.28 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 a_229_368.t1 C.t0 a_498_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_498_368.t1 C.t1 a_229_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_701_368.t0 A.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1736 ps=1.43 w=1.12 l=0.15
X6 a_229_368.t3 a_27_392.t3 Y.t7 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t8 a_27_392.t4 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1469 ps=1.16 w=0.74 l=0.15
X8 Y.t6 a_27_392.t5 a_229_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X9 VGND.t3 A.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=2.08 as=0.12395 ps=1.075 w=0.74 l=0.15
X10 VGND.t4 D_N.t1 a_27_392.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1469 pd=1.16 as=0.1824 ps=1.85 w=0.64 l=0.15
X11 Y.t1 C.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1998 ps=1.28 w=0.74 l=0.15
X12 Y.t0 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12395 pd=1.075 as=0.26825 ps=1.465 w=0.74 l=0.15
X13 Y.t5 B.t1 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1369 pd=1.11 as=0.148 ps=1.14 w=0.74 l=0.15
X14 VGND.t2 C.t3 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.148 pd=1.14 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VGND.t5 B.t2 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.26825 pd=1.465 as=0.1369 ps=1.11 w=0.74 l=0.15
X16 VPWR.t1 A.t3 a_701_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_701_368.t2 B.t3 a_498_368.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B.n0 B.t3 344.606
R1 B.n1 B.t0 226.809
R2 B.n2 B.t1 209.16
R3 B.n0 B.t2 196.013
R4 B.n2 B 153.637
R5 B.n4 B.n3 152
R6 B.n3 B.n2 49.6611
R7 B.n3 B.n1 10.955
R8 B.n4 B 8.48422
R9 B B.n4 5.80515
R10 B.n1 B.n0 2.19141
R11 a_701_368.n1 a_701_368.t3 448.33
R12 a_701_368.t0 a_701_368.n1 294.255
R13 a_701_368.n1 a_701_368.n0 207.946
R14 a_701_368.n0 a_701_368.t1 26.3844
R15 a_701_368.n0 a_701_368.t2 26.3844
R16 a_498_368.n1 a_498_368.n0 979.997
R17 a_498_368.n0 a_498_368.t0 26.3844
R18 a_498_368.n0 a_498_368.t1 26.3844
R19 a_498_368.t2 a_498_368.n1 26.3844
R20 a_498_368.n1 a_498_368.t3 26.3844
R21 VPB.t0 VPB.t8 515.861
R22 VPB.t2 VPB.t6 515.861
R23 VPB VPB.t2 257.93
R24 VPB.t5 VPB.t1 234.946
R25 VPB.t7 VPB.t5 229.839
R26 VPB.t8 VPB.t7 229.839
R27 VPB.t4 VPB.t0 229.839
R28 VPB.t3 VPB.t4 229.839
R29 VPB.t6 VPB.t3 229.839
R30 D_N.n0 D_N.t1 268.313
R31 D_N.n0 D_N.t0 225.202
R32 D_N D_N.n0 154.522
R33 a_27_392.n0 a_27_392.t3 300.325
R34 a_27_392.t1 a_27_392.n5 277.921
R35 a_27_392.n2 a_27_392.t5 261.62
R36 a_27_392.n3 a_27_392.t4 164.464
R37 a_27_392.n4 a_27_392.n1 162.363
R38 a_27_392.n0 a_27_392.t2 154.24
R39 a_27_392.n4 a_27_392.n3 152
R40 a_27_392.n5 a_27_392.t0 141.343
R41 a_27_392.n5 a_27_392.n4 44.5585
R42 a_27_392.n3 a_27_392.n2 35.7853
R43 a_27_392.n2 a_27_392.n1 13.8763
R44 a_27_392.n1 a_27_392.n0 13.146
R45 VPWR.n1 VPWR.n0 322.839
R46 VPWR.n1 VPWR.t2 257.553
R47 VPWR.n0 VPWR.t0 28.1434
R48 VPWR.n0 VPWR.t1 26.3844
R49 VPWR VPWR.n1 0.191868
R50 Y.n4 Y.n0 454.332
R51 Y.n8 Y.n7 185
R52 Y.n9 Y.n8 185
R53 Y.n6 Y.n5 180.393
R54 Y.n3 Y.n2 163.782
R55 Y.n3 Y.n1 95.0012
R56 Y.n8 Y.t4 34.0546
R57 Y.n2 Y.t9 34.0546
R58 Y.n6 Y.n4 32.377
R59 Y.n5 Y.t3 31.6221
R60 Y.n0 Y.t7 26.3844
R61 Y.n0 Y.t6 26.3844
R62 Y.n8 Y.t5 25.9464
R63 Y.n4 Y.n3 24.7808
R64 Y.n5 Y.t0 22.7032
R65 Y.n1 Y.t2 22.7032
R66 Y.n1 Y.t1 22.7032
R67 Y.n2 Y.t8 22.7032
R68 Y.n9 Y 12.6066
R69 Y.n7 Y.n6 5.04292
R70 Y.n7 Y 4.84898
R71 Y Y.n9 1.74595
R72 VGND.n14 VGND.n13 211.183
R73 VGND.n6 VGND.n5 185
R74 VGND.n8 VGND.n7 185
R75 VGND.n20 VGND.n19 185
R76 VGND.n9 VGND.t3 168.427
R77 VGND.n1 VGND.n0 114.885
R78 VGND.n7 VGND.n6 72.1627
R79 VGND.n19 VGND.t1 49.46
R80 VGND.n0 VGND.t4 39.3755
R81 VGND.n19 VGND.t8 38.1086
R82 VGND.n22 VGND.n21 36.1417
R83 VGND.n0 VGND.t7 35.7861
R84 VGND.n13 VGND.t2 34.0546
R85 VGND.n13 VGND.t6 30.8113
R86 VGND.n18 VGND.n3 29.9148
R87 VGND.n12 VGND.n11 27.6485
R88 VGND.n14 VGND.n12 24.8476
R89 VGND.n7 VGND.t0 22.7032
R90 VGND.n6 VGND.t5 22.7032
R91 VGND.n14 VGND.n3 22.5887
R92 VGND.n21 VGND.n20 10.1295
R93 VGND.n24 VGND.n1 9.96261
R94 VGND.n23 VGND.n22 9.3005
R95 VGND.n21 VGND.n2 9.3005
R96 VGND.n18 VGND.n17 9.3005
R97 VGND.n16 VGND.n3 9.3005
R98 VGND.n15 VGND.n14 9.3005
R99 VGND.n12 VGND.n4 9.3005
R100 VGND.n11 VGND.n10 9.3005
R101 VGND.n22 VGND.n1 9.03579
R102 VGND.n9 VGND.n8 7.16793
R103 VGND.n8 VGND.n5 6.51021
R104 VGND.n20 VGND.n18 2.80342
R105 VGND.n10 VGND.n9 0.58252
R106 VGND.n11 VGND.n5 0.366214
R107 VGND VGND.n24 0.163644
R108 VGND.n24 VGND.n23 0.144205
R109 VGND.n10 VGND.n4 0.122949
R110 VGND.n15 VGND.n4 0.122949
R111 VGND.n16 VGND.n15 0.122949
R112 VGND.n17 VGND.n16 0.122949
R113 VGND.n17 VGND.n2 0.122949
R114 VGND.n23 VGND.n2 0.122949
R115 VNB.t5 VNB.t0 2021
R116 VNB.t8 VNB.t1 1593.7
R117 VNB VNB.t4 1455.12
R118 VNB.t4 VNB.t7 1316.54
R119 VNB.t2 VNB.t6 1270.34
R120 VNB.t6 VNB.t5 1201.05
R121 VNB.t7 VNB.t8 1154.86
R122 VNB.t0 VNB.t3 1120.21
R123 VNB.t1 VNB.t2 993.177
R124 C.n0 C.t0 233.381
R125 C.n1 C.t1 226.809
R126 C.n1 C.t2 199.666
R127 C.n0 C.t3 196.013
R128 C.n3 C.n2 152
R129 C.n2 C.n0 49.6611
R130 C.n3 C 12.0563
R131 C.n2 C.n1 9.49444
R132 C C.n3 2.23306
R133 a_229_368.t1 a_229_368.n1 686.431
R134 a_229_368.n1 a_229_368.t2 297.844
R135 a_229_368.n1 a_229_368.n0 287.964
R136 a_229_368.n0 a_229_368.t0 26.3844
R137 a_229_368.n0 a_229_368.t3 26.3844
R138 A.n0 A.t0 226.809
R139 A.n1 A.t3 226.809
R140 A.n0 A.t1 198.204
R141 A.n1 A.t2 197.475
R142 A.n5 A.n4 152
R143 A.n3 A.n2 152
R144 A.n4 A.n3 49.6611
R145 A.n4 A.n0 10.955
R146 A.n2 A 10.2703
R147 A A.n5 8.18655
R148 A.n3 A.n1 6.57323
R149 A.n5 A 6.10283
R150 A.n2 A 4.0191
C0 VGND B 0.038477f
C1 C VPWR 0.015083f
C2 B A 0.072002f
C3 VGND A 0.065334f
C4 C Y 0.209391f
C5 B VPWR 0.018209f
C6 VGND VPWR 0.093146f
C7 A VPWR 0.042696f
C8 B Y 0.151604f
C9 VPB C 0.067634f
C10 VGND Y 0.660592f
C11 A Y 0.087023f
C12 VPB B 0.093995f
C13 D_N C 0.004474f
C14 VGND VPB 0.011279f
C15 VPWR Y 0.01538f
C16 VPB A 0.069537f
C17 VGND D_N 0.015835f
C18 VPB VPWR 0.151437f
C19 D_N VPWR 0.052921f
C20 VPB Y 0.009192f
C21 D_N Y 7.98e-19
C22 VPB D_N 0.063104f
C23 C B 0.036473f
C24 VGND C 0.031382f
C25 VGND VNB 0.71819f
C26 Y VNB 0.045934f
C27 VPWR VNB 0.543893f
C28 A VNB 0.258364f
C29 B VNB 0.244444f
C30 C VNB 0.197741f
C31 D_N VNB 0.162343f
C32 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4b_1 VNB VPB VPWR VGND Y D_N A B C
X0 Y.t0 C.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1591 ps=1.17 w=0.74 l=0.15
X1 VPWR.t0 D_N.t0 a_57_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2177 pd=1.54 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 a_344_368.t0 B.t0 a_260_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.1512 ps=1.39 w=1.12 l=0.15
X3 a_446_368.t0 C.t1 a_344_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2016 ps=1.48 w=1.12 l=0.15
X4 a_260_368.t1 A.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.2177 ps=1.54 w=1.12 l=0.15
X5 VGND.t1 D_N.t1 a_57_368.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.13925 pd=1.16 as=0.15675 ps=1.67 w=0.55 l=0.15
X6 Y.t1 a_57_368.t2 a_446_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.4648 pd=3.07 as=0.2352 ps=1.54 w=1.12 l=0.15
X7 Y.t4 A.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.13925 ps=1.16 w=0.74 l=0.15
X8 VGND.t2 a_57_368.t3 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VGND.t3 B.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1591 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 C.n0 C.t1 250.909
R1 C.n0 C.t0 220.113
R2 C C.n0 156.614
R3 VGND.n3 VGND.t2 248.095
R4 VGND.n1 VGND.n0 210.018
R5 VGND.n5 VGND.n4 208.079
R6 VGND.n0 VGND.t1 45.8187
R7 VGND.n0 VGND.t4 39.2753
R8 VGND.n7 VGND.n6 36.1417
R9 VGND.n4 VGND.t0 35.6762
R10 VGND.n4 VGND.t3 34.0546
R11 VGND.n9 VGND.n1 12.9744
R12 VGND.n5 VGND.n3 10.1204
R13 VGND.n6 VGND.n2 9.3005
R14 VGND.n8 VGND.n7 9.3005
R15 VGND.n6 VGND.n5 8.28285
R16 VGND.n7 VGND.n1 6.02403
R17 VGND.n3 VGND.n2 0.654227
R18 VGND VGND.n9 0.163644
R19 VGND.n9 VGND.n8 0.144205
R20 VGND.n8 VGND.n2 0.122949
R21 Y Y.n0 589.324
R22 Y.n5 Y.n0 585
R23 Y.n4 Y.n0 585
R24 Y.n3 Y.n1 152.911
R25 Y.n3 Y.n2 101.71
R26 Y Y.n3 96.0717
R27 Y.n0 Y.t1 47.4916
R28 Y.n1 Y.t3 22.7032
R29 Y.n1 Y.t4 22.7032
R30 Y.n2 Y.t2 22.7032
R31 Y.n2 Y.t0 22.7032
R32 Y Y.n4 10.5519
R33 Y Y.n5 9.51401
R34 Y.n5 Y 3.28699
R35 Y.n4 Y 2.24915
R36 VNB VNB.t1 1547.51
R37 VNB.t3 VNB.t0 1339.63
R38 VNB.t1 VNB.t4 1316.54
R39 VNB.t0 VNB.t2 993.177
R40 VNB.t4 VNB.t3 993.177
R41 D_N.n0 D_N.t0 270.188
R42 D_N.n0 D_N.t1 173.52
R43 D_N D_N.n0 154.25
R44 a_57_368.t0 a_57_368.n0 387.56
R45 a_57_368.n0 a_57_368.n1 332.767
R46 a_57_368.n0 a_57_368.t1 294.753
R47 a_57_368.n1 a_57_368.t2 250.909
R48 a_57_368.n1 a_57_368.t3 220.113
R49 VPWR VPWR.n0 343.911
R50 VPWR.n0 VPWR.t0 63.3219
R51 VPWR.n0 VPWR.t1 29.6087
R52 VPB VPB.t0 334.543
R53 VPB.t2 VPB.t4 291.13
R54 VPB.t0 VPB.t3 291.13
R55 VPB.t1 VPB.t2 260.485
R56 VPB.t3 VPB.t1 214.517
R57 B.n0 B.t0 250.909
R58 B.n0 B.t1 220.113
R59 B B.n0 154.828
R60 a_260_368.t0 a_260_368.t1 47.4916
R61 a_344_368.t0 a_344_368.t1 63.3219
R62 a_446_368.t0 a_446_368.t1 73.8755
R63 A.n0 A.t0 250.909
R64 A.n0 A.t1 220.113
R65 A A.n0 154.522
C0 Y A 0.012261f
C1 VPWR C 0.008208f
C2 D_N B 4.43e-19
C3 VGND VPB 0.007954f
C4 D_N Y 0.006816f
C5 VPWR VGND 0.054715f
C6 D_N C 1.91e-19
C7 VGND A 0.025753f
C8 Y B 0.04658f
C9 D_N VGND 0.020993f
C10 B C 0.085884f
C11 Y C 0.049952f
C12 VGND B 0.012912f
C13 Y VGND 0.335421f
C14 VGND C 0.014419f
C15 VPWR VPB 0.096033f
C16 VPB A 0.035637f
C17 D_N VPB 0.039133f
C18 VPWR A 0.017281f
C19 VPWR D_N 0.010859f
C20 VPB B 0.031819f
C21 VPWR B 0.011286f
C22 D_N A 0.056066f
C23 Y VPB 0.016734f
C24 VPWR Y 0.057162f
C25 A B 0.095516f
C26 VPB C 0.033998f
C27 VGND VNB 0.464994f
C28 Y VNB 0.109537f
C29 D_N VNB 0.166249f
C30 VPWR VNB 0.360086f
C31 C VNB 0.102898f
C32 B VNB 0.102837f
C33 A VNB 0.106126f
C34 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4_4 VNB VPB VPWR VGND Y A B C D
X0 a_496_368.t5 C.t0 a_27_368.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_27_368.t2 D.t0 Y.t7 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_879_368.t3 A.t0 VPWR.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3 VGND.t5 C.t1 Y.t9 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.444 ps=1.94 w=0.74 l=0.15
X4 VPWR.t3 A.t1 a_879_368.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=1.45 w=0.74 l=0.15
X6 a_879_368.t4 B.t0 a_496_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_496_368.t1 B.t1 a_879_368.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X8 Y.t6 D.t1 a_27_368.t7 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t8 C.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.444 pd=1.94 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 a_27_368.t0 D.t2 Y.t5 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t3 D.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.4329 pd=1.91 as=0.2442 ps=2.14 w=0.74 l=0.15
X12 VGND.t1 B.t2 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.8621 pd=3.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t2 A.t2 a_879_368.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VGND.t2 D.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.4329 ps=1.91 w=0.74 l=0.15
X15 a_496_368.t6 B.t3 a_879_368.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X16 a_879_368.t7 B.t4 a_496_368.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_879_368.t0 A.t3 VPWR.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=1.45 as=0.8621 ps=3.07 w=0.74 l=0.15
X19 Y.t4 D.t5 a_27_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X20 Y.t0 B.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X21 a_27_368.t5 C.t3 a_496_368.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_496_368.t3 C.t4 a_27_368.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_27_368.t3 C.t5 a_496_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 C.n0 C.t3 232.184
R1 C.n2 C.t4 226.809
R2 C.n3 C.t5 226.809
R3 C.n4 C.t0 226.809
R4 C.n4 C.t2 202.587
R5 C.n0 C.t1 196.013
R6 C C.n1 155.126
R7 C.n10 C.n9 152
R8 C.n8 C.n7 152
R9 C.n6 C.n5 152
R10 C.n9 C.n8 49.6611
R11 C.n2 C.n1 46.0096
R12 C.n5 C.n3 37.246
R13 C.n5 C.n4 28.4823
R14 C.n1 C.n0 13.146
R15 C.n8 C.n3 12.4157
R16 C.n7 C.n6 10.1214
R17 C.n10 C 7.29352
R18 C C.n10 6.99585
R19 C.n9 C.n2 3.65202
R20 C.n7 C 2.82841
R21 C.n6 C 1.34003
R22 a_27_368.n1 a_27_368.t5 430.988
R23 a_27_368.n4 a_27_368.t1 390.623
R24 a_27_368.n5 a_27_368.n4 305.998
R25 a_27_368.n1 a_27_368.n0 300.08
R26 a_27_368.n3 a_27_368.n2 183.916
R27 a_27_368.n4 a_27_368.n3 92.5131
R28 a_27_368.n3 a_27_368.n1 82.9171
R29 a_27_368.n2 a_27_368.t6 26.3844
R30 a_27_368.n2 a_27_368.t2 26.3844
R31 a_27_368.n0 a_27_368.t4 26.3844
R32 a_27_368.n0 a_27_368.t3 26.3844
R33 a_27_368.n5 a_27_368.t7 26.3844
R34 a_27_368.t0 a_27_368.n5 26.3844
R35 a_496_368.n2 a_496_368.n0 347.824
R36 a_496_368.n5 a_496_368.n4 346.411
R37 a_496_368.n4 a_496_368.n3 303.495
R38 a_496_368.n2 a_496_368.n1 303.401
R39 a_496_368.n4 a_496_368.n2 85.0829
R40 a_496_368.n0 a_496_368.t0 26.3844
R41 a_496_368.n0 a_496_368.t1 26.3844
R42 a_496_368.n1 a_496_368.t7 26.3844
R43 a_496_368.n1 a_496_368.t6 26.3844
R44 a_496_368.n3 a_496_368.t4 26.3844
R45 a_496_368.n3 a_496_368.t3 26.3844
R46 a_496_368.n5 a_496_368.t2 26.3844
R47 a_496_368.t5 a_496_368.n5 26.3844
R48 VPB.t7 VPB.t9 515.861
R49 VPB VPB.t3 283.469
R50 VPB.t14 VPB.t15 280.914
R51 VPB.t13 VPB.t11 280.914
R52 VPB.t12 VPB.t4 255.376
R53 VPB.t10 VPB.t1 240.054
R54 VPB.t11 VPB.t14 229.839
R55 VPB.t0 VPB.t13 229.839
R56 VPB.t1 VPB.t0 229.839
R57 VPB.t9 VPB.t10 229.839
R58 VPB.t6 VPB.t7 229.839
R59 VPB.t5 VPB.t6 229.839
R60 VPB.t8 VPB.t5 229.839
R61 VPB.t4 VPB.t8 229.839
R62 VPB.t2 VPB.t12 229.839
R63 VPB.t3 VPB.t2 229.839
R64 D.n0 D.t0 240.361
R65 D.n2 D.t1 226.809
R66 D.n3 D.t2 226.809
R67 D.n4 D.t5 226.809
R68 D.n4 D.t3 198.204
R69 D.n0 D.t4 196.013
R70 D D.n1 155.423
R71 D.n10 D.n9 152
R72 D.n8 D.n7 152
R73 D.n6 D.n5 152
R74 D.n9 D.n8 49.6611
R75 D.n5 D.n3 46.0096
R76 D.n2 D.n1 37.246
R77 D.n1 D.n0 21.9096
R78 D.n5 D.n4 19.7187
R79 D.n9 D.n2 12.4157
R80 D.n7 D.n6 10.1214
R81 D.n10 D 7.5912
R82 D D.n10 6.69817
R83 D.n8 D.n3 3.65202
R84 D.n7 D 2.53073
R85 D.n6 D 1.63771
R86 Y.n2 Y.n0 346.632
R87 Y.n2 Y.n1 299.952
R88 Y.n6 Y.n5 153.624
R89 Y.n10 Y.n9 92.5005
R90 Y.n8 Y.n4 92.5005
R91 Y.n7 Y.n6 92.5005
R92 Y.n15 Y.n14 92.5005
R93 Y.n13 Y.n3 92.5005
R94 Y.n12 Y.n11 92.5005
R95 Y.n8 Y.n7 80.2708
R96 Y.n13 Y.n12 76.2167
R97 Y.n9 Y.n8 68.9194
R98 Y.n14 Y.n13 68.1086
R99 Y Y.n2 65.49
R100 Y.n11 Y.n10 54.4572
R101 Y.n0 Y.t6 35.1791
R102 Y Y.n15 28.136
R103 Y.n0 Y.t7 26.3844
R104 Y.n1 Y.t5 26.3844
R105 Y.n1 Y.t4 26.3844
R106 Y.n12 Y.t2 22.7032
R107 Y.n14 Y.t3 22.7032
R108 Y.n7 Y.t9 22.7032
R109 Y.n9 Y.t8 22.7032
R110 Y.n5 Y.t1 22.7032
R111 Y.n5 Y.t0 22.7032
R112 Y.n6 Y.n4 7.63423
R113 Y.n11 Y.n3 7.24869
R114 Y.n10 Y.n4 6.55472
R115 Y.n15 Y.n3 6.47761
R116 A.n2 A.t1 390.128
R117 A.n5 A.t0 269.925
R118 A.n7 A.t2 240.197
R119 A.n3 A.t3 240.197
R120 A.n2 A.n1 179.947
R121 A.n5 A.n4 179.947
R122 A.n6 A.n0 152
R123 A A.n8 79.1892
R124 A.n7 A.n6 44.549
R125 A.n8 A.n3 33.3172
R126 A.n8 A.n7 25.6895
R127 A.n6 A.n5 13.146
R128 A.n0 A 12.0894
R129 A.n3 A.n2 2.19141
R130 A A.n0 1.56494
R131 VPWR.n2 VPWR.n1 322.423
R132 VPWR.n2 VPWR.n0 322.043
R133 VPWR.n0 VPWR.t1 35.1791
R134 VPWR.n0 VPWR.t3 35.1791
R135 VPWR.n1 VPWR.t0 35.1791
R136 VPWR.n1 VPWR.t2 35.1791
R137 VPWR VPWR.n2 2.05607
R138 a_879_368.n1 a_879_368.t6 440.801
R139 a_879_368.n1 a_879_368.n0 300.08
R140 a_879_368.t3 a_879_368.n5 279.959
R141 a_879_368.n3 a_879_368.n2 205.282
R142 a_879_368.n5 a_879_368.n4 203.458
R143 a_879_368.n3 a_879_368.n1 52.3299
R144 a_879_368.n5 a_879_368.n3 50.4476
R145 a_879_368.n0 a_879_368.t5 28.1434
R146 a_879_368.n0 a_879_368.t7 28.1434
R147 a_879_368.n2 a_879_368.t2 26.3844
R148 a_879_368.n2 a_879_368.t4 26.3844
R149 a_879_368.n4 a_879_368.t1 26.3844
R150 a_879_368.n4 a_879_368.t0 26.3844
R151 VGND.n18 VGND.t3 241.183
R152 VGND.n5 VGND.n4 211.183
R153 VGND.n12 VGND.n11 211.183
R154 VGND.n6 VGND.t1 108.689
R155 VGND.n9 VGND.n3 36.1417
R156 VGND.n10 VGND.n9 36.1417
R157 VGND.n16 VGND.n1 36.1417
R158 VGND.n17 VGND.n16 36.1417
R159 VGND.n4 VGND.t0 34.0546
R160 VGND.n11 VGND.t4 34.0546
R161 VGND.n12 VGND.n10 30.1181
R162 VGND.n4 VGND.t5 22.7032
R163 VGND.n11 VGND.t2 22.7032
R164 VGND.n18 VGND.n17 20.7064
R165 VGND.n12 VGND.n1 17.3181
R166 VGND.n5 VGND.n3 12.0476
R167 VGND.n19 VGND.n18 9.3005
R168 VGND.n17 VGND.n0 9.3005
R169 VGND.n16 VGND.n15 9.3005
R170 VGND.n14 VGND.n1 9.3005
R171 VGND.n13 VGND.n12 9.3005
R172 VGND.n10 VGND.n2 9.3005
R173 VGND.n9 VGND.n8 9.3005
R174 VGND.n7 VGND.n3 9.3005
R175 VGND.n6 VGND.n5 7.35284
R176 VGND.n7 VGND.n6 0.393893
R177 VGND.n8 VGND.n7 0.122949
R178 VGND.n8 VGND.n2 0.122949
R179 VGND.n13 VGND.n2 0.122949
R180 VGND.n14 VGND.n13 0.122949
R181 VGND.n15 VGND.n14 0.122949
R182 VGND.n15 VGND.n0 0.122949
R183 VGND.n19 VGND.n0 0.122949
R184 VGND VGND.n19 0.0617245
R185 VNB.t4 VNB.t5 3118.11
R186 VNB.t3 VNB.t2 3048.82
R187 VNB VNB.t3 1247.24
R188 VNB.t5 VNB.t0 1154.86
R189 VNB.t2 VNB.t4 1154.86
R190 VNB.t0 VNB.t1 993.177
R191 B.n1 B.t0 246.526
R192 B.n2 B.t1 226.809
R193 B.n3 B.t4 226.809
R194 B.n8 B.t3 226.809
R195 B.n4 B.t5 209.16
R196 B.n7 B.t2 196.013
R197 B.n1 B.n0 152
R198 B.n14 B.n13 152
R199 B.n12 B.n11 152
R200 B.n10 B.n9 152
R201 B.n7 B.n6 152
R202 B.n5 B.n4 152
R203 B.n13 B.n12 49.6611
R204 B.n7 B.n4 49.6611
R205 B.n2 B.n1 46.0096
R206 B.n9 B.n3 34.3247
R207 B.n9 B.n8 31.4035
R208 B.n8 B.n7 18.2581
R209 B.n12 B.n3 15.3369
R210 B.n0 B 11.7586
R211 B.n11 B.n10 10.1214
R212 B.n6 B 9.37724
R213 B.n5 B 9.07957
R214 B B.n14 7.5912
R215 B.n14 B 6.69817
R216 B B.n5 5.2098
R217 B.n6 B 4.91213
R218 B.n13 B.n2 3.65202
R219 B.n11 B 3.42376
R220 B B.n0 2.53073
R221 B.n10 B 0.744686
C0 C B 0.076635f
C1 D Y 0.382992f
C2 C A 4.65e-20
C3 VPB VPWR 0.183052f
C4 C Y 0.163531f
C5 D VPWR 0.023325f
C6 B A 0.057605f
C7 VPB VGND 0.01083f
C8 D VGND 0.041352f
C9 C VPWR 0.027061f
C10 B Y 0.23547f
C11 A Y 0.09577f
C12 B VPWR 0.031028f
C13 C VGND 0.038024f
C14 A VPWR 0.075421f
C15 B VGND 0.04942f
C16 A VGND 0.081824f
C17 Y VPWR 0.032542f
C18 Y VGND 1.06134f
C19 VPB D 0.140908f
C20 VPWR VGND 0.137597f
C21 VPB C 0.139088f
C22 VPB B 0.176315f
C23 D C 0.070646f
C24 VPB A 0.148479f
C25 VPB Y 0.010837f
C26 D A 2.27e-20
C27 VGND VNB 1.03916f
C28 VPWR VNB 0.780665f
C29 Y VNB 0.129705f
C30 A VNB 0.41918f
C31 B VNB 0.400584f
C32 C VNB 0.340808f
C33 D VNB 0.37065f
C34 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4_2 VNB VPB VPWR VGND C A B D Y
X0 a_490_368.t2 A.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_116_368.t2 C.t0 a_27_368.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t0 A.t1 a_490_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2184 ps=1.51 w=1.12 l=0.15
X3 Y.t4 D.t0 a_116_368.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.182 pd=1.445 as=0.1764 ps=1.435 w=1.12 l=0.15
X4 VGND.t3 C.t1 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1184 ps=1.06 w=0.74 l=0.15
X5 Y.t2 D.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.3329 ps=3 w=0.74 l=0.15
X6 VGND.t1 A.t2 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_490_368.t0 B.t0 a_27_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1848 ps=1.45 w=1.12 l=0.15
X8 a_27_368.t2 C.t2 a_116_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X10 a_116_368.t0 D.t2 Y.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.182 ps=1.445 w=1.12 l=0.15
X11 a_27_368.t1 B.t2 a_490_368.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n1 A.t0 276.955
R1 A.n0 A.t1 263.81
R2 A A.n1 161.067
R3 A.n0 A.t2 154.24
R4 A.n1 A.n0 48.2005
R5 VPWR VPWR.n0 611.568
R6 VPWR.n0 VPWR.t1 26.3844
R7 VPWR.n0 VPWR.t0 26.3844
R8 a_490_368.n1 a_490_368.n0 646.279
R9 a_490_368.n0 a_490_368.t1 35.1791
R10 a_490_368.n0 a_490_368.t0 33.4201
R11 a_490_368.n1 a_490_368.t3 26.3844
R12 a_490_368.t2 a_490_368.n1 26.3844
R13 VPB.t0 VPB.t2 275.807
R14 VPB VPB.t5 257.93
R15 VPB.t4 VPB.t0 245.161
R16 VPB.t7 VPB.t1 242.608
R17 VPB.t5 VPB.t7 237.5
R18 VPB.t3 VPB.t6 229.839
R19 VPB.t2 VPB.t3 229.839
R20 VPB.t1 VPB.t4 229.839
R21 C C.t0 520.183
R22 C.n0 C.t2 258.942
R23 C.n0 C.t1 210.474
R24 C.n1 C.n0 160.922
R25 C.n1 C 16.6962
R26 C C.n1 3.89615
R27 C.n1 C 3.29747
R28 a_27_368.n0 a_27_368.t1 545.159
R29 a_27_368.n0 a_27_368.t3 350.3
R30 a_27_368.n1 a_27_368.n0 195.115
R31 a_27_368.t0 a_27_368.n1 31.6612
R32 a_27_368.n1 a_27_368.t2 26.3844
R33 a_116_368.n1 a_116_368.n0 1207.4
R34 a_116_368.n1 a_116_368.t3 28.1434
R35 a_116_368.t2 a_116_368.n1 27.2639
R36 a_116_368.n0 a_116_368.t1 26.3844
R37 a_116_368.n0 a_116_368.t0 26.3844
R38 D D.n1 501.894
R39 D.n1 D.t0 274.74
R40 D.n0 D.t2 269.652
R41 D.n0 D.t1 145.153
R42 D.n1 D.n0 66.1856
R43 Y Y.n0 587.4
R44 Y Y.n3 189.397
R45 Y.n3 Y.n1 155.799
R46 Y.n3 Y.n2 95.742
R47 Y.n2 Y.t2 29.1897
R48 Y.n0 Y.t3 29.0228
R49 Y.n0 Y.t4 28.1434
R50 Y.n2 Y.t5 22.7032
R51 Y.n1 Y.t1 22.7032
R52 Y.n1 Y.t0 22.7032
R53 VGND.n6 VGND.n0 369.139
R54 VGND.n4 VGND.n3 210.018
R55 VGND.n7 VGND.n6 185
R56 VGND.n2 VGND.t1 143.519
R57 VGND.n6 VGND.t2 38.8915
R58 VGND.n3 VGND.t0 34.0546
R59 VGND.n3 VGND.t3 34.0546
R60 VGND.n5 VGND.n4 27.8593
R61 VGND.n7 VGND.n5 25.6719
R62 VGND.n9 VGND.n8 9.3005
R63 VGND.n5 VGND.n1 9.3005
R64 VGND.n10 VGND.n0 8.42306
R65 VGND.n8 VGND.n0 8.03554
R66 VGND.n4 VGND.n2 6.55159
R67 VGND.n2 VGND.n1 0.50072
R68 VGND.n8 VGND.n7 0.280792
R69 VGND VGND.n10 0.160812
R70 VGND.n10 VGND.n9 0.147
R71 VGND.n9 VGND.n1 0.122949
R72 VNB VNB.t2 3372.18
R73 VNB.t3 VNB.t0 1316.54
R74 VNB.t2 VNB.t3 1085.56
R75 VNB.t0 VNB.t1 993.177
R76 B B.n0 272.339
R77 B.n0 B.t0 258.942
R78 B.n4 B.t2 256.428
R79 B.n0 B.t1 210.474
R80 B.n5 B.n4 152
R81 B.n3 B.n2 152
R82 B.n3 B.n1 114.257
R83 B.n4 B.n3 33.4454
R84 B.n2 B 11.055
R85 B.n5 B 9.89141
R86 B B.n1 7.43094
R87 B.n1 B 6.49682
R88 B B.n5 4.46111
R89 B.n2 B 3.29747
C0 C B 0.085493f
C1 A Y 0.010402f
C2 D B 0.004048f
C3 A VPWR 0.026531f
C4 A VGND 0.058416f
C5 Y VPWR 0.010509f
C6 A VPB 0.057476f
C7 Y VGND 0.355987f
C8 A C 0.001747f
C9 Y VPB 0.009593f
C10 VPWR VGND 0.067701f
C11 VPWR VPB 0.101227f
C12 A D 4.07e-19
C13 Y C 0.299837f
C14 Y D 0.100699f
C15 A B 0.233762f
C16 VGND VPB 0.005596f
C17 VPWR C 0.02029f
C18 VGND C 0.021974f
C19 VPWR D 0.01124f
C20 Y B 0.060231f
C21 VPB C 0.065459f
C22 VPWR B 0.028059f
C23 VGND D 0.089216f
C24 VPB D 0.062331f
C25 VGND B 0.119301f
C26 C D 0.168398f
C27 VPB B 0.083008f
C28 VGND VNB 0.544815f
C29 VPWR VNB 0.424689f
C30 Y VNB 0.089445f
C31 A VNB 0.175226f
C32 B VNB 0.438919f
C33 D VNB 0.368654f
C34 C VNB 0.203785f
C35 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor4_1 VNB VPB VPWR VGND Y D C B A
X0 Y.t0 D.t0 a_342_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X1 VGND.t1 B.t0 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1924 pd=1.26 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t2 C.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1924 ps=1.26 w=0.74 l=0.15
X3 Y.t4 A.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X4 a_228_368.t1 B.t1 a_144_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.1512 ps=1.39 w=1.12 l=0.15
X5 a_144_368.t1 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 a_342_368.t0 C.t1 a_228_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.2352 ps=1.54 w=1.12 l=0.15
X7 VGND.t0 D.t1 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.23225 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 D.n0 D.t0 250.909
R1 D.n0 D.t1 220.113
R2 D D.n0 158.102
R3 a_342_368.t0 a_342_368.t1 73.8755
R4 Y Y.n0 588.077
R5 Y.n4 Y.n0 290.363
R6 Y.n3 Y.n1 162.103
R7 Y.n4 Y.n3 108.48
R8 Y.n3 Y.n2 101.71
R9 Y.n0 Y.t0 26.3844
R10 Y.n1 Y.t3 22.7032
R11 Y.n1 Y.t4 22.7032
R12 Y.n2 Y.t1 22.7032
R13 Y.n2 Y.t2 22.7032
R14 Y Y.n4 9.81567
R15 VPB VPB.t0 329.435
R16 VPB.t1 VPB.t2 291.13
R17 VPB.t3 VPB.t1 291.13
R18 VPB.t0 VPB.t3 214.517
R19 B.n0 B.t1 250.909
R20 B.n0 B.t0 220.113
R21 B B.n0 154.447
R22 VGND.n3 VGND.t0 241.319
R23 VGND.n2 VGND.n1 211.183
R24 VGND.n7 VGND.t3 145.03
R25 VGND.n1 VGND.t2 50.2708
R26 VGND.n6 VGND.n5 36.1417
R27 VGND.n1 VGND.t1 34.0546
R28 VGND.n3 VGND.n2 17.6341
R29 VGND.n8 VGND.n7 9.3005
R30 VGND.n5 VGND.n4 9.3005
R31 VGND.n6 VGND.n0 9.3005
R32 VGND.n7 VGND.n6 8.28285
R33 VGND.n5 VGND.n2 0.753441
R34 VGND.n4 VGND.n3 0.667728
R35 VGND.n4 VGND.n0 0.122949
R36 VGND.n8 VGND.n0 0.122949
R37 VGND VGND.n8 0.0617245
R38 VNB.t1 VNB.t2 1547.51
R39 VNB VNB.t3 1524.41
R40 VNB.t2 VNB.t0 993.177
R41 VNB.t3 VNB.t1 993.177
R42 C.n0 C.t1 250.909
R43 C.n0 C.t0 220.113
R44 C C.n0 154.522
R45 A.n0 A.t1 276.767
R46 A.n0 A.t0 169.389
R47 A A.n0 159.612
R48 a_144_368.t0 a_144_368.t1 47.4916
R49 a_228_368.t0 a_228_368.t1 73.8755
R50 VPWR VPWR.t0 256.74
C0 C VPWR 0.016108f
C1 D VPWR 0.011278f
C2 A VGND 0.05525f
C3 VGND VPB 0.007525f
C4 Y VGND 0.330614f
C5 B VGND 0.015873f
C6 C VGND 0.013638f
C7 A VPB 0.044137f
C8 A Y 0.009149f
C9 Y VPB 0.025359f
C10 D VGND 0.014116f
C11 A B 0.081019f
C12 B VPB 0.036802f
C13 B Y 0.063295f
C14 VPWR VGND 0.050518f
C15 A C 2.53e-19
C16 C VPB 0.036913f
C17 C Y 0.063905f
C18 B C 0.105574f
C19 A D 1.49e-19
C20 D VPB 0.039039f
C21 D Y 0.117332f
C22 A VPWR 0.04734f
C23 B D 0.001655f
C24 VPWR VPB 0.090802f
C25 VPWR Y 0.067628f
C26 B VPWR 0.087703f
C27 C D 0.093486f
C28 VGND VNB 0.442654f
C29 Y VNB 0.114573f
C30 VPWR VNB 0.355318f
C31 D VNB 0.133428f
C32 C VNB 0.105202f
C33 B VNB 0.112937f
C34 A VNB 0.175904f
C35 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3b_4 VNB VPB VPWR VGND Y A B C_N
X0 Y.t7 a_468_264.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 VPWR.t2 C_N.t0 a_468_264.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X2 a_468_264.t1 C_N.t1 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.231 ps=1.555 w=0.84 l=0.15
X3 VGND.t5 A.t0 Y.t9 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=1.29 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t6 A.t1 Y.t10 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 VGND.t0 B.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_126_368# B.t1 a_27_368.t7 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.495 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_27_368.t6 B.t2 a_126_368# VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR A a_126_368# VPB sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t6 a_468_264.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 a_126_368# A.t2 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X11 a_126_368# A.t3 VPWR.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 Y.t14 A.t4 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2035 ps=1.29 w=0.74 l=0.15
X13 VPWR.t4 A.t5 a_126_368# VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y.t11 B.t3 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.2442 ps=2.14 w=0.74 l=0.15
X15 Y.t12 B.t4 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 VGND.t2 a_468_264.t5 Y.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t1 a_468_264.t6 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_27_368.t3 a_468_264.t7 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t2 a_468_264.t8 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 VGND.t10 B.t5 Y.t13 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.11285 ps=1.045 w=0.74 l=0.15
X21 a_126_368# B.t6 a_27_368.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X22 a_27_368.t1 a_468_264.t9 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 Y.t8 a_468_264.t10 a_27_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_27_368.t4 B.t7 a_126_368# VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.21 ps=1.495 w=1.12 l=0.15
X25 Y.t15 A.t6 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X26 a_468_264.t2 C_N.t2 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.6771 pd=3.31 as=0.1295 ps=1.09 w=0.74 l=0.15
R0 a_468_264.n13 a_468_264.n12 307.411
R1 a_468_264.n4 a_468_264.t10 244.335
R2 a_468_264.n1 a_468_264.t7 234.841
R3 a_468_264.n8 a_468_264.t8 234.841
R4 a_468_264.n3 a_468_264.t9 234.841
R5 a_468_264.n12 a_468_264.n11 213.946
R6 a_468_264.n1 a_468_264.t5 197.328
R7 a_468_264.n9 a_468_264.t4 186.374
R8 a_468_264.n4 a_468_264.t3 186.374
R9 a_468_264.n2 a_468_264.t6 186.374
R10 a_468_264.n6 a_468_264.n5 165.189
R11 a_468_264.n7 a_468_264.n6 152
R12 a_468_264.n9 a_468_264.n0 152
R13 a_468_264.n11 a_468_264.n10 152
R14 a_468_264.n12 a_468_264.t2 150.008
R15 a_468_264.n10 a_468_264.n9 49.6611
R16 a_468_264.n5 a_468_264.n4 36.5157
R17 a_468_264.n8 a_468_264.n7 35.7853
R18 a_468_264.t0 a_468_264.n13 35.1791
R19 a_468_264.n13 a_468_264.t1 35.1791
R20 a_468_264.n7 a_468_264.n2 23.3702
R21 a_468_264.n5 a_468_264.n3 19.7187
R22 a_468_264.n9 a_468_264.n8 13.8763
R23 a_468_264.n11 a_468_264.n0 13.1884
R24 a_468_264.n6 a_468_264.n0 13.1884
R25 a_468_264.n3 a_468_264.n2 6.57323
R26 a_468_264.n10 a_468_264.n1 2.19141
R27 VGND.n24 VGND.n2 211.183
R28 VGND.n17 VGND.n5 210.018
R29 VGND.n20 VGND.n19 210.018
R30 VGND.n13 VGND.n12 205.559
R31 VGND.n10 VGND.n9 199.331
R32 VGND.n26 VGND.t8 157.612
R33 VGND.n8 VGND.n7 122.692
R34 VGND.n9 VGND.t11 44.5951
R35 VGND.n9 VGND.t5 44.5951
R36 VGND.n7 VGND.t7 34.0546
R37 VGND.n12 VGND.t12 34.0546
R38 VGND.n12 VGND.t2 34.0546
R39 VGND.n5 VGND.t3 34.0546
R40 VGND.n19 VGND.t0 34.0546
R41 VGND.n2 VGND.t9 34.0546
R42 VGND.n2 VGND.t10 34.0546
R43 VGND.n20 VGND.n1 32.7534
R44 VGND.n11 VGND.n10 31.2476
R45 VGND.n25 VGND.n24 29.7417
R46 VGND.n13 VGND.n4 28.2358
R47 VGND.n18 VGND.n17 25.224
R48 VGND.n7 VGND.t6 22.7032
R49 VGND.n5 VGND.t1 22.7032
R50 VGND.n19 VGND.t4 22.7032
R51 VGND.n17 VGND.n4 22.2123
R52 VGND.n26 VGND.n25 20.7064
R53 VGND.n13 VGND.n11 19.2005
R54 VGND.n24 VGND.n1 17.6946
R55 VGND.n20 VGND.n18 14.6829
R56 VGND.n27 VGND.n26 9.3005
R57 VGND.n11 VGND.n6 9.3005
R58 VGND.n14 VGND.n13 9.3005
R59 VGND.n15 VGND.n4 9.3005
R60 VGND.n17 VGND.n16 9.3005
R61 VGND.n18 VGND.n3 9.3005
R62 VGND.n21 VGND.n20 9.3005
R63 VGND.n22 VGND.n1 9.3005
R64 VGND.n24 VGND.n23 9.3005
R65 VGND.n25 VGND.n0 9.3005
R66 VGND.n10 VGND.n8 5.29514
R67 VGND.n8 VGND.n6 0.44172
R68 VGND.n14 VGND.n6 0.122949
R69 VGND.n15 VGND.n14 0.122949
R70 VGND.n16 VGND.n15 0.122949
R71 VGND.n16 VGND.n3 0.122949
R72 VGND.n21 VGND.n3 0.122949
R73 VGND.n22 VGND.n21 0.122949
R74 VGND.n23 VGND.n22 0.122949
R75 VGND.n23 VGND.n0 0.122949
R76 VGND.n27 VGND.n0 0.122949
R77 VGND VGND.n27 0.0617245
R78 Y.n2 Y.n0 631.081
R79 Y.n2 Y.n1 585
R80 Y.n5 Y.n4 174.263
R81 Y.n9 Y.n7 156.904
R82 Y.n12 Y.n6 101.391
R83 Y.n5 Y.n3 97.8322
R84 Y.n9 Y.n8 96.6686
R85 Y.n11 Y.n10 96.6686
R86 Y.n12 Y.n11 61.4793
R87 Y.n11 Y.n9 50.4476
R88 Y Y.n2 38.701
R89 Y.n7 Y.t10 34.0546
R90 Y.n13 Y.n12 33.5882
R91 Y Y.n13 27.8266
R92 Y.n4 Y.t11 26.7573
R93 Y.n1 Y.t1 26.3844
R94 Y.n1 Y.t8 26.3844
R95 Y.n0 Y.t3 26.3844
R96 Y.n0 Y.t2 26.3844
R97 Y.n4 Y.t13 22.7032
R98 Y.n3 Y.t0 22.7032
R99 Y.n3 Y.t12 22.7032
R100 Y.n10 Y.t5 22.7032
R101 Y.n10 Y.t6 22.7032
R102 Y.n7 Y.t14 22.7032
R103 Y.n8 Y.t9 22.7032
R104 Y.n8 Y.t15 22.7032
R105 Y.n6 Y.t4 22.7032
R106 Y.n6 Y.t7 22.7032
R107 Y.n13 Y.n5 6.4005
R108 VNB.t5 VNB.t11 1616.8
R109 VNB.t2 VNB.t12 1316.54
R110 VNB.t10 VNB.t9 1316.54
R111 VNB VNB.t8 1247.24
R112 VNB.t6 VNB.t7 1154.86
R113 VNB.t11 VNB.t6 1154.86
R114 VNB.t1 VNB.t3 1154.86
R115 VNB.t0 VNB.t4 1154.86
R116 VNB.t8 VNB.t10 1050.92
R117 VNB.t12 VNB.t5 993.177
R118 VNB.t3 VNB.t2 993.177
R119 VNB.t4 VNB.t1 993.177
R120 VNB.t9 VNB.t0 993.177
R121 C_N.n1 C_N.t0 216.845
R122 C_N.n0 C_N.t2 187.981
R123 C_N.n0 C_N.t1 160.399
R124 C_N C_N.n1 158.788
R125 C_N.n1 C_N.n0 18.2986
R126 VPWR.n9 VPWR.t0 838.082
R127 VPWR.n4 VPWR.t2 368.798
R128 VPWR.n7 VPWR.n2 315.349
R129 VPWR.n3 VPWR.t1 286.628
R130 VPWR.n7 VPWR.n6 27.8593
R131 VPWR.n2 VPWR.t3 26.3844
R132 VPWR.n2 VPWR.t4 26.3844
R133 VPWR.n9 VPWR.n8 23.3417
R134 VPWR.n8 VPWR.n7 19.577
R135 VPWR.n6 VPWR.n3 18.824
R136 VPWR.n6 VPWR.n5 9.3005
R137 VPWR.n7 VPWR.n1 9.3005
R138 VPWR.n8 VPWR.n0 9.3005
R139 VPWR.n10 VPWR.n9 7.16774
R140 VPWR.n4 VPWR.n3 6.90183
R141 VPWR VPWR.n10 1.13494
R142 VPWR.n5 VPWR.n4 0.606651
R143 VPWR.n10 VPWR.n0 0.157082
R144 VPWR.n5 VPWR.n1 0.122949
R145 VPWR.n1 VPWR.n0 0.122949
R146 VPB.t9 VPB.t6 528.63
R147 VPB.t3 VPB.t4 515.861
R148 VPB VPB.t11 283.469
R149 VPB.t5 VPB.t12 268.146
R150 VPB.t6 VPB.t7 229.839
R151 VPB.t10 VPB.t9 229.839
R152 VPB.t4 VPB.t10 229.839
R153 VPB.t2 VPB.t3 229.839
R154 VPB.t1 VPB.t2 229.839
R155 VPB.t0 VPB.t1 229.839
R156 VPB.t12 VPB.t0 229.839
R157 VPB.t8 VPB.t5 229.839
R158 VPB.t11 VPB.t8 229.839
R159 A.n2 A.n1 276.205
R160 A.n13 A.t3 261.62
R161 A.n3 A.t5 261.62
R162 A.n5 A.t2 261.62
R163 A.n4 A.t6 180.531
R164 A.n8 A.n4 165.189
R165 A.n6 A.t0 154.24
R166 A.n11 A.t4 154.24
R167 A.n2 A.t1 154.24
R168 A.n15 A.n14 152
R169 A.n12 A.n0 152
R170 A.n10 A.n9 152
R171 A.n8 A.n7 152
R172 A.n7 A.n3 43.0884
R173 A.n14 A.n13 40.1672
R174 A.n11 A.n10 39.4369
R175 A.n5 A.n4 27.0217
R176 A A.n15 16.6793
R177 A.n15 A.n0 13.1884
R178 A.n9 A.n0 13.1884
R179 A.n9 A.n8 13.1884
R180 A.n14 A.n2 13.146
R181 A.n7 A.n6 13.146
R182 A.n12 A.n11 10.2247
R183 A.n13 A.n12 9.49444
R184 A.n6 A.n5 9.49444
R185 A.n10 A.n3 6.57323
R186 B.n0 B.t7 226.809
R187 B.n3 B.t1 226.809
R188 B.n10 B.t2 226.809
R189 B.n4 B.t6 226.809
R190 B.n4 B.t3 198.204
R191 B.n0 B.t0 198.204
R192 B.n9 B.t5 196.013
R193 B.n2 B.t4 196.013
R194 B B.n1 153.637
R195 B.n12 B.n11 152
R196 B.n8 B.n7 152
R197 B.n6 B.n5 152
R198 B.n8 B.n5 49.6611
R199 B.n1 B.n0 48.2005
R200 B.n11 B.n10 44.549
R201 B.n11 B.n3 21.1793
R202 B.n3 B.n2 16.0672
R203 B.n6 B 14.14
R204 B.n2 B.n1 12.4157
R205 B.n5 B.n4 10.955
R206 B.n7 B 9.97259
R207 B B.n12 8.48422
R208 B.n12 B 5.80515
R209 B.n7 B 4.31678
R210 B.n9 B.n8 3.65202
R211 B.n10 B.n9 1.46111
R212 B B.n6 0.149337
R213 a_27_368.t3 a_27_368.n5 871.107
R214 a_27_368.n3 a_27_368.n2 585
R215 a_27_368.n5 a_27_368.n4 585
R216 a_27_368.n1 a_27_368.n0 305.901
R217 a_27_368.n1 a_27_368.t5 303.455
R218 a_27_368.n3 a_27_368.n1 65.2554
R219 a_27_368.n5 a_27_368.n3 53.5848
R220 a_27_368.n4 a_27_368.t2 26.3844
R221 a_27_368.n4 a_27_368.t1 26.3844
R222 a_27_368.n2 a_27_368.t0 26.3844
R223 a_27_368.n2 a_27_368.t4 26.3844
R224 a_27_368.n0 a_27_368.t7 26.3844
R225 a_27_368.n0 a_27_368.t6 26.3844
C0 VPWR a_126_368# 0.379458f
C1 a_126_368# C_N 4.62e-19
C2 VPB B 0.144553f
C3 VPB VGND 0.010413f
C4 VPB A 0.147214f
C5 B VGND 0.098492f
C6 VPB Y 0.010084f
C7 A VGND 0.099797f
C8 B Y 0.217669f
C9 VPB VPWR 0.204685f
C10 VPB C_N 0.073208f
C11 Y VGND 0.920112f
C12 A Y 0.184591f
C13 B VPWR 0.025888f
C14 VPB a_126_368# 0.013547f
C15 VPWR VGND 0.124895f
C16 C_N VGND 0.018764f
C17 A VPWR 0.075615f
C18 A C_N 0.079326f
C19 B a_126_368# 0.163886f
C20 a_126_368# VGND 0.009012f
C21 Y VPWR 0.021363f
C22 Y C_N 2.4e-19
C23 A a_126_368# 0.056279f
C24 VPWR C_N 0.032278f
C25 Y a_126_368# 0.170951f
C26 VGND VNB 0.922761f
C27 C_N VNB 0.204546f
C28 VPWR VNB 0.729758f
C29 Y VNB 0.056122f
C30 A VNB 0.459472f
C31 B VNB 0.455587f
C32 VPB VNB 1.79899f
C33 a_126_368# VNB 0.008642f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nor3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3b_2 VNB VPB VPWR VGND A B Y C_N
X0 VPWR.t2 A.t0 a_495_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_495_368.t1 A.t1 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
X2 VGND.t3 C_N.t0 a_27_392.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1469 pd=1.16 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 VGND.t4 A.t2 Y.t6 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=2.09 as=0.1221 ps=1.07 w=0.74 l=0.15
X4 VGND.t1 a_27_392.t2 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2664 pd=1.46 as=0.10915 ps=1.035 w=0.74 l=0.15
X5 Y.t5 A.t3 VGND.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.3108 ps=1.58 w=0.74 l=0.15
X6 Y.t7 B.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2664 ps=1.46 w=0.74 l=0.15
X7 a_227_368.t3 B.t1 a_495_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Y.t0 a_27_392.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1469 ps=1.16 w=0.74 l=0.15
X9 a_495_368.t3 B.t2 a_227_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_227_368.t1 a_27_392.t4 Y.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VGND.t2 B.t3 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3108 pd=1.58 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VPWR.t0 C_N.t1 a_27_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X13 Y.t2 a_27_392.t5 a_227_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
R0 A.n0 A.t0 229
R1 A.n1 A.t1 226.809
R2 A.n1 A.t3 202.587
R3 A.n0 A.t2 196.013
R4 A.n5 A.n4 152
R5 A.n3 A.n2 152
R6 A.n4 A.n3 49.6611
R7 A.n4 A.n0 13.146
R8 A.n2 A 10.1214
R9 A A.n5 8.33538
R10 A.n5 A 5.95399
R11 A.n2 A 4.16794
R12 A.n3 A.n1 0.730803
R13 a_495_368.n1 a_495_368.n0 594.696
R14 a_495_368.n0 a_495_368.t2 26.3844
R15 a_495_368.n0 a_495_368.t1 26.3844
R16 a_495_368.t0 a_495_368.n1 26.3844
R17 a_495_368.n1 a_495_368.t3 26.3844
R18 VPWR.n4 VPWR.t1 342.878
R19 VPWR.n3 VPWR.t2 262.353
R20 VPWR.n12 VPWR.t0 251.91
R21 VPWR.n6 VPWR.n5 36.1417
R22 VPWR.n6 VPWR.n1 36.1417
R23 VPWR.n10 VPWR.n1 36.1417
R24 VPWR.n11 VPWR.n10 36.1417
R25 VPWR.n5 VPWR.n4 25.6005
R26 VPWR.n12 VPWR.n11 23.3417
R27 VPWR.n5 VPWR.n2 9.3005
R28 VPWR.n7 VPWR.n6 9.3005
R29 VPWR.n8 VPWR.n1 9.3005
R30 VPWR.n10 VPWR.n9 9.3005
R31 VPWR.n11 VPWR.n0 9.3005
R32 VPWR.n13 VPWR.n12 7.25439
R33 VPWR.n4 VPWR.n3 6.56006
R34 VPWR.n3 VPWR.n2 0.625092
R35 VPWR VPWR.n13 0.157727
R36 VPWR.n13 VPWR.n0 0.150046
R37 VPWR.n7 VPWR.n2 0.122949
R38 VPWR.n8 VPWR.n7 0.122949
R39 VPWR.n9 VPWR.n8 0.122949
R40 VPWR.n9 VPWR.n0 0.122949
R41 VPB.t3 VPB.t4 510.753
R42 VPB.t2 VPB.t1 510.753
R43 VPB VPB.t2 255.376
R44 VPB.t4 VPB.t5 229.839
R45 VPB.t6 VPB.t3 229.839
R46 VPB.t0 VPB.t6 229.839
R47 VPB.t1 VPB.t0 229.839
R48 C_N.n0 C_N.t0 267.267
R49 C_N.n0 C_N.t1 235.936
R50 C_N C_N.n0 153.745
R51 a_27_392.n0 a_27_392.t4 333.904
R52 a_27_392.t1 a_27_392.n3 294.481
R53 a_27_392.n1 a_27_392.t5 261.62
R54 a_27_392.n3 a_27_392.n2 201.159
R55 a_27_392.n2 a_27_392.t3 168.846
R56 a_27_392.n0 a_27_392.t2 154.24
R57 a_27_392.n3 a_27_392.t0 143.913
R58 a_27_392.n2 a_27_392.n1 48.2005
R59 a_27_392.n1 a_27_392.n0 2.19141
R60 VGND.n9 VGND.n8 185
R61 VGND.n7 VGND.n6 185
R62 VGND.n11 VGND.n1 185
R63 VGND.n13 VGND.n12 185
R64 VGND.n5 VGND.t4 167.632
R65 VGND.n20 VGND.n19 115.66
R66 VGND.n8 VGND.n7 90.8113
R67 VGND.n12 VGND.n11 71.3518
R68 VGND.n19 VGND.t3 39.3755
R69 VGND.n19 VGND.t0 35.7861
R70 VGND.n18 VGND.n17 29.6318
R71 VGND.n13 VGND.n10 26.0484
R72 VGND.n12 VGND.t6 22.7032
R73 VGND.n11 VGND.t1 22.7032
R74 VGND.n7 VGND.t5 22.7032
R75 VGND.n8 VGND.t2 22.7032
R76 VGND.n10 VGND.n9 19.4119
R77 VGND.n20 VGND.n18 18.824
R78 VGND.n18 VGND.n0 9.3005
R79 VGND.n17 VGND.n16 9.3005
R80 VGND.n15 VGND.n14 9.3005
R81 VGND.n10 VGND.n2 9.3005
R82 VGND.n4 VGND.n3 9.3005
R83 VGND.n14 VGND.n1 8.03554
R84 VGND.n21 VGND.n20 7.44972
R85 VGND.n6 VGND.n3 7.03676
R86 VGND.n6 VGND.n5 6.9507
R87 VGND.n9 VGND.n3 1.34787
R88 VGND.n17 VGND.n1 0.934807
R89 VGND.n5 VGND.n4 0.626959
R90 VGND.n14 VGND.n13 0.187361
R91 VGND VGND.n21 0.160299
R92 VGND.n21 VGND.n0 0.147507
R93 VGND.n4 VGND.n2 0.122949
R94 VGND.n15 VGND.n2 0.122949
R95 VGND.n16 VGND.n15 0.122949
R96 VGND.n16 VGND.n0 0.122949
R97 VNB.t2 VNB.t4 2286.61
R98 VNB.t1 VNB.t6 2009.45
R99 VNB.t3 VNB.t0 1316.54
R100 VNB VNB.t3 1154.86
R101 VNB.t4 VNB.t5 1108.66
R102 VNB.t0 VNB.t1 1027.82
R103 VNB.t6 VNB.t2 993.177
R104 Y.n4 Y.n0 367.49
R105 Y.n3 Y.n2 197.655
R106 Y Y.n5 110.162
R107 Y.n3 Y.n1 96.6047
R108 Y.n2 Y.t6 30.8113
R109 Y.n0 Y.t3 26.3844
R110 Y.n0 Y.t2 26.3844
R111 Y.n5 Y.t1 25.1356
R112 Y.n1 Y.t4 22.7032
R113 Y.n1 Y.t7 22.7032
R114 Y.n5 Y.t0 22.7032
R115 Y.n2 Y.t5 22.7032
R116 Y Y.n3 18.6672
R117 Y.n4 Y 12.4449
R118 Y Y.n4 4.62272
R119 B.n0 B.t1 226.809
R120 B.n2 B.t2 226.809
R121 B.n2 B.t0 198.204
R122 B.n1 B.t3 196.013
R123 B B.n0 192.208
R124 B B.n3 159.888
R125 B.n3 B.n2 54.0429
R126 B.n3 B.n1 6.57323
R127 B.n1 B.n0 5.11262
R128 a_227_368.n0 a_227_368.t3 383.305
R129 a_227_368.n0 a_227_368.t0 279.81
R130 a_227_368.n1 a_227_368.n0 213.232
R131 a_227_368.n1 a_227_368.t2 26.3844
R132 a_227_368.t1 a_227_368.n1 26.3844
C0 A VPB 0.076238f
C1 Y VGND 0.515785f
C2 VPWR VPB 0.150208f
C3 B A 0.058858f
C4 C_N VPWR 0.050846f
C5 Y VPB 0.007215f
C6 B VPWR 0.013856f
C7 C_N Y 0.007219f
C8 A VPWR 0.06979f
C9 B Y 0.103351f
C10 A Y 0.074766f
C11 VPWR Y 0.011358f
C12 VGND VPB 0.010087f
C13 C_N VGND 0.017353f
C14 B VGND 0.036085f
C15 C_N VPB 0.056645f
C16 A VGND 0.067592f
C17 B VPB 0.083043f
C18 VPWR VGND 0.079707f
C19 VGND VNB 0.610109f
C20 Y VNB 0.034173f
C21 VPWR VNB 0.499003f
C22 A VNB 0.262188f
C23 B VNB 0.234873f
C24 C_N VNB 0.155263f
C25 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2bb2a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2a_1 VNB VPB VPWR VGND B2 A2_N X B1 A1_N
X0 VPWR.t0 a_83_260.t3 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2278 pd=1.555 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_588_74.t1 a_233_384.t3 a_83_260.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X2 VGND.t1 a_83_260.t4 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.18895 pd=1.275 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_233_384.t0 A2_N.t0 a_253_94.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0768 ps=0.88 w=0.64 l=0.15
X4 VPWR.t3 A2_N.t1 a_233_384.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.4767 pd=1.975 as=0.1491 ps=1.195 w=0.84 l=0.15
X5 a_233_384.t1 A1_N.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1491 pd=1.195 as=0.2278 ps=1.555 w=0.84 l=0.15
X6 VGND.t0 B2.t0 a_588_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1216 pd=1.02 as=0.0896 ps=0.92 w=0.64 l=0.15
X7 a_83_260.t2 a_233_384.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1724 pd=1.36 as=0.4767 ps=1.975 w=0.84 l=0.15
X8 VPWR.t4 B1.t0 a_693_384.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X9 a_588_74.t2 B1.t1 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1216 ps=1.02 w=0.64 l=0.15
X10 a_253_94.t1 A1_N.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.18895 ps=1.275 w=0.64 l=0.15
X11 a_693_384.t1 B2.t1 a_83_260.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.1724 ps=1.36 w=1 l=0.15
R0 a_83_260.n2 a_83_260.n1 403.67
R1 a_83_260.n1 a_83_260.n0 357.144
R2 a_83_260.n0 a_83_260.t3 263.589
R3 a_83_260.n0 a_83_260.t4 203.339
R4 a_83_260.n1 a_83_260.t1 124.865
R5 a_83_260.n2 a_83_260.t2 46.9053
R6 a_83_260.t0 a_83_260.n2 33.9999
R7 X.n1 X 589.444
R8 X.n1 X.n0 585
R9 X.n2 X.n1 585
R10 X X.t0 205.94
R11 X.n1 X.t1 26.3844
R12 X X.n2 11.9116
R13 X X.n0 10.3116
R14 X X.n0 2.84494
R15 X.n2 X 1.24494
R16 VPWR.n8 VPWR.n2 585
R17 VPWR.n10 VPWR.n9 585
R18 VPWR.n7 VPWR.n6 585
R19 VPWR.n5 VPWR.t4 260.313
R20 VPWR.n16 VPWR.n1 225.375
R21 VPWR.n9 VPWR.n7 98.5005
R22 VPWR.n9 VPWR.n8 97.3279
R23 VPWR.n1 VPWR.t2 57.4585
R24 VPWR.n1 VPWR.t0 36.3318
R25 VPWR.n7 VPWR.t1 35.1791
R26 VPWR.n8 VPWR.t3 35.1791
R27 VPWR.n15 VPWR.n14 34.5909
R28 VPWR.n6 VPWR.n5 32.017
R29 VPWR.n16 VPWR.n15 19.2005
R30 VPWR.n4 VPWR.n3 9.3005
R31 VPWR.n12 VPWR.n11 9.3005
R32 VPWR.n14 VPWR.n13 9.3005
R33 VPWR.n15 VPWR.n0 9.3005
R34 VPWR.n17 VPWR.n16 7.43488
R35 VPWR.n10 VPWR.n4 5.37252
R36 VPWR.n11 VPWR.n2 4.51034
R37 VPWR.n14 VPWR.n2 1.85749
R38 VPWR.n11 VPWR.n10 0.995319
R39 VPWR.n5 VPWR.n3 0.541527
R40 VPWR.n6 VPWR.n4 0.199464
R41 VPWR VPWR.n17 0.160103
R42 VPWR.n17 VPWR.n0 0.1477
R43 VPWR.n12 VPWR.n3 0.122949
R44 VPWR.n13 VPWR.n12 0.122949
R45 VPWR.n13 VPWR.n0 0.122949
R46 VPB.t4 VPB.t2 656.317
R47 VPB.t1 VPB.t3 298.791
R48 VPB.t2 VPB.t0 260.485
R49 VPB.t3 VPB.t4 257.93
R50 VPB VPB.t1 257.93
R51 VPB.t0 VPB.t5 214.517
R52 a_233_384.n2 a_233_384.n1 640.929
R53 a_233_384.n0 a_233_384.t4 350.692
R54 a_233_384.n1 a_233_384.n0 252.549
R55 a_233_384.n1 a_233_384.t0 248.746
R56 a_233_384.n0 a_233_384.t3 128.534
R57 a_233_384.n2 a_233_384.t2 48.0779
R58 a_233_384.t1 a_233_384.n2 35.1791
R59 a_588_74.n0 a_588_74.t2 290.526
R60 a_588_74.t0 a_588_74.n0 26.2505
R61 a_588_74.n0 a_588_74.t1 26.2505
R62 VNB.t3 VNB.t2 2967.98
R63 VNB.t1 VNB.t5 1582.15
R64 VNB.t0 VNB.t4 1224.15
R65 VNB VNB.t1 1166.4
R66 VNB.t2 VNB.t0 993.177
R67 VNB.t5 VNB.t3 900.788
R68 VGND.n2 VGND.n0 212.868
R69 VGND.n2 VGND.n1 103.019
R70 VGND.n1 VGND.t3 49.4014
R71 VGND.n0 VGND.t0 39.3755
R72 VGND.n1 VGND.t1 37.994
R73 VGND.n0 VGND.t2 31.8755
R74 VGND VGND.n2 0.22228
R75 A2_N.n0 A2_N.t0 229.754
R76 A2_N.n0 A2_N.t1 205.922
R77 A2_N A2_N.n0 154.744
R78 a_253_94.t0 a_253_94.t1 45.0005
R79 A1_N.n0 A1_N.t0 219.31
R80 A1_N.n0 A1_N.t1 208.429
R81 A1_N A1_N.n0 153.28
R82 B2.n0 B2.t1 298.572
R83 B2.n0 B2.t0 181.554
R84 B2.n1 B2.n0 152
R85 B2 B2.n1 12.0247
R86 B2.n1 B2 6.59444
R87 B1.n0 B1.t0 306.741
R88 B1.n0 B1.t1 174.558
R89 B1 B1.n0 157.237
R90 a_693_384.t0 a_693_384.t1 53.1905
C0 VPB B2 0.040511f
C1 VGND X 0.090049f
C2 X B2 1.28e-20
C3 VPB B1 0.044048f
C4 VGND B2 0.01609f
C5 VPB A1_N 0.045631f
C6 VPB VPWR 0.151746f
C7 VGND B1 0.01647f
C8 VPB A2_N 0.044804f
C9 X A1_N 0.006642f
C10 B2 B1 0.09866f
C11 X VPWR 0.127235f
C12 VGND A1_N 0.014252f
C13 X A2_N 2.83e-19
C14 VGND VPWR 0.072821f
C15 VGND A2_N 0.005566f
C16 VPWR B2 0.025277f
C17 VPWR B1 0.043291f
C18 VPWR A1_N 0.022731f
C19 A1_N A2_N 0.095484f
C20 VPWR A2_N 0.016003f
C21 VPB X 0.016174f
C22 VGND VPB 0.009673f
C23 VGND VNB 0.534984f
C24 A2_N VNB 0.102833f
C25 A1_N VNB 0.107194f
C26 B1 VNB 0.176456f
C27 B2 VNB 0.116631f
C28 VPWR VNB 0.465606f
C29 X VNB 0.112581f
C30 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2bb2a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2a_2 VNB VPB VPWR VGND A1_N A2_N X B1 B2
X0 X.t1 a_201_392.t3 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.320525 ps=1.795 w=1.12 l=0.15
X1 a_270_48.t1 A2_N.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.23 as=0.253325 ps=1.58 w=0.84 l=0.15
X2 X.t3 a_201_392.t4 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1453 ps=1.155 w=0.74 l=0.15
X3 a_117_392.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X4 VPWR.t2 A1_N.t0 a_270_48.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.320525 pd=1.795 as=0.1638 ps=1.23 w=0.84 l=0.15
X5 VGND.t1 B1.t1 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VGND.t3 a_201_392.t5 X.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_201_392.t0 a_270_48.t3 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 a_27_74.t0 B2.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_201_392.t2 B2.t1 a_117_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t1 a_270_48.t4 a_201_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.253325 pd=1.58 as=0.18 ps=1.36 w=1 l=0.15
X11 VGND.t2 A1_N.t1 a_500_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1453 pd=1.155 as=0.0768 ps=0.88 w=0.64 l=0.15
X12 a_500_74.t1 A2_N.t1 a_270_48.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X13 VPWR.t4 a_201_392.t6 X.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 a_201_392.n4 a_201_392.n3 396.312
R1 a_201_392.n3 a_201_392.t0 287.161
R2 a_201_392.n0 a_201_392.t6 239.589
R3 a_201_392.n2 a_201_392.t3 238.858
R4 a_201_392.n1 a_201_392.t4 181.554
R5 a_201_392.n0 a_201_392.t5 181.554
R6 a_201_392.n3 a_201_392.n2 166.607
R7 a_201_392.n1 a_201_392.n0 62.8066
R8 a_201_392.n4 a_201_392.t2 41.3705
R9 a_201_392.t1 a_201_392.n4 29.5505
R10 a_201_392.n2 a_201_392.n1 2.19141
R11 VPWR.n2 VPWR.n1 646.715
R12 VPWR.n6 VPWR.n5 622.431
R13 VPWR.n4 VPWR.t4 266.272
R14 VPWR.n14 VPWR.t0 251.91
R15 VPWR.n5 VPWR.t2 79.7386
R16 VPWR.n1 VPWR.t3 69.185
R17 VPWR.n5 VPWR.t5 41.3484
R18 VPWR.n13 VPWR.n12 36.1417
R19 VPWR.n8 VPWR.n7 36.1417
R20 VPWR.n1 VPWR.t1 35.2195
R21 VPWR.n12 VPWR.n2 28.9887
R22 VPWR.n14 VPWR.n13 20.3299
R23 VPWR.n8 VPWR.n2 16.5652
R24 VPWR.n7 VPWR.n6 14.024
R25 VPWR.n6 VPWR.n4 9.42285
R26 VPWR.n7 VPWR.n3 9.3005
R27 VPWR.n9 VPWR.n8 9.3005
R28 VPWR.n10 VPWR.n2 9.3005
R29 VPWR.n12 VPWR.n11 9.3005
R30 VPWR.n13 VPWR.n0 9.3005
R31 VPWR.n15 VPWR.n14 9.3005
R32 VPWR.n4 VPWR.n3 0.526566
R33 VPWR.n9 VPWR.n3 0.122949
R34 VPWR.n10 VPWR.n9 0.122949
R35 VPWR.n11 VPWR.n10 0.122949
R36 VPWR.n11 VPWR.n0 0.122949
R37 VPWR.n15 VPWR.n0 0.122949
R38 VPWR VPWR.n15 0.0617245
R39 X.n2 X 589.639
R40 X.n2 X.n0 585
R41 X.n3 X.n2 585
R42 X X.n1 159.54
R43 X.n2 X.t0 26.3844
R44 X.n2 X.t1 26.3844
R45 X.n1 X.t2 22.7032
R46 X.n1 X.t3 22.7032
R47 X X.n3 12.4295
R48 X X.n0 10.7599
R49 X X.n0 2.96862
R50 X.n3 X 1.29905
R51 VPB.t2 VPB.t6 377.957
R52 VPB.t1 VPB.t3 329.435
R53 VPB.t3 VPB.t2 275.807
R54 VPB.t4 VPB.t1 260.485
R55 VPB VPB.t0 260.485
R56 VPB.t6 VPB.t5 229.839
R57 VPB.t0 VPB.t4 214.517
R58 A2_N.n0 A2_N.t1 284.38
R59 A2_N.n0 A2_N.t0 205.922
R60 A2_N A2_N.n0 155.298
R61 a_270_48.n2 a_270_48.n1 639.619
R62 a_270_48.n1 a_270_48.t2 270.447
R63 a_270_48.n0 a_270_48.t3 246.429
R64 a_270_48.n0 a_270_48.t4 231.167
R65 a_270_48.n1 a_270_48.n0 152
R66 a_270_48.t0 a_270_48.n2 45.7326
R67 a_270_48.n2 a_270_48.t1 45.7326
R68 VGND.n2 VGND.t3 178.791
R69 VGND.n4 VGND.n3 115.29
R70 VGND.n12 VGND.n11 115.066
R71 VGND.n3 VGND.t4 44.2236
R72 VGND.n5 VGND.n1 36.1417
R73 VGND.n9 VGND.n1 36.1417
R74 VGND.n10 VGND.n9 36.1417
R75 VGND.n3 VGND.t2 30.0005
R76 VGND.n12 VGND.n10 24.4711
R77 VGND.n11 VGND.t0 22.7032
R78 VGND.n11 VGND.t1 22.7032
R79 VGND.n5 VGND.n4 18.4476
R80 VGND.n10 VGND.n0 9.3005
R81 VGND.n9 VGND.n8 9.3005
R82 VGND.n7 VGND.n1 9.3005
R83 VGND.n6 VGND.n5 9.3005
R84 VGND.n13 VGND.n12 7.19894
R85 VGND.n4 VGND.n2 6.98414
R86 VGND.n6 VGND.n2 0.550243
R87 VGND VGND.n13 0.156997
R88 VGND.n13 VGND.n0 0.150766
R89 VGND.n7 VGND.n6 0.122949
R90 VGND.n8 VGND.n7 0.122949
R91 VGND.n8 VGND.n0 0.122949
R92 VNB.t1 VNB.t4 2309.71
R93 VNB.t3 VNB.t6 1304.99
R94 VNB.t0 VNB.t1 1154.86
R95 VNB VNB.t2 1143.31
R96 VNB.t6 VNB.t5 993.177
R97 VNB.t2 VNB.t0 993.177
R98 VNB.t4 VNB.t3 900.788
R99 B1.n0 B1.t1 252.248
R100 B1.n0 B1.t0 235.159
R101 B1 B1.n0 161.697
R102 a_117_392.t0 a_117_392.t1 53.1905
R103 A1_N.n0 A1_N.t1 274.649
R104 A1_N.n0 A1_N.t0 204.225
R105 A1_N A1_N.n0 157.625
R106 a_27_74.n0 a_27_74.t2 318.83
R107 a_27_74.n0 a_27_74.t1 34.0546
R108 a_27_74.t0 a_27_74.n0 22.7032
R109 B2.n0 B2.t0 252.248
R110 B2.n0 B2.t1 236.983
R111 B2 B2.n0 157.43
R112 a_500_74.t0 a_500_74.t1 45.0005
C0 A1_N VPB 0.051612f
C1 X VPB 0.00599f
C2 VGND VPB 0.010443f
C3 A2_N VPWR 0.009592f
C4 A1_N VPWR 0.011844f
C5 VGND B1 0.018446f
C6 VGND B2 0.018647f
C7 X VPWR 0.1544f
C8 VGND VPWR 0.082548f
C9 VPB B1 0.046675f
C10 A2_N A1_N 0.095087f
C11 VPB B2 0.040383f
C12 A2_N X 2.16e-19
C13 VPB VPWR 0.14493f
C14 B1 B2 0.091816f
C15 A2_N VGND 0.006192f
C16 A1_N X 0.002239f
C17 B1 VPWR 0.055202f
C18 A1_N VGND 0.018535f
C19 B2 VPWR 0.022104f
C20 X VGND 0.150106f
C21 A2_N VPB 0.050766f
C22 VGND VNB 0.572731f
C23 X VNB 0.030015f
C24 A1_N VNB 0.11327f
C25 A2_N VNB 0.13385f
C26 VPWR VNB 0.506976f
C27 B2 VNB 0.101655f
C28 B1 VNB 0.150332f
C29 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2bb2a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2a_4 VNB VPB VPWR VGND X B2 B1 A2_N A1_N
X0 a_41_392.t2 B2.t0 a_310_392.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X1 a_310_392.t4 B2.t1 a_41_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X2 a_41_392.t0 B1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X3 VPWR.t2 a_476_48.t3 a_310_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2583 pd=1.73 as=0.1554 ps=1.21 w=0.84 l=0.15
X4 X.t7 a_310_392.t6 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.2709 ps=1.73 w=1.12 l=0.15
X5 a_27_74.t1 a_476_48.t4 a_310_392.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2048 pd=1.92 as=0.1008 ps=0.955 w=0.64 l=0.15
X6 X.t3 a_310_392.t7 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.15725 pd=1.165 as=0.1693 ps=1.23 w=0.74 l=0.15
X7 a_476_48.t2 A2_N.t0 VPWR.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2583 ps=1.73 w=0.84 l=0.15
X8 a_27_74.t5 B2.t2 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0992 pd=0.95 as=0.112 ps=0.99 w=0.64 l=0.15
X9 VGND.t1 B1.t1 a_27_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.1824 ps=1.85 w=0.64 l=0.15
X10 X.t6 a_310_392.t8 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.196 ps=1.47 w=1.12 l=0.15
X11 VPWR.t0 B1.t2 a_41_392.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X12 VGND.t2 A1_N.t0 a_835_94.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1693 pd=1.23 as=0.0768 ps=0.88 w=0.64 l=0.15
X13 VGND.t7 a_310_392.t9 X.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t6 a_310_392.t10 X.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.1708 ps=1.425 w=1.12 l=0.15
X15 VGND.t3 B2.t3 a_27_74.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 VPWR.t5 a_310_392.t11 X.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.224 ps=1.52 w=1.12 l=0.15
X17 X.t1 a_310_392.t12 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 a_310_392.t2 a_476_48.t5 VPWR.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1554 pd=1.21 as=0.2478 ps=2.27 w=0.84 l=0.15
X19 a_310_392.t3 a_476_48.t6 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1008 pd=0.955 as=0.0992 ps=0.95 w=0.64 l=0.15
X20 a_27_74.t2 B1.t3 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1344 ps=1.06 w=0.64 l=0.15
X21 a_835_94.t1 A2_N.t1 a_476_48.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1952 ps=1.89 w=0.64 l=0.15
X22 VPWR.t4 A1_N.t1 a_476_48.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2709 pd=1.73 as=0.126 ps=1.14 w=0.84 l=0.15
X23 VGND.t5 a_310_392.t13 X.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.15725 ps=1.165 w=0.74 l=0.15
R0 B2.n4 B2.t2 247.136
R1 B2.n1 B2.t3 244.214
R2 B2.n1 B2.t1 215.805
R3 B2.n3 B2.t0 212.883
R4 B2.n5 B2.n4 152
R5 B2.n2 B2.n0 152
R6 B2.n3 B2.n2 42.3581
R7 B2.n2 B2.n1 20.449
R8 B2.n5 B2.n0 13.1884
R9 B2.n4 B2.n3 7.30353
R10 B2 B2.n5 3.87929
R11 B2.n0 B2 1.55202
R12 a_310_392.n12 a_310_392.n11 585
R13 a_310_392.n13 a_310_392.n12 404.834
R14 a_310_392.n10 a_310_392.n2 402.053
R15 a_310_392.n4 a_310_392.t10 329.902
R16 a_310_392.n0 a_310_392.t8 261.62
R17 a_310_392.n1 a_310_392.t11 261.62
R18 a_310_392.n7 a_310_392.t6 261.62
R19 a_310_392.n12 a_310_392.n10 225.416
R20 a_310_392.n4 a_310_392.t9 174.323
R21 a_310_392.n5 a_310_392.n3 165.189
R22 a_310_392.n7 a_310_392.t7 156.431
R23 a_310_392.n1 a_310_392.t13 154.24
R24 a_310_392.n0 a_310_392.t12 154.24
R25 a_310_392.n9 a_310_392.n8 152
R26 a_310_392.n6 a_310_392.n3 152
R27 a_310_392.n0 a_310_392.n4 100.052
R28 a_310_392.n11 a_310_392.t0 50.4231
R29 a_310_392.n8 a_310_392.n6 49.6611
R30 a_310_392.n5 a_310_392.n0 44.549
R31 a_310_392.n11 a_310_392.t2 36.3517
R32 a_310_392.n2 a_310_392.t1 32.813
R33 a_310_392.n13 a_310_392.t5 29.5505
R34 a_310_392.t4 a_310_392.n13 29.5505
R35 a_310_392.n1 a_310_392.n5 28.4823
R36 a_310_392.n2 a_310_392.t3 26.2505
R37 a_310_392.n6 a_310_392.n1 21.1793
R38 a_310_392.n9 a_310_392.n3 13.1884
R39 a_310_392.n8 a_310_392.n7 10.955
R40 a_310_392.n10 a_310_392.n9 8.53383
R41 a_41_392.t2 a_41_392.n1 395.264
R42 a_41_392.n1 a_41_392.t3 294.043
R43 a_41_392.n1 a_41_392.n0 189.115
R44 a_41_392.n0 a_41_392.t1 29.5505
R45 a_41_392.n0 a_41_392.t0 29.5505
R46 VPB.t5 VPB.t1 515.861
R47 VPB.t2 VPB.t9 316.668
R48 VPB.t0 VPB.t10 316.668
R49 VPB VPB.t11 293.683
R50 VPB.t9 VPB.t6 280.914
R51 VPB.t1 VPB.t0 265.591
R52 VPB.t6 VPB.t8 255.376
R53 VPB.t8 VPB.t7 232.393
R54 VPB.t10 VPB.t2 229.839
R55 VPB.t4 VPB.t5 229.839
R56 VPB.t3 VPB.t4 229.839
R57 VPB.t11 VPB.t3 229.839
R58 B1.n1 B1.t0 263.762
R59 B1.n4 B1.t2 263.762
R60 B1.n1 B1.t3 189.606
R61 B1.n6 B1.n5 184.864
R62 B1.n5 B1.t1 183.161
R63 B1.n2 B1 159.906
R64 B1.n3 B1.n0 152
R65 B1.n3 B1.n2 49.6611
R66 B1.n5 B1.n4 11.6853
R67 B1.n2 B1.n1 10.955
R68 B1.n6 B1.n0 8.53383
R69 B1.n4 B1.n3 5.11262
R70 B1 B1.n6 2.88677
R71 B1 B1.n0 0.627951
R72 VPWR.n19 VPWR.n5 786.356
R73 VPWR.n21 VPWR.t3 783.755
R74 VPWR.n13 VPWR.n12 742.111
R75 VPWR.n27 VPWR.n1 331.5
R76 VPWR.n8 VPWR.t6 264.7
R77 VPWR.n10 VPWR.n9 221.766
R78 VPWR.n12 VPWR.t4 65.6672
R79 VPWR.n5 VPWR.t9 55.1136
R80 VPWR.n5 VPWR.t2 55.1136
R81 VPWR.n25 VPWR.n2 36.1417
R82 VPWR.n26 VPWR.n25 36.1417
R83 VPWR.n20 VPWR.n19 36.1417
R84 VPWR.n18 VPWR.n6 36.1417
R85 VPWR.n14 VPWR.n11 36.1417
R86 VPWR.n9 VPWR.t7 35.1791
R87 VPWR.n12 VPWR.t8 34.0942
R88 VPWR.n27 VPWR.n26 30.1181
R89 VPWR.n1 VPWR.t1 29.5505
R90 VPWR.n1 VPWR.t0 29.5505
R91 VPWR.n21 VPWR.n2 28.9887
R92 VPWR.n9 VPWR.t5 26.3844
R93 VPWR.n21 VPWR.n20 18.4476
R94 VPWR.n11 VPWR.n10 17.6946
R95 VPWR.n28 VPWR.n27 13.7273
R96 VPWR.n19 VPWR.n18 11.2946
R97 VPWR.n11 VPWR.n7 9.3005
R98 VPWR.n15 VPWR.n14 9.3005
R99 VPWR.n16 VPWR.n6 9.3005
R100 VPWR.n18 VPWR.n17 9.3005
R101 VPWR.n19 VPWR.n4 9.3005
R102 VPWR.n20 VPWR.n3 9.3005
R103 VPWR.n22 VPWR.n21 9.3005
R104 VPWR.n23 VPWR.n2 9.3005
R105 VPWR.n25 VPWR.n24 9.3005
R106 VPWR.n26 VPWR.n0 9.3005
R107 VPWR.n13 VPWR.n6 8.28285
R108 VPWR.n10 VPWR.n8 6.96039
R109 VPWR.n14 VPWR.n13 3.01226
R110 VPWR.n8 VPWR.n7 0.594857
R111 VPWR VPWR.n28 0.163644
R112 VPWR.n28 VPWR.n0 0.144205
R113 VPWR.n15 VPWR.n7 0.122949
R114 VPWR.n16 VPWR.n15 0.122949
R115 VPWR.n17 VPWR.n16 0.122949
R116 VPWR.n17 VPWR.n4 0.122949
R117 VPWR.n4 VPWR.n3 0.122949
R118 VPWR.n22 VPWR.n3 0.122949
R119 VPWR.n23 VPWR.n22 0.122949
R120 VPWR.n24 VPWR.n23 0.122949
R121 VPWR.n24 VPWR.n0 0.122949
R122 a_476_48.n8 a_476_48.n7 636.634
R123 a_476_48.n7 a_476_48.t0 241.835
R124 a_476_48.n1 a_476_48.t6 233.924
R125 a_476_48.n5 a_476_48.t3 211.643
R126 a_476_48.n2 a_476_48.t4 196.013
R127 a_476_48.n3 a_476_48.t5 195.21
R128 a_476_48.n1 a_476_48.n0 165.77
R129 a_476_48.n4 a_476_48.n0 152
R130 a_476_48.n6 a_476_48.n5 152
R131 a_476_48.n5 a_476_48.n4 49.6611
R132 a_476_48.n2 a_476_48.n1 38.7066
R133 a_476_48.t1 a_476_48.n8 35.1791
R134 a_476_48.n8 a_476_48.t2 35.1791
R135 a_476_48.n6 a_476_48.n0 13.1884
R136 a_476_48.n4 a_476_48.n3 10.955
R137 a_476_48.n7 a_476_48.n6 9.30959
R138 a_476_48.n3 a_476_48.n2 2.19141
R139 X.n4 X.n2 261.149
R140 X.n4 X.n3 210.702
R141 X.n0 X 197.607
R142 X.n1 X.n0 185
R143 X.n6 X.n5 96.0198
R144 X.n2 X.t4 35.1791
R145 X.n2 X.t7 35.1791
R146 X.n0 X.t3 34.8654
R147 X.n0 X.t0 34.0546
R148 X.n6 X.n4 33.231
R149 X.n3 X.t5 27.2639
R150 X.n3 X.t6 26.3844
R151 X.n5 X.t2 22.7032
R152 X.n5 X.t1 22.7032
R153 X X.n6 18.8389
R154 X.n7 X 17.6005
R155 X X.n7 8.0005
R156 X.n7 X.n1 1.74595
R157 X.n1 X 1.74595
R158 a_27_74.t1 a_27_74.n3 254.286
R159 a_27_74.n1 a_27_74.t3 191.244
R160 a_27_74.n3 a_27_74.n2 185
R161 a_27_74.n1 a_27_74.n0 98.4905
R162 a_27_74.n3 a_27_74.n1 32.207
R163 a_27_74.n2 a_27_74.t0 29.063
R164 a_27_74.n2 a_27_74.t5 29.063
R165 a_27_74.n0 a_27_74.t4 26.2505
R166 a_27_74.n0 a_27_74.t2 26.2505
R167 VNB.t1 VNB.t2 2725.46
R168 VNB.t5 VNB.t11 1478.22
R169 VNB.t11 VNB.t8 1328.08
R170 VNB.t4 VNB.t3 1316.54
R171 VNB.t8 VNB.t9 1154.86
R172 VNB.t6 VNB.t7 1154.86
R173 VNB VNB.t4 1143.31
R174 VNB.t0 VNB.t1 1074.02
R175 VNB.t7 VNB.t0 1062.47
R176 VNB.t9 VNB.t10 993.177
R177 VNB.t3 VNB.t6 993.177
R178 VNB.t2 VNB.t5 900.788
R179 VGND.n24 VGND.n23 206.333
R180 VGND.n8 VGND.n7 205.752
R181 VGND.n21 VGND.n2 205.171
R182 VGND.n11 VGND.n10 200.171
R183 VGND.n6 VGND.t7 161.433
R184 VGND.n10 VGND.t2 45.938
R185 VGND.n10 VGND.t8 42.3486
R186 VGND.n2 VGND.t3 39.3755
R187 VGND.n23 VGND.t0 39.3755
R188 VGND.n23 VGND.t1 39.3755
R189 VGND.n15 VGND.n4 36.1417
R190 VGND.n16 VGND.n15 36.1417
R191 VGND.n17 VGND.n16 36.1417
R192 VGND.n17 VGND.n1 36.1417
R193 VGND.n11 VGND.n4 34.6358
R194 VGND.n7 VGND.t6 34.0546
R195 VGND.n11 VGND.n9 33.1299
R196 VGND.n22 VGND.n21 31.2476
R197 VGND.n2 VGND.t4 26.2505
R198 VGND.n7 VGND.t5 22.7032
R199 VGND.n24 VGND.n22 19.2005
R200 VGND.n9 VGND.n8 17.6946
R201 VGND.n21 VGND.n1 16.1887
R202 VGND.n22 VGND.n0 9.3005
R203 VGND.n21 VGND.n20 9.3005
R204 VGND.n19 VGND.n1 9.3005
R205 VGND.n18 VGND.n17 9.3005
R206 VGND.n16 VGND.n3 9.3005
R207 VGND.n15 VGND.n14 9.3005
R208 VGND.n13 VGND.n4 9.3005
R209 VGND.n9 VGND.n5 9.3005
R210 VGND.n25 VGND.n24 7.43488
R211 VGND.n8 VGND.n6 6.96039
R212 VGND.n12 VGND.n11 4.62059
R213 VGND.n6 VGND.n5 0.594857
R214 VGND.n12 VGND.n5 0.184273
R215 VGND.n13 VGND.n12 0.184273
R216 VGND VGND.n25 0.160103
R217 VGND.n25 VGND.n0 0.1477
R218 VGND.n14 VGND.n13 0.122949
R219 VGND.n14 VGND.n3 0.122949
R220 VGND.n18 VGND.n3 0.122949
R221 VGND.n19 VGND.n18 0.122949
R222 VGND.n20 VGND.n19 0.122949
R223 VGND.n20 VGND.n0 0.122949
R224 A2_N.n0 A2_N.t0 205.922
R225 A2_N.n0 A2_N.t1 204.048
R226 A2_N A2_N.n0 154.377
R227 A1_N.n0 A1_N.t1 205.922
R228 A1_N.n0 A1_N.t0 204.048
R229 A1_N A1_N.n0 155.126
R230 a_835_94.t0 a_835_94.t1 45.0005
C0 B2 VGND 0.028012f
C1 VPWR X 0.384921f
C2 B2 VPWR 0.013222f
C3 VPB A1_N 0.037927f
C4 VPWR VGND 0.129855f
C5 A2_N X 2.68e-19
C6 A2_N VGND 0.005918f
C7 A1_N X 0.001916f
C8 VPWR A2_N 0.005602f
C9 A1_N VGND 0.014323f
C10 VPWR A1_N 0.008166f
C11 A2_N A1_N 0.093395f
C12 VPB B1 0.100247f
C13 VPB X 0.013755f
C14 VPB B2 0.093104f
C15 VPB VGND 0.015264f
C16 VPB VPWR 0.229995f
C17 B1 B2 0.088579f
C18 B1 VGND 0.034198f
C19 B2 X 6.37e-20
C20 X VGND 0.280971f
C21 VPB A2_N 0.035261f
C22 B1 VPWR 0.032136f
C23 VGND VNB 0.877532f
C24 X VNB 0.038851f
C25 A1_N VNB 0.107488f
C26 A2_N VNB 0.109958f
C27 VPWR VNB 0.709385f
C28 B2 VNB 0.220678f
C29 B1 VNB 0.310246f
C30 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2bb2ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2ai_1 VNB VPB VPWR VGND Y B2 A1_N B1 A2_N
X0 a_131_383.t1 A1_N.t0 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2898 ps=2.37 w=0.84 l=0.15
X1 a_397_74.t1 B1.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_114_74.t0 A1_N.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 a_131_383.t2 A2_N.t0 a_114_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0768 ps=0.88 w=0.64 l=0.15
X4 VGND.t0 B2.t0 a_397_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 a_397_74.t2 a_131_383.t3 Y.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VPWR.t1 A2_N.t1 a_131_383.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.371 pd=1.865 as=0.126 ps=1.14 w=0.84 l=0.15
X7 a_490_368.t1 B2.t1 Y.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t2 B1.t1 a_490_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1848 ps=1.45 w=1.12 l=0.15
X9 Y.t2 a_131_383.t4 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.371 ps=1.865 w=1.12 l=0.15
R0 A1_N.n0 A1_N.t0 262.923
R1 A1_N.n0 A1_N.t1 174.558
R2 A1_N A1_N.n0 157.237
R3 VPWR.n5 VPWR.t3 404.202
R4 VPWR.n1 VPWR.t2 265.072
R5 VPWR.n3 VPWR.n2 148.514
R6 VPWR.n2 VPWR.t1 81.8078
R7 VPWR.n2 VPWR.t0 69.1735
R8 VPWR.n4 VPWR.n3 31.624
R9 VPWR.n5 VPWR.n4 18.824
R10 VPWR.n4 VPWR.n0 9.3005
R11 VPWR.n6 VPWR.n5 9.3005
R12 VPWR.n3 VPWR.n1 4.12254
R13 VPWR.n1 VPWR.n0 0.237326
R14 VPWR.n6 VPWR.n0 0.122949
R15 VPWR VPWR.n6 0.0617245
R16 a_131_383.n2 a_131_383.n1 339.887
R17 a_131_383.n0 a_131_383.t4 229
R18 a_131_383.n1 a_131_383.n0 208.233
R19 a_131_383.n0 a_131_383.t3 196.013
R20 a_131_383.n1 a_131_383.t2 167.921
R21 a_131_383.t0 a_131_383.n2 35.1791
R22 a_131_383.n2 a_131_383.t1 35.1791
R23 VPB.t0 VPB.t4 457.125
R24 VPB VPB.t2 296.238
R25 VPB.t3 VPB.t1 245.161
R26 VPB.t4 VPB.t3 229.839
R27 VPB.t2 VPB.t0 229.839
R28 B1.n0 B1.t1 256.428
R29 B1.n0 B1.t0 196.178
R30 B1 B1.n0 156.462
R31 VGND.n1 VGND.n0 229.38
R32 VGND.n1 VGND.t2 158.5
R33 VGND.n0 VGND.t1 22.7032
R34 VGND.n0 VGND.t0 22.7032
R35 VGND VGND.n1 0.100891
R36 a_397_74.n0 a_397_74.t1 395.452
R37 a_397_74.n0 a_397_74.t2 34.0546
R38 a_397_74.t0 a_397_74.n0 22.7032
R39 VNB.t3 VNB.t4 2367.45
R40 VNB.t4 VNB.t0 1154.86
R41 VNB VNB.t2 1143.31
R42 VNB.t0 VNB.t1 993.177
R43 VNB.t2 VNB.t3 900.788
R44 a_114_74.t0 a_114_74.t1 45.0005
R45 A2_N.n0 A2_N.t1 286.95
R46 A2_N A2_N.n0 164.024
R47 A2_N.n0 A2_N.t0 162.274
R48 B2.n0 B2.t1 264.298
R49 B2.n0 B2.t0 204.048
R50 B2 B2.n0 156.4
R51 Y Y.n0 588.516
R52 Y.n2 Y.n0 585
R53 Y.n1 Y.n0 585
R54 Y.n1 Y.t1 221.077
R55 Y.n0 Y.t0 26.3844
R56 Y.n0 Y.t2 26.3844
R57 Y Y.n2 6.33017
R58 Y Y.n1 5.76753
R59 Y.n2 Y 4.07962
R60 a_490_368.t0 a_490_368.t1 58.0451
C0 VPWR Y 0.17791f
C1 Y VGND 0.038334f
C2 VPWR VGND 0.059461f
C3 VPB B2 0.033263f
C4 VPB B1 0.04372f
C5 A1_N VPB 0.051178f
C6 B2 B1 0.107731f
C7 A2_N VPB 0.041751f
C8 Y VPB 0.007318f
C9 VPWR VPB 0.125844f
C10 VGND VPB 0.007335f
C11 Y B2 0.058408f
C12 VPWR B2 0.021451f
C13 A1_N A2_N 0.099529f
C14 Y B1 0.005681f
C15 VGND B2 0.014304f
C16 VPWR B1 0.046406f
C17 VGND B1 0.01532f
C18 VPWR A1_N 0.03939f
C19 A2_N Y 0.001601f
C20 A1_N VGND 0.047354f
C21 VPWR A2_N 0.018449f
C22 A2_N VGND 0.022389f
C23 VGND VNB 0.469982f
C24 Y VNB 0.019767f
C25 A2_N VNB 0.12636f
C26 A1_N VNB 0.179486f
C27 VPWR VNB 0.429241f
C28 B1 VNB 0.168215f
C29 B2 VNB 0.104589f
C30 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2bb2ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2ai_2 VNB VPB VPWR VGND B2 A2_N Y B1 A1_N
X0 VPWR.t5 A1_N.t0 a_133_387.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2709 pd=1.665 as=0.1723 ps=1.33 w=0.84 l=0.15
X1 VPWR.t7 a_133_387.t6 Y.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1764 ps=1.435 w=1.12 l=0.15
X2 a_796_368.t1 B2.t0 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t0 B2.t1 a_796_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t2 B1.t0 a_796_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_133_387.t3 A2_N.t0 a_134_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1136 pd=0.995 as=0.0896 ps=0.92 w=0.64 l=0.15
X6 a_796_368.t3 B1.t1 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2184 ps=1.51 w=1.12 l=0.15
X7 a_518_74.t5 a_133_387.t7 Y.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_134_74.t3 A1_N.t1 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2272 ps=1.99 w=0.64 l=0.15
X9 a_518_74.t3 B1.t2 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10915 ps=1.035 w=0.74 l=0.15
X10 a_518_74.t1 B2.t2 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 Y.t3 a_133_387.t8 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.2709 ps=1.665 w=1.12 l=0.15
X12 Y.t5 a_133_387.t9 a_518_74.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 VPWR.t0 A2_N.t1 a_133_387.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.232925 pd=1.555 as=0.126 ps=1.14 w=0.84 l=0.15
X14 VGND.t2 B1.t3 a_518_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1147 ps=1.05 w=0.74 l=0.15
X15 a_133_387.t1 A2_N.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1723 pd=1.33 as=0.232925 ps=1.555 w=0.84 l=0.15
X16 a_134_74.t0 A2_N.t3 a_133_387.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1136 ps=0.995 w=0.64 l=0.15
X17 VGND.t0 B2.t3 a_518_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1221 ps=1.07 w=0.74 l=0.15
X18 a_133_387.t4 A1_N.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.3801 ps=2.86 w=0.84 l=0.15
X19 VGND.t4 A1_N.t3 a_134_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 A1_N.n2 A1_N.n0 404.599
R1 A1_N.n1 A1_N.t2 235.944
R2 A1_N.n0 A1_N.t3 219.416
R3 A1_N.n1 A1_N.t1 211.309
R4 A1_N.n0 A1_N.t0 205.922
R5 A1_N A1_N.n1 156.147
R6 A1_N A1_N.n2 2.78311
R7 A1_N.n2 A1_N 1.80332
R8 a_133_387.n6 a_133_387.n0 625.284
R9 a_133_387.n7 a_133_387.n6 585
R10 a_133_387.n3 a_133_387.t8 539.038
R11 a_133_387.n5 a_133_387.n3 268.512
R12 a_133_387.n1 a_133_387.t6 246.892
R13 a_133_387.n5 a_133_387.n4 201.129
R14 a_133_387.n1 a_133_387.t7 182.317
R15 a_133_387.n2 a_133_387.t9 179.947
R16 a_133_387.n2 a_133_387.n1 65.5841
R17 a_133_387.n0 a_133_387.t5 57.5459
R18 a_133_387.n6 a_133_387.n5 52.5622
R19 a_133_387.n4 a_133_387.t2 40.313
R20 a_133_387.n0 a_133_387.t1 38.0274
R21 a_133_387.t0 a_133_387.n7 35.1791
R22 a_133_387.n7 a_133_387.t4 35.1791
R23 a_133_387.n3 a_133_387.n2 32.3972
R24 a_133_387.n4 a_133_387.t3 26.2505
R25 VPWR.n17 VPWR.t4 865.899
R26 VPWR.n15 VPWR.n2 670.581
R27 VPWR.n8 VPWR.n7 315.349
R28 VPWR.n6 VPWR.t2 265.139
R29 VPWR.n10 VPWR.n5 233.226
R30 VPWR.n5 VPWR.t5 91.8365
R31 VPWR.n2 VPWR.t1 55.1136
R32 VPWR.n2 VPWR.t0 55.1136
R33 VPWR.n14 VPWR.n3 36.1417
R34 VPWR.n7 VPWR.t3 36.0585
R35 VPWR.n16 VPWR.n15 35.0123
R36 VPWR.n7 VPWR.t7 32.5407
R37 VPWR.n5 VPWR.t6 30.3299
R38 VPWR.n10 VPWR.n3 25.977
R39 VPWR.n9 VPWR.n8 25.6005
R40 VPWR.n10 VPWR.n9 21.4593
R41 VPWR.n17 VPWR.n16 20.7064
R42 VPWR.n15 VPWR.n14 12.424
R43 VPWR.n9 VPWR.n4 9.3005
R44 VPWR.n11 VPWR.n10 9.3005
R45 VPWR.n12 VPWR.n3 9.3005
R46 VPWR.n14 VPWR.n13 9.3005
R47 VPWR.n15 VPWR.n1 9.3005
R48 VPWR.n16 VPWR.n0 9.3005
R49 VPWR.n18 VPWR.n17 9.3005
R50 VPWR.n8 VPWR.n6 7.03002
R51 VPWR.n6 VPWR.n4 0.172977
R52 VPWR.n11 VPWR.n4 0.122949
R53 VPWR.n12 VPWR.n11 0.122949
R54 VPWR.n13 VPWR.n12 0.122949
R55 VPWR.n13 VPWR.n1 0.122949
R56 VPWR.n1 VPWR.n0 0.122949
R57 VPWR.n18 VPWR.n0 0.122949
R58 VPWR VPWR.n18 0.0617245
R59 VPB.t7 VPB.t8 354.974
R60 VPB.t1 VPB.t2 316.668
R61 VPB VPB.t6 301.344
R62 VPB.t2 VPB.t7 278.361
R63 VPB.t9 VPB.t5 275.807
R64 VPB.t8 VPB.t9 237.5
R65 VPB.t3 VPB.t4 229.839
R66 VPB.t0 VPB.t3 229.839
R67 VPB.t5 VPB.t0 229.839
R68 VPB.t6 VPB.t1 229.839
R69 Y.n2 Y.n1 392.608
R70 Y.n2 Y.n0 200.391
R71 Y.n4 Y.n3 185
R72 Y.n0 Y.t4 29.0228
R73 Y.n0 Y.t3 26.3844
R74 Y.n1 Y.t1 26.3844
R75 Y.n1 Y.t0 26.3844
R76 Y.n3 Y.t2 22.7032
R77 Y.n3 Y.t5 22.7032
R78 Y Y.n4 15.5107
R79 Y Y.n2 6.24004
R80 Y.n4 Y 0.883259
R81 B2.n0 B2.t0 261.62
R82 B2.n1 B2.t1 261.62
R83 B2 B2.n2 158.788
R84 B2.n1 B2.t2 156.431
R85 B2.n0 B2.t3 156.431
R86 B2.n2 B2.n0 43.0884
R87 B2.n2 B2.n1 22.6399
R88 a_796_368.n1 a_796_368.n0 553.654
R89 a_796_368.n0 a_796_368.t0 26.3844
R90 a_796_368.n0 a_796_368.t3 26.3844
R91 a_796_368.n1 a_796_368.t2 26.3844
R92 a_796_368.t1 a_796_368.n1 26.3844
R93 B1.n1 B1.t1 250.909
R94 B1.n0 B1.t0 250.909
R95 B1 B1.n1 247.954
R96 B1.n1 B1.t3 220.113
R97 B1.n0 B1.t2 220.113
R98 B1.n2 B1.n0 158.995
R99 B1 B1.n2 4.16794
R100 B1.n2 B1 1.12991
R101 A2_N.n0 A2_N.t0 244.798
R102 A2_N.n1 A2_N.t3 242.607
R103 A2_N.n2 A2_N.t2 199.349
R104 A2_N.n0 A2_N.t1 181.821
R105 A2_N A2_N.n2 154.102
R106 A2_N.n1 A2_N.n0 71.5702
R107 A2_N.n2 A2_N.n1 1.46111
R108 a_134_74.n1 a_134_74.n0 344.798
R109 a_134_74.n0 a_134_74.t2 26.2505
R110 a_134_74.n0 a_134_74.t0 26.2505
R111 a_134_74.t1 a_134_74.n1 26.2505
R112 a_134_74.n1 a_134_74.t3 26.2505
R113 VNB.t6 VNB.t8 2286.61
R114 VNB VNB.t7 1374.28
R115 VNB.t1 VNB.t0 1166.4
R116 VNB.t4 VNB.t3 1154.86
R117 VNB.t3 VNB.t2 1108.66
R118 VNB.t9 VNB.t4 1062.47
R119 VNB.t2 VNB.t5 1027.82
R120 VNB.t8 VNB.t9 993.177
R121 VNB.t0 VNB.t6 993.177
R122 VNB.t7 VNB.t1 993.177
R123 a_518_74.t4 a_518_74.n3 286.658
R124 a_518_74.n1 a_518_74.t3 186.786
R125 a_518_74.n1 a_518_74.n0 96.0666
R126 a_518_74.n3 a_518_74.n2 89.0748
R127 a_518_74.n3 a_518_74.n1 64.7247
R128 a_518_74.n2 a_518_74.t5 27.5681
R129 a_518_74.n0 a_518_74.t0 26.7573
R130 a_518_74.n0 a_518_74.t1 26.7573
R131 a_518_74.n2 a_518_74.t2 22.7032
R132 VGND.n12 VGND.t4 243.743
R133 VGND.n7 VGND.n4 209.677
R134 VGND.n6 VGND.n5 206.333
R135 VGND.n18 VGND.t5 155.126
R136 VGND.n10 VGND.n3 36.1417
R137 VGND.n11 VGND.n10 36.1417
R138 VGND.n16 VGND.n1 36.1417
R139 VGND.n17 VGND.n16 36.1417
R140 VGND.n5 VGND.t2 34.0546
R141 VGND.n12 VGND.n1 30.1181
R142 VGND.n6 VGND.n3 27.1064
R143 VGND.n4 VGND.t3 24.3248
R144 VGND.n4 VGND.t0 23.514
R145 VGND.n5 VGND.t1 22.7032
R146 VGND.n12 VGND.n11 22.5887
R147 VGND.n18 VGND.n17 18.4476
R148 VGND.n19 VGND.n18 9.3005
R149 VGND.n8 VGND.n3 9.3005
R150 VGND.n10 VGND.n9 9.3005
R151 VGND.n11 VGND.n2 9.3005
R152 VGND.n13 VGND.n12 9.3005
R153 VGND.n14 VGND.n1 9.3005
R154 VGND.n16 VGND.n15 9.3005
R155 VGND.n17 VGND.n0 9.3005
R156 VGND.n7 VGND.n6 6.49467
R157 VGND.n8 VGND.n7 0.585239
R158 VGND.n9 VGND.n8 0.122949
R159 VGND.n9 VGND.n2 0.122949
R160 VGND.n13 VGND.n2 0.122949
R161 VGND.n14 VGND.n13 0.122949
R162 VGND.n15 VGND.n14 0.122949
R163 VGND.n15 VGND.n0 0.122949
R164 VGND.n19 VGND.n0 0.122949
R165 VGND VGND.n19 0.0617245
C0 B2 VPB 0.0559f
C1 VGND VPB 0.009793f
C2 A1_N VPB 0.120167f
C3 B2 VPWR 0.011835f
C4 VGND VPWR 0.095552f
C5 A2_N VPB 0.092108f
C6 A1_N VPWR 0.247418f
C7 B1 VPB 0.075577f
C8 Y VPB 0.007432f
C9 A2_N VPWR 0.01821f
C10 VGND B2 0.0294f
C11 B1 VPWR 0.052465f
C12 Y VPWR 0.238959f
C13 VGND A1_N 0.064063f
C14 VGND A2_N 0.012283f
C15 B1 B2 0.199837f
C16 VGND B1 0.03104f
C17 B2 Y 0.024088f
C18 A1_N A2_N 0.166374f
C19 VGND Y 0.012423f
C20 A1_N Y 0.006837f
C21 B1 A2_N 8.67e-20
C22 A2_N Y 4.04e-19
C23 B1 Y 0.122979f
C24 VPB VPWR 0.183491f
C25 VGND VNB 0.721282f
C26 Y VNB 0.011711f
C27 A2_N VNB 0.216584f
C28 A1_N VNB 0.339001f
C29 B2 VNB 0.199528f
C30 B1 VNB 0.264768f
C31 VPWR VNB 0.592533f
C32 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21a_1 VNB VPB VPWR VGND X A2 B1 A1
X0 VGND.t1 A2.t0 a_320_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 VPWR.t1 a_83_244.t3 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.334825 pd=1.765 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VGND.t0 a_83_244.t4 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_320_74.t2 A1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 a_320_74.t0 B1.t0 a_83_244.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X5 a_376_387.t1 A2.t1 a_83_244.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.1703 ps=1.355 w=1 l=0.15
X6 a_83_244.t1 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1703 pd=1.355 as=0.334825 ps=1.765 w=0.84 l=0.15
X7 VPWR.t2 A1.t1 a_376_387.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.21 ps=1.42 w=1 l=0.15
R0 A2.n0 A2.t0 266.707
R1 A2.n0 A2.t1 231.629
R2 A2 A2.n0 159.452
R3 a_320_74.n0 a_320_74.t2 300.832
R4 a_320_74.n0 a_320_74.t1 26.2505
R5 a_320_74.t0 a_320_74.n0 26.2505
R6 VGND.n1 VGND.n0 213.268
R7 VGND.n1 VGND.t0 143.971
R8 VGND.n0 VGND.t2 26.2505
R9 VGND.n0 VGND.t1 26.2505
R10 VGND VGND.n1 0.242346
R11 VNB.t1 VNB.t0 2379
R12 VNB VNB.t1 1143.31
R13 VNB.t2 VNB.t3 993.177
R14 VNB.t0 VNB.t2 993.177
R15 a_83_244.n2 a_83_244.n1 380.702
R16 a_83_244.n0 a_83_244.t3 279.293
R17 a_83_244.n1 a_83_244.t0 178.959
R18 a_83_244.n0 a_83_244.t4 171.913
R19 a_83_244.n1 a_83_244.n0 152
R20 a_83_244.t2 a_83_244.n2 44.5535
R21 a_83_244.n2 a_83_244.t1 35.1791
R22 X.n1 X 589.85
R23 X.n1 X.n0 585
R24 X.n2 X.n1 585
R25 X.t1 X.n3 279.738
R26 X.n4 X.t1 279.738
R27 X.n1 X.t0 26.3844
R28 X.n4 X 16.6405
R29 X.n2 X 12.9944
R30 X.n3 X 12.5445
R31 X.n0 X 11.249
R32 X.n3 X 6.4005
R33 X.n0 X 3.10353
R34 X X.n4 2.3045
R35 X X.n2 1.35808
R36 VPWR.n4 VPWR.n3 599.198
R37 VPWR.n1 VPWR.n0 589.914
R38 VPWR.n2 VPWR.n0 585
R39 VPWR.n5 VPWR.t2 260.019
R40 VPWR.n3 VPWR.n2 51.5957
R41 VPWR.n2 VPWR.t0 35.1791
R42 VPWR.n1 VPWR.t1 22.3123
R43 VPWR.n3 VPWR.n1 19.9985
R44 VPWR.n5 VPWR.n4 15.6988
R45 VPWR.n4 VPWR.n0 8.15625
R46 VPWR VPWR.n5 0.267443
R47 VPB.t1 VPB.t0 406.048
R48 VPB.t3 VPB.t2 291.13
R49 VPB.t0 VPB.t3 257.93
R50 VPB VPB.t1 257.93
R51 A1.n0 A1.t1 263.459
R52 A1.n0 A1.t0 213.118
R53 A1 A1.n0 156.462
R54 B1.n0 B1.t0 221.575
R55 B1.n0 B1.t1 205.922
R56 B1 B1.n0 157.923
R57 a_376_387.t0 a_376_387.t1 82.7405
C0 B1 VPB 0.054477f
C1 B1 X 0.00111f
C2 A1 VPWR 0.054557f
C3 VGND VPB 0.007554f
C4 A2 VPB 0.046063f
C5 B1 VPWR 0.014938f
C6 VGND X 0.079552f
C7 A2 X 2.97e-20
C8 A1 B1 5.11e-19
C9 VGND VPWR 0.048911f
C10 A2 VPWR 0.026028f
C11 A1 VGND 0.017826f
C12 A2 A1 0.097805f
C13 B1 VGND 0.013448f
C14 A2 B1 0.074603f
C15 A2 VGND 0.017095f
C16 VPB X 0.012691f
C17 VPB VPWR 0.09628f
C18 A1 VPB 0.051741f
C19 X VPWR 0.098555f
C20 VGND VNB 0.393445f
C21 B1 VNB 0.142106f
C22 A1 VNB 0.181119f
C23 A2 VNB 0.110427f
C24 VPWR VNB 0.343911f
C25 X VNB 0.110492f
C26 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21a_2 VNB VPB VPWR VGND A1 A2 B1 X
X0 X.t3 a_244_368.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2931 ps=1.66 w=1.12 l=0.15
X1 X.t1 a_244_368.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X2 a_244_368.t0 A2.t0 a_160_368.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X3 a_160_368.t0 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X4 a_244_368.t1 B1.t0 a_54_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.12025 ps=1.065 w=0.74 l=0.15
X5 VPWR.t3 B1.t1 a_244_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2931 pd=1.66 as=0.21 ps=1.42 w=1 l=0.15
X6 VGND.t3 A1.t1 a_54_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1702 pd=1.2 as=0.2627 ps=2.19 w=0.74 l=0.15
X7 a_54_74.t2 A2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.1702 ps=1.2 w=0.74 l=0.15
X8 VPWR.t0 a_244_368.t5 X.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VGND.t0 a_244_368.t6 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_244_368.n0 a_244_368.t6 282.762
R1 a_244_368.n2 a_244_368.t3 272.574
R2 a_244_368.n4 a_244_368.n3 268.12
R3 a_244_368.n1 a_244_368.t5 260.012
R4 a_244_368.n0 a_244_368.t4 152.637
R5 a_244_368.n3 a_244_368.n2 152
R6 a_244_368.n3 a_244_368.t1 143.201
R7 a_244_368.n2 a_244_368.n1 56.2338
R8 a_244_368.t0 a_244_368.n4 53.1905
R9 a_244_368.n4 a_244_368.t2 29.5505
R10 a_244_368.n1 a_244_368.n0 7.03871
R11 VPWR.n4 VPWR.t0 358.962
R12 VPWR.n9 VPWR.t2 256.668
R13 VPWR.n3 VPWR.n2 221.764
R14 VPWR.n2 VPWR.t3 66.9805
R15 VPWR.n7 VPWR.n1 36.1417
R16 VPWR.n8 VPWR.n7 36.1417
R17 VPWR.n2 VPWR.t1 33.8013
R18 VPWR.n3 VPWR.n1 21.4593
R19 VPWR.n10 VPWR.n9 16.4534
R20 VPWR.n5 VPWR.n1 9.3005
R21 VPWR.n7 VPWR.n6 9.3005
R22 VPWR.n8 VPWR.n0 9.3005
R23 VPWR.n4 VPWR.n3 6.88087
R24 VPWR.n9 VPWR.n8 4.14168
R25 VPWR.n5 VPWR.n4 0.513127
R26 VPWR.n6 VPWR.n5 0.122949
R27 VPWR.n6 VPWR.n0 0.122949
R28 VPWR.n10 VPWR.n0 0.122949
R29 VPWR VPWR.n10 0.0617245
R30 X X.n0 232.231
R31 X.n3 X.n2 185
R32 X.n2 X.n1 185
R33 X.n0 X.t2 26.3844
R34 X.n0 X.t3 26.3844
R35 X.n2 X.t0 22.7032
R36 X.n2 X.t1 22.7032
R37 X.n1 X 12.6066
R38 X X.n3 9.50353
R39 X.n3 X 4.84898
R40 X.n1 X 1.74595
R41 VPB VPB.t3 370.296
R42 VPB.t4 VPB.t2 352.42
R43 VPB.t0 VPB.t4 291.13
R44 VPB.t2 VPB.t1 229.839
R45 VPB.t3 VPB.t0 214.517
R46 VGND.n7 VGND.n6 198.593
R47 VGND.n2 VGND.t0 178.799
R48 VGND.n1 VGND.t1 149.984
R49 VGND.n6 VGND.t2 39.7302
R50 VGND.n5 VGND.n4 36.1417
R51 VGND.n6 VGND.t3 34.8654
R52 VGND.n7 VGND.n5 33.5064
R53 VGND.n4 VGND.n1 22.9652
R54 VGND.n5 VGND.n0 9.3005
R55 VGND.n4 VGND.n3 9.3005
R56 VGND.n2 VGND.n1 6.74444
R57 VGND.n8 VGND.n7 4.77522
R58 VGND.n3 VGND.n2 0.585372
R59 VGND VGND.n8 0.237916
R60 VGND.n8 VGND.n0 0.192318
R61 VGND.n3 VGND.n0 0.122949
R62 VNB.t4 VNB.t1 2609.97
R63 VNB VNB.t3 1616.8
R64 VNB.t3 VNB.t2 1408.92
R65 VNB.t2 VNB.t4 1097.11
R66 VNB.t1 VNB.t0 993.177
R67 A2.n0 A2.t0 266.44
R68 A2.n0 A2.t1 178.34
R69 A2 A2.n0 158.788
R70 a_160_368.t0 a_160_368.t1 53.1905
R71 A1.n0 A1.t0 246.31
R72 A1.n0 A1.t1 154.24
R73 A1.n1 A1.n0 97.0285
R74 A1 A1.n1 10.4704
R75 A1.n1 A1 5.75841
R76 B1.n0 B1.t1 266.44
R77 B1.n0 B1.t0 178.34
R78 B1 B1.n0 158.746
R79 a_54_74.t0 a_54_74.n0 288.976
R80 a_54_74.n0 a_54_74.t2 30.0005
R81 a_54_74.n0 a_54_74.t1 22.7032
C0 VPWR X 0.229443f
C1 VPB A2 0.031519f
C2 VPWR VGND 0.070156f
C3 A1 A2 0.081856f
C4 B1 VPWR 0.014055f
C5 X VGND 0.168711f
C6 B1 X 8.31e-19
C7 B1 VGND 0.014685f
C8 VPB VPWR 0.157617f
C9 A1 VPWR 0.050364f
C10 VPB X 0.011329f
C11 VPB VGND 0.017878f
C12 A2 VPWR 0.017503f
C13 VPB B1 0.036446f
C14 A1 VGND 0.01847f
C15 A2 VGND 0.015369f
C16 A2 B1 0.080588f
C17 VPB A1 0.055163f
C18 VGND VNB 0.534676f
C19 X VNB 0.040572f
C20 VPWR VNB 0.45911f
C21 B1 VNB 0.114438f
C22 A2 VNB 0.106469f
C23 A1 VNB 0.194835f
C24 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21a_4 VNB VPB VPWR VGND A1 A2 B1 X
X0 VPWR.t2 A1.t0 a_116_387.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.185 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X1 X.t7 a_216_387.t6 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 a_116_387.t1 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X3 a_27_125.t5 A2.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1136 ps=0.995 w=0.64 l=0.15
X4 a_216_387.t1 B1.t0 a_27_125.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 a_216_387.t0 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1596 pd=1.22 as=0.185 ps=1.39 w=0.84 l=0.15
X6 X.t3 a_216_387.t7 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X7 VGND.t4 a_216_387.t8 X.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 X.t5 a_216_387.t9 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11655 ps=1.055 w=0.74 l=0.15
X9 VPWR.t4 a_216_387.t10 X.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t6 a_216_387.t11 X.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_116_387.t3 A2.t1 a_216_387.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X12 VGND.t0 A2.t2 a_27_125.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.07 as=0.0896 ps=0.92 w=0.64 l=0.15
X13 a_216_387.t2 A2.t3 a_116_387.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X14 a_27_125.t3 B1.t2 a_216_387.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2336 pd=2.01 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 VGND.t2 A1.t2 a_27_125.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1136 pd=0.995 as=0.1824 ps=1.85 w=0.64 l=0.15
X16 VPWR.t5 a_216_387.t12 X.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X17 X.t0 a_216_387.t13 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2807 ps=1.7 w=1.12 l=0.15
X18 a_27_125.t1 A1.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1376 ps=1.07 w=0.64 l=0.15
X19 VPWR.t7 B1.t3 a_216_387.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2807 pd=1.7 as=0.1596 ps=1.22 w=0.84 l=0.15
R0 A1.t3 A1.t2 930.26
R1 A1.t2 A1.t1 450.938
R2 A1.n0 A1.t0 231.629
R3 A1.n0 A1.t3 184.768
R4 A1 A1.n0 156.394
R5 a_116_387.n1 a_116_387.n0 570.744
R6 a_116_387.n0 a_116_387.t3 39.4005
R7 a_116_387.n1 a_116_387.t1 39.4005
R8 a_116_387.n0 a_116_387.t2 29.5505
R9 a_116_387.t0 a_116_387.n1 29.5505
R10 VPWR.n15 VPWR.n3 618.939
R11 VPWR.n5 VPWR.n4 608.067
R12 VPWR.n6 VPWR.t4 264.243
R13 VPWR.n21 VPWR.t1 252.982
R14 VPWR.n8 VPWR.n7 221.766
R15 VPWR.n4 VPWR.t6 69.6583
R16 VPWR.n4 VPWR.t7 60.9767
R17 VPWR.n3 VPWR.t0 44.56
R18 VPWR.n3 VPWR.t2 43.6235
R19 VPWR.n19 VPWR.n1 36.1417
R20 VPWR.n20 VPWR.n19 36.1417
R21 VPWR.n14 VPWR.n13 36.1417
R22 VPWR.n7 VPWR.t3 35.1791
R23 VPWR.n7 VPWR.t5 35.1791
R24 VPWR.n9 VPWR.n5 35.0123
R25 VPWR.n15 VPWR.n1 28.9887
R26 VPWR.n21 VPWR.n20 20.7064
R27 VPWR.n15 VPWR.n14 18.4476
R28 VPWR.n9 VPWR.n8 17.6946
R29 VPWR.n10 VPWR.n9 9.3005
R30 VPWR.n11 VPWR.n5 9.3005
R31 VPWR.n13 VPWR.n12 9.3005
R32 VPWR.n14 VPWR.n2 9.3005
R33 VPWR.n16 VPWR.n15 9.3005
R34 VPWR.n17 VPWR.n1 9.3005
R35 VPWR.n19 VPWR.n18 9.3005
R36 VPWR.n20 VPWR.n0 9.3005
R37 VPWR.n22 VPWR.n21 9.3005
R38 VPWR.n8 VPWR.n6 6.96039
R39 VPWR.n13 VPWR.n5 1.12991
R40 VPWR.n10 VPWR.n6 0.594857
R41 VPWR.n11 VPWR.n10 0.122949
R42 VPWR.n12 VPWR.n11 0.122949
R43 VPWR.n12 VPWR.n2 0.122949
R44 VPWR.n16 VPWR.n2 0.122949
R45 VPWR.n17 VPWR.n16 0.122949
R46 VPWR.n18 VPWR.n17 0.122949
R47 VPWR.n18 VPWR.n0 0.122949
R48 VPWR.n22 VPWR.n0 0.122949
R49 VPWR VPWR.n22 0.0617245
R50 VPB.t9 VPB.t8 372.849
R51 VPB.t7 VPB.t5 280.914
R52 VPB.t3 VPB.t0 275.807
R53 VPB.t0 VPB.t9 270.7
R54 VPB VPB.t2 257.93
R55 VPB.t4 VPB.t3 255.376
R56 VPB.t2 VPB.t1 255.376
R57 VPB.t5 VPB.t6 229.839
R58 VPB.t8 VPB.t7 229.839
R59 VPB.t1 VPB.t4 229.839
R60 a_216_387.n16 a_216_387.n15 388.046
R61 a_216_387.n15 a_216_387.n14 300.514
R62 a_216_387.n9 a_216_387.t12 261.62
R63 a_216_387.n10 a_216_387.t13 261.62
R64 a_216_387.n3 a_216_387.t10 205.387
R65 a_216_387.n5 a_216_387.t7 205.387
R66 a_216_387.n11 a_216_387.n10 173.179
R67 a_216_387.n7 a_216_387.n6 163.606
R68 a_216_387.n3 a_216_387.t11 161.177
R69 a_216_387.n4 a_216_387.t9 154.24
R70 a_216_387.n1 a_216_387.t6 154.24
R71 a_216_387.n2 a_216_387.t8 154.24
R72 a_216_387.n1 a_216_387.n0 152
R73 a_216_387.n8 a_216_387.n7 152
R74 a_216_387.n13 a_216_387.n12 150.891
R75 a_216_387.n15 a_216_387.n13 74.9181
R76 a_216_387.n14 a_216_387.t5 51.5957
R77 a_216_387.n6 a_216_387.n2 37.9763
R78 a_216_387.n14 a_216_387.t0 37.5243
R79 a_216_387.n1 a_216_387.n9 37.246
R80 a_216_387.n4 a_216_387.n3 33.0264
R81 a_216_387.n16 a_216_387.t3 29.5505
R82 a_216_387.t2 a_216_387.n16 29.5505
R83 a_216_387.n10 a_216_387.n1 28.4823
R84 a_216_387.n12 a_216_387.t4 26.2505
R85 a_216_387.n12 a_216_387.t1 26.2505
R86 a_216_387.n6 a_216_387.n5 13.146
R87 a_216_387.n9 a_216_387.n8 12.4157
R88 a_216_387.n8 a_216_387.n2 11.6853
R89 a_216_387.n7 a_216_387.n0 11.6058
R90 a_216_387.n11 a_216_387.n0 11.6058
R91 a_216_387.n5 a_216_387.n4 7.14124
R92 a_216_387.n13 a_216_387.n11 4.0965
R93 VGND.n16 VGND.n2 214.868
R94 VGND.n19 VGND.n18 214.422
R95 VGND.n6 VGND.n5 202.535
R96 VGND.n7 VGND.t6 170.607
R97 VGND.n10 VGND.t5 144.959
R98 VGND.n2 VGND.t0 41.2505
R99 VGND.n2 VGND.t1 39.3755
R100 VGND.n18 VGND.t2 39.3755
R101 VGND.n12 VGND.n11 36.1417
R102 VGND.n12 VGND.n1 36.1417
R103 VGND.n11 VGND.n10 33.1299
R104 VGND.n18 VGND.t3 27.188
R105 VGND.n17 VGND.n16 27.1064
R106 VGND.n5 VGND.t7 25.9464
R107 VGND.n6 VGND.n4 25.6005
R108 VGND.n5 VGND.t4 25.1356
R109 VGND.n10 VGND.n4 20.3299
R110 VGND.n16 VGND.n1 20.3299
R111 VGND.n19 VGND.n17 18.824
R112 VGND.n17 VGND.n0 9.3005
R113 VGND.n16 VGND.n15 9.3005
R114 VGND.n14 VGND.n1 9.3005
R115 VGND.n13 VGND.n12 9.3005
R116 VGND.n11 VGND.n3 9.3005
R117 VGND.n10 VGND.n9 9.3005
R118 VGND.n8 VGND.n4 9.3005
R119 VGND.n20 VGND.n19 7.43488
R120 VGND.n7 VGND.n6 6.26985
R121 VGND.n8 VGND.n7 0.733933
R122 VGND VGND.n20 0.160103
R123 VGND.n20 VGND.n0 0.1477
R124 VGND.n9 VGND.n8 0.122949
R125 VGND.n9 VGND.n3 0.122949
R126 VGND.n13 VGND.n3 0.122949
R127 VGND.n14 VGND.n13 0.122949
R128 VGND.n15 VGND.n14 0.122949
R129 VGND.n15 VGND.n0 0.122949
R130 X.n5 X.n3 261.149
R131 X.n5 X.n4 210.702
R132 X.n2 X.n1 158.627
R133 X.n2 X.n0 98.1558
R134 X.n6 X.n2 47.0802
R135 X.n4 X.t2 26.3844
R136 X.n4 X.t3 26.3844
R137 X.n3 X.t1 26.3844
R138 X.n3 X.t0 26.3844
R139 X.n0 X.t4 22.7032
R140 X.n0 X.t5 22.7032
R141 X.n1 X.t6 22.7032
R142 X.n1 X.t7 22.7032
R143 X X.n6 16.1396
R144 X.n6 X.n5 2.13383
R145 VNB.t5 VNB.t9 2471.39
R146 VNB.t1 VNB.t2 1339.63
R147 VNB.t3 VNB.t4 1166.4
R148 VNB VNB.t3 1143.31
R149 VNB.t8 VNB.t7 1074.02
R150 VNB.t7 VNB.t6 993.177
R151 VNB.t9 VNB.t8 993.177
R152 VNB.t0 VNB.t5 993.177
R153 VNB.t2 VNB.t0 993.177
R154 VNB.t4 VNB.t1 993.177
R155 A2.n0 A2.t1 211.179
R156 A2.n2 A2.t3 207.529
R157 A2.n3 A2.t0 160.667
R158 A2.n0 A2.t2 160.667
R159 A2 A2.n1 160.597
R160 A2 A2.n3 156.394
R161 A2.n2 A2.n1 48.9308
R162 A2.n1 A2.n0 13.146
R163 A2.n3 A2.n2 0.730803
R164 a_27_125.n1 a_27_125.t3 312.486
R165 a_27_125.t2 a_27_125.n3 186.942
R166 a_27_125.n3 a_27_125.n2 100.754
R167 a_27_125.n1 a_27_125.n0 89.3175
R168 a_27_125.n3 a_27_125.n1 60.671
R169 a_27_125.n0 a_27_125.t0 26.2505
R170 a_27_125.n0 a_27_125.t1 26.2505
R171 a_27_125.n2 a_27_125.t4 26.2505
R172 a_27_125.n2 a_27_125.t5 26.2505
R173 B1.n4 B1.t3 192.776
R174 B1.n1 B1.t1 181.821
R175 B1.n1 B1.t0 168.701
R176 B1.n3 B1.t2 160.667
R177 B1.n5 B1.n4 152
R178 B1.n2 B1.n0 152
R179 B1.n3 B1.n2 37.9763
R180 B1.n2 B1.n1 16.7975
R181 B1.n5 B1.n0 16.4231
R182 B1.n4 B1.n3 11.6853
R183 B1 B1.n5 4.10616
R184 B1.n0 B1 2.6571
C0 VPB X 0.013999f
C1 VPB A2 0.076691f
C2 A1 X 1.06e-19
C3 VPB VGND 0.009705f
C4 A1 A2 0.144992f
C5 VPB VPWR 0.178525f
C6 A1 VGND 0.093608f
C7 X VGND 0.296014f
C8 A1 VPWR 0.042184f
C9 VPB B1 0.094226f
C10 A2 VGND 0.023451f
C11 VPWR X 0.44459f
C12 A2 VPWR 0.011489f
C13 A1 B1 0.07292f
C14 VPWR VGND 0.097724f
C15 B1 X 0.001704f
C16 B1 VGND 0.011396f
C17 VPWR B1 0.030394f
C18 VPB A1 0.080689f
C19 VGND VNB 0.744028f
C20 X VNB 0.04606f
C21 B1 VNB 0.189902f
C22 VPWR VNB 0.615471f
C23 A2 VNB 0.173963f
C24 A1 VNB 0.424116f
C25 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o21ai_1 VNB VPB VPWR VGND Y B1 A2 A1
X0 a_27_74.t2 A2.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3361 ps=1.68 w=0.74 l=0.15
X1 VGND.t0 A1.t0 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.3361 pd=1.68 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 Y.t1 B1.t0 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t2 A2.t1 a_162_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2828 pd=1.625 as=0.1512 ps=1.39 w=1.12 l=0.15
X4 a_162_368.t1 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.4648 ps=3.07 w=1.12 l=0.15
X5 VPWR.t0 B1.t1 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2828 ps=1.625 w=1.12 l=0.15
R0 A2.n0 A2.t1 245.972
R1 A2.n0 A2.t0 215.178
R2 A2 A2.n0 155.423
R3 VGND VGND.n0 157.105
R4 VGND.n0 VGND.t1 61.6221
R5 VGND.n0 VGND.t0 61.6221
R6 a_27_74.n0 a_27_74.t1 406.166
R7 a_27_74.t0 a_27_74.n0 22.7032
R8 a_27_74.n0 a_27_74.t2 22.7032
R9 VNB.t1 VNB.t2 2101.84
R10 VNB VNB.t1 1143.31
R11 VNB.t2 VNB.t0 993.177
R12 A1.n0 A1.t1 296.673
R13 A1 A1.n0 175.466
R14 A1.n0 A1.t0 154.24
R15 B1.n0 B1.t1 250.909
R16 B1.n0 B1.t0 220.113
R17 B1.n1 B1.n0 152
R18 B1.n1 B1 8.63306
R19 B1 B1.n1 5.65631
R20 Y Y.n0 586.952
R21 Y.n2 Y.n0 585
R22 Y.n1 Y.n0 585
R23 Y.n1 Y.t1 286.558
R24 Y.n0 Y.t0 62.4425
R25 Y.n0 Y.t2 26.3844
R26 Y Y.n2 3.5127
R27 Y Y.n1 3.2005
R28 Y.n2 Y 2.26391
R29 a_162_368.t0 a_162_368.t1 47.4916
R30 VPB VPB.t2 375.404
R31 VPB.t1 VPB.t0 334.543
R32 VPB.t2 VPB.t1 214.517
R33 VPWR.n0 VPWR.t1 274.452
R34 VPWR.n0 VPWR.t0 255.597
R35 VPWR VPWR.n0 0.157417
C0 B1 VPWR 0.059725f
C1 B1 Y 0.086644f
C2 B1 VPB 0.043237f
C3 VPWR Y 0.256431f
C4 B1 VGND 0.011733f
C5 VPWR VPB 0.095144f
C6 VPWR VGND 0.041766f
C7 VPWR A1 0.032709f
C8 B1 A2 0.091515f
C9 Y VPB 0.011264f
C10 Y VGND 0.058046f
C11 Y A1 0.060002f
C12 VGND VPB 0.007526f
C13 VPWR A2 0.005067f
C14 VPB A1 0.047622f
C15 Y A2 0.125472f
C16 VGND A1 0.015265f
C17 VPB A2 0.037595f
C18 VGND A2 0.013236f
C19 A1 A2 0.048992f
C20 VGND VNB 0.319948f
C21 Y VNB 0.072494f
C22 VPWR VNB 0.34592f
C23 B1 VNB 0.153851f
C24 A2 VNB 0.114332f
C25 A1 VNB 0.183536f
C26 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__o2bb2ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2ai_4 VNB VPB VPWR VGND Y A2_N A1_N B1 B2
X0 VPWR.t8 A2_N.t0 a_114_368.t7 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_857_74.t10 a_114_368.t12 Y.t11 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_114_368.t6 A2_N.t1 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_857_74.t9 a_114_368.t13 Y.t10 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t9 B1.t0 a_857_74.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VPWR.t6 A2_N.t2 a_114_368.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_114_368.t4 A2_N.t3 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VGND.t11 B2.t0 a_857_74.t11 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t0 A1_N.t0 a_114_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_114_368.t1 A1_N.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_114_368.t8 A2_N.t4 a_27_74.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_857_74.t4 B1.t1 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VPWR.t3 A1_N.t2 a_114_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t0 A1_N.t3 a_27_74.t7 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 Y.t9 a_114_368.t14 a_857_74.t8 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_857_74.t6 B2.t1 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 a_1215_368.t3 B1.t2 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_27_74.t2 A2_N.t5 a_114_368.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.13875 pd=1.115 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VPWR.t2 B1.t3 a_1215_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t8 a_114_368.t15 a_857_74.t7 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X20 a_1215_368.t1 B1.t4 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_114_368.t11 A2_N.t6 a_27_74.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.13875 ps=1.115 w=0.74 l=0.15
X22 VPWR.t11 B1.t5 a_1215_368.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_27_74.t6 A1_N.t4 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_1215_368.t7 B2.t2 Y.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 Y.t7 a_114_368.t16 VPWR.t15 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 Y.t1 B2.t3 a_1215_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 VGND.t4 B2.t4 a_857_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VPWR.t14 a_114_368.t17 Y.t6 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 VPWR.t13 a_114_368.t18 Y.t5 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_1215_368.t5 B2.t5 Y.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X31 a_114_368.t3 A1_N.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X32 a_857_74.t0 B1.t6 VGND.t7 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X33 Y.t3 B2.t6 a_1215_368.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X34 a_27_74.t5 A1_N.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X35 VGND.t3 A1_N.t7 a_27_74.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1073 ps=1.03 w=0.74 l=0.15
X36 a_27_74.t0 A2_N.t7 a_114_368.t9 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.12025 ps=1.065 w=0.74 l=0.15
X37 a_857_74.t3 B2.t7 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X38 VGND.t6 B1.t7 a_857_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X39 Y.t4 a_114_368.t19 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A2_N.n0 A2_N.t0 303.699
R1 A2_N.n1 A2_N.t1 226.809
R2 A2_N.n4 A2_N.t2 226.809
R3 A2_N.n5 A2_N.t3 226.809
R4 A2_N.n0 A2_N.t7 207.03
R5 A2_N.n5 A2_N.t4 195.746
R6 A2_N.n7 A2_N.t5 186.374
R7 A2_N.n2 A2_N.t6 186.374
R8 A2_N.n6 A2_N 156.912
R9 A2_N A2_N.n3 153.042
R10 A2_N.n9 A2_N.n8 152
R11 A2_N.n1 A2_N.n0 98.8105
R12 A2_N.n4 A2_N.n3 43.5144
R13 A2_N.n7 A2_N.n6 35.4811
R14 A2_N.n3 A2_N.n2 14.7283
R15 A2_N.n6 A2_N.n5 12.7199
R16 A2_N.n8 A2_N.n7 10.0422
R17 A2_N A2_N.n9 9.07957
R18 A2_N.n9 A2_N 5.2098
R19 A2_N.n2 A2_N.n1 2.00883
R20 A2_N.n8 A2_N.n4 2.00883
R21 a_114_368.n6 a_114_368.t12 345.255
R22 a_114_368.n15 a_114_368.t19 261.252
R23 a_114_368.n22 a_114_368.n21 246.312
R24 a_114_368.n3 a_114_368.n1 246.114
R25 a_114_368.n7 a_114_368.t18 240.197
R26 a_114_368.n5 a_114_368.t16 240.197
R27 a_114_368.n14 a_114_368.t17 240.197
R28 a_114_368.n18 a_114_368.n0 203.394
R29 a_114_368.n20 a_114_368.n19 203.394
R30 a_114_368.n23 a_114_368.n22 203.394
R31 a_114_368.n3 a_114_368.n2 194.115
R32 a_114_368.n12 a_114_368.t15 179.947
R33 a_114_368.n8 a_114_368.t13 179.947
R34 a_114_368.n6 a_114_368.t14 174.704
R35 a_114_368.n10 a_114_368.n9 165.189
R36 a_114_368.n16 a_114_368.n15 152
R37 a_114_368.n13 a_114_368.n4 152
R38 a_114_368.n11 a_114_368.n10 152
R39 a_114_368.n15 a_114_368.n14 44.549
R40 a_114_368.n20 a_114_368.n18 42.9181
R41 a_114_368.n22 a_114_368.n20 42.9181
R42 a_114_368.n12 a_114_368.n11 40.1672
R43 a_114_368.n2 a_114_368.t11 30.0005
R44 a_114_368.n17 a_114_368.n16 28.3157
R45 a_114_368.n18 a_114_368.n17 27.7795
R46 a_114_368.n9 a_114_368.n7 27.0217
R47 a_114_368.n9 a_114_368.n8 27.0217
R48 a_114_368.n21 a_114_368.t2 26.3844
R49 a_114_368.n21 a_114_368.t3 26.3844
R50 a_114_368.n0 a_114_368.t7 26.3844
R51 a_114_368.n0 a_114_368.t6 26.3844
R52 a_114_368.n19 a_114_368.t5 26.3844
R53 a_114_368.n19 a_114_368.t4 26.3844
R54 a_114_368.t0 a_114_368.n23 26.3844
R55 a_114_368.n23 a_114_368.t1 26.3844
R56 a_114_368.n2 a_114_368.t9 22.7032
R57 a_114_368.n1 a_114_368.t10 22.7032
R58 a_114_368.n1 a_114_368.t8 22.7032
R59 a_114_368.n7 a_114_368.n6 17.3833
R60 a_114_368.n10 a_114_368.n4 13.1884
R61 a_114_368.n16 a_114_368.n4 13.1884
R62 a_114_368.n8 a_114_368.n5 11.6853
R63 a_114_368.n17 a_114_368.n3 11.3817
R64 a_114_368.n11 a_114_368.n5 10.955
R65 a_114_368.n13 a_114_368.n12 9.49444
R66 a_114_368.n14 a_114_368.n13 5.11262
R67 VPWR.n8 VPWR.t13 342.784
R68 VPWR.n12 VPWR.n11 336.163
R69 VPWR.n26 VPWR.n7 334.173
R70 VPWR.n44 VPWR.n1 331.5
R71 VPWR.n38 VPWR.n37 331.5
R72 VPWR.n35 VPWR.n4 331.5
R73 VPWR.n14 VPWR.n13 321.661
R74 VPWR.n46 VPWR.t4 257.433
R75 VPWR.n29 VPWR.n28 243.916
R76 VPWR.n30 VPWR.n27 36.1417
R77 VPWR.n34 VPWR.n5 36.1417
R78 VPWR.n39 VPWR.n36 36.1417
R79 VPWR.n43 VPWR.n2 36.1417
R80 VPWR.n15 VPWR.n10 36.1417
R81 VPWR.n19 VPWR.n10 36.1417
R82 VPWR.n20 VPWR.n19 36.1417
R83 VPWR.n21 VPWR.n20 36.1417
R84 VPWR.n25 VPWR.n8 35.0123
R85 VPWR.n45 VPWR.n44 33.8829
R86 VPWR.n38 VPWR.n2 29.3652
R87 VPWR.n15 VPWR.n14 28.2358
R88 VPWR.n46 VPWR.n45 27.4829
R89 VPWR.n1 VPWR.t1 26.3844
R90 VPWR.n1 VPWR.t3 26.3844
R91 VPWR.n37 VPWR.t5 26.3844
R92 VPWR.n37 VPWR.t0 26.3844
R93 VPWR.n4 VPWR.t7 26.3844
R94 VPWR.n4 VPWR.t6 26.3844
R95 VPWR.n28 VPWR.t12 26.3844
R96 VPWR.n28 VPWR.t8 26.3844
R97 VPWR.n7 VPWR.t15 26.3844
R98 VPWR.n7 VPWR.t14 26.3844
R99 VPWR.n13 VPWR.t10 26.3844
R100 VPWR.n13 VPWR.t11 26.3844
R101 VPWR.n11 VPWR.t9 26.3844
R102 VPWR.n11 VPWR.t2 26.3844
R103 VPWR.n36 VPWR.n35 24.8476
R104 VPWR.n26 VPWR.n25 20.3299
R105 VPWR.n29 VPWR.n5 20.3299
R106 VPWR.n27 VPWR.n26 15.8123
R107 VPWR.n30 VPWR.n29 15.8123
R108 VPWR.n21 VPWR.n8 12.424
R109 VPWR.n35 VPWR.n34 11.2946
R110 VPWR.n16 VPWR.n15 9.3005
R111 VPWR.n17 VPWR.n10 9.3005
R112 VPWR.n19 VPWR.n18 9.3005
R113 VPWR.n20 VPWR.n9 9.3005
R114 VPWR.n22 VPWR.n21 9.3005
R115 VPWR.n23 VPWR.n8 9.3005
R116 VPWR.n25 VPWR.n24 9.3005
R117 VPWR.n27 VPWR.n6 9.3005
R118 VPWR.n31 VPWR.n30 9.3005
R119 VPWR.n32 VPWR.n5 9.3005
R120 VPWR.n34 VPWR.n33 9.3005
R121 VPWR.n36 VPWR.n3 9.3005
R122 VPWR.n40 VPWR.n39 9.3005
R123 VPWR.n41 VPWR.n2 9.3005
R124 VPWR.n43 VPWR.n42 9.3005
R125 VPWR.n45 VPWR.n0 9.3005
R126 VPWR.n47 VPWR.n46 9.3005
R127 VPWR.n14 VPWR.n12 6.807
R128 VPWR.n39 VPWR.n38 6.77697
R129 VPWR.n44 VPWR.n43 2.25932
R130 VPWR.n16 VPWR.n12 0.50363
R131 VPWR.n17 VPWR.n16 0.122949
R132 VPWR.n18 VPWR.n17 0.122949
R133 VPWR.n18 VPWR.n9 0.122949
R134 VPWR.n22 VPWR.n9 0.122949
R135 VPWR.n23 VPWR.n22 0.122949
R136 VPWR.n24 VPWR.n23 0.122949
R137 VPWR.n24 VPWR.n6 0.122949
R138 VPWR.n31 VPWR.n6 0.122949
R139 VPWR.n32 VPWR.n31 0.122949
R140 VPWR.n33 VPWR.n32 0.122949
R141 VPWR.n33 VPWR.n3 0.122949
R142 VPWR.n40 VPWR.n3 0.122949
R143 VPWR.n41 VPWR.n40 0.122949
R144 VPWR.n42 VPWR.n41 0.122949
R145 VPWR.n42 VPWR.n0 0.122949
R146 VPWR.n47 VPWR.n0 0.122949
R147 VPWR VPWR.n47 0.0617245
R148 VPB.t17 VPB.t8 505.646
R149 VPB VPB.t4 252.823
R150 VPB.t2 VPB.t13 229.839
R151 VPB.t14 VPB.t2 229.839
R152 VPB.t15 VPB.t14 229.839
R153 VPB.t5 VPB.t15 229.839
R154 VPB.t6 VPB.t5 229.839
R155 VPB.t7 VPB.t6 229.839
R156 VPB.t8 VPB.t7 229.839
R157 VPB.t19 VPB.t17 229.839
R158 VPB.t18 VPB.t19 229.839
R159 VPB.t16 VPB.t18 229.839
R160 VPB.t12 VPB.t16 229.839
R161 VPB.t11 VPB.t12 229.839
R162 VPB.t10 VPB.t11 229.839
R163 VPB.t9 VPB.t10 229.839
R164 VPB.t0 VPB.t9 229.839
R165 VPB.t1 VPB.t0 229.839
R166 VPB.t3 VPB.t1 229.839
R167 VPB.t4 VPB.t3 229.839
R168 Y.n5 Y.n3 341.385
R169 Y.n5 Y.n4 298.467
R170 Y.n9 Y.n7 260.13
R171 Y.n2 Y.n0 231.329
R172 Y.n9 Y.n8 229.512
R173 Y.n2 Y.n1 191.965
R174 Y.n6 Y.n5 62.1299
R175 Y.n6 Y.n2 53.6476
R176 Y.n7 Y.t6 26.3844
R177 Y.n7 Y.t4 26.3844
R178 Y.n3 Y.t0 26.3844
R179 Y.n3 Y.t1 26.3844
R180 Y.n4 Y.t2 26.3844
R181 Y.n4 Y.t3 26.3844
R182 Y.n8 Y.t5 26.3844
R183 Y.n8 Y.t7 26.3844
R184 Y.n1 Y.t11 22.7032
R185 Y.n1 Y.t9 22.7032
R186 Y.n0 Y.t10 22.7032
R187 Y.n0 Y.t8 22.7032
R188 Y Y.n6 7.8005
R189 Y Y.n9 5.56264
R190 a_857_74.n1 a_857_74.t7 212.715
R191 a_857_74.n3 a_857_74.t0 203.258
R192 a_857_74.n1 a_857_74.n0 195.918
R193 a_857_74.n3 a_857_74.n2 104.579
R194 a_857_74.n5 a_857_74.n4 104.579
R195 a_857_74.n7 a_857_74.n6 104.579
R196 a_857_74.n8 a_857_74.n1 87.0504
R197 a_857_74.n9 a_857_74.n8 84.741
R198 a_857_74.n8 a_857_74.n7 76.5092
R199 a_857_74.n5 a_857_74.n3 51.9534
R200 a_857_74.n7 a_857_74.n5 51.2005
R201 a_857_74.n2 a_857_74.t1 22.7032
R202 a_857_74.n2 a_857_74.t4 22.7032
R203 a_857_74.n4 a_857_74.t5 22.7032
R204 a_857_74.n4 a_857_74.t6 22.7032
R205 a_857_74.n6 a_857_74.t2 22.7032
R206 a_857_74.n6 a_857_74.t3 22.7032
R207 a_857_74.n0 a_857_74.t8 22.7032
R208 a_857_74.n0 a_857_74.t9 22.7032
R209 a_857_74.n9 a_857_74.t11 22.7032
R210 a_857_74.t10 a_857_74.n9 22.7032
R211 VNB.t8 VNB.t15 2286.61
R212 VNB.t10 VNB.t9 1212.6
R213 VNB.t1 VNB.t0 1154.86
R214 VNB.t6 VNB.t14 1154.86
R215 VNB.t19 VNB.t7 1154.86
R216 VNB VNB.t2 1143.31
R217 VNB.t9 VNB.t8 1097.11
R218 VNB.t4 VNB.t5 1016.27
R219 VNB.t12 VNB.t1 993.177
R220 VNB.t13 VNB.t12 993.177
R221 VNB.t14 VNB.t13 993.177
R222 VNB.t7 VNB.t6 993.177
R223 VNB.t18 VNB.t19 993.177
R224 VNB.t16 VNB.t18 993.177
R225 VNB.t17 VNB.t16 993.177
R226 VNB.t15 VNB.t17 993.177
R227 VNB.t11 VNB.t10 993.177
R228 VNB.t3 VNB.t11 993.177
R229 VNB.t5 VNB.t3 993.177
R230 VNB.t2 VNB.t4 993.177
R231 B1.n11 B1.t2 226.809
R232 B1.n9 B1.t3 226.809
R233 B1.n1 B1.t4 226.809
R234 B1.n2 B1.t5 204.048
R235 B1.n2 B1.t0 197.474
R236 B1.n4 B1.t1 196.013
R237 B1.n11 B1.t6 196.013
R238 B1.n8 B1.t7 196.013
R239 B1.n12 B1.n11 165.145
R240 B1.n10 B1.n0 152
R241 B1.n7 B1.n6 152
R242 B1.n5 B1.n4 152
R243 B1.n3 B1 152
R244 B1.n4 B1.n3 49.6611
R245 B1.n7 B1.n1 45.2793
R246 B1.n11 B1.n10 36.5157
R247 B1.n10 B1.n9 29.2126
R248 B1.n8 B1.n7 13.146
R249 B1.n3 B1.n2 11.6853
R250 B1.n12 B1.n0 10.1214
R251 B1.n5 B1 10.1214
R252 B1.n6 B1 8.33538
R253 B1.n9 B1.n8 7.30353
R254 B1.n6 B1 5.95399
R255 B1.n4 B1.n1 4.38232
R256 B1 B1.n5 4.16794
R257 B1 B1.n12 2.3819
R258 B1 B1.n0 1.78655
R259 VGND.n13 VGND.n10 215.841
R260 VGND.n12 VGND.n11 210.213
R261 VGND.n16 VGND.n9 210.213
R262 VGND.n19 VGND.n18 210.213
R263 VGND.n35 VGND.n2 208.079
R264 VGND.n38 VGND.n37 208.079
R265 VGND.n23 VGND.n6 36.1417
R266 VGND.n24 VGND.n23 36.1417
R267 VGND.n25 VGND.n24 36.1417
R268 VGND.n25 VGND.n4 36.1417
R269 VGND.n29 VGND.n4 36.1417
R270 VGND.n30 VGND.n29 36.1417
R271 VGND.n31 VGND.n30 36.1417
R272 VGND.n31 VGND.n1 36.1417
R273 VGND.n10 VGND.t6 34.0546
R274 VGND.n9 VGND.t10 34.0546
R275 VGND.n18 VGND.t5 34.0546
R276 VGND.n19 VGND.n6 31.2476
R277 VGND.n35 VGND.n1 31.2476
R278 VGND.n17 VGND.n16 28.9887
R279 VGND.n12 VGND.n8 26.7299
R280 VGND.n38 VGND.n36 24.4711
R281 VGND.n10 VGND.t7 22.7032
R282 VGND.n11 VGND.t8 22.7032
R283 VGND.n11 VGND.t9 22.7032
R284 VGND.n9 VGND.t4 22.7032
R285 VGND.n18 VGND.t11 22.7032
R286 VGND.n2 VGND.t1 22.7032
R287 VGND.n2 VGND.t3 22.7032
R288 VGND.n37 VGND.t2 22.7032
R289 VGND.n37 VGND.t0 22.7032
R290 VGND.n16 VGND.n8 18.4476
R291 VGND.n19 VGND.n17 16.1887
R292 VGND.n36 VGND.n35 16.1887
R293 VGND.n14 VGND.n8 9.3005
R294 VGND.n16 VGND.n15 9.3005
R295 VGND.n17 VGND.n7 9.3005
R296 VGND.n20 VGND.n19 9.3005
R297 VGND.n21 VGND.n6 9.3005
R298 VGND.n23 VGND.n22 9.3005
R299 VGND.n24 VGND.n5 9.3005
R300 VGND.n26 VGND.n25 9.3005
R301 VGND.n27 VGND.n4 9.3005
R302 VGND.n29 VGND.n28 9.3005
R303 VGND.n30 VGND.n3 9.3005
R304 VGND.n32 VGND.n31 9.3005
R305 VGND.n33 VGND.n1 9.3005
R306 VGND.n35 VGND.n34 9.3005
R307 VGND.n36 VGND.n0 9.3005
R308 VGND.n39 VGND.n38 7.19894
R309 VGND.n13 VGND.n12 6.53914
R310 VGND.n14 VGND.n13 0.568152
R311 VGND VGND.n39 0.156997
R312 VGND.n39 VGND.n0 0.150766
R313 VGND.n15 VGND.n14 0.122949
R314 VGND.n15 VGND.n7 0.122949
R315 VGND.n20 VGND.n7 0.122949
R316 VGND.n21 VGND.n20 0.122949
R317 VGND.n22 VGND.n21 0.122949
R318 VGND.n22 VGND.n5 0.122949
R319 VGND.n26 VGND.n5 0.122949
R320 VGND.n27 VGND.n26 0.122949
R321 VGND.n28 VGND.n27 0.122949
R322 VGND.n28 VGND.n3 0.122949
R323 VGND.n32 VGND.n3 0.122949
R324 VGND.n33 VGND.n32 0.122949
R325 VGND.n34 VGND.n33 0.122949
R326 VGND.n34 VGND.n0 0.122949
R327 B2.n0 B2.t2 226.809
R328 B2.n2 B2.t3 226.809
R329 B2.n10 B2.t5 226.809
R330 B2.n4 B2.t6 226.809
R331 B2.n4 B2.t0 206.238
R332 B2.n0 B2.t1 197.475
R333 B2.n9 B2.t7 196.013
R334 B2.n3 B2.t4 196.013
R335 B2 B2.n1 155.572
R336 B2.n12 B2.n11 152
R337 B2.n8 B2.n7 152
R338 B2.n6 B2.n5 152
R339 B2.n8 B2.n5 49.6611
R340 B2.n1 B2.n0 45.2793
R341 B2.n11 B2.n10 36.5157
R342 B2.n11 B2.n3 23.3702
R343 B2.n2 B2.n1 20.449
R344 B2.n9 B2.n8 10.2247
R345 B2.n7 B2.n6 10.1214
R346 B2.n12 B2 7.74003
R347 B2 B2.n12 6.54934
R348 B2.n3 B2.n2 5.84292
R349 B2.n10 B2.n9 2.92171
R350 B2.n5 B2.n4 2.92171
R351 B2.n7 B2 2.3819
R352 B2.n6 B2 1.78655
R353 A1_N.n0 A1_N.t0 234.112
R354 A1_N.n11 A1_N.t1 226.809
R355 A1_N.n2 A1_N.t2 226.809
R356 A1_N.n5 A1_N.t5 226.809
R357 A1_N.n5 A1_N.t3 196.013
R358 A1_N.n3 A1_N.t6 196.013
R359 A1_N.n10 A1_N.t7 196.013
R360 A1_N.n0 A1_N.t4 196.013
R361 A1_N.n5 A1_N.n4 164.416
R362 A1_N A1_N.n1 157.209
R363 A1_N.n13 A1_N.n12 152
R364 A1_N.n9 A1_N.n8 152
R365 A1_N.n7 A1_N.n6 152
R366 A1_N.n12 A1_N.n1 49.6611
R367 A1_N.n10 A1_N.n9 40.1672
R368 A1_N.n6 A1_N.n5 37.246
R369 A1_N.n6 A1_N.n3 25.5611
R370 A1_N.n9 A1_N.n2 21.1793
R371 A1_N.n8 A1_N.n7 10.1214
R372 A1_N.n13 A1_N 9.37724
R373 A1_N.n4 A1_N 7.5912
R374 A1_N.n4 A1_N 6.69817
R375 A1_N.n12 A1_N.n11 5.11262
R376 A1_N A1_N.n13 4.91213
R377 A1_N.n11 A1_N.n10 4.38232
R378 A1_N.n1 A1_N.n0 3.65202
R379 A1_N.n7 A1_N 3.42376
R380 A1_N.n3 A1_N.n2 2.92171
R381 A1_N.n8 A1_N 0.744686
R382 a_27_74.n1 a_27_74.t0 209.173
R383 a_27_74.n3 a_27_74.t7 204.012
R384 a_27_74.n1 a_27_74.n0 185
R385 a_27_74.n3 a_27_74.n2 109.109
R386 a_27_74.n5 a_27_74.n4 84.741
R387 a_27_74.n4 a_27_74.n1 83.5077
R388 a_27_74.n4 a_27_74.n3 77.2621
R389 a_27_74.n0 a_27_74.t2 34.0546
R390 a_27_74.n0 a_27_74.t1 26.7573
R391 a_27_74.n2 a_27_74.t4 23.514
R392 a_27_74.n2 a_27_74.t5 23.514
R393 a_27_74.t3 a_27_74.n5 22.7032
R394 a_27_74.n5 a_27_74.t6 22.7032
R395 a_1215_368.n2 a_1215_368.t4 384.327
R396 a_1215_368.n2 a_1215_368.n1 309.351
R397 a_1215_368.t3 a_1215_368.n5 272.635
R398 a_1215_368.n5 a_1215_368.n4 203.333
R399 a_1215_368.n3 a_1215_368.n0 185.442
R400 a_1215_368.n3 a_1215_368.n2 85.4811
R401 a_1215_368.n5 a_1215_368.n3 74.5074
R402 a_1215_368.n0 a_1215_368.t0 26.3844
R403 a_1215_368.n0 a_1215_368.t7 26.3844
R404 a_1215_368.n1 a_1215_368.t6 26.3844
R405 a_1215_368.n1 a_1215_368.t5 26.3844
R406 a_1215_368.n4 a_1215_368.t2 26.3844
R407 a_1215_368.n4 a_1215_368.t1 26.3844
C0 VPWR A1_N 0.091516f
C1 Y VPB 0.024828f
C2 VGND VPB 0.011574f
C3 B1 B2 0.077258f
C4 VPWR A2_N 0.05743f
C5 VPWR B2 0.026347f
C6 VGND A1_N 0.073434f
C7 Y A2_N 3.01e-19
C8 B1 VPWR 0.078242f
C9 VGND A2_N 0.024938f
C10 Y B2 0.245978f
C11 B1 Y 3.69e-19
C12 VGND B2 0.069775f
C13 B1 VGND 0.072519f
C14 VPWR Y 0.431638f
C15 VPWR VGND 0.163479f
C16 VPB A1_N 0.14625f
C17 Y VGND 0.02396f
C18 VPB A2_N 0.130441f
C19 VPB B2 0.143425f
C20 A1_N A2_N 0.088517f
C21 B1 VPB 0.146283f
C22 VPWR VPB 0.269034f
C23 VGND VNB 1.12783f
C24 Y VNB 0.019188f
C25 VPWR VNB 0.956096f
C26 B1 VNB 0.458611f
C27 B2 VNB 0.408651f
C28 A2_N VNB 0.407927f
C29 A1_N VNB 0.454632f
C30 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_1 VNB VPB VPWR VGND
C0 VPB VGND 0.006682f
C1 VPB VPWR 0.025145f
C2 VGND VPWR 0.010643f
C3 VGND VNB 0.11882f
C4 VPWR VNB 0.100356f
C5 VPB VNB 0.191952f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_2 VNB VPB VPWR VGND
C0 VPWR VPB 0.046866f
C1 VGND VPB 0.013363f
C2 VGND VPWR 0.021287f
C3 VGND VNB 0.184043f
C4 VPWR VNB 0.150541f
C5 VPB VNB 0.299088f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_4 VNB VPB VPWR VGND
C0 VGND VPWR 0.042573f
C1 VPB VGND 0.026726f
C2 VPB VPWR 0.090307f
C3 VGND VNB 0.31449f
C4 VPWR VNB 0.250909f
C5 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_8 VNB VPB VPWR VGND
C0 VGND VPB 0.053452f
C1 VPB VPWR 0.177189f
C2 VGND VPWR 0.085146f
C3 VGND VNB 0.575383f
C4 VPWR VNB 0.451646f
C5 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_diode_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_diode_2 VNB VPB VPWR VGND
C0 VPB VPWR 0.040116f
C1 VPB VGND 0.006237f
C2 VPWR VGND 0.033971f
C3 VGND VNB 0.214225f
C4 VPWR VNB 0.178751f
C5 VPB VNB 0.299088f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_2 VNB VPB VPWR VGND
C0 VPWR VPB 0.046866f
C1 VGND VPB 0.013363f
C2 VGND VPWR 0.021287f
C3 VGND VNB 0.184043f
C4 VPWR VNB 0.150541f
C5 VPB VNB 0.299088f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_diode_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_diode_4 VNB VPB VPWR VGND
C0 VPB VPWR 0.063062f
C1 VPWR VGND 0.074126f
C2 VPB VGND 0.008898f
C3 VGND VNB 0.328699f
C4 VPWR VNB 0.270417f
C5 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_4 VNB VPB VPWR VGND
C0 VGND VPWR 0.042573f
C1 VPB VGND 0.026726f
C2 VPB VPWR 0.090307f
C3 VGND VNB 0.31449f
C4 VPWR VNB 0.250909f
C5 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_diode_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_diode_8 VNB VPB VPWR VGND
C0 VPWR VPB 0.108195f
C1 VGND VPB 0.013547f
C2 VPWR VGND 0.151209f
C3 VGND VNB 0.56393f
C4 VPWR VNB 0.460891f
C5 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fill_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fill_8 VNB VPB VPWR VGND
C0 VGND VPB 0.053452f
C1 VPB VPWR 0.177189f
C2 VGND VPWR 0.085146f
C3 VGND VNB 0.575383f
C4 VPWR VNB 0.451646f
C5 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ha_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ha_1 VNB VPB VPWR VGND B SUM COUT A
X0 VPWR.t0 a_83_260.t3 SUM.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3562 pd=1.815 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 COUT.t0 a_239_294.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1245 ps=1.09 w=0.74 l=0.15
X2 a_305_130.t2 a_239_294.t4 a_83_260.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1726 ps=1.85 w=0.64 l=0.15
X3 a_305_130.t1 A.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.125525 ps=1.065 w=0.64 l=0.15
X4 VGND.t0 a_83_260.t4 SUM.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.19515 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 VGND.t1 B.t0 a_305_130.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.125525 pd=1.065 as=0.0896 ps=0.92 w=0.64 l=0.15
X6 COUT.t1 a_239_294.t5 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2051 ps=1.52 w=1.12 l=0.15
X7 VPWR.t1 A.t1 a_239_294.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.126 ps=1.14 w=0.84 l=0.15
X8 a_239_294.t1 B.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.3047 ps=1.675 w=0.84 l=0.15
X9 a_386_392.t1 B.t2 a_83_260.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.1703 ps=1.355 w=1 l=0.15
X10 VGND.t4 A.t2 a_695_119.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1245 pd=1.09 as=0.0672 ps=0.85 w=0.64 l=0.15
X11 a_83_260.t0 a_239_294.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1703 pd=1.355 as=0.3562 ps=1.815 w=0.84 l=0.15
X12 VPWR.t5 A.t3 a_386_392.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3047 pd=1.675 as=0.21 ps=1.42 w=1 l=0.15
X13 a_695_119.t1 B.t3 a_239_294.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1824 ps=1.85 w=0.64 l=0.15
R0 a_83_260.n2 a_83_260.n1 695.098
R1 a_83_260.n0 a_83_260.t3 258.272
R2 a_83_260.n1 a_83_260.t2 247.841
R3 a_83_260.n0 a_83_260.t4 198.023
R4 a_83_260.n1 a_83_260.n0 152
R5 a_83_260.t1 a_83_260.n2 44.5535
R6 a_83_260.n2 a_83_260.t0 35.1791
R7 SUM.n1 SUM 589.85
R8 SUM.n1 SUM.n0 585
R9 SUM.n2 SUM.n1 585
R10 SUM.t1 SUM.n3 279.738
R11 SUM.n4 SUM.t1 279.738
R12 SUM.n1 SUM.t0 26.3844
R13 SUM.n2 SUM 12.9944
R14 SUM.n4 SUM 12.6066
R15 SUM.n0 SUM 11.249
R16 SUM.n3 SUM 10.6672
R17 SUM.n3 SUM 4.84898
R18 SUM.n0 SUM 3.10353
R19 SUM SUM.n4 1.74595
R20 SUM SUM.n2 1.35808
R21 VPWR.n11 VPWR.n10 585
R22 VPWR.n5 VPWR.n4 323.406
R23 VPWR.n3 VPWR.n2 138.37
R24 VPWR.n10 VPWR.t2 83.2565
R25 VPWR.n2 VPWR.t3 73.4067
R26 VPWR.n2 VPWR.t5 70.1253
R27 VPWR.n10 VPWR.t0 53.9524
R28 VPWR.n4 VPWR.t1 46.9053
R29 VPWR.n4 VPWR.t4 42.7253
R30 VPWR.n8 VPWR.n1 36.1417
R31 VPWR.n9 VPWR.n8 35.8489
R32 VPWR.n3 VPWR.n1 24.4711
R33 VPWR.n12 VPWR.n11 10.8486
R34 VPWR.n6 VPWR.n1 9.3005
R35 VPWR.n8 VPWR.n7 9.3005
R36 VPWR.n9 VPWR.n0 9.3005
R37 VPWR.n11 VPWR.n9 4.68547
R38 VPWR.n5 VPWR.n3 3.85859
R39 VPWR.n6 VPWR.n5 0.443135
R40 VPWR VPWR.n12 0.160989
R41 VPWR.n12 VPWR.n0 0.146825
R42 VPWR.n7 VPWR.n6 0.122949
R43 VPWR.n7 VPWR.n0 0.122949
R44 VPB.n0 VPB 1588.44
R45 VPB VPB.n1 952.731
R46 VPB.t2 VPB.t0 431.587
R47 VPB.t6 VPB.n0 373.995
R48 VPB.t4 VPB.t6 311.207
R49 VPB.t1 VPB.t5 280.914
R50 VPB.t0 VPB 257.93
R51 VPB.t3 VPB.t1 229.839
R52 VPB.n1 VPB.t2 201.748
R53 VPB.n0 VPB.t3 71.5059
R54 VPB.n1 VPB.t4 60.058
R55 a_239_294.n4 a_239_294.n3 308.255
R56 a_239_294.n3 a_239_294.n0 306.457
R57 a_239_294.n1 a_239_294.t5 250.909
R58 a_239_294.n0 a_239_294.t6 205.922
R59 a_239_294.n0 a_239_294.t4 184.768
R60 a_239_294.n1 a_239_294.t3 179.947
R61 a_239_294.n2 a_239_294.n1 177.406
R62 a_239_294.n2 a_239_294.t2 158.343
R63 a_239_294.t0 a_239_294.n4 35.1791
R64 a_239_294.n4 a_239_294.t1 35.1791
R65 a_239_294.n3 a_239_294.n2 25.7215
R66 VGND.n8 VGND.t0 237.845
R67 VGND.n2 VGND.n1 214.075
R68 VGND.n4 VGND.n3 129.725
R69 VGND.n1 VGND.t2 42.3444
R70 VGND.n7 VGND.n6 36.1417
R71 VGND.n3 VGND.t3 35.7861
R72 VGND.n3 VGND.t4 26.2505
R73 VGND.n8 VGND.n7 24.4711
R74 VGND.n1 VGND.t1 23.6423
R75 VGND.n6 VGND.n2 18.824
R76 VGND.n7 VGND.n0 9.3005
R77 VGND.n6 VGND.n5 9.3005
R78 VGND.n9 VGND.n8 7.46433
R79 VGND.n4 VGND.n2 7.29889
R80 VGND.n5 VGND.n4 0.168939
R81 VGND VGND.n9 0.160491
R82 VGND.n9 VGND.n0 0.147317
R83 VGND.n5 VGND.n0 0.122949
R84 COUT COUT.n0 588.952
R85 COUT.n2 COUT.n0 585
R86 COUT.n1 COUT.n0 585
R87 COUT COUT.t0 192.887
R88 COUT.n0 COUT.t1 26.3844
R89 COUT COUT.n1 9.64001
R90 COUT COUT.n2 8.69186
R91 COUT.n2 COUT 3.00297
R92 COUT.n1 COUT 2.05482
R93 VNB.t2 VNB.t3 2286.61
R94 VNB.t0 VNB.t4 2205.77
R95 VNB.t1 VNB.t2 1224.15
R96 VNB.t6 VNB.t5 1154.86
R97 VNB VNB.t0 1143.31
R98 VNB.t4 VNB.t1 993.177
R99 VNB.t3 VNB.t6 831.496
R100 a_305_130.n0 a_305_130.t1 373.613
R101 a_305_130.t0 a_305_130.n0 26.2505
R102 a_305_130.n0 a_305_130.t2 26.2505
R103 A.n0 A.t2 552.982
R104 A.t2 A.t1 504.226
R105 A.t0 A.t3 438.889
R106 A.n0 A.t0 156.046
R107 A A.n0 153.851
R108 B.n0 B.t3 259.022
R109 B.n0 B.t1 246.161
R110 B.n1 B.t2 231.629
R111 B B.n1 205.721
R112 B.n1 B.t0 184.768
R113 B B.n0 155.88
R114 a_386_392.t0 a_386_392.t1 82.7405
R115 a_695_119.t0 a_695_119.t1 39.3755
C0 VPWR B 0.038468f
C1 VGND VPB 0.008997f
C2 COUT VPB 0.017555f
C3 VGND B 0.028946f
C4 VPWR A 0.039811f
C5 VPWR SUM 0.069681f
C6 VGND A 0.161013f
C7 VGND SUM 0.075536f
C8 COUT A 0.004048f
C9 VPB B 0.103036f
C10 VPB A 0.082084f
C11 VPB SUM 0.012825f
C12 B A 0.172988f
C13 VPWR VGND 0.080869f
C14 B SUM 5.22e-20
C15 VPWR COUT 0.120537f
C16 A SUM 1.22e-19
C17 VGND COUT 0.093924f
C18 VPWR VPB 0.132722f
C19 COUT VNB 0.108431f
C20 VGND VNB 0.624679f
C21 VPWR VNB 0.463736f
C22 SUM VNB 0.110576f
C23 A VNB 0.398161f
C24 B VNB 0.219964f
C25 VPB VNB 1.13652f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ha_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ha_2 VNB VPB VPWR VGND B A SUM COUT
X0 COUT.t1 a_27_74.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t6 a_391_388.t3 SUM.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t1 a_27_74.t4 COUT.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_27_74.t1 B.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X4 VPWR.t3 a_27_74.t5 a_391_388.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.38685 pd=1.855 as=0.495 ps=1.99 w=1 l=0.15
X5 SUM.t0 a_391_388.t4 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.38685 ps=1.855 w=1.12 l=0.15
X6 SUM.t3 a_391_388.t5 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1962 ps=2.05 w=0.74 l=0.15
X7 COUT.t3 a_27_74.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_114_74.t1 B.t1 a_27_74.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 VGND.t1 a_27_74.t7 COUT.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VGND.t6 B.t2 a_278_74.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.19515 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VGND.t0 A.t0 a_114_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.0888 ps=0.98 w=0.74 l=0.15
X12 VGND.t4 a_391_388.t6 SUM.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X13 a_278_74.t0 a_27_74.t8 a_391_388.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2011 pd=2.05 as=0.201625 ps=2.05 w=0.74 l=0.15
X14 VPWR.t0 A.t1 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.17925 pd=1.375 as=0.15 ps=1.3 w=1 l=0.15
X15 a_278_74.t1 A.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_391_388.t2 B.t3 a_307_388.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.495 pd=1.99 as=0.135 ps=1.27 w=1 l=0.15
X17 a_307_388.t1 A.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.17925 ps=1.375 w=1 l=0.15
R0 a_27_74.n5 a_27_74.n4 649.754
R1 a_27_74.n3 a_27_74.n0 518.116
R2 a_27_74.n2 a_27_74.t5 274.74
R3 a_27_74.n1 a_27_74.t3 243.294
R4 a_27_74.n0 a_27_74.t4 240.197
R5 a_27_74.n1 a_27_74.t6 179.947
R6 a_27_74.n0 a_27_74.t7 179.947
R7 a_27_74.n4 a_27_74.t2 179.204
R8 a_27_74.n2 a_27_74.t8 173.52
R9 a_27_74.n4 a_27_74.n3 111.812
R10 a_27_74.n3 a_27_74.n2 106.312
R11 a_27_74.n0 a_27_74.n1 62.8066
R12 a_27_74.t0 a_27_74.n5 29.5505
R13 a_27_74.n5 a_27_74.t1 29.5505
R14 VPWR.n8 VPWR.t1 872.976
R15 VPWR.n24 VPWR.t5 843.596
R16 VPWR.n7 VPWR.n6 605.946
R17 VPWR.n22 VPWR.n2 603.452
R18 VPWR.n13 VPWR.n12 588.629
R19 VPWR.n15 VPWR.n14 585
R20 VPWR.n14 VPWR.n13 78.0588
R21 VPWR.n17 VPWR.n3 36.1417
R22 VPWR.n21 VPWR.n3 36.1417
R23 VPWR.n2 VPWR.t4 34.2662
R24 VPWR.n17 VPWR.n16 33.8265
R25 VPWR.n2 VPWR.t0 33.3958
R26 VPWR.n14 VPWR.t3 29.5505
R27 VPWR.n6 VPWR.t2 26.3844
R28 VPWR.n6 VPWR.t6 26.3844
R29 VPWR.n11 VPWR.n7 25.224
R30 VPWR.n23 VPWR.n22 22.2123
R31 VPWR.n22 VPWR.n21 21.0829
R32 VPWR.n13 VPWR.t7 20.7211
R33 VPWR.n24 VPWR.n23 20.7064
R34 VPWR.n12 VPWR.n11 20.5681
R35 VPWR.n11 VPWR.n10 9.3005
R36 VPWR.n9 VPWR.n5 9.3005
R37 VPWR.n16 VPWR.n4 9.3005
R38 VPWR.n18 VPWR.n17 9.3005
R39 VPWR.n19 VPWR.n3 9.3005
R40 VPWR.n21 VPWR.n20 9.3005
R41 VPWR.n22 VPWR.n1 9.3005
R42 VPWR.n23 VPWR.n0 9.3005
R43 VPWR.n25 VPWR.n24 9.3005
R44 VPWR.n8 VPWR.n7 6.50549
R45 VPWR.n15 VPWR.n5 6.18281
R46 VPWR.n16 VPWR.n15 2.17737
R47 VPWR.n12 VPWR.n5 1.3937
R48 VPWR.n10 VPWR.n8 0.686474
R49 VPWR.n10 VPWR.n9 0.122949
R50 VPWR.n9 VPWR.n4 0.122949
R51 VPWR.n18 VPWR.n4 0.122949
R52 VPWR.n19 VPWR.n18 0.122949
R53 VPWR.n20 VPWR.n19 0.122949
R54 VPWR.n20 VPWR.n1 0.122949
R55 VPWR.n1 VPWR.n0 0.122949
R56 VPWR.n25 VPWR.n0 0.122949
R57 VPWR VPWR.n25 0.0617245
R58 COUT.n1 COUT.n0 650.141
R59 COUT.n2 COUT.n1 185
R60 COUT.n3 COUT.n2 185
R61 COUT.n0 COUT.t0 26.3844
R62 COUT.n0 COUT.t1 26.3844
R63 COUT.n2 COUT.t2 22.7032
R64 COUT.n2 COUT.t3 22.7032
R65 COUT.n3 COUT 12.6066
R66 COUT.n1 COUT 4.84898
R67 COUT COUT.n3 1.74595
R68 VPB.t5 VPB.t1 582.259
R69 VPB.t1 VPB.t8 452.017
R70 VPB.t0 VPB.t4 257.93
R71 VPB VPB.t6 257.93
R72 VPB.t3 VPB.t2 229.839
R73 VPB.t7 VPB.t3 229.839
R74 VPB.t8 VPB.t7 229.839
R75 VPB.t6 VPB.t0 229.839
R76 VPB.t4 VPB.t5 214.517
R77 a_391_388.n6 a_391_388.n5 644.091
R78 a_391_388.n5 a_391_388.t1 273.961
R79 a_391_388.n1 a_391_388.t3 261.62
R80 a_391_388.n0 a_391_388.t4 261.62
R81 a_391_388.n4 a_391_388.n3 170.654
R82 a_391_388.n6 a_391_388.t2 165.481
R83 a_391_388.n1 a_391_388.t6 161.482
R84 a_391_388.n2 a_391_388.t5 154.24
R85 a_391_388.n4 a_391_388.n0 95.2419
R86 a_391_388.n3 a_391_388.n2 35.055
R87 a_391_388.t0 a_391_388.n6 29.5505
R88 a_391_388.n3 a_391_388.n1 27.752
R89 a_391_388.n5 a_391_388.n4 10.3536
R90 a_391_388.n2 a_391_388.n0 2.92171
R91 SUM.n2 SUM.n1 585
R92 SUM SUM.n0 279.183
R93 SUM.n0 SUM.t2 26.7573
R94 SUM.n0 SUM.t3 26.7573
R95 SUM.n1 SUM.t1 26.3844
R96 SUM.n1 SUM.t0 26.3844
R97 SUM SUM.n2 12.6176
R98 SUM.n2 SUM 4.93764
R99 B.n0 B.t0 273.786
R100 B.n1 B.t3 231.629
R101 B.n1 B.t2 230.825
R102 B.n2 B.n0 210.742
R103 B.n0 B.t1 202.671
R104 B B.n1 195.704
R105 B.n2 B 27.2005
R106 B B.n2 3.5205
R107 VGND.n14 VGND.t6 231.453
R108 VGND.n8 VGND.t5 231.453
R109 VGND.n4 VGND.n3 212.137
R110 VGND.n17 VGND.n16 204.976
R111 VGND.n5 VGND.t1 178.81
R112 VGND.n9 VGND.n1 36.1417
R113 VGND.n13 VGND.n1 36.1417
R114 VGND.n9 VGND.n8 32.0005
R115 VGND.n17 VGND.n15 31.2476
R116 VGND.n7 VGND.n4 28.2358
R117 VGND.n3 VGND.t2 22.7032
R118 VGND.n3 VGND.t4 22.7032
R119 VGND.n16 VGND.t3 22.7032
R120 VGND.n16 VGND.t0 22.7032
R121 VGND.n8 VGND.n7 15.4358
R122 VGND.n15 VGND.n0 9.3005
R123 VGND.n13 VGND.n12 9.3005
R124 VGND.n11 VGND.n1 9.3005
R125 VGND.n10 VGND.n9 9.3005
R126 VGND.n8 VGND.n2 9.3005
R127 VGND.n7 VGND.n6 9.3005
R128 VGND.n15 VGND.n14 8.65932
R129 VGND.n5 VGND.n4 6.79022
R130 VGND.n18 VGND.n17 6.66636
R131 VGND.n14 VGND.n13 2.63579
R132 VGND.n6 VGND.n5 0.5771
R133 VGND VGND.n18 0.267138
R134 VGND.n18 VGND.n0 0.163541
R135 VGND.n6 VGND.n2 0.122949
R136 VGND.n10 VGND.n2 0.122949
R137 VGND.n11 VGND.n10 0.122949
R138 VGND.n12 VGND.n11 0.122949
R139 VGND.n12 VGND.n0 0.122949
R140 VNB.t7 VNB.t1 2748.56
R141 VNB.t1 VNB.t6 2286.61
R142 VNB VNB.t8 1143.31
R143 VNB.t6 VNB.t5 1108.66
R144 VNB.t3 VNB.t2 993.177
R145 VNB.t5 VNB.t3 993.177
R146 VNB.t4 VNB.t7 993.177
R147 VNB.t0 VNB.t4 993.177
R148 VNB.t8 VNB.t0 900.788
R149 a_114_74.t0 a_114_74.t1 38.9194
R150 a_278_74.n1 a_278_74.n0 519.528
R151 a_278_74.n2 a_278_74.n1 67.2005
R152 a_278_74.n0 a_278_74.t2 22.7032
R153 a_278_74.n0 a_278_74.t1 22.7032
R154 a_278_74.n1 a_278_74.t0 18.5827
R155 A.n0 A.t3 238.292
R156 A.n1 A.t0 225.213
R157 A.n0 A.t2 212.081
R158 A.n1 A.t1 207.529
R159 A A.n2 156.268
R160 A.n2 A.n1 36.1505
R161 A.n2 A.n0 12.0505
R162 a_307_388.t0 a_307_388.t1 53.1905
C0 SUM COUT 0.096605f
C1 VPWR VGND 0.09838f
C2 COUT VPB 0.002506f
C3 SUM VGND 0.05545f
C4 VGND VPB 0.01085f
C5 COUT VGND 0.132153f
C6 B A 0.184763f
C7 B VPWR 0.166917f
C8 B SUM 1.58e-20
C9 B VPB 0.108543f
C10 B COUT 8.25e-21
C11 A VPWR 0.033519f
C12 B VGND 0.028262f
C13 A VPB 0.076762f
C14 VPWR SUM 0.023642f
C15 VPWR VPB 0.164877f
C16 VPWR COUT 0.013188f
C17 A VGND 0.031091f
C18 SUM VPB 0.004763f
C19 VGND VNB 0.741142f
C20 COUT VNB 0.011811f
C21 SUM VNB 0.013209f
C22 VPWR VNB 0.571346f
C23 A VNB 0.193799f
C24 B VNB 0.307672f
C25 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__maj3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__maj3_1 VNB VPB VPWR VGND A B X C
X0 a_84_74.t3 B.t0 a_226_384.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_406_384.t1 B.t1 a_84_74.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X2 a_598_384.t1 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X3 a_226_384.t0 A.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.1934 ps=1.475 w=1 l=0.15
X4 VGND.t0 C.t0 a_403_136.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
X5 a_84_74.t1 C.t1 a_595_136.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1733 pd=1.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 a_403_136.t1 B.t2 a_84_74.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1222 ps=1.08 w=0.64 l=0.15
X7 a_595_136.t1 A.t2 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0864 pd=0.91 as=0.1344 ps=1.06 w=0.64 l=0.15
X8 VGND.t1 a_84_74.t6 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1389 pd=1.135 as=0.2081 ps=2.05 w=0.74 l=0.15
X9 VPWR.t1 a_84_74.t7 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.3304 ps=2.83 w=1.12 l=0.15
X10 a_84_74.t2 B.t3 a_223_120.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1222 pd=1.08 as=0.0768 ps=0.88 w=0.64 l=0.15
X11 a_223_120.t1 A.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1389 ps=1.135 w=0.64 l=0.15
X12 VPWR.t0 C.t2 a_406_384.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X13 a_84_74.t0 C.t3 a_598_384.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
R0 B.n0 B.t1 209.72
R1 B.n1 B.t0 207.529
R2 B.n1 B.t3 170.453
R3 B B.n2 166.811
R4 B.n0 B.t2 138.173
R5 B.n2 B.n0 61.346
R6 B.n2 B.n1 6.57323
R7 a_226_384.t0 a_226_384.t1 53.1905
R8 a_84_74.t0 a_84_74.n5 340.596
R9 a_84_74.n3 a_84_74.t1 319.877
R10 a_84_74.n0 a_84_74.t7 250.548
R11 a_84_74.n2 a_84_74.n0 223.374
R12 a_84_74.n5 a_84_74.n4 210.905
R13 a_84_74.n0 a_84_74.t6 177.981
R14 a_84_74.n2 a_84_74.n1 98.8784
R15 a_84_74.n5 a_84_74.n3 51.9534
R16 a_84_74.n1 a_84_74.t5 42.0902
R17 a_84_74.n4 a_84_74.t3 35.4605
R18 a_84_74.n4 a_84_74.t4 29.5505
R19 a_84_74.n1 a_84_74.t2 23.133
R20 a_84_74.n3 a_84_74.n2 12.8005
R21 VPB VPB.t6 280.914
R22 VPB.t0 VPB.t2 275.807
R23 VPB.t6 VPB.t3 257.93
R24 VPB.t5 VPB.t4 245.161
R25 VPB.t2 VPB.t1 214.517
R26 VPB.t4 VPB.t0 214.517
R27 VPB.t3 VPB.t5 214.517
R28 a_406_384.t0 a_406_384.t1 53.1905
R29 A.n0 A.t3 759.953
R30 A.t3 A.t1 453.616
R31 A.t2 A.t0 432.193
R32 A A.n0 180.649
R33 A.n0 A.t2 162.274
R34 VPWR.n2 VPWR.n0 319.214
R35 VPWR.n2 VPWR.n1 229.377
R36 VPWR.n0 VPWR.t2 39.4005
R37 VPWR.n0 VPWR.t0 37.4305
R38 VPWR.n1 VPWR.t1 36.2945
R39 VPWR.n1 VPWR.t3 30.5355
R40 VPWR VPWR.n2 0.217021
R41 a_598_384.t0 a_598_384.t1 53.1905
R42 C.n0 C.t3 231.629
R43 C.n1 C.t2 229.619
R44 C C.n0 184.72
R45 C.n0 C.t1 162.274
R46 C C.n1 155.84
R47 C.n1 C.t0 154.643
R48 a_403_136.t0 a_403_136.t1 45.0005
R49 VGND.n2 VGND.n1 264.442
R50 VGND.n2 VGND.n0 216.863
R51 VGND.n0 VGND.t1 39.5361
R52 VGND.n1 VGND.t2 39.3755
R53 VGND.n1 VGND.t0 39.3755
R54 VGND.n0 VGND.t3 30.938
R55 VGND VGND.n2 0.235935
R56 VNB.t1 VNB.t6 1316.54
R57 VNB.t4 VNB.t5 1258.79
R58 VNB.t2 VNB.t3 1177.95
R59 VNB VNB.t4 1143.31
R60 VNB.t6 VNB.t0 970.08
R61 VNB.t3 VNB.t1 900.788
R62 VNB.t5 VNB.t2 900.788
R63 a_595_136.t0 a_595_136.t1 50.6255
R64 X X.n0 588.952
R65 X.n2 X.n0 585
R66 X.n1 X.n0 585
R67 X X.t0 177.417
R68 X.n0 X.t1 26.3844
R69 X X.n1 9.64001
R70 X X.n2 8.69186
R71 X.n2 X 3.00297
R72 X.n1 X 2.05482
R73 a_223_120.t0 a_223_120.t1 45.0005
C0 VPB VPWR 0.109434f
C1 VPB C 0.08299f
C2 X VPWR 0.131851f
C3 VPB A 0.061787f
C4 VPB VGND 0.007908f
C5 VPB B 0.073192f
C6 X A 0.002596f
C7 X VGND 0.06879f
C8 VPWR C 0.034079f
C9 X B 0.003396f
C10 VPWR A 0.041004f
C11 A C 0.135088f
C12 VPWR VGND 0.061917f
C13 C VGND 0.019846f
C14 VPWR B 0.038008f
C15 A VGND 0.252486f
C16 B C 0.058958f
C17 A B 0.100842f
C18 B VGND 0.017031f
C19 VPB X 0.018055f
C20 VGND VNB 0.498255f
C21 C VNB 0.212639f
C22 B VNB 0.164573f
C23 A VNB 0.454494f
C24 VPWR VNB 0.390409f
C25 X VNB 0.105759f
C26 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__maj3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__maj3_2 VNB VPB VPWR VGND B C X A
X0 a_790_368.t1 A.t0 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2184 ps=1.525 w=1 l=0.15
X1 X.t1 a_87_264.t6 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t2 C.t0 a_584_347.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.525 as=0.155 ps=1.31 w=1 l=0.15
X3 a_413_74.t1 A.t1 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.33115 ps=1.635 w=0.74 l=0.15
X4 VPWR.t0 a_87_264.t7 X.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.4032 pd=1.885 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_87_264.t3 C.t1 a_793_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6 VGND.t0 a_87_264.t8 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.33115 pd=1.635 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 X.t2 a_87_264.t9 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8 a_393_368.t1 A.t2 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.186675 pd=1.46 as=0.4032 ps=1.885 w=1 l=0.15
X9 a_87_264.t0 B.t0 a_413_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.0888 ps=0.98 w=0.74 l=0.15
X10 VGND.t2 C.t2 a_577_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1665 pd=1.19 as=0.1221 ps=1.07 w=0.74 l=0.15
X11 a_584_347.t0 B.t1 a_87_264.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.31 as=0.15 ps=1.3 w=1 l=0.15
X12 a_87_264.t2 B.t2 a_393_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.186675 ps=1.46 w=1 l=0.15
X13 a_577_74.t0 B.t3 a_87_264.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_793_74.t1 A.t3 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1665 ps=1.19 w=0.74 l=0.15
X15 a_87_264.t1 C.t3 a_790_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
R0 A.t2 A.t0 1075.4
R1 A.t0 A.t3 506.101
R2 A.n0 A.t2 242.339
R3 A A.n0 196.764
R4 A.n0 A.t1 168.846
R5 VPWR.n2 VPWR.n1 326.168
R6 VPWR.n6 VPWR.t1 259.171
R7 VPWR.n4 VPWR.n3 139.466
R8 VPWR.n3 VPWR.t3 69.3402
R9 VPWR.n3 VPWR.t0 65.6186
R10 VPWR.n1 VPWR.t2 56.6157
R11 VPWR.n1 VPWR.t4 28.8981
R12 VPWR.n5 VPWR.n4 27.4829
R13 VPWR.n6 VPWR.n5 25.224
R14 VPWR.n5 VPWR.n0 9.3005
R15 VPWR.n7 VPWR.n6 9.3005
R16 VPWR.n4 VPWR.n2 4.07289
R17 VPWR.n2 VPWR.n0 0.213523
R18 VPWR.n7 VPWR.n0 0.122949
R19 VPWR VPWR.n7 0.0617245
R20 a_790_368.t0 a_790_368.t1 53.1905
R21 VPB.n0 VPB 1953.63
R22 VPB VPB.n1 906.49
R23 VPB.n1 VPB.t0 459.678
R24 VPB.t1 VPB 268.146
R25 VPB.t4 VPB.n0 251.399
R26 VPB.t6 VPB.t3 244.149
R27 VPB.t0 VPB.t1 229.839
R28 VPB.t5 VPB.t4 222.393
R29 VPB.t3 VPB.t5 217.558
R30 VPB.t7 VPB.t2 214.517
R31 VPB.n0 VPB.t7 12.4188
R32 VPB.n1 VPB.t6 3.72599
R33 a_87_264.t1 a_87_264.n7 352.272
R34 a_87_264.n7 a_87_264.n0 292.5
R35 a_87_264.n2 a_87_264.t3 266.197
R36 a_87_264.n6 a_87_264.n5 246.329
R37 a_87_264.n5 a_87_264.t7 234.841
R38 a_87_264.n3 a_87_264.t9 234.841
R39 a_87_264.n3 a_87_264.t6 187.834
R40 a_87_264.n4 a_87_264.t8 186.374
R41 a_87_264.n2 a_87_264.n1 92.5005
R42 a_87_264.n6 a_87_264.n2 62.7049
R43 a_87_264.n4 a_87_264.n3 61.346
R44 a_87_264.n0 a_87_264.t4 29.5505
R45 a_87_264.n0 a_87_264.t2 29.5505
R46 a_87_264.n1 a_87_264.t5 22.7032
R47 a_87_264.n1 a_87_264.t0 22.7032
R48 a_87_264.n7 a_87_264.n6 9.06385
R49 a_87_264.n5 a_87_264.n4 4.38232
R50 VGND.n7 VGND.n6 205.262
R51 VGND.n3 VGND.n1 185
R52 VGND.n2 VGND.n1 185
R53 VGND.n10 VGND.t1 171.77
R54 VGND.n5 VGND.n4 74.5346
R55 VGND.n6 VGND.t3 36.487
R56 VGND.n6 VGND.t2 36.487
R57 VGND.n4 VGND.n3 35.9339
R58 VGND.n4 VGND.n2 35.9339
R59 VGND.n2 VGND.t4 33.2437
R60 VGND.n9 VGND.n8 26.7299
R61 VGND.n10 VGND.n9 25.224
R62 VGND.n3 VGND.t0 22.7032
R63 VGND.n11 VGND.n10 9.3005
R64 VGND.n9 VGND.n0 9.3005
R65 VGND.n8 VGND.n5 8.97828
R66 VGND.n5 VGND.n1 6.04494
R67 VGND.n8 VGND.n7 4.05562
R68 VGND.n7 VGND.n0 0.216105
R69 VGND.n11 VGND.n0 0.122949
R70 VGND VGND.n11 0.0617245
R71 X.n2 X 589.444
R72 X.n2 X.n0 585
R73 X.n3 X.n2 585
R74 X X.n1 159.339
R75 X.n2 X.t3 26.3844
R76 X.n2 X.t2 26.3844
R77 X.n1 X.t0 22.7032
R78 X.n1 X.t1 22.7032
R79 X X.n3 11.9116
R80 X X.n0 10.3116
R81 X X.n0 2.84494
R82 X.n3 X 1.24494
R83 VNB VNB.n0 4583.33
R84 VNB.n0 VNB.t1 2148.03
R85 VNB.t4 VNB.t6 1466.67
R86 VNB.t2 VNB 1189.5
R87 VNB.t5 VNB.t4 1173.33
R88 VNB.t0 VNB.t5 1051.11
R89 VNB.t1 VNB.t2 993.177
R90 VNB.t6 VNB.t3 953.333
R91 VNB.t7 VNB.t0 953.333
R92 VNB.n0 VNB.t7 281.111
R93 C.n0 C.t3 245.018
R94 C.n1 C.t0 231.629
R95 C.n0 C.t1 204.048
R96 C.n1 C.t2 186.374
R97 C C.n0 182.191
R98 C C.n1 155.231
R99 a_584_347.t0 a_584_347.t1 61.0705
R100 a_413_74.t0 a_413_74.t1 38.9194
R101 a_793_74.t0 a_793_74.t1 38.9194
R102 a_393_368.n0 a_393_368.t1 45.8843
R103 a_393_368.n1 a_393_368.n0 40.8873
R104 a_393_368.n0 a_393_368.t0 26.9849
R105 B.n0 B.t1 212.641
R106 B.n1 B.t2 207.529
R107 B.n1 B.t0 164.464
R108 B.n0 B.t3 162.274
R109 B B.n2 67.3122
R110 B.n2 B.n1 32.0985
R111 B.n2 B.n0 21.7022
R112 a_577_74.t0 a_577_74.t1 53.514
C0 C VPB 0.071671f
C1 B A 0.075758f
C2 X VPWR 0.212737f
C3 C A 0.133217f
C4 B VPWR 0.012715f
C5 VGND VPB 0.011066f
C6 VGND A 0.059897f
C7 C VPWR 0.028848f
C8 VGND VPWR 0.091441f
C9 X B 1.16e-19
C10 VPB A 0.260499f
C11 X VGND 0.158809f
C12 B C 0.086393f
C13 VPB VPWR 0.140874f
C14 B VGND 0.017533f
C15 A VPWR 0.108468f
C16 C VGND 0.031022f
C17 X VPB 0.006114f
C18 B VPB 0.06247f
C19 X A 0.004782f
C20 VGND VNB 0.626989f
C21 C VNB 0.250483f
C22 B VNB 0.168283f
C23 X VNB 0.031408f
C24 VPWR VNB 0.51029f
C25 A VNB 0.298721f
C26 VPB VNB 1.18075f
.ends

* NGSPICE file created from sky130_fd_sc_hs__maj3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__maj3_4 VNB VPB VPWR VGND C B X A
X0 VGND.t2 A.t0 a_114_125.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
X1 VPWR.t8 a_219_392.t12 X.t2 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_906_78.t1 A.t1 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.133125 pd=1.205 as=0.112 ps=0.99 w=0.64 l=0.15
X3 X.t1 a_219_392.t13 VPWR.t7 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t6 a_219_392.t14 X.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 X.t3 a_219_392.t15 VPWR.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1934 ps=1.475 w=1.12 l=0.15
X6 a_219_392.t5 C.t0 a_906_78.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.133125 ps=1.205 w=0.64 l=0.15
X7 VPWR.t4 C.t1 a_501_392.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X8 a_504_125.t1 C.t2 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1088 pd=0.98 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 a_219_392.t6 C.t3 a_905_392# VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X10 VPWR A a_905_392# VPB sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.15 ps=1.3 w=1 l=0.15
X11 a_219_392.t2 B.t0 a_114_125.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.174875 ps=1.315 w=0.64 l=0.15
X12 VGND.t8 C.t4 a_504_125.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.162075 ps=1.32 w=0.64 l=0.15
X13 a_114_125.t2 B.t1 a_219_392.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X14 a_905_392# A.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.21 ps=1.42 w=1 l=0.15
X15 a_905_392# C.t5 a_219_392.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X16 X.t7 a_219_392.t16 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.12945 ps=1.1 w=0.74 l=0.15
X17 a_501_392.t0 B.t2 a_219_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X18 a_906_78.t2 C.t6 a_219_392.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X19 a_119_392.t1 A.t3 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X20 X.t6 a_219_392.t17 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 a_114_125.t0 A.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.174875 pd=1.315 as=0.1824 ps=1.85 w=0.64 l=0.15
X22 a_219_392.t10 B.t3 a_504_125.t3 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1088 ps=0.98 w=0.64 l=0.15
X23 VGND.t0 A.t5 a_906_78.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.0896 ps=0.92 w=0.64 l=0.15
X24 VGND.t6 a_219_392.t18 X.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1962 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 a_219_392.t11 B.t4 a_501_392.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X26 VPWR.t2 A.t6 a_119_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X27 a_501_392.t1 C.t7 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.18 ps=1.36 w=1 l=0.15
X28 VGND.t7 a_219_392.t19 X.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1184 ps=1.06 w=0.74 l=0.15
X29 a_119_392.t3 B.t5 a_219_392.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X30 a_219_392.t8 B.t6 a_119_392.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X31 a_504_125.t2 B.t7 a_219_392.t9 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.162075 pd=1.32 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 A.t0 A.t4 931.867
R1 A.t1 A.t5 798.514
R2 A.t5 A.n0 463.553
R3 A.t4 A.t3 455.519
R4 A A.n1 329.067
R5 A.n1 A.t1 268.313
R6 A.n2 A.t6 231.629
R7 A.n1 A.t2 231.629
R8 A.n2 A.t0 192.8
R9 A A.n2 156.268
R10 a_114_125.n1 a_114_125.n0 482.296
R11 a_114_125.n1 a_114_125.t3 41.2505
R12 a_114_125.t0 a_114_125.n1 41.2505
R13 a_114_125.n0 a_114_125.t2 39.3755
R14 a_114_125.n0 a_114_125.t1 26.2505
R15 VGND.n8 VGND.t6 243.413
R16 VGND.n26 VGND.n3 237.329
R17 VGND.n10 VGND.n9 210.988
R18 VGND.n20 VGND.n19 205.752
R19 VGND.n33 VGND.t1 162.518
R20 VGND.n13 VGND.n12 129.95
R21 VGND.n12 VGND.t0 41.0701
R22 VGND.n19 VGND.t3 39.3755
R23 VGND.n17 VGND.n6 36.1417
R24 VGND.n18 VGND.n17 36.1417
R25 VGND.n24 VGND.n4 36.1417
R26 VGND.n25 VGND.n24 36.1417
R27 VGND.n27 VGND.n1 36.1417
R28 VGND.n31 VGND.n1 36.1417
R29 VGND.n32 VGND.n31 36.1417
R30 VGND.n13 VGND.n6 32.7534
R31 VGND.n26 VGND.n25 30.8711
R32 VGND.n20 VGND.n4 30.4946
R33 VGND.n11 VGND.n10 28.2358
R34 VGND.n19 VGND.t8 26.2505
R35 VGND.n3 VGND.t9 26.2505
R36 VGND.n3 VGND.t2 26.2505
R37 VGND.n9 VGND.t5 22.7032
R38 VGND.n9 VGND.t7 22.7032
R39 VGND.n12 VGND.t4 21.1849
R40 VGND.n13 VGND.n11 20.7064
R41 VGND.n33 VGND.n32 20.7064
R42 VGND.n20 VGND.n18 16.9417
R43 VGND.n34 VGND.n33 9.3005
R44 VGND.n11 VGND.n7 9.3005
R45 VGND.n14 VGND.n13 9.3005
R46 VGND.n15 VGND.n6 9.3005
R47 VGND.n17 VGND.n16 9.3005
R48 VGND.n18 VGND.n5 9.3005
R49 VGND.n21 VGND.n20 9.3005
R50 VGND.n22 VGND.n4 9.3005
R51 VGND.n24 VGND.n23 9.3005
R52 VGND.n25 VGND.n2 9.3005
R53 VGND.n28 VGND.n27 9.3005
R54 VGND.n29 VGND.n1 9.3005
R55 VGND.n31 VGND.n30 9.3005
R56 VGND.n32 VGND.n0 9.3005
R57 VGND.n10 VGND.n8 6.26985
R58 VGND.n27 VGND.n26 5.27109
R59 VGND.n8 VGND.n7 0.733933
R60 VGND.n14 VGND.n7 0.122949
R61 VGND.n15 VGND.n14 0.122949
R62 VGND.n16 VGND.n15 0.122949
R63 VGND.n16 VGND.n5 0.122949
R64 VGND.n21 VGND.n5 0.122949
R65 VGND.n22 VGND.n21 0.122949
R66 VGND.n23 VGND.n22 0.122949
R67 VGND.n23 VGND.n2 0.122949
R68 VGND.n28 VGND.n2 0.122949
R69 VGND.n29 VGND.n28 0.122949
R70 VGND.n30 VGND.n29 0.122949
R71 VGND.n30 VGND.n0 0.122949
R72 VGND.n34 VGND.n0 0.122949
R73 VGND VGND.n34 0.0617245
R74 VNB.t14 VNB.t10 1362.73
R75 VNB.t1 VNB.t9 1362.73
R76 VNB.t0 VNB.t5 1177.95
R77 VNB.t2 VNB.t12 1177.95
R78 VNB.t10 VNB.t2 1154.86
R79 VNB.t4 VNB.t3 1154.86
R80 VNB VNB.t1 1143.31
R81 VNB.t13 VNB.t15 1131.76
R82 VNB.t5 VNB.t8 1085.56
R83 VNB.t6 VNB.t7 993.177
R84 VNB.t8 VNB.t6 993.177
R85 VNB.t11 VNB.t0 993.177
R86 VNB.t12 VNB.t11 993.177
R87 VNB.t15 VNB.t14 993.177
R88 VNB.t3 VNB.t13 993.177
R89 VNB.t9 VNB.t4 993.177
R90 a_219_392.n16 a_219_392.n15 585
R91 a_219_392.n2 a_219_392.n0 336.531
R92 a_219_392.n19 a_219_392.n17 306.159
R93 a_219_392.n21 a_219_392.n20 295.856
R94 a_219_392.n19 a_219_392.n18 294.236
R95 a_219_392.n12 a_219_392.t15 228.148
R96 a_219_392.n6 a_219_392.t13 228.148
R97 a_219_392.n9 a_219_392.t14 228.148
R98 a_219_392.n4 a_219_392.t12 206.715
R99 a_219_392.n7 a_219_392.n3 165.189
R100 a_219_392.n4 a_219_392.t18 156.424
R101 a_219_392.n11 a_219_392.t16 154.24
R102 a_219_392.n8 a_219_392.t19 154.24
R103 a_219_392.n5 a_219_392.t17 154.24
R104 a_219_392.n13 a_219_392.n12 152
R105 a_219_392.n10 a_219_392.n3 152
R106 a_219_392.n20 a_219_392.n16 128.572
R107 a_219_392.n20 a_219_392.n19 121.828
R108 a_219_392.n2 a_219_392.n1 90.4996
R109 a_219_392.n5 a_219_392.n4 60.6205
R110 a_219_392.n11 a_219_392.n10 45.2793
R111 a_219_392.n16 a_219_392.n14 41.2308
R112 a_219_392.n21 a_219_392.t11 39.4005
R113 a_219_392.n14 a_219_392.n2 32.9542
R114 a_219_392.n14 a_219_392.n13 32.1944
R115 a_219_392.n7 a_219_392.n6 32.1338
R116 a_219_392.n18 a_219_392.t7 29.5505
R117 a_219_392.n18 a_219_392.t8 29.5505
R118 a_219_392.n15 a_219_392.t3 29.5505
R119 a_219_392.n15 a_219_392.t6 29.5505
R120 a_219_392.t1 a_219_392.n21 29.5505
R121 a_219_392.n8 a_219_392.n7 26.2914
R122 a_219_392.n17 a_219_392.t0 26.2505
R123 a_219_392.n17 a_219_392.t2 26.2505
R124 a_219_392.n1 a_219_392.t4 26.2505
R125 a_219_392.n1 a_219_392.t5 26.2505
R126 a_219_392.n0 a_219_392.t9 26.2505
R127 a_219_392.n0 a_219_392.t10 26.2505
R128 a_219_392.n10 a_219_392.n9 16.0672
R129 a_219_392.n13 a_219_392.n3 13.1884
R130 a_219_392.n9 a_219_392.n8 7.30353
R131 a_219_392.n6 a_219_392.n5 4.38232
R132 a_219_392.n12 a_219_392.n11 4.38232
R133 X.n2 X.n1 261.877
R134 X.n2 X.n0 210.614
R135 X.n5 X.n4 185
R136 X.n5 X.n3 159.456
R137 X X.n2 62.6747
R138 X X.n5 33.4082
R139 X.n3 X.t7 29.1897
R140 X.n0 X.t2 26.3844
R141 X.n0 X.t1 26.3844
R142 X.n1 X.t0 26.3844
R143 X.n1 X.t3 26.3844
R144 X.n4 X.t5 22.7032
R145 X.n4 X.t6 22.7032
R146 X.n3 X.t4 22.7032
R147 VPWR.n25 VPWR.n3 615.032
R148 VPWR.n19 VPWR.n6 608.662
R149 VPWR.n11 VPWR.n10 324.702
R150 VPWR.n13 VPWR.t5 269.568
R151 VPWR.n31 VPWR.t0 260.733
R152 VPWR.n9 VPWR.t8 256.671
R153 VPWR.n6 VPWR.t1 43.3405
R154 VPWR.n3 VPWR.t3 40.3855
R155 VPWR.n6 VPWR.t4 39.4005
R156 VPWR.n29 VPWR.n1 36.1417
R157 VPWR.n30 VPWR.n29 36.1417
R158 VPWR.n23 VPWR.n4 36.1417
R159 VPWR.n24 VPWR.n23 36.1417
R160 VPWR.n17 VPWR.n7 36.1417
R161 VPWR.n18 VPWR.n17 36.1417
R162 VPWR.n13 VPWR.n7 31.624
R163 VPWR.n12 VPWR.n11 31.2476
R164 VPWR.n3 VPWR.t2 30.5355
R165 VPWR.n19 VPWR.n4 29.3652
R166 VPWR.n25 VPWR.n1 28.6123
R167 VPWR.n10 VPWR.t7 26.3844
R168 VPWR.n10 VPWR.t6 26.3844
R169 VPWR.n31 VPWR.n30 25.6005
R170 VPWR.n25 VPWR.n24 24.0946
R171 VPWR.n13 VPWR.n12 21.8358
R172 VPWR.n19 VPWR.n18 18.0711
R173 VPWR.n12 VPWR.n8 9.3005
R174 VPWR.n14 VPWR.n13 9.3005
R175 VPWR.n15 VPWR.n7 9.3005
R176 VPWR.n17 VPWR.n16 9.3005
R177 VPWR.n18 VPWR.n5 9.3005
R178 VPWR.n20 VPWR.n19 9.3005
R179 VPWR.n21 VPWR.n4 9.3005
R180 VPWR.n23 VPWR.n22 9.3005
R181 VPWR.n24 VPWR.n2 9.3005
R182 VPWR.n26 VPWR.n25 9.3005
R183 VPWR.n27 VPWR.n1 9.3005
R184 VPWR.n29 VPWR.n28 9.3005
R185 VPWR.n30 VPWR.n0 9.3005
R186 VPWR.n32 VPWR.n31 9.3005
R187 VPWR.n11 VPWR.n9 6.50549
R188 VPWR.n9 VPWR.n8 0.686474
R189 VPWR.n14 VPWR.n8 0.122949
R190 VPWR.n15 VPWR.n14 0.122949
R191 VPWR.n16 VPWR.n15 0.122949
R192 VPWR.n16 VPWR.n5 0.122949
R193 VPWR.n20 VPWR.n5 0.122949
R194 VPWR.n21 VPWR.n20 0.122949
R195 VPWR.n22 VPWR.n21 0.122949
R196 VPWR.n22 VPWR.n2 0.122949
R197 VPWR.n26 VPWR.n2 0.122949
R198 VPWR.n27 VPWR.n26 0.122949
R199 VPWR.n28 VPWR.n27 0.122949
R200 VPWR.n28 VPWR.n0 0.122949
R201 VPWR.n32 VPWR.n0 0.122949
R202 VPWR VPWR.n32 0.0617245
R203 VPB.t4 VPB.t11 487.769
R204 VPB.t6 VPB.t2 291.13
R205 VPB VPB.t1 265.591
R206 VPB.t0 VPB.t5 260.485
R207 VPB.t3 VPB.t6 255.376
R208 VPB.t10 VPB.t3 255.376
R209 VPB.t1 VPB.t9 255.376
R210 VPB.t13 VPB.t14 229.839
R211 VPB.t12 VPB.t13 229.839
R212 VPB.t11 VPB.t12 229.839
R213 VPB.t7 VPB.t4 229.839
R214 VPB.t2 VPB.t7 229.839
R215 VPB.t5 VPB.t10 229.839
R216 VPB.t8 VPB.t0 229.839
R217 VPB.t9 VPB.t8 229.839
R218 a_906_78.n1 a_906_78.n0 466.406
R219 a_906_78.n1 a_906_78.t3 49.6449
R220 a_906_78.n0 a_906_78.t0 26.2505
R221 a_906_78.n0 a_906_78.t2 26.2505
R222 a_906_78.t1 a_906_78.n1 21.4851
R223 C.t4 C.t2 853.14
R224 C.t2 C.t7 457.632
R225 C.n3 C.t1 255.69
R226 C.n4 C.n2 239.308
R227 C.n3 C.t4 236.411
R228 C.n1 C.t3 217.023
R229 C.n0 C.t5 207.529
R230 C.n0 C.t6 186.089
R231 C.n1 C.t0 178.34
R232 C.n4 C.n3 152
R233 C.n2 C.n0 43.0884
R234 C.n2 C.n1 13.146
R235 C C.n4 7.34659
R236 a_501_392.n1 a_501_392.n0 1241.39
R237 a_501_392.n1 a_501_392.t0 39.4005
R238 a_501_392.n0 a_501_392.t3 29.5505
R239 a_501_392.n0 a_501_392.t1 29.5505
R240 a_501_392.t2 a_501_392.n1 29.5505
R241 a_504_125.n1 a_504_125.n0 454.568
R242 a_504_125.n0 a_504_125.t2 61.9565
R243 a_504_125.n0 a_504_125.t0 34.688
R244 a_504_125.n1 a_504_125.t3 31.8755
R245 a_504_125.t1 a_504_125.n1 31.8755
R246 B B.n6 245.087
R247 B.n1 B.t4 241
R248 B.n5 B.t6 240.27
R249 B.n0 B.t2 235.57
R250 B.n4 B.t5 232.968
R251 B.n3 B.n2 152
R252 B.n4 B.t1 144.746
R253 B.n0 B.t7 138.173
R254 B.n1 B.t3 138.173
R255 B.n5 B.t0 138.173
R256 B.n2 B.n0 59.8853
R257 B.n6 B.n5 31.4035
R258 B.n6 B.n4 24.8308
R259 B B.n3 8.90485
R260 B.n2 B.n1 2.92171
R261 B.n3 B 1.78137
R262 a_119_392.n1 a_119_392.n0 943.856
R263 a_119_392.n1 a_119_392.t2 39.4005
R264 a_119_392.n0 a_119_392.t0 29.5505
R265 a_119_392.n0 a_119_392.t3 29.5505
R266 a_119_392.t1 a_119_392.n1 29.5505
C0 B C 0.194293f
C1 A VPWR 0.076821f
C2 VGND X 0.202158f
C3 B VPWR 0.025078f
C4 C VPWR 0.048082f
C5 a_905_392# VPB 0.006783f
C6 VGND VPB 0.014188f
C7 a_905_392# A 0.011009f
C8 VGND A 0.158343f
C9 X VPB 0.012918f
C10 VGND B 0.050107f
C11 X A 0.002319f
C12 a_905_392# C 0.024483f
C13 X B 6.41e-21
C14 VGND C 0.08557f
C15 a_905_392# VPWR 0.162651f
C16 VGND VPWR 0.143571f
C17 VPB A 0.176766f
C18 X VPWR 0.426813f
C19 VPB B 0.153706f
C20 A B 0.296311f
C21 VPB C 0.148889f
C22 VPB VPWR 0.225293f
C23 A C 0.447343f
C24 VGND a_905_392# 0.002795f
C25 X VNB 0.057792f
C26 VGND VNB 0.976318f
C27 VPWR VNB 0.825249f
C28 C VNB 0.55436f
C29 B VNB 0.333277f
C30 A VNB 0.783982f
C31 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2_1 VNB VPB VPWR VGND X S A0 A1
X0 VGND.t2 a_27_112.t2 a_443_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.20905 pd=1.305 as=0.2997 ps=1.55 w=0.74 l=0.15
X1 VPWR.t3 S.t0 a_27_112.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 X.t1 a_304_74.t4 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2557 ps=1.59 w=1.12 l=0.15
X3 VPWR.t0 a_27_112.t3 a_524_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2557 pd=1.59 as=0.21 ps=1.42 w=1 l=0.15
X4 a_304_74.t0 A1.t0 a_226_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.20165 pd=1.285 as=0.0888 ps=0.98 w=0.74 l=0.15
X5 X.t0 a_304_74.t5 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.20905 ps=1.305 w=0.74 l=0.15
X6 a_223_368.t1 S.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.4075 pd=1.815 as=0.1853 ps=1.385 w=1 l=0.15
X7 a_304_74.t2 A0.t0 a_223_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.4075 ps=1.815 w=1 l=0.15
X8 a_443_74.t1 A0.t1 a_304_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=1.55 as=0.20165 ps=1.285 w=0.74 l=0.15
X9 a_524_368.t0 A1.t1 a_304_74.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.195 ps=1.39 w=1 l=0.15
X10 a_226_74.t1 S.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.144575 ps=1.15 w=0.74 l=0.15
X11 VGND.t1 S.t3 a_27_112.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.144575 pd=1.15 as=0.15675 ps=1.67 w=0.55 l=0.15
R0 a_27_112.t1 a_27_112.n1 783.771
R1 a_27_112.t1 a_27_112.n2 718.559
R2 a_27_112.n1 a_27_112.n0 497.986
R3 a_27_112.n2 a_27_112.t0 292.997
R4 a_27_112.n0 a_27_112.t3 239.661
R5 a_27_112.n0 a_27_112.t2 210.474
R6 a_27_112.n2 a_27_112.n1 3.29747
R7 a_443_74.t0 a_443_74.t1 131.351
R8 VGND.n2 VGND.n0 216.272
R9 VGND.n2 VGND.n1 120.71
R10 VGND.n0 VGND.t2 46.2167
R11 VGND.n0 VGND.t3 45.4059
R12 VGND.n1 VGND.t1 42.8374
R13 VGND.n1 VGND.t0 32.2699
R14 VGND VGND.n2 0.204724
R15 VNB.t5 VNB.t3 2217.32
R16 VNB.t3 VNB.t4 1651.44
R17 VNB.t2 VNB.t5 1605.25
R18 VNB.t1 VNB.t0 1293.44
R19 VNB VNB.t1 1143.31
R20 VNB.t0 VNB.t2 900.788
R21 S.n0 S.t1 207.529
R22 S.n0 S.t2 198.204
R23 S.n1 S.t0 181.821
R24 S.n1 S.t3 166.947
R25 S S.n2 154.522
R26 S.n2 S.n0 54.0429
R27 S.n2 S.n1 24.1005
R28 VPWR.n2 VPWR.n1 622.521
R29 VPWR.n2 VPWR.n0 229.951
R30 VPWR.n1 VPWR.t3 55.1136
R31 VPWR.n0 VPWR.t0 53.1905
R32 VPWR.n0 VPWR.t1 35.2408
R33 VPWR.n1 VPWR.t2 30.4598
R34 VPWR VPWR.n2 0.202943
R35 VPB.t4 VPB.t2 492.877
R36 VPB.t1 VPB.t3 316.668
R37 VPB.t0 VPB.t1 291.13
R38 VPB.t2 VPB.t0 275.807
R39 VPB.t5 VPB.t4 273.253
R40 VPB VPB.t5 257.93
R41 a_304_74.n3 a_304_74.n2 486.913
R42 a_304_74.n2 a_304_74.n0 301.521
R43 a_304_74.n0 a_304_74.t4 264.298
R44 a_304_74.n0 a_304_74.t5 204.048
R45 a_304_74.n2 a_304_74.n1 185
R46 a_304_74.t1 a_304_74.n3 47.2805
R47 a_304_74.n1 a_304_74.t3 44.5951
R48 a_304_74.n1 a_304_74.t0 43.7843
R49 a_304_74.n3 a_304_74.t2 29.5505
R50 X.n1 X 588.636
R51 X.n1 X.n0 585
R52 X.n2 X.n1 585
R53 X X.t0 205.1
R54 X.n1 X.t1 26.3844
R55 X X.n2 9.74595
R56 X X.n0 8.43686
R57 X X.n0 2.32777
R58 X.n2 X 1.01868
R59 a_524_368.t0 a_524_368.t1 82.7405
R60 A1 A1.t1 425.228
R61 A1.n0 A1.t0 419
R62 A1.n0 A1 12.2187
R63 A1 A1.n0 2.13383
R64 a_226_74.t0 a_226_74.t1 38.9194
R65 a_223_368.t0 a_223_368.t1 160.555
R66 A0.n0 A0.t0 266.44
R67 A0.n0 A0.t1 178.34
R68 A0 A0.n0 157.744
C0 VPB X 0.019138f
C1 VPB VPWR 0.120525f
C2 S A1 0.040558f
C3 VPB VGND 0.007976f
C4 S X 7.35e-20
C5 A0 A1 0.169224f
C6 S VPWR 0.029088f
C7 S VGND 0.053687f
C8 A0 VPWR 0.005355f
C9 A0 VGND 0.006604f
C10 A1 VPWR 0.008123f
C11 A1 VGND 0.018598f
C12 VPWR X 0.145606f
C13 X VGND 0.076208f
C14 VPWR VGND 0.070402f
C15 VPB S 0.082896f
C16 VPB A0 0.036036f
C17 VPB A1 0.046616f
C18 S A0 0.008407f
C19 VGND VNB 0.551037f
C20 X VNB 0.112862f
C21 VPWR VNB 0.436357f
C22 A1 VNB 0.16319f
C23 A0 VNB 0.112787f
C24 S VNB 0.240566f
C25 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ha_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ha_4 VNB VPB VPWR SUM VGND COUT B A
X0 a_435_99.t3 A.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.175875 pd=1.425 as=0.126 ps=1.14 w=0.84 l=0.15
X1 VPWR.t8 a_294_392.t6 SUM.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3136 ps=1.68 w=1.12 l=0.15
X2 VPWR.t9 B.t0 a_435_99.t4 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.222525 ps=1.58 w=0.84 l=0.15
X3 a_27_125.t5 B.t1 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0992 pd=0.95 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 a_27_125.t3 a_435_99.t6 a_294_392.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2144 pd=1.95 as=0.1024 ps=0.96 w=0.64 l=0.15
X5 VPWR.t4 A.t1 a_435_99.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.273 pd=1.63 as=0.175875 ps=1.425 w=0.84 l=0.15
X6 a_27_392.t3 B.t2 a_294_392.t4 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.15 ps=1.3 w=1 l=0.15
X7 VGND.t2 a_294_392.t7 SUM.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.14985 ps=1.145 w=0.74 l=0.15
X8 a_435_99.t5 B.t3 VPWR.t10 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.222525 pd=1.58 as=0.126 ps=1.14 w=0.84 l=0.15
X9 a_707_119.t1 A.t2 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.176 pd=1.83 as=0.112 ps=0.99 w=0.64 l=0.15
X10 a_294_392.t5 B.t4 a_27_392.t2 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR.t0 a_435_99.t7 a_294_392.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X12 VPWR.t11 a_435_99.t8 COUT.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2576 ps=1.58 w=1.12 l=0.15
X13 a_27_392.t1 A.t3 VPWR.t7 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X14 a_294_392.t2 a_435_99.t9 VPWR.t12 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2394 ps=2.25 w=0.84 l=0.15
X15 SUM.t1 a_294_392.t8 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.14985 pd=1.145 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 COUT.t4 a_435_99.t10 VPWR.t13 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2576 pd=1.58 as=0.273 ps=1.63 w=1.12 l=0.15
X17 VGND.t6 A.t4 a_707_119.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.112 ps=0.99 w=0.64 l=0.15
X18 a_294_392.t1 a_435_99.t11 a_27_125.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.0992 ps=0.95 w=0.64 l=0.15
X19 a_435_99.t1 B.t5 a_707_119.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1856 ps=1.86 w=0.64 l=0.15
X20 VGND.t0 a_294_392.t9 SUM.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VGND.t5 A.t5 a_27_125.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0912 pd=0.925 as=0.1824 ps=1.85 w=0.64 l=0.15
X22 a_27_125.t0 A.t6 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0912 ps=0.925 w=0.64 l=0.15
X23 VGND.t8 a_435_99.t12 COUT.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VPWR.t6 A.t7 a_27_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.285 ps=2.57 w=1 l=0.15
X25 a_707_119.t2 B.t6 a_435_99.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X26 SUM.t5 a_294_392.t10 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=1.68 as=0.168 ps=1.42 w=1.12 l=0.15
X27 VGND.t7 a_435_99.t13 COUT.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VPWR.t2 a_294_392.t11 SUM.t4 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 SUM.t3 a_294_392.t12 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X30 VPWR.t14 a_435_99.t14 COUT.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X31 VGND.t9 B.t7 a_27_125.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X32 COUT.t2 a_435_99.t15 VPWR.t15 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.t6 A.t4 1687
R1 A.n1 A.t0 254.404
R2 A.n2 A.t3 213.98
R3 A.n3 A.t7 211.544
R4 A.n0 A.t1 197.385
R5 A.n2 A.t6 163.881
R6 A.n3 A.t5 163.881
R7 A.n5 A.n4 152
R8 A.n0 A.t2 126.927
R9 A.t4 A.n1 126.927
R10 A.n1 A.n0 75.313
R11 A.n4 A.n3 33.5944
R12 A.n4 A.n2 29.9429
R13 A.n5 A 15.1278
R14 A A.n5 3.49141
R15 VPWR.n36 VPWR.t12 790.742
R16 VPWR.n28 VPWR.n9 631.946
R17 VPWR.n34 VPWR.n5 613.703
R18 VPWR.n7 VPWR.n6 607.692
R19 VPWR.n23 VPWR.n12 606.333
R20 VPWR.n21 VPWR.n13 606.333
R21 VPWR.n17 VPWR.t8 349.466
R22 VPWR.n42 VPWR.n1 323.925
R23 VPWR.n16 VPWR.n15 315.812
R24 VPWR.n9 VPWR.t4 70.3576
R25 VPWR.n40 VPWR.n2 36.1417
R26 VPWR.n41 VPWR.n40 36.1417
R27 VPWR.n27 VPWR.n10 36.1417
R28 VPWR.n20 VPWR.n14 36.1417
R29 VPWR.n9 VPWR.t13 35.8187
R30 VPWR.n5 VPWR.t10 35.1791
R31 VPWR.n5 VPWR.t0 35.1791
R32 VPWR.n6 VPWR.t5 35.1791
R33 VPWR.n6 VPWR.t9 35.1791
R34 VPWR.n29 VPWR.n28 33.8829
R35 VPWR.n23 VPWR.n22 32.7534
R36 VPWR.n42 VPWR.n41 29.7417
R37 VPWR.n1 VPWR.t7 29.5505
R38 VPWR.n1 VPWR.t6 29.5505
R39 VPWR.n34 VPWR.n33 28.2358
R40 VPWR.n12 VPWR.t15 26.3844
R41 VPWR.n12 VPWR.t11 26.3844
R42 VPWR.n13 VPWR.t3 26.3844
R43 VPWR.n13 VPWR.t14 26.3844
R44 VPWR.n15 VPWR.t1 26.3844
R45 VPWR.n15 VPWR.t2 26.3844
R46 VPWR.n33 VPWR.n7 26.3534
R47 VPWR.n36 VPWR.n2 23.7181
R48 VPWR.n36 VPWR.n35 23.7181
R49 VPWR.n29 VPWR.n7 21.0829
R50 VPWR.n35 VPWR.n34 19.2005
R51 VPWR.n23 VPWR.n10 14.6829
R52 VPWR.n17 VPWR.n16 12.8919
R53 VPWR.n22 VPWR.n21 10.1652
R54 VPWR.n18 VPWR.n14 9.3005
R55 VPWR.n20 VPWR.n19 9.3005
R56 VPWR.n22 VPWR.n11 9.3005
R57 VPWR.n24 VPWR.n23 9.3005
R58 VPWR.n25 VPWR.n10 9.3005
R59 VPWR.n27 VPWR.n26 9.3005
R60 VPWR.n28 VPWR.n8 9.3005
R61 VPWR.n30 VPWR.n29 9.3005
R62 VPWR.n31 VPWR.n7 9.3005
R63 VPWR.n33 VPWR.n32 9.3005
R64 VPWR.n34 VPWR.n4 9.3005
R65 VPWR.n35 VPWR.n3 9.3005
R66 VPWR.n37 VPWR.n36 9.3005
R67 VPWR.n38 VPWR.n2 9.3005
R68 VPWR.n40 VPWR.n39 9.3005
R69 VPWR.n41 VPWR.n0 9.3005
R70 VPWR.n43 VPWR.n42 7.23624
R71 VPWR.n16 VPWR.n14 5.64756
R72 VPWR.n28 VPWR.n27 4.14168
R73 VPWR.n21 VPWR.n20 1.12991
R74 VPWR.n18 VPWR.n17 0.537576
R75 VPWR VPWR.n43 0.157488
R76 VPWR.n43 VPWR.n0 0.150282
R77 VPWR.n19 VPWR.n18 0.122949
R78 VPWR.n19 VPWR.n11 0.122949
R79 VPWR.n24 VPWR.n11 0.122949
R80 VPWR.n25 VPWR.n24 0.122949
R81 VPWR.n26 VPWR.n25 0.122949
R82 VPWR.n26 VPWR.n8 0.122949
R83 VPWR.n30 VPWR.n8 0.122949
R84 VPWR.n31 VPWR.n30 0.122949
R85 VPWR.n32 VPWR.n31 0.122949
R86 VPWR.n32 VPWR.n4 0.122949
R87 VPWR.n4 VPWR.n3 0.122949
R88 VPWR.n37 VPWR.n3 0.122949
R89 VPWR.n38 VPWR.n37 0.122949
R90 VPWR.n39 VPWR.n38 0.122949
R91 VPWR.n39 VPWR.n0 0.122949
R92 a_435_99.n19 a_435_99.n18 660.562
R93 a_435_99.n21 a_435_99.n20 629.931
R94 a_435_99.n14 a_435_99.t11 277.2
R95 a_435_99.n11 a_435_99.t10 249.886
R96 a_435_99.n3 a_435_99.t14 234.841
R97 a_435_99.n5 a_435_99.t15 234.841
R98 a_435_99.n8 a_435_99.t8 234.841
R99 a_435_99.n3 a_435_99.t12 200.195
R100 a_435_99.n16 a_435_99.t7 190.974
R101 a_435_99.n10 a_435_99.n1 186.374
R102 a_435_99.n7 a_435_99.t13 186.374
R103 a_435_99.n4 a_435_99.n2 186.374
R104 a_435_99.n15 a_435_99.t9 181.821
R105 a_435_99.n17 a_435_99.n16 180.898
R106 a_435_99.n6 a_435_99.n0 165.189
R107 a_435_99.n12 a_435_99.n11 152
R108 a_435_99.n9 a_435_99.n0 152
R109 a_435_99.n14 a_435_99.t6 124.796
R110 a_435_99.n17 a_435_99.n13 113.724
R111 a_435_99.n23 a_435_99.n22 78.0571
R112 a_435_99.n18 a_435_99.t4 72.6962
R113 a_435_99.n20 a_435_99.n19 67.8771
R114 a_435_99.n4 a_435_99.n3 51.852
R115 a_435_99.n20 a_435_99.n12 51.2005
R116 a_435_99.n16 a_435_99.n15 45.76
R117 a_435_99.n6 a_435_99.n5 40.1672
R118 a_435_99.n18 a_435_99.t5 38.01
R119 a_435_99.n21 a_435_99.t2 34.55
R120 a_435_99.n22 a_435_99.t3 32.253
R121 a_435_99.n22 a_435_99.n21 31.2703
R122 a_435_99.n11 a_435_99.n10 27.752
R123 a_435_99.n13 a_435_99.t0 26.2505
R124 a_435_99.n13 a_435_99.t1 26.2505
R125 a_435_99.n15 a_435_99.n14 25.7458
R126 a_435_99.n9 a_435_99.n8 24.1005
R127 a_435_99.n10 a_435_99.n9 21.9096
R128 a_435_99.n8 a_435_99.n7 16.7975
R129 a_435_99.n5 a_435_99.n4 13.8763
R130 a_435_99.n12 a_435_99.n0 13.1884
R131 a_435_99.n7 a_435_99.n6 8.76414
R132 a_435_99.n19 a_435_99.n17 4.84944
R133 VPB.t15 VPB.t10 520.968
R134 VPB.t0 VPB.t13 362.635
R135 VPB.t5 VPB.t9 337.098
R136 VPB.t9 VPB.t11 311.56
R137 VPB.t16 VPB.t14 309.005
R138 VPB.t6 VPB.t5 268.146
R139 VPB VPB.t3 252.823
R140 VPB.t1 VPB.t0 229.839
R141 VPB.t2 VPB.t1 229.839
R142 VPB.t8 VPB.t2 229.839
R143 VPB.t7 VPB.t8 229.839
R144 VPB.t11 VPB.t7 229.839
R145 VPB.t14 VPB.t6 229.839
R146 VPB.t12 VPB.t16 229.839
R147 VPB.t10 VPB.t12 229.839
R148 VPB.t17 VPB.t15 229.839
R149 VPB.t4 VPB.t17 229.839
R150 VPB.t3 VPB.t4 229.839
R151 a_294_392.n20 a_294_392.n19 585
R152 a_294_392.n19 a_294_392.n18 409.781
R153 a_294_392.n2 a_294_392.n1 363.759
R154 a_294_392.n16 a_294_392.t12 242.875
R155 a_294_392.n5 a_294_392.t6 237.032
R156 a_294_392.n4 a_294_392.t10 234.841
R157 a_294_392.n13 a_294_392.t11 234.841
R158 a_294_392.n16 a_294_392.n15 186.374
R159 a_294_392.n12 a_294_392.t9 186.374
R160 a_294_392.n7 a_294_392.t8 186.374
R161 a_294_392.n6 a_294_392.t7 186.374
R162 a_294_392.n9 a_294_392.n5 166.159
R163 a_294_392.n18 a_294_392.n17 152
R164 a_294_392.n14 a_294_392.n3 152
R165 a_294_392.n11 a_294_392.n10 152
R166 a_294_392.n9 a_294_392.n8 152
R167 a_294_392.n2 a_294_392.n0 148.857
R168 a_294_392.n17 a_294_392.n14 53.3126
R169 a_294_392.n12 a_294_392.n11 51.1217
R170 a_294_392.n8 a_294_392.n6 45.2793
R171 a_294_392.n8 a_294_392.n7 35.7853
R172 a_294_392.t3 a_294_392.n20 35.1791
R173 a_294_392.n20 a_294_392.t2 35.1791
R174 a_294_392.n0 a_294_392.t1 33.7505
R175 a_294_392.n1 a_294_392.t4 29.5505
R176 a_294_392.n1 a_294_392.t5 29.5505
R177 a_294_392.n0 a_294_392.t0 26.2505
R178 a_294_392.n19 a_294_392.n2 25.9884
R179 a_294_392.n10 a_294_392.n9 15.3217
R180 a_294_392.n10 a_294_392.n3 15.3217
R181 a_294_392.n18 a_294_392.n3 14.1581
R182 a_294_392.n7 a_294_392.n4 12.4157
R183 a_294_392.n11 a_294_392.n4 9.49444
R184 a_294_392.n6 a_294_392.n5 8.03383
R185 a_294_392.n13 a_294_392.n12 5.11262
R186 a_294_392.n17 a_294_392.n16 2.92171
R187 a_294_392.n14 a_294_392.n13 1.46111
R188 SUM.n6 SUM.n5 230.814
R189 SUM.n1 SUM.t0 201.816
R190 SUM.n4 SUM.n3 201.362
R191 SUM.n1 SUM.n0 100.547
R192 SUM.n2 SUM.n1 91.5627
R193 SUM.n3 SUM.t5 52.7684
R194 SUM.n3 SUM.t6 45.7326
R195 SUM.n0 SUM.t1 34.0546
R196 SUM.n0 SUM.t2 31.6221
R197 SUM.n5 SUM.t4 26.3844
R198 SUM.n5 SUM.t3 26.3844
R199 SUM.n4 SUM.n2 23.2732
R200 SUM.n6 SUM.n4 13.9641
R201 SUM SUM.n6 10.0101
R202 SUM SUM.n2 9.3467
R203 B.n2 B.n1 953.321
R204 B.n1 B.t0 345.166
R205 B.n0 B.t6 335.793
R206 B.n1 B.t3 250.105
R207 B.t3 B.n0 239.929
R208 B.n0 B.t5 197.62
R209 B.n2 B.t2 186.107
R210 B.n4 B.t4 186.107
R211 B.n4 B.t7 168.671
R212 B.n3 B.t1 163.881
R213 B.n6 B.n5 152
R214 B.n5 B.n4 37.9934
R215 B B.n6 13.3823
R216 B.n5 B.n3 6.80521
R217 B.n3 B.n2 6.23815
R218 B.n6 B 5.23686
R219 VGND.n7 VGND.t8 295.558
R220 VGND.n16 VGND.t7 295.558
R221 VGND.n8 VGND.t2 241.192
R222 VGND.n36 VGND.n35 224.68
R223 VGND.n39 VGND.n38 224.68
R224 VGND.n10 VGND.n9 207.498
R225 VGND.n23 VGND.n22 124.478
R226 VGND.n22 VGND.t6 39.3755
R227 VGND.n24 VGND.n3 36.1417
R228 VGND.n28 VGND.n3 36.1417
R229 VGND.n29 VGND.n28 36.1417
R230 VGND.n30 VGND.n29 36.1417
R231 VGND.n30 VGND.n1 36.1417
R232 VGND.n34 VGND.n1 36.1417
R233 VGND.n9 VGND.t0 34.0546
R234 VGND.n11 VGND.n7 32.377
R235 VGND.n39 VGND.n37 30.4946
R236 VGND.n21 VGND.n5 30.1181
R237 VGND.n24 VGND.n23 29.3652
R238 VGND.n38 VGND.t4 27.188
R239 VGND.n22 VGND.t3 26.2505
R240 VGND.n35 VGND.t10 26.2505
R241 VGND.n35 VGND.t9 26.2505
R242 VGND.n38 VGND.t5 26.2505
R243 VGND.n16 VGND.n15 24.8476
R244 VGND.n17 VGND.n5 23.3417
R245 VGND.n9 VGND.t1 22.7032
R246 VGND.n17 VGND.n16 22.5887
R247 VGND.n23 VGND.n21 18.0711
R248 VGND.n37 VGND.n36 15.8123
R249 VGND.n15 VGND.n7 15.0593
R250 VGND.n11 VGND.n10 12.8005
R251 VGND.n37 VGND.n0 9.3005
R252 VGND.n34 VGND.n33 9.3005
R253 VGND.n32 VGND.n1 9.3005
R254 VGND.n31 VGND.n30 9.3005
R255 VGND.n29 VGND.n2 9.3005
R256 VGND.n28 VGND.n27 9.3005
R257 VGND.n26 VGND.n3 9.3005
R258 VGND.n25 VGND.n24 9.3005
R259 VGND.n23 VGND.n4 9.3005
R260 VGND.n12 VGND.n11 9.3005
R261 VGND.n13 VGND.n7 9.3005
R262 VGND.n15 VGND.n14 9.3005
R263 VGND.n16 VGND.n6 9.3005
R264 VGND.n18 VGND.n17 9.3005
R265 VGND.n19 VGND.n5 9.3005
R266 VGND.n21 VGND.n20 9.3005
R267 VGND.n40 VGND.n39 7.19894
R268 VGND.n10 VGND.n8 7.12592
R269 VGND.n36 VGND.n34 1.50638
R270 VGND.n12 VGND.n8 0.599569
R271 VGND VGND.n40 0.156997
R272 VGND.n40 VGND.n0 0.150766
R273 VGND.n13 VGND.n12 0.122949
R274 VGND.n14 VGND.n13 0.122949
R275 VGND.n14 VGND.n6 0.122949
R276 VGND.n18 VGND.n6 0.122949
R277 VGND.n19 VGND.n18 0.122949
R278 VGND.n20 VGND.n19 0.122949
R279 VGND.n20 VGND.n4 0.122949
R280 VGND.n25 VGND.n4 0.122949
R281 VGND.n26 VGND.n25 0.122949
R282 VGND.n27 VGND.n26 0.122949
R283 VGND.n27 VGND.n2 0.122949
R284 VGND.n31 VGND.n2 0.122949
R285 VGND.n32 VGND.n31 0.122949
R286 VGND.n33 VGND.n32 0.122949
R287 VGND.n33 VGND.n0 0.122949
R288 COUT.n2 COUT.n0 617
R289 COUT.n2 COUT.n1 585
R290 COUT.n3 COUT.t1 282.913
R291 COUT.n3 COUT.t0 181.299
R292 COUT.n0 COUT.t4 53.6478
R293 COUT.n0 COUT.t5 27.2639
R294 COUT.n1 COUT.t3 26.3844
R295 COUT.n1 COUT.t2 26.3844
R296 COUT COUT.n3 7.6063
R297 COUT COUT.n2 1.29905
R298 VNB.n0 VNB 11098.2
R299 VNB VNB.n1 8523.5
R300 VNB.t6 VNB.t7 3233.6
R301 VNB.t8 VNB.t0 1986.35
R302 VNB.t7 VNB.t8 1986.35
R303 VNB.n1 VNB.t10 1905.51
R304 VNB.t1 VNB.t2 1281.89
R305 VNB.t0 VNB.t1 1154.86
R306 VNB.t5 VNB.t6 1154.86
R307 VNB.t4 VNB 1143.31
R308 VNB.t12 VNB.n0 1142.08
R309 VNB.t10 VNB.t9 1085.56
R310 VNB.t9 VNB.t14 1062.47
R311 VNB.t13 VNB.t12 1033.88
R312 VNB.t3 VNB.t4 1004.72
R313 VNB.t14 VNB.t11 993.177
R314 VNB.t11 VNB.t3 993.177
R315 VNB.n1 VNB.t13 853.553
R316 VNB.n0 VNB.t5 29.4516
R317 a_27_125.n1 a_27_125.t3 224.637
R318 a_27_125.t1 a_27_125.n3 184.076
R319 a_27_125.n3 a_27_125.n2 100.871
R320 a_27_125.n1 a_27_125.n0 89.2272
R321 a_27_125.n3 a_27_125.n1 55.5811
R322 a_27_125.n0 a_27_125.t2 31.8755
R323 a_27_125.n0 a_27_125.t5 26.2505
R324 a_27_125.n2 a_27_125.t4 26.2505
R325 a_27_125.n2 a_27_125.t0 26.2505
R326 a_27_392.n0 a_27_392.t3 408.207
R327 a_27_392.n0 a_27_392.t0 304.64
R328 a_27_392.n1 a_27_392.n0 187.346
R329 a_27_392.n1 a_27_392.t2 29.5505
R330 a_27_392.t1 a_27_392.n1 29.5505
R331 a_707_119.t1 a_707_119.n1 230.558
R332 a_707_119.n1 a_707_119.t3 218.279
R333 a_707_119.n1 a_707_119.n0 89.2272
R334 a_707_119.n0 a_707_119.t2 39.3755
R335 a_707_119.n0 a_707_119.t0 26.2505
C0 VPWR VPB 0.270959f
C1 B COUT 5.75e-20
C2 VPB A 0.188468f
C3 VPWR A 0.060623f
C4 VGND VPB 0.015017f
C5 B SUM 2.85e-19
C6 VPWR VGND 0.142873f
C7 COUT VPB 0.006592f
C8 VGND A 0.18421f
C9 VPWR COUT 0.044117f
C10 SUM VPB 0.022145f
C11 COUT A 8.94e-19
C12 VPWR SUM 0.391252f
C13 VGND COUT 0.195627f
C14 SUM A 5.26e-19
C15 VGND SUM 0.329708f
C16 COUT SUM 0.018187f
C17 B VPB 0.493329f
C18 B VPWR 0.145786f
C19 B A 0.187524f
C20 B VGND 0.030482f
C21 SUM VNB 0.084084f
C22 COUT VNB 0.017775f
C23 VGND VNB 1.1907f
C24 VPWR VNB 0.928702f
C25 B VNB 0.418703f
C26 A VNB 0.884773f
C27 VPB VNB 2.34601f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2_4 VNB VPB VPWR VGND Y B A
X0 Y.t7 A.t0 a_27_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X1 Y.t0 B.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.6216 pd=2.23 as=0.336 ps=2.84 w=1.12 l=0.15
X2 VPWR.t1 A.t1 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.7532 ps=2.465 w=1.12 l=0.15
X3 Y.t6 A.t2 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.15355 pd=1.155 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 Y.t3 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.7532 pd=2.465 as=0.196 ps=1.47 w=1.12 l=0.15
X5 VGND.t3 B.t1 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_27_74.t3 A.t4 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1147 ps=1.05 w=0.74 l=0.15
X7 VPWR.t2 B.t2 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.6216 ps=2.23 w=1.12 l=0.15
X8 a_27_74.t1 B.t3 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_27_74.t2 A.t5 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2442 pd=2.14 as=0.15355 ps=1.155 w=0.74 l=0.15
X10 a_27_74.t7 B.t4 VGND.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VGND.t0 B.t5 a_27_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t1 226.809
R1 A.n3 A.t3 226.809
R2 A.n3 A.t0 198.204
R3 A.n0 A.t5 198.204
R4 A.n2 A.t4 196.013
R5 A.n8 A.t2 196.013
R6 A A.n1 155.423
R7 A.n10 A.n9 152
R8 A.n7 A.n6 152
R9 A.n5 A.n4 152
R10 A.n9 A.n1 49.6611
R11 A.n4 A.n3 49.6611
R12 A.n8 A.n7 38.7066
R13 A.n7 A.n2 34.3247
R14 A.n1 A.n0 19.7187
R15 A.n4 A.n2 15.3369
R16 A.n9 A.n8 10.955
R17 A.n6 A.n5 10.1214
R18 A.n10 A 7.5912
R19 A A.n10 6.69817
R20 A.n6 A 2.53073
R21 A.n5 A 1.63771
R22 a_27_74.n2 a_27_74.t2 283.353
R23 a_27_74.t0 a_27_74.n5 210.411
R24 a_27_74.n2 a_27_74.n1 185
R25 a_27_74.n5 a_27_74.n0 103.65
R26 a_27_74.n4 a_27_74.n3 87.0786
R27 a_27_74.n5 a_27_74.n4 75.8546
R28 a_27_74.n4 a_27_74.n2 74.0928
R29 a_27_74.n1 a_27_74.t3 34.0546
R30 a_27_74.n3 a_27_74.t5 29.1897
R31 a_27_74.n3 a_27_74.t1 22.7032
R32 a_27_74.n1 a_27_74.t4 22.7032
R33 a_27_74.n0 a_27_74.t6 22.7032
R34 a_27_74.n0 a_27_74.t7 22.7032
R35 Y.n11 Y.n9 251.626
R36 Y.n3 Y.n1 195
R37 Y.n5 Y.n4 195
R38 Y.n6 Y.n0 195
R39 Y.n8 Y.n7 195
R40 Y.n11 Y.n10 185
R41 Y.n3 Y.n2 98.8947
R42 Y.n2 Y.t0 80.0499
R43 Y.n2 Y.t1 77.7787
R44 Y.n6 Y.n5 62.4425
R45 Y.n7 Y.n6 60.6835
R46 Y.n5 Y.n1 60.6835
R47 Y Y.n8 46.9492
R48 Y.n10 Y.t6 37.2978
R49 Y Y.n11 30.1314
R50 Y.n10 Y.t4 30.0005
R51 Y.n9 Y.t7 27.5681
R52 Y.n7 Y.t2 26.3844
R53 Y.n1 Y.t3 26.3844
R54 Y.n9 Y.t5 22.7032
R55 Y.n4 Y.n0 4.41215
R56 Y.n8 Y.n0 4.28788
R57 Y.n4 Y.n3 4.28788
R58 VNB.t4 VNB.t2 1304.99
R59 VNB.t3 VNB.t4 1154.86
R60 VNB VNB.t0 1143.31
R61 VNB.t1 VNB.t5 1085.56
R62 VNB.t5 VNB.t3 1062.47
R63 VNB.t6 VNB.t1 993.177
R64 VNB.t7 VNB.t6 993.177
R65 VNB.t0 VNB.t7 993.177
R66 B.n0 B.t2 226.809
R67 B.n3 B.t0 226.809
R68 B.n3 B.t1 198.204
R69 B.n0 B.t3 198.204
R70 B.n7 B.t5 196.013
R71 B.n2 B.t4 196.013
R72 B.n5 B.n4 165.189
R73 B.n5 B.n1 152
R74 B.n9 B.n8 152
R75 B.n7 B.n6 152
R76 B.n8 B.n7 49.6611
R77 B.n7 B.n1 49.6611
R78 B.n4 B.n2 36.5157
R79 B.n4 B.n3 24.1005
R80 B.n2 B.n1 13.146
R81 B B.n9 11.3121
R82 B.n8 B.n0 10.955
R83 B.n6 B 7.14469
R84 B.n6 B 7.14469
R85 B B.n5 3.60867
R86 B.n9 B 2.97724
R87 VPWR.n4 VPWR.t1 358.829
R88 VPWR.n3 VPWR.n2 316.259
R89 VPWR.n9 VPWR.t3 250.651
R90 VPWR.n7 VPWR.n1 36.1417
R91 VPWR.n8 VPWR.n7 36.1417
R92 VPWR.n2 VPWR.t0 35.1791
R93 VPWR.n2 VPWR.t2 26.3844
R94 VPWR.n9 VPWR.n8 20.7064
R95 VPWR.n3 VPWR.n1 11.2946
R96 VPWR.n5 VPWR.n1 9.3005
R97 VPWR.n7 VPWR.n6 9.3005
R98 VPWR.n8 VPWR.n0 9.3005
R99 VPWR.n10 VPWR.n9 9.3005
R100 VPWR.n4 VPWR.n3 7.63859
R101 VPWR.n5 VPWR.n4 0.161319
R102 VPWR.n6 VPWR.n5 0.122949
R103 VPWR.n6 VPWR.n0 0.122949
R104 VPWR.n10 VPWR.n0 0.122949
R105 VPWR VPWR.n10 0.0617245
R106 VPB.t0 VPB.t1 763.576
R107 VPB.t3 VPB.t2 643.548
R108 VPB VPB.t3 260.485
R109 VPB.t2 VPB.t0 255.376
R110 VGND.n2 VGND.n0 214.661
R111 VGND.n2 VGND.n1 214.655
R112 VGND.n0 VGND.t2 22.7032
R113 VGND.n0 VGND.t0 22.7032
R114 VGND.n1 VGND.t1 22.7032
R115 VGND.n1 VGND.t3 22.7032
R116 VGND VGND.n2 0.597443
C0 Y VGND 0.031583f
C1 VPB Y 0.027359f
C2 B Y 0.169794f
C3 VPB VGND 0.007548f
C4 B VGND 0.069379f
C5 A Y 0.383629f
C6 VPB B 0.122713f
C7 A VGND 0.024408f
C8 VPWR Y 0.614609f
C9 VPB A 0.133753f
C10 VPWR VGND 0.069325f
C11 VPB VPWR 0.134016f
C12 B A 0.099561f
C13 B VPWR 0.05101f
C14 A VPWR 0.039892f
C15 VGND VNB 0.516664f
C16 Y VNB 0.07344f
C17 VPWR VNB 0.490387f
C18 A VNB 0.404593f
C19 B VNB 0.391908f
C20 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2_2 VNB VPB VPWR VGND Y B A
X0 VPWR.t1 A.t0 Y.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t1 A.t1 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t2 A.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X3 Y.t5 B.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4 VGND.t1 B.t1 a_27_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 VPWR.t2 B.t2 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_27_74.t3 B.t3 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X7 a_27_74.t0 A.t3 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=2.09 as=0.1221 ps=1.07 w=0.74 l=0.15
R0 A.n0 A.t0 226.809
R1 A.n1 A.t2 226.809
R2 A.n1 A.t1 198.204
R3 A.n0 A.t3 198.204
R4 A A.n2 154.522
R5 A.n2 A.n1 33.5944
R6 A.n2 A.n0 32.1338
R7 Y.n2 Y.n1 270.894
R8 Y Y.n3 220.093
R9 Y.n2 Y.n0 208.897
R10 Y Y.n2 55.4399
R11 Y.n3 Y.t0 30.8113
R12 Y.n0 Y.t3 26.3844
R13 Y.n0 Y.t2 26.3844
R14 Y.n1 Y.t4 26.3844
R15 Y.n1 Y.t5 26.3844
R16 Y.n3 Y.t1 22.7032
R17 VPWR.n1 VPWR.t1 348.793
R18 VPWR.n3 VPWR.n2 315.928
R19 VPWR.n5 VPWR.t3 259.171
R20 VPWR.n2 VPWR.t0 28.1434
R21 VPWR.n2 VPWR.t2 26.3844
R22 VPWR.n5 VPWR.n4 26.3534
R23 VPWR.n4 VPWR.n3 22.5887
R24 VPWR.n4 VPWR.n0 9.3005
R25 VPWR.n6 VPWR.n5 9.3005
R26 VPWR.n3 VPWR.n1 6.65145
R27 VPWR.n1 VPWR.n0 0.677131
R28 VPWR.n6 VPWR.n0 0.122949
R29 VPWR VPWR.n6 0.0617245
R30 VPB VPB.t3 260.485
R31 VPB.t2 VPB.t0 234.946
R32 VPB.t0 VPB.t1 229.839
R33 VPB.t3 VPB.t2 229.839
R34 a_27_74.n0 a_27_74.t0 300.735
R35 a_27_74.n0 a_27_74.t2 233.084
R36 a_27_74.n1 a_27_74.n0 84.741
R37 a_27_74.t1 a_27_74.n1 22.7032
R38 a_27_74.n1 a_27_74.t3 22.7032
R39 VNB VNB.t2 1143.31
R40 VNB.t1 VNB.t0 1108.66
R41 VNB.t2 VNB.t3 1108.66
R42 VNB.t3 VNB.t1 993.177
R43 B.n0 B.t2 226.809
R44 B.n1 B.t0 226.809
R45 B.n1 B.t1 198.204
R46 B.n0 B.t3 198.204
R47 B.n3 B.n2 152
R48 B.n2 B.n1 37.9763
R49 B.n2 B.n0 27.752
R50 B B.n3 10.2703
R51 B.n3 B 4.0191
R52 VGND VGND.n0 214.124
R53 VGND.n0 VGND.t0 30.8113
R54 VGND.n0 VGND.t1 22.7032
C0 B A 0.09794f
C1 B VPWR 0.040599f
C2 B VPB 0.065844f
C3 B Y 0.087085f
C4 A VPWR 0.039637f
C5 A VPB 0.063501f
C6 B VGND 0.036647f
C7 A Y 0.15934f
C8 VPWR VPB 0.085694f
C9 A VGND 0.012584f
C10 VPWR Y 0.377948f
C11 Y VPB 0.012275f
C12 VPWR VGND 0.040991f
C13 VGND VPB 0.005423f
C14 Y VGND 0.01404f
C15 VGND VNB 0.319892f
C16 Y VNB 0.074709f
C17 VPWR VNB 0.33234f
C18 A VNB 0.220242f
C19 B VNB 0.238522f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2_1 VNB VPB VPWR VGND B Y A
X0 a_117_74.t0 B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VPWR.t1 A.t0 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t1 A.t1 a_117_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3 Y.t0 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
R0 B.n0 B.t1 278.188
R1 B.n0 B.t0 170.81
R2 B B.n0 158.788
R3 VGND VGND.t0 166.618
R4 a_117_74.t0 a_117_74.t1 38.9194
R5 VNB VNB.t0 1177.95
R6 VNB.t0 VNB.t1 900.788
R7 A.n0 A.t0 277.214
R8 A.n0 A.t1 169.834
R9 A A.n0 158.788
R10 Y.n1 Y 591.957
R11 Y.n1 Y.n0 585
R12 Y.n2 Y.n1 585
R13 Y Y.t1 168.683
R14 Y.n1 Y.t2 26.3844
R15 Y.n1 Y.t0 26.3844
R16 Y Y.n2 18.644
R17 Y Y.n0 16.1396
R18 Y Y.n0 4.45267
R19 Y.n2 Y 1.94833
R20 VPWR.n0 VPWR.t1 256.714
R21 VPWR.n0 VPWR.t0 256.543
R22 VPWR VPWR.n0 0.625604
R23 VPB VPB.t0 252.823
R24 VPB.t0 VPB.t1 229.839
C0 Y VPB 0.006523f
C1 VPWR B 0.051044f
C2 VGND VPB 0.004689f
C3 Y B 0.055465f
C4 VPWR A 0.050796f
C5 VGND B 0.052533f
C6 Y A 0.097251f
C7 VGND A 0.014967f
C8 VPWR Y 0.224451f
C9 VPWR VGND 0.027464f
C10 Y VGND 0.081749f
C11 VPB B 0.039081f
C12 VPB A 0.040249f
C13 B A 0.061674f
C14 VPWR VPB 0.064491f
C15 VGND VNB 0.257375f
C16 Y VNB 0.064463f
C17 VPWR VNB 0.267241f
C18 A VNB 0.169029f
C19 B VNB 0.165458f
C20 VPB VNB 0.406224f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux4_4 VNB VPB VPWR VGND S1 A0 A1 A2 A3 S0 X
X0 VPWR.t4 S0.t0 a_758_306.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_509_392.t7 S1.t0 a_2199_74.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X2 a_1465_377.t1 S0.t1 a_1191_121# VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X3 VGND.t3 A2.t0 a_1278_121.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 a_116_392.t1 A1.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X5 a_509_392.t0 a_2489_347.t1 a_2199_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.224 ps=1.34 w=0.64 l=0.15
X6 a_1285_377# a_758_306.t2 a_1191_121# VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X7 a_2199_74.t1 a_2489_347.t2 a_1191_121# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.175 ps=1.35 w=1 l=0.15
X8 a_2199_74.t5 S1.t1 a_1191_121# VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.224 pd=1.34 as=0.166175 ps=1.255 w=0.64 l=0.15
X9 a_1278_121.t3 a_758_306.t3 a_1191_121# VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X10 VGND.t9 A3.t0 a_1450_121.t3 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X11 a_509_392.t9 a_758_306.t4 a_116_392.t3 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X12 a_1450_121.t2 A3.t1 VGND.t11 VNB.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X13 X.t5 a_2199_74.t8 VPWR.t7 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2044 ps=1.485 w=1.12 l=0.15
X14 a_116_392.t2 a_758_306.t5 a_509_392.t8 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1625 ps=1.325 w=1 l=0.15
X15 VPWR.t10 A3.t2 a_1285_377# VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X16 X.t2 a_2199_74.t9 VGND.t6 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VPWR.t5 A0.t0 a_296_392.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X18 a_1278_121.t0 A2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2887 ps=2.39 w=0.64 l=0.15
X19 VPWR.t2 A2.t2 a_1465_377.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.27525 pd=1.715 as=0.15 ps=1.3 w=1 l=0.15
X20 a_1465_377.t2 A2.t3 VPWR.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.44815 ps=3.23 w=1 l=0.15
X21 a_1191_121# a_758_306.t6 a_1278_121.t2 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X22 a_1191_121# a_2489_347.t3 a_2199_74.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X23 a_299_126.t1 A0.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1104 ps=0.985 w=0.64 l=0.15
X24 a_509_392.t3 S0.t2 a_114_126.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.104 ps=0.965 w=0.64 l=0.15
X25 a_509_392.t5 S0.t3 a_296_392.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.1625 ps=1.325 w=1 l=0.15
X26 VGND.t8 a_2199_74.t10 X.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 a_1285_377# A3.t3 VPWR.t11 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.27525 ps=1.715 w=1 l=0.15
X28 VPWR.t8 a_2199_74.t11 X.t4 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X29 a_296_392.t2 S0.t4 a_509_392.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.31 ps=2.62 w=1 l=0.15
X30 a_114_126.t2 S0.t5 a_509_392.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.31625 ps=2.58 w=0.64 l=0.15
X31 X.t0 a_2199_74.t12 VGND.t7 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=1.32 w=0.74 l=0.15
X32 a_296_392.t0 A0.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X33 VGND.t1 A0.t3 a_299_126.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.3525 pd=2.83 as=0.0896 ps=0.92 w=0.64 l=0.15
X34 a_1450_121.t1 S0.t6 a_1191_121# VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X35 VPWR.t1 A1.t1 a_116_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X36 a_2199_74.t6 S1.t2 a_509_392.t6 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X37 a_299_126.t3 a_758_306.t7 a_509_392.t11 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X38 a_2199_74.t3 a_2489_347.t4 a_509_392.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X39 VGND.t5 A1.t2 a_114_126.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1104 pd=0.985 as=0.0896 ps=0.92 w=0.64 l=0.15
X40 a_1191_121# S0.t7 a_1450_121.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2336 pd=2.01 as=0.0896 ps=0.92 w=0.64 l=0.15
X41 VPWR.t9 a_2199_74.t13 X.t3 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X42 a_114_126.t0 A1.t3 VGND.t10 VNB.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X43 a_509_392.t10 a_758_306.t8 a_299_126.t2 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X44 a_1191_121# S1.t3 a_2199_74.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.166175 pd=1.255 as=0.1824 ps=1.85 w=0.64 l=0.15
X45 VGND.t4 S0.t8 a_758_306.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X46 VPWR.t12 S1.t4 a_2489_347.t0 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.2044 pd=1.485 as=0.3696 ps=2.9 w=1.12 l=0.15
R0 S0.n10 S0.n1 1312.94
R1 S0.n1 S0.n0 594.467
R2 S0.t8 S0.t0 502.351
R3 S0.t2 S0.t3 456.265
R4 S0.t5 S0.t4 456.265
R5 S0.n0 S0.t5 364.714
R6 S0.n0 S0.t2 212.081
R7 S0.n3 S0.n2 207.529
R8 S0.n5 S0.t1 207.529
R9 S0.n5 S0.t6 164.02
R10 S0.n1 S0.t8 155.847
R11 S0.n11 S0.n10 152
R12 S0.n9 S0.n8 152
R13 S0.n7 S0.n6 152
R14 S0.n4 S0.t7 151.028
R15 S0.n10 S0.n9 49.6611
R16 S0.n6 S0.n5 30.6732
R17 S0.n6 S0.n4 21.1793
R18 S0.n9 S0.n3 14.6066
R19 S0.n4 S0.n3 13.8763
R20 S0.n8 S0.n7 12.8005
R21 S0.n11 S0 11.4829
R22 S0 S0.n11 6.58874
R23 S0.n7 S0 3.95344
R24 S0.n8 S0 1.31815
R25 a_758_306.t0 a_758_306.n9 252.774
R26 a_758_306.n9 a_758_306.n0 244.309
R27 a_758_306.n8 a_758_306.t5 243.797
R28 a_758_306.n0 a_758_306.t4 239.661
R29 a_758_306.n2 a_758_306.n1 223.595
R30 a_758_306.n4 a_758_306.t2 215.561
R31 a_758_306.n6 a_758_306.n5 168.798
R32 a_758_306.n7 a_758_306.t1 167.262
R33 a_758_306.n6 a_758_306.n3 165.189
R34 a_758_306.n8 a_758_306.t7 160.667
R35 a_758_306.n0 a_758_306.t8 160.667
R36 a_758_306.n5 a_758_306.t3 141.387
R37 a_758_306.n2 a_758_306.t6 141.387
R38 a_758_306.n0 a_758_306.n8 78.2118
R39 a_758_306.n7 a_758_306.n6 69.2711
R40 a_758_306.n3 a_758_306.n2 29.9429
R41 a_758_306.n4 a_758_306.n3 27.752
R42 a_758_306.n5 a_758_306.n4 5.11262
R43 a_758_306.n9 a_758_306.n7 1.71596
R44 VPWR.n43 VPWR.t6 905.35
R45 VPWR.n3 VPWR.t5 848.437
R46 VPWR.n41 VPWR.n40 644.101
R47 VPWR.n34 VPWR.t10 361.14
R48 VPWR.n19 VPWR.t8 359.074
R49 VPWR.n20 VPWR.t9 351.639
R50 VPWR.n68 VPWR.n2 323.158
R51 VPWR.n70 VPWR.t3 260.599
R52 VPWR.n55 VPWR.t4 250.081
R53 VPWR.n22 VPWR.n18 223.696
R54 VPWR.n40 VPWR.t11 47.2805
R55 VPWR.n40 VPWR.t2 47.2805
R56 VPWR.n57 VPWR.n56 36.1417
R57 VPWR.n57 VPWR.n5 36.1417
R58 VPWR.n61 VPWR.n5 36.1417
R59 VPWR.n62 VPWR.n61 36.1417
R60 VPWR.n63 VPWR.n62 36.1417
R61 VPWR.n49 VPWR.n48 36.1417
R62 VPWR.n50 VPWR.n49 36.1417
R63 VPWR.n50 VPWR.n8 36.1417
R64 VPWR.n54 VPWR.n8 36.1417
R65 VPWR.n44 VPWR.n42 36.1417
R66 VPWR.n26 VPWR.n16 36.1417
R67 VPWR.n27 VPWR.n26 36.1417
R68 VPWR.n28 VPWR.n27 36.1417
R69 VPWR.n28 VPWR.n14 36.1417
R70 VPWR.n32 VPWR.n14 36.1417
R71 VPWR.n33 VPWR.n32 36.1417
R72 VPWR.n35 VPWR.n33 36.1417
R73 VPWR.n39 VPWR.n12 36.1417
R74 VPWR.n18 VPWR.t7 35.1791
R75 VPWR.n48 VPWR.n10 32.3937
R76 VPWR.n22 VPWR.n21 31.2476
R77 VPWR.n2 VPWR.t0 29.5505
R78 VPWR.n2 VPWR.t1 29.5505
R79 VPWR.n18 VPWR.t12 29.0228
R80 VPWR.n69 VPWR.n68 28.2358
R81 VPWR.n67 VPWR.n3 27.4829
R82 VPWR.n56 VPWR.n55 27.1064
R83 VPWR.n70 VPWR.n69 26.7299
R84 VPWR.n63 VPWR.n3 25.977
R85 VPWR.n68 VPWR.n67 25.224
R86 VPWR.n44 VPWR.n43 22.0115
R87 VPWR.n21 VPWR.n20 21.4593
R88 VPWR.n55 VPWR.n54 20.3299
R89 VPWR.n35 VPWR.n34 18.824
R90 VPWR.n34 VPWR.n12 17.3181
R91 VPWR.n22 VPWR.n16 16.1887
R92 VPWR.n41 VPWR.n39 13.1184
R93 VPWR.n21 VPWR.n17 9.3005
R94 VPWR.n23 VPWR.n22 9.3005
R95 VPWR.n24 VPWR.n16 9.3005
R96 VPWR.n26 VPWR.n25 9.3005
R97 VPWR.n27 VPWR.n15 9.3005
R98 VPWR.n29 VPWR.n28 9.3005
R99 VPWR.n30 VPWR.n14 9.3005
R100 VPWR.n32 VPWR.n31 9.3005
R101 VPWR.n33 VPWR.n13 9.3005
R102 VPWR.n36 VPWR.n35 9.3005
R103 VPWR.n37 VPWR.n12 9.3005
R104 VPWR.n39 VPWR.n38 9.3005
R105 VPWR.n42 VPWR.n11 9.3005
R106 VPWR.n45 VPWR.n44 9.3005
R107 VPWR.n46 VPWR.n10 9.3005
R108 VPWR.n48 VPWR.n47 9.3005
R109 VPWR.n49 VPWR.n9 9.3005
R110 VPWR.n51 VPWR.n50 9.3005
R111 VPWR.n52 VPWR.n8 9.3005
R112 VPWR.n54 VPWR.n53 9.3005
R113 VPWR.n55 VPWR.n7 9.3005
R114 VPWR.n56 VPWR.n6 9.3005
R115 VPWR.n58 VPWR.n57 9.3005
R116 VPWR.n59 VPWR.n5 9.3005
R117 VPWR.n61 VPWR.n60 9.3005
R118 VPWR.n62 VPWR.n4 9.3005
R119 VPWR.n64 VPWR.n63 9.3005
R120 VPWR.n65 VPWR.n3 9.3005
R121 VPWR.n67 VPWR.n66 9.3005
R122 VPWR.n68 VPWR.n1 9.3005
R123 VPWR.n69 VPWR.n0 9.3005
R124 VPWR.n71 VPWR.n70 9.3005
R125 VPWR.n42 VPWR.n41 7.09488
R126 VPWR.n20 VPWR.n19 7.03723
R127 VPWR.n43 VPWR.n10 2.41828
R128 VPWR.n19 VPWR.n17 0.600107
R129 VPWR.n23 VPWR.n17 0.122949
R130 VPWR.n24 VPWR.n23 0.122949
R131 VPWR.n25 VPWR.n24 0.122949
R132 VPWR.n25 VPWR.n15 0.122949
R133 VPWR.n29 VPWR.n15 0.122949
R134 VPWR.n30 VPWR.n29 0.122949
R135 VPWR.n31 VPWR.n30 0.122949
R136 VPWR.n31 VPWR.n13 0.122949
R137 VPWR.n36 VPWR.n13 0.122949
R138 VPWR.n37 VPWR.n36 0.122949
R139 VPWR.n38 VPWR.n37 0.122949
R140 VPWR.n38 VPWR.n11 0.122949
R141 VPWR.n45 VPWR.n11 0.122949
R142 VPWR.n46 VPWR.n45 0.122949
R143 VPWR.n47 VPWR.n46 0.122949
R144 VPWR.n47 VPWR.n9 0.122949
R145 VPWR.n51 VPWR.n9 0.122949
R146 VPWR.n52 VPWR.n51 0.122949
R147 VPWR.n53 VPWR.n52 0.122949
R148 VPWR.n53 VPWR.n7 0.122949
R149 VPWR.n7 VPWR.n6 0.122949
R150 VPWR.n58 VPWR.n6 0.122949
R151 VPWR.n59 VPWR.n58 0.122949
R152 VPWR.n60 VPWR.n59 0.122949
R153 VPWR.n60 VPWR.n4 0.122949
R154 VPWR.n64 VPWR.n4 0.122949
R155 VPWR.n65 VPWR.n64 0.122949
R156 VPWR.n66 VPWR.n65 0.122949
R157 VPWR.n66 VPWR.n1 0.122949
R158 VPWR.n1 VPWR.n0 0.122949
R159 VPWR.n71 VPWR.n0 0.122949
R160 VPWR VPWR.n71 0.0617245
R161 VPB.t10 VPB.t13 789.114
R162 VPB.t5 VPB.t22 646.102
R163 VPB.t20 VPB.t7 618.011
R164 VPB.t12 VPB.t8 523.521
R165 VPB.t11 VPB.t16 515.861
R166 VPB.t15 VPB.t11 515.861
R167 VPB.t19 VPB.t18 485.216
R168 VPB.t16 VPB.t10 459.678
R169 VPB.t2 VPB.t21 321.774
R170 VPB.t22 VPB.t17 263.038
R171 VPB VPB.t4 257.93
R172 VPB.t6 VPB.t5 255.376
R173 VPB.t3 VPB.t6 255.376
R174 VPB.t7 VPB.t3 255.376
R175 VPB.t0 VPB.t12 255.376
R176 VPB.t9 VPB.t14 242.608
R177 VPB.t8 VPB.t9 242.608
R178 VPB.t17 VPB.t19 229.839
R179 VPB.t21 VPB.t20 229.839
R180 VPB.t13 VPB.t2 229.839
R181 VPB.t14 VPB.t15 229.839
R182 VPB.t1 VPB.t0 229.839
R183 VPB.t4 VPB.t1 229.839
R184 S1.n5 S1.n1 325.897
R185 S1.n4 S1.t2 281.168
R186 S1.n2 S1.t0 281.168
R187 S1.n1 S1.t4 272.062
R188 S1.n2 S1.t3 204.339
R189 S1 S1.n4 201.008
R190 S1.n3 S1.t1 162.274
R191 S1.n1 S1.n0 154.24
R192 S1.n3 S1.n2 59.8853
R193 S1.n4 S1.n3 13.146
R194 S1 S1.n5 4.14168
R195 S1.n5 S1 0.760896
R196 a_2199_74.n19 a_2199_74.t7 317.235
R197 a_2199_74.n18 a_2199_74.t1 300.916
R198 a_2199_74.n18 a_2199_74.n17 288.351
R199 a_2199_74.n12 a_2199_74.t8 282.481
R200 a_2199_74.n5 a_2199_74.t11 240.197
R201 a_2199_74.n9 a_2199_74.n3 240.197
R202 a_2199_74.n11 a_2199_74.t13 240.197
R203 a_2199_74.n20 a_2199_74.t4 211.25
R204 a_2199_74.n5 a_2199_74.t10 193.093
R205 a_2199_74.n22 a_2199_74.n21 185
R206 a_2199_74.n16 a_2199_74.n0 185
R207 a_2199_74.n10 a_2199_74.n2 179.947
R208 a_2199_74.n12 a_2199_74.t12 179.947
R209 a_2199_74.n4 a_2199_74.t9 179.947
R210 a_2199_74.n7 a_2199_74.n6 165.189
R211 a_2199_74.n14 a_2199_74.n13 152
R212 a_2199_74.n10 a_2199_74.n1 152
R213 a_2199_74.n8 a_2199_74.n7 152
R214 a_2199_74.n15 a_2199_74.n14 150.006
R215 a_2199_74.n15 a_2199_74.t3 130.536
R216 a_2199_74.n19 a_2199_74.n18 72.0568
R217 a_2199_74.n22 a_2199_74.n0 65.6255
R218 a_2199_74.n21 a_2199_74.n20 60.9848
R219 a_2199_74.n20 a_2199_74.n19 58.0354
R220 a_2199_74.n16 a_2199_74.n15 56.2339
R221 a_2199_74.n10 a_2199_74.n9 46.7399
R222 a_2199_74.n17 a_2199_74.t6 39.4005
R223 a_2199_74.n0 a_2199_74.t0 39.3755
R224 a_2199_74.n6 a_2199_74.n4 36.5157
R225 a_2199_74.n17 a_2199_74.t2 29.5505
R226 a_2199_74.n11 a_2199_74.n10 26.2914
R227 a_2199_74.t5 a_2199_74.n22 26.2505
R228 a_2199_74.n13 a_2199_74.n11 23.3702
R229 a_2199_74.n7 a_2199_74.n1 13.1884
R230 a_2199_74.n14 a_2199_74.n1 13.1884
R231 a_2199_74.n6 a_2199_74.n5 13.146
R232 a_2199_74.n8 a_2199_74.n4 13.146
R233 a_2199_74.n13 a_2199_74.n12 13.146
R234 a_2199_74.n21 a_2199_74.n16 12.2745
R235 a_2199_74.n9 a_2199_74.n8 2.92171
R236 a_509_392.n2 a_509_392.t4 864.72
R237 a_509_392.n9 a_509_392.n8 592.564
R238 a_509_392.n5 a_509_392.t2 415.664
R239 a_509_392.n8 a_509_392.n0 290.373
R240 a_509_392.n3 a_509_392.t9 218.837
R241 a_509_392.n5 a_509_392.n4 218.506
R242 a_509_392.n2 a_509_392.n1 209.275
R243 a_509_392.n6 a_509_392.t10 125.135
R244 a_509_392.n6 a_509_392.n5 73.3428
R245 a_509_392.n7 a_509_392.n6 69.532
R246 a_509_392.n3 a_509_392.n2 61.1633
R247 a_509_392.t7 a_509_392.n9 39.4005
R248 a_509_392.n1 a_509_392.t5 34.4755
R249 a_509_392.n1 a_509_392.t8 29.5505
R250 a_509_392.n9 a_509_392.t6 29.5505
R251 a_509_392.n4 a_509_392.t11 26.2505
R252 a_509_392.n4 a_509_392.t3 26.2505
R253 a_509_392.n0 a_509_392.t1 26.2505
R254 a_509_392.n0 a_509_392.t0 26.2505
R255 a_509_392.n8 a_509_392.n7 24.9278
R256 a_509_392.n7 a_509_392.n3 15.4798
R257 a_1465_377.t1 a_1465_377.n0 1389.24
R258 a_1465_377.n0 a_1465_377.t0 29.5505
R259 a_1465_377.n0 a_1465_377.t2 29.5505
R260 A2.n4 A2.t3 283.479
R261 A2.n2 A2.t2 263.762
R262 A2.n1 A2.t0 199.958
R263 A2.n3 A2.t1 183.161
R264 A2.n1 A2.n0 152
R265 A2.n5 A2.n4 152
R266 A2.n3 A2.n2 42.3581
R267 A2.n5 A2.n0 8.45099
R268 A2.n2 A2.n1 3.65202
R269 A2.n4 A2.n3 3.65202
R270 A2 A2.n5 3.35584
R271 A2.n0 A2 0.124772
R272 a_1278_121.n1 a_1278_121.n0 577.172
R273 a_1278_121.n0 a_1278_121.t1 26.2505
R274 a_1278_121.n0 a_1278_121.t0 26.2505
R275 a_1278_121.t2 a_1278_121.n1 26.2505
R276 a_1278_121.n1 a_1278_121.t3 26.2505
R277 VGND.n62 VGND.t1 414.019
R278 VGND.n42 VGND.t2 308.827
R279 VGND.n17 VGND.t6 239.703
R280 VGND.n16 VGND.t8 238.587
R281 VGND.n36 VGND.n35 213.161
R282 VGND.n5 VGND.t4 164.077
R283 VGND.n34 VGND.t9 160.042
R284 VGND.n15 VGND.t7 156.047
R285 VGND.n69 VGND.n68 142.571
R286 VGND.n69 VGND.t10 124.615
R287 VGND.n70 VGND.n69 47.0773
R288 VGND.n22 VGND.n21 36.1417
R289 VGND.n23 VGND.n22 36.1417
R290 VGND.n23 VGND.n13 36.1417
R291 VGND.n27 VGND.n13 36.1417
R292 VGND.n28 VGND.n27 36.1417
R293 VGND.n29 VGND.n28 36.1417
R294 VGND.n29 VGND.n11 36.1417
R295 VGND.n33 VGND.n11 36.1417
R296 VGND.n41 VGND.n9 36.1417
R297 VGND.n44 VGND.n43 36.1417
R298 VGND.n44 VGND.n7 36.1417
R299 VGND.n48 VGND.n7 36.1417
R300 VGND.n49 VGND.n48 36.1417
R301 VGND.n50 VGND.n49 36.1417
R302 VGND.n55 VGND.n54 36.1417
R303 VGND.n56 VGND.n55 36.1417
R304 VGND.n56 VGND.n3 36.1417
R305 VGND.n60 VGND.n3 36.1417
R306 VGND.n61 VGND.n60 36.1417
R307 VGND.n66 VGND.n1 36.1417
R308 VGND.n67 VGND.n66 36.1417
R309 VGND.n37 VGND.n34 34.2593
R310 VGND.n68 VGND.t0 32.813
R311 VGND.n68 VGND.t5 31.8755
R312 VGND.n18 VGND.n17 28.2358
R313 VGND.n70 VGND.n67 26.7299
R314 VGND.n35 VGND.t11 26.2505
R315 VGND.n35 VGND.t3 26.2505
R316 VGND.n54 VGND.n5 25.224
R317 VGND.n62 VGND.n61 24.8476
R318 VGND.n18 VGND.n15 24.0946
R319 VGND.n62 VGND.n1 22.5887
R320 VGND.n50 VGND.n5 22.2123
R321 VGND.n34 VGND.n33 19.2005
R322 VGND.n21 VGND.n15 12.0476
R323 VGND.n37 VGND.n36 11.6711
R324 VGND.n43 VGND.n42 11.4201
R325 VGND.n71 VGND.n70 9.3005
R326 VGND.n19 VGND.n18 9.3005
R327 VGND.n21 VGND.n20 9.3005
R328 VGND.n22 VGND.n14 9.3005
R329 VGND.n24 VGND.n23 9.3005
R330 VGND.n25 VGND.n13 9.3005
R331 VGND.n27 VGND.n26 9.3005
R332 VGND.n28 VGND.n12 9.3005
R333 VGND.n30 VGND.n29 9.3005
R334 VGND.n31 VGND.n11 9.3005
R335 VGND.n33 VGND.n32 9.3005
R336 VGND.n34 VGND.n10 9.3005
R337 VGND.n38 VGND.n37 9.3005
R338 VGND.n39 VGND.n9 9.3005
R339 VGND.n41 VGND.n40 9.3005
R340 VGND.n43 VGND.n8 9.3005
R341 VGND.n45 VGND.n44 9.3005
R342 VGND.n46 VGND.n7 9.3005
R343 VGND.n48 VGND.n47 9.3005
R344 VGND.n49 VGND.n6 9.3005
R345 VGND.n51 VGND.n50 9.3005
R346 VGND.n52 VGND.n5 9.3005
R347 VGND.n54 VGND.n53 9.3005
R348 VGND.n55 VGND.n4 9.3005
R349 VGND.n57 VGND.n56 9.3005
R350 VGND.n58 VGND.n3 9.3005
R351 VGND.n60 VGND.n59 9.3005
R352 VGND.n61 VGND.n2 9.3005
R353 VGND.n63 VGND.n62 9.3005
R354 VGND.n64 VGND.n1 9.3005
R355 VGND.n66 VGND.n65 9.3005
R356 VGND.n67 VGND.n0 9.3005
R357 VGND.n42 VGND.n41 8.40834
R358 VGND.n17 VGND.n16 6.70714
R359 VGND.n36 VGND.n9 5.64756
R360 VGND.n19 VGND.n16 0.645862
R361 VGND.n20 VGND.n19 0.122949
R362 VGND.n20 VGND.n14 0.122949
R363 VGND.n24 VGND.n14 0.122949
R364 VGND.n25 VGND.n24 0.122949
R365 VGND.n26 VGND.n25 0.122949
R366 VGND.n26 VGND.n12 0.122949
R367 VGND.n30 VGND.n12 0.122949
R368 VGND.n31 VGND.n30 0.122949
R369 VGND.n32 VGND.n31 0.122949
R370 VGND.n32 VGND.n10 0.122949
R371 VGND.n38 VGND.n10 0.122949
R372 VGND.n39 VGND.n38 0.122949
R373 VGND.n40 VGND.n39 0.122949
R374 VGND.n40 VGND.n8 0.122949
R375 VGND.n45 VGND.n8 0.122949
R376 VGND.n46 VGND.n45 0.122949
R377 VGND.n47 VGND.n46 0.122949
R378 VGND.n47 VGND.n6 0.122949
R379 VGND.n51 VGND.n6 0.122949
R380 VGND.n52 VGND.n51 0.122949
R381 VGND.n53 VGND.n52 0.122949
R382 VGND.n53 VGND.n4 0.122949
R383 VGND.n57 VGND.n4 0.122949
R384 VGND.n58 VGND.n57 0.122949
R385 VGND.n59 VGND.n58 0.122949
R386 VGND.n59 VGND.n2 0.122949
R387 VGND.n63 VGND.n2 0.122949
R388 VGND.n64 VGND.n63 0.122949
R389 VGND.n65 VGND.n64 0.122949
R390 VGND.n65 VGND.n0 0.122949
R391 VGND.n71 VGND.n0 0.122949
R392 VGND VGND.n71 0.0617245
R393 VNB.t5 VNB.t14 4134.38
R394 VNB.t7 VNB.t2 3118.11
R395 VNB.t1 VNB.t9 2656.17
R396 VNB.t21 VNB.t11 2563.78
R397 VNB.t6 VNB.t20 2286.61
R398 VNB.t17 VNB.t6 2286.61
R399 VNB.t14 VNB.t16 1986.35
R400 VNB.t12 VNB.t4 1963.25
R401 VNB.t11 VNB.t12 1362.73
R402 VNB.t13 VNB.t0 1143.31
R403 VNB VNB.t22 1143.31
R404 VNB.t9 VNB.t10 1097.11
R405 VNB.t16 VNB.t15 993.177
R406 VNB.t4 VNB.t5 993.177
R407 VNB.t23 VNB.t21 993.177
R408 VNB.t3 VNB.t23 993.177
R409 VNB.t2 VNB.t3 993.177
R410 VNB.t8 VNB.t7 993.177
R411 VNB.t19 VNB.t8 993.177
R412 VNB.t20 VNB.t19 993.177
R413 VNB.t18 VNB.t17 993.177
R414 VNB.t10 VNB.t18 993.177
R415 VNB.t0 VNB.t1 993.177
R416 VNB.t22 VNB.t13 993.177
R417 A1.n0 A1.t1 217.266
R418 A1.n2 A1.t0 212.883
R419 A1.n4 A1.n3 168.067
R420 A1.n3 A1.t3 160.667
R421 A1.n0 A1.t2 160.667
R422 A1 A1.n1 155.492
R423 A1.n2 A1.n1 32.1338
R424 A1.n1 A1.n0 29.2126
R425 A1 A1.n4 9.69747
R426 A1.n4 A1 8.92171
R427 A1.n3 A1.n2 1.46111
R428 a_116_392.n1 a_116_392.n0 787.687
R429 a_116_392.n0 a_116_392.t3 29.5505
R430 a_116_392.n0 a_116_392.t2 29.5505
R431 a_116_392.n1 a_116_392.t0 29.5505
R432 a_116_392.t1 a_116_392.n1 29.5505
R433 a_2489_347.t0 a_2489_347.n2 442.974
R434 a_2489_347.n2 a_2489_347.t4 257.61
R435 a_2489_347.n0 a_2489_347.t3 252.924
R436 a_2489_347.n0 a_2489_347.t1 250.641
R437 a_2489_347.n1 a_2489_347.t2 184.768
R438 a_2489_347.n1 a_2489_347.n0 27.8752
R439 a_2489_347.n2 a_2489_347.n1 15.0993
R440 A3.n2 A3.t1 251.37
R441 A3.n0 A3.t0 226.696
R442 A3.n0 A3.t2 214.881
R443 A3.n2 A3.t3 214.222
R444 A3 A3.n1 152.388
R445 A3.n4 A3.n3 152
R446 A3.n3 A3.n1 49.6611
R447 A3 A3.n4 12.8005
R448 A3.n1 A3.n0 10.9788
R449 A3.n4 A3 5.81868
R450 A3.n3 A3.n2 4.38232
R451 a_1450_121.n1 a_1450_121.n0 469.649
R452 a_1450_121.n0 a_1450_121.t3 26.2505
R453 a_1450_121.n0 a_1450_121.t2 26.2505
R454 a_1450_121.n1 a_1450_121.t0 26.2505
R455 a_1450_121.t1 a_1450_121.n1 26.2505
R456 X.n1 X.n0 254.282
R457 X.n1 X.t4 233.983
R458 X.n3 X.t0 196.274
R459 X.n3 X.n2 102.019
R460 X X.n1 38.8097
R461 X X.n3 29.5125
R462 X.n0 X.t3 26.3844
R463 X.n0 X.t5 26.3844
R464 X.n2 X.t1 22.7032
R465 X.n2 X.t2 22.7032
R466 A0.n1 A0.t2 209.72
R467 A0.n0 A0.t0 207.529
R468 A0 A0.n0 198.089
R469 A0.n4 A0.t3 167.094
R470 A0.n1 A0.t1 167.094
R471 A0.n5 A0.n4 152
R472 A0.n3 A0.n2 152
R473 A0.n4 A0.n3 49.6611
R474 A0.n2 A0 15.3217
R475 A0.n3 A0.n1 13.146
R476 A0.n5 A0 9.89141
R477 A0 A0.n5 8.72777
R478 A0.n4 A0.n0 8.03383
R479 A0.n2 A0 3.29747
R480 a_296_392.n1 a_296_392.n0 682.574
R481 a_296_392.n1 a_296_392.t0 39.4005
R482 a_296_392.n0 a_296_392.t3 34.4755
R483 a_296_392.n0 a_296_392.t2 29.5505
R484 a_296_392.t1 a_296_392.n1 29.5505
R485 a_299_126.n1 a_299_126.n0 457.125
R486 a_299_126.n0 a_299_126.t2 26.2505
R487 a_299_126.n0 a_299_126.t3 26.2505
R488 a_299_126.n1 a_299_126.t0 26.2505
R489 a_299_126.t1 a_299_126.n1 26.2505
R490 a_114_126.n1 a_114_126.n0 547.537
R491 a_114_126.n0 a_114_126.t3 34.688
R492 a_114_126.n0 a_114_126.t2 26.2505
R493 a_114_126.t1 a_114_126.n1 26.2505
R494 a_114_126.n1 a_114_126.t0 26.2505
C0 S0 VGND 0.17201f
C1 A3 a_1191_121# 0.109133f
C2 A2 a_1285_377# 0.019332f
C3 VPB VPWR 0.447531f
C4 A3 S1 0.019709f
C5 S0 X 6.08e-20
C6 A2 VGND 0.022766f
C7 A3 a_1285_377# 0.022776f
C8 S1 a_1191_121# 0.029549f
C9 a_1191_121# a_1285_377# 0.226151f
C10 VPB A1 0.089697f
C11 A3 VGND 0.040441f
C12 VGND a_1191_121# 0.272306f
C13 VPB A0 0.107707f
C14 VPWR A1 0.059104f
C15 S1 VGND 0.028579f
C16 VPB S0 0.219412f
C17 VPWR A0 0.03418f
C18 S1 X 1.92e-19
C19 VPWR S0 0.0429f
C20 VPB A2 0.091736f
C21 A1 A0 0.079935f
C22 VGND X 0.306569f
C23 VPWR A2 0.015375f
C24 VPB A3 0.08761f
C25 A1 S0 2.71e-20
C26 VPB a_1191_121# 0.075309f
C27 VPWR A3 0.015847f
C28 A0 S0 0.021477f
C29 VPB S1 0.159692f
C30 VPWR a_1191_121# 0.463618f
C31 VPB a_1285_377# 0.029289f
C32 VPB VGND 0.024389f
C33 VPWR S1 0.038753f
C34 VPWR a_1285_377# 0.451157f
C35 S0 A2 0.060155f
C36 VPWR VGND 0.149686f
C37 VPB X 0.016934f
C38 A0 a_1191_121# 1.21e-20
C39 S0 a_1191_121# 0.209976f
C40 VPWR X 0.45187f
C41 A1 VGND 0.10844f
C42 A2 A3 0.082686f
C43 S0 a_1285_377# 0.020539f
C44 A2 a_1191_121# 0.082952f
C45 A0 VGND 0.042844f
C46 X VNB 0.069926f
C47 VGND VNB 1.90515f
C48 S1 VNB 0.479905f
C49 A3 VNB 0.227743f
C50 A2 VNB 0.227348f
C51 S0 VNB 1.20927f
C52 A0 VNB 0.220905f
C53 A1 VNB 0.231687f
C54 VPWR VNB 1.5237f
C55 VPB VNB 3.83458f
C56 a_1191_121# VNB 0.072457f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux4_2 VNB VPB VPWR VGND X A0 A1 A3 S1 S0 A2
X0 a_1047_74.t0 a_31_94.t2 a_909_74.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2886 pd=1.52 as=0.1998 ps=1.28 w=0.74 l=0.15
X1 a_264_392.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.45 pd=1.9 as=0.225 ps=1.45 w=1 l=0.15
X2 a_840_392.t0 A3.t0 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.36 pd=1.72 as=0.27 ps=1.54 w=1 l=0.15
X3 VGND.t1 A0.t0 a_507_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=1.28 as=0.2886 ps=1.52 w=0.74 l=0.15
X4 a_333_74.t2 a_31_94.t3 a_264_392.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.285 pd=1.57 as=0.45 ps=1.9 w=1 l=0.15
X5 VPWR.t3 A2.t0 a_1152_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t4 S1.t0 a_1500_94.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3849 pd=1.855 as=0.425 ps=2.85 w=1 l=0.15
X7 X.t1 a_1429_74.t3 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3849 ps=1.855 w=1.12 l=0.15
X8 a_1152_392.t0 S0.t0 a_909_74.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.27 ps=1.54 w=1 l=0.15
X9 a_255_74.t0 A1.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.18545 ps=1.275 w=0.74 l=0.15
X10 VGND.t5 A2.t1 a_1047_74.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.2886 ps=1.52 w=0.74 l=0.15
X11 VPWR.t2 A0.t1 a_618_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.27 pd=1.54 as=0.135 ps=1.27 w=1 l=0.15
X12 a_333_74.t0 a_1500_94.t2 a_1429_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151475 ps=1.325 w=0.74 l=0.15
X13 VGND.t3 S0.t1 a_31_94.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.18545 pd=1.275 as=0.1824 ps=1.85 w=0.64 l=0.15
X14 a_618_392.t0 S0.t2 a_333_74.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.285 ps=1.57 w=1 l=0.15
X15 a_909_74.t5 S0.t3 a_831_74.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=1.28 as=0.0888 ps=0.98 w=0.74 l=0.15
X16 a_1429_74.t1 S1.t1 a_909_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.151475 pd=1.325 as=0.2072 ps=2.04 w=0.74 l=0.15
X17 VGND.t4 S1.t2 a_1500_94.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.25105 pd=1.48 as=0.276725 ps=2.15 w=0.64 l=0.15
X18 a_909_74.t2 a_31_94.t4 a_840_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.27 pd=1.54 as=0.36 ps=1.72 w=1 l=0.15
X19 a_831_74.t1 A3.t1 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1998 ps=1.28 w=0.74 l=0.15
X20 a_507_74.t1 a_31_94.t5 a_333_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2886 pd=1.52 as=0.2664 ps=1.46 w=0.74 l=0.15
X21 VGND.t6 a_1429_74.t4 X.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_909_74.t1 a_1500_94.t3 a_1429_74.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.15 ps=1.3 w=1 l=0.15
X23 VPWR.t1 S0.t4 a_31_94.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.45 as=0.295 ps=2.59 w=1 l=0.15
X24 a_333_74.t4 S0.t5 a_255_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2664 pd=1.46 as=0.0888 ps=0.98 w=0.74 l=0.15
R0 a_31_94.n3 a_31_94.t1 292.101
R1 a_31_94.n1 a_31_94.t5 265.392
R2 a_31_94.n0 a_31_94.t2 255.46
R3 a_31_94.t0 a_31_94.n3 241.308
R4 a_31_94.n1 a_31_94.t3 236.983
R5 a_31_94.n0 a_31_94.t4 236.619
R6 a_31_94.n2 a_31_94.n1 180.5
R7 a_31_94.n2 a_31_94.n0 179.206
R8 a_31_94.n3 a_31_94.n2 10.9135
R9 a_909_74.n3 a_909_74.n0 755.437
R10 a_909_74.n3 a_909_74.n2 334.969
R11 a_909_74.t1 a_909_74.n3 325.312
R12 a_909_74.n2 a_909_74.n1 213.696
R13 a_909_74.n2 a_909_74.t0 119.361
R14 a_909_74.n0 a_909_74.t4 53.1905
R15 a_909_74.n0 a_909_74.t2 53.1905
R16 a_909_74.n1 a_909_74.t5 50.2708
R17 a_909_74.n1 a_909_74.t3 37.2978
R18 a_1047_74.t0 a_1047_74.t1 126.487
R19 VNB.t6 VNB.t11 3048.82
R20 VNB.t1 VNB.t6 2621.52
R21 VNB.t9 VNB.t4 2263.52
R22 VNB.t8 VNB.t9 2148.03
R23 VNB.t7 VNB.t3 2148.03
R24 VNB.t10 VNB.t7 2009.45
R25 VNB.t12 VNB.t8 1593.7
R26 VNB.t3 VNB.t0 1593.7
R27 VNB.t5 VNB.t2 1582.15
R28 VNB VNB.t5 1189.5
R29 VNB.t4 VNB.t1 1166.4
R30 VNB.t0 VNB.t12 900.788
R31 VNB.t2 VNB.t10 900.788
R32 a_1429_74.t2 a_1429_74.n5 1030
R33 a_1429_74.n5 a_1429_74.n1 386.498
R34 a_1429_74.n4 a_1429_74.n3 238.386
R35 a_1429_74.n0 a_1429_74.t3 226.809
R36 a_1429_74.n5 a_1429_74.n0 207.504
R37 a_1429_74.n4 a_1429_74.t4 154.24
R38 a_1429_74.n0 a_1429_74.n2 154.24
R39 a_1429_74.n0 a_1429_74.n4 67.6266
R40 a_1429_74.n1 a_1429_74.t0 41.6348
R41 a_1429_74.n1 a_1429_74.t1 22.7032
R42 X.n1 X 589.572
R43 X.n1 X.n0 585
R44 X.n2 X.n1 585
R45 X.t0 X.n3 281.43
R46 X.n4 X.t0 281.43
R47 X.n1 X.t1 26.3844
R48 X.n2 X 12.2519
R49 X.n0 X 10.6062
R50 X.n3 X 9.89141
R51 X.n4 X 7.56414
R52 X X.n4 6.78838
R53 X.n3 X 4.46111
R54 X.n0 X 2.92621
R55 X X.n2 1.2805
R56 VPWR.n10 VPWR.t3 835.754
R57 VPWR.n5 VPWR.n4 315.928
R58 VPWR.n9 VPWR.n8 252.917
R59 VPWR.n28 VPWR.n1 222.359
R60 VPWR.n8 VPWR.t4 115.246
R61 VPWR.n4 VPWR.t6 53.1905
R62 VPWR.n4 VPWR.t2 53.1905
R63 VPWR.n1 VPWR.t0 49.2505
R64 VPWR.n1 VPWR.t1 39.4005
R65 VPWR.n21 VPWR.n20 36.1417
R66 VPWR.n22 VPWR.n21 36.1417
R67 VPWR.n22 VPWR.n2 36.1417
R68 VPWR.n26 VPWR.n2 36.1417
R69 VPWR.n27 VPWR.n26 36.1417
R70 VPWR.n11 VPWR.n7 36.1417
R71 VPWR.n15 VPWR.n7 36.1417
R72 VPWR.n16 VPWR.n15 36.1417
R73 VPWR.n17 VPWR.n16 36.1417
R74 VPWR.n8 VPWR.t5 25.5754
R75 VPWR.n11 VPWR.n10 12.424
R76 VPWR.n29 VPWR.n28 10.3391
R77 VPWR.n17 VPWR.n5 10.1652
R78 VPWR.n12 VPWR.n11 9.3005
R79 VPWR.n13 VPWR.n7 9.3005
R80 VPWR.n15 VPWR.n14 9.3005
R81 VPWR.n16 VPWR.n6 9.3005
R82 VPWR.n18 VPWR.n17 9.3005
R83 VPWR.n20 VPWR.n19 9.3005
R84 VPWR.n21 VPWR.n3 9.3005
R85 VPWR.n23 VPWR.n22 9.3005
R86 VPWR.n24 VPWR.n2 9.3005
R87 VPWR.n26 VPWR.n25 9.3005
R88 VPWR.n27 VPWR.n0 9.3005
R89 VPWR.n28 VPWR.n27 8.65932
R90 VPWR.n10 VPWR.n9 7.61447
R91 VPWR.n20 VPWR.n5 1.12991
R92 VPWR VPWR.n29 0.163644
R93 VPWR.n12 VPWR.n9 0.150248
R94 VPWR.n29 VPWR.n0 0.144205
R95 VPWR.n13 VPWR.n12 0.122949
R96 VPWR.n14 VPWR.n13 0.122949
R97 VPWR.n14 VPWR.n6 0.122949
R98 VPWR.n18 VPWR.n6 0.122949
R99 VPWR.n19 VPWR.n18 0.122949
R100 VPWR.n19 VPWR.n3 0.122949
R101 VPWR.n23 VPWR.n3 0.122949
R102 VPWR.n24 VPWR.n23 0.122949
R103 VPWR.n25 VPWR.n24 0.122949
R104 VPWR.n25 VPWR.n0 0.122949
R105 VPB.n0 VPB 4226.48
R106 VPB VPB.n1 3729.83
R107 VPB.t7 VPB.t0 536.29
R108 VPB.t8 VPB.t10 452.017
R109 VPB.t6 VPB.t11 444.356
R110 VPB.n1 VPB.t4 411.156
R111 VPB.t5 VPB.n0 369.745
R112 VPB.t2 VPB.t7 367.743
R113 VPB.n1 VPB.t5 367.046
R114 VPB.t9 VPB.t6 352.42
R115 VPB.t11 VPB.t3 352.42
R116 VPB.t1 VPB 329.435
R117 VPB.t0 VPB.t1 306.452
R118 VPB.n0 VPB.t8 229.839
R119 VPB.t4 VPB.t9 214.517
R120 VPB.t3 VPB.t2 214.517
R121 A1.n0 A1.t1 252.248
R122 A1.n0 A1.t0 237.143
R123 A1 A1.n0 153.319
R124 a_264_392.t0 a_264_392.t1 177.3
R125 A3.n0 A3.t1 252.248
R126 A3.n0 A3.t0 239.833
R127 A3 A3.n0 153.319
R128 a_840_392.t0 a_840_392.t1 141.84
R129 A0.n0 A0.t1 236.983
R130 A0.n0 A0.t0 215.44
R131 A0 A0.n0 153.358
R132 a_507_74.t0 a_507_74.t1 126.487
R133 VGND.n7 VGND.t5 301.404
R134 VGND.n11 VGND.t4 255.41
R135 VGND.n12 VGND.t6 183.728
R136 VGND.n1 VGND.n0 115.835
R137 VGND.n33 VGND.n32 108.447
R138 VGND.n0 VGND.t3 73.8826
R139 VGND.n32 VGND.t2 57.5681
R140 VGND.n12 VGND.n11 39.4932
R141 VGND.n15 VGND.n14 36.1417
R142 VGND.n16 VGND.n15 36.1417
R143 VGND.n16 VGND.n9 36.1417
R144 VGND.n20 VGND.n9 36.1417
R145 VGND.n21 VGND.n20 36.1417
R146 VGND.n22 VGND.n21 36.1417
R147 VGND.n26 VGND.n25 36.1417
R148 VGND.n27 VGND.n26 36.1417
R149 VGND.n27 VGND.n5 36.1417
R150 VGND.n31 VGND.n5 36.1417
R151 VGND.n34 VGND.n3 36.1417
R152 VGND.n38 VGND.n3 36.1417
R153 VGND.n39 VGND.n38 36.1417
R154 VGND.n40 VGND.n39 36.1417
R155 VGND.n32 VGND.t1 30.0005
R156 VGND.n34 VGND.n33 24.4711
R157 VGND.n0 VGND.t0 21.1849
R158 VGND.n42 VGND.n1 15.2332
R159 VGND.n33 VGND.n31 11.6711
R160 VGND.n25 VGND.n7 10.5417
R161 VGND.n41 VGND.n40 9.3005
R162 VGND.n39 VGND.n2 9.3005
R163 VGND.n38 VGND.n37 9.3005
R164 VGND.n36 VGND.n3 9.3005
R165 VGND.n35 VGND.n34 9.3005
R166 VGND.n33 VGND.n4 9.3005
R167 VGND.n31 VGND.n30 9.3005
R168 VGND.n29 VGND.n5 9.3005
R169 VGND.n28 VGND.n27 9.3005
R170 VGND.n26 VGND.n6 9.3005
R171 VGND.n25 VGND.n24 9.3005
R172 VGND.n23 VGND.n22 9.3005
R173 VGND.n21 VGND.n8 9.3005
R174 VGND.n20 VGND.n19 9.3005
R175 VGND.n18 VGND.n9 9.3005
R176 VGND.n17 VGND.n16 9.3005
R177 VGND.n15 VGND.n10 9.3005
R178 VGND.n14 VGND.n13 9.3005
R179 VGND.n40 VGND.n1 3.76521
R180 VGND.n13 VGND.n12 2.17006
R181 VGND.n14 VGND.n11 1.88285
R182 VGND.n22 VGND.n7 0.753441
R183 VGND VGND.n42 0.163644
R184 VGND.n42 VGND.n41 0.144205
R185 VGND.n13 VGND.n10 0.122949
R186 VGND.n17 VGND.n10 0.122949
R187 VGND.n18 VGND.n17 0.122949
R188 VGND.n19 VGND.n18 0.122949
R189 VGND.n19 VGND.n8 0.122949
R190 VGND.n23 VGND.n8 0.122949
R191 VGND.n24 VGND.n23 0.122949
R192 VGND.n24 VGND.n6 0.122949
R193 VGND.n28 VGND.n6 0.122949
R194 VGND.n29 VGND.n28 0.122949
R195 VGND.n30 VGND.n29 0.122949
R196 VGND.n30 VGND.n4 0.122949
R197 VGND.n35 VGND.n4 0.122949
R198 VGND.n36 VGND.n35 0.122949
R199 VGND.n37 VGND.n36 0.122949
R200 VGND.n37 VGND.n2 0.122949
R201 VGND.n41 VGND.n2 0.122949
R202 a_333_74.n1 a_333_74.t0 666.299
R203 a_333_74.n1 a_333_74.n0 270.142
R204 a_333_74.n2 a_333_74.n1 195
R205 a_333_74.n0 a_333_74.t4 67.2978
R206 a_333_74.n2 a_333_74.t2 57.1305
R207 a_333_74.t1 a_333_74.n2 55.1605
R208 a_333_74.n0 a_333_74.t3 49.46
R209 A2.n0 A2.t0 298.572
R210 A2.n0 A2.t1 178.34
R211 A2.n1 A2.n0 152
R212 A2 A2.n1 5.80515
R213 A2.n1 A2 5.2098
R214 a_1152_392.t0 a_1152_392.t1 53.1905
R215 S1.t1 S1.t2 893.308
R216 S1.t2 S1.t0 458.971
R217 S1.n1 S1.t1 252.248
R218 S1.n1 S1.n0 236.983
R219 S1 S1.n1 163.249
R220 a_1500_94.t1 a_1500_94.n1 660.734
R221 a_1500_94.n1 a_1500_94.t0 254.406
R222 a_1500_94.n0 a_1500_94.t3 212.883
R223 a_1500_94.n0 a_1500_94.t2 156.431
R224 a_1500_94.n1 a_1500_94.n0 137.923
R225 S0.n1 S0.t0 476.776
R226 S0.n2 S0.t2 408.894
R227 S0.n3 S0.t5 361.481
R228 S0.n1 S0.t3 330.341
R229 S0.n0 S0.t4 298.572
R230 S0.n3 S0.n2 173.512
R231 S0.n0 S0.t1 162.274
R232 S0 S0.n0 153.212
R233 S0.n2 S0.n1 101.93
R234 S0 S0.n3 56.146
R235 a_255_74.t0 a_255_74.t1 38.9194
R236 a_618_392.t0 a_618_392.t1 53.1905
R237 a_831_74.t0 a_831_74.t1 38.9194
C0 A2 S1 0.024569f
C1 A0 A3 0.079046f
C2 A2 VPWR 0.013201f
C3 VPB A2 0.044815f
C4 A2 VGND 0.015006f
C5 S1 VPWR 0.014502f
C6 VPB S1 0.087277f
C7 S0 A2 0.0982f
C8 S1 VGND 0.052691f
C9 VPB VPWR 0.284296f
C10 S0 S1 4.52e-20
C11 VPWR VGND 0.104693f
C12 S1 X 5.35e-19
C13 VPB VGND 0.020253f
C14 S0 VPWR 0.046519f
C15 VPWR X 0.22134f
C16 VPB S0 0.166933f
C17 A1 VPWR 0.032817f
C18 VPB X 0.006636f
C19 S0 VGND 0.339652f
C20 VGND X 0.159022f
C21 VPB A1 0.053284f
C22 A1 VGND 0.014959f
C23 A0 VPWR 0.010139f
C24 VPB A0 0.04157f
C25 S0 A1 0.159898f
C26 A0 VGND 0.019934f
C27 A3 VPWR 0.012331f
C28 S0 A0 0.123291f
C29 VPB A3 0.050925f
C30 A3 VGND 0.013699f
C31 S0 A3 0.089338f
C32 X VNB 0.024518f
C33 VGND VNB 1.26292f
C34 VPWR VNB 1.00209f
C35 S1 VNB 0.430804f
C36 A2 VNB 0.125123f
C37 A3 VNB 0.105202f
C38 A0 VNB 0.114103f
C39 A1 VNB 0.10812f
C40 S0 VNB 0.488342f
C41 VPB VNB 2.42543f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux4_1 VNB VPB VPWR VGND S0 A3 A2 A1 A0 S1 X
X0 a_342_74.t3 a_27_74.t2 a_264_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
X1 a_450_74.t0 S0.t0 a_342_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.24 pd=1.39 as=0.1248 ps=1.03 w=0.64 l=0.15
X2 VGND.t1 A1.t0 a_450_74.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1728 pd=1.18 as=0.24 ps=1.39 w=0.64 l=0.15
X3 a_768_74.t0 A2.t0 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1728 ps=1.18 w=0.64 l=0.15
X4 VGND.t4 A3.t0 a_979_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0768 ps=0.88 w=0.64 l=0.15
X5 a_1338_125# S1.t0 a_846_74# VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.454475 ps=3.19 w=0.64 l=0.15
X6 a_846_74# S0.t1 a_763_341.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.4275 pd=1.855 as=0.197625 ps=1.585 w=1 l=0.15
X7 VGND.t2 S0.t2 a_27_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.192 pd=1.24 as=0.1824 ps=1.85 w=0.64 l=0.15
X8 VPWR.t2 S1.t1 a_1396_99.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.336275 pd=1.76 as=0.345 ps=2.69 w=1 l=0.15
X9 X a_1338_125# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3472 pd=2.86 as=0.336275 ps=1.76 w=1.12 l=0.15
X10 a_342_74.t4 a_1396_99.t1 a_1338_125# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0928 ps=0.93 w=0.64 l=0.15
X11 X.t0 a_1338_125# VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1469 ps=1.16 w=0.74 l=0.15
X12 a_763_341.t0 A2.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.197625 pd=1.585 as=0.2756 ps=1.75 w=1 l=0.15
X13 a_264_74.t0 A0.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.192 ps=1.24 w=0.64 l=0.15
X14 a_537_341.t1 a_27_74.t3 a_342_74.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X15 a_255_341.t1 A0.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.405 pd=1.81 as=0.2293 ps=1.57 w=1 l=0.15
X16 a_846_74# a_27_74.t4 a_768_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.155 as=0.0768 ps=0.88 w=0.64 l=0.15
X17 a_342_74.t0 S0.t3 a_255_341.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.405 ps=1.81 w=1 l=0.15
X18 VPWR.t4 A1.t1 a_537_341.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2756 pd=1.75 as=0.18 ps=1.36 w=1 l=0.15
X19 VPWR.t5 S0.t4 a_27_74.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2293 pd=1.57 as=0.295 ps=2.59 w=1 l=0.15
X20 a_979_74.t1 S0.t5 a_846_74# VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1648 ps=1.155 w=0.64 l=0.15
X21 VPWR.t0 A3.t1 a_1065_387.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1065_387.t1 a_27_74.t5 a_846_74# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.4275 ps=1.855 w=1 l=0.15
R0 a_27_74.n0 a_27_74.t5 456.401
R1 a_27_74.n1 a_27_74.t3 421.673
R2 a_27_74.n2 a_27_74.t2 359.18
R3 a_27_74.n0 a_27_74.t4 314.274
R4 a_27_74.t0 a_27_74.n3 304.865
R5 a_27_74.n2 a_27_74.n1 139.957
R6 a_27_74.n3 a_27_74.t1 135.66
R7 a_27_74.n1 a_27_74.n0 100.802
R8 a_27_74.n3 a_27_74.n2 88.0946
R9 a_264_74.t0 a_264_74.t1 45.0005
R10 a_342_74.n1 a_342_74.t4 742.106
R11 a_342_74.n1 a_342_74.n0 254.529
R12 a_342_74.n2 a_342_74.n1 192.305
R13 a_342_74.n0 a_342_74.t3 46.8755
R14 a_342_74.n2 a_342_74.t2 29.5505
R15 a_342_74.t0 a_342_74.n2 29.5505
R16 a_342_74.n0 a_342_74.t1 26.2505
R17 VNB VNB.n0 9839.37
R18 VNB.t7 VNB.t6 4561.68
R19 VNB.t8 VNB.t11 3245.14
R20 VNB.t9 VNB.t2 2237.29
R21 VNB.t1 VNB.t3 1864.41
R22 VNB.t10 VNB.t9 1715.25
R23 VNB.t2 VNB.t5 1342.37
R24 VNB.n0 VNB.t0 1293.44
R25 VNB.t3 VNB 1230.51
R26 VNB.t11 VNB.t7 1016.27
R27 VNB.t4 VNB.t10 969.492
R28 VNB.t5 VNB.t1 969.492
R29 VNB.t0 VNB.t8 900.788
R30 VNB.n0 VNB.t4 261.017
R31 S0.n0 S0.t1 834.396
R32 S0.t4 S0.n0 686.314
R33 S0.t1 S0.t5 638.169
R34 S0.t3 S0.t0 457.632
R35 S0.n0 S0.t3 283.844
R36 S0.n1 S0.t4 265.769
R37 S0.n1 S0.t2 190.792
R38 S0 S0.n1 158.919
R39 a_450_74.t0 a_450_74.t1 140.625
R40 A1.n0 A1.t1 231.629
R41 A1.n0 A1.t0 192.8
R42 A1 A1.n0 159.758
R43 VGND.n23 VGND.n22 203.052
R44 VGND.n14 VGND.n13 185
R45 VGND.n5 VGND.t3 163.743
R46 VGND.n6 VGND.t4 150.758
R47 VGND.n22 VGND.t2 60.938
R48 VGND.n22 VGND.t0 51.563
R49 VGND.n13 VGND.t5 50.6255
R50 VGND.n13 VGND.t1 50.6255
R51 VGND.n8 VGND.n7 36.1417
R52 VGND.n8 VGND.n3 36.1417
R53 VGND.n16 VGND.n15 36.1417
R54 VGND.n16 VGND.n1 36.1417
R55 VGND.n20 VGND.n1 36.1417
R56 VGND.n21 VGND.n20 36.1417
R57 VGND.n12 VGND.n3 29.407
R58 VGND.n7 VGND.n6 16.5652
R59 VGND.n21 VGND.n0 9.3005
R60 VGND.n20 VGND.n19 9.3005
R61 VGND.n18 VGND.n1 9.3005
R62 VGND.n17 VGND.n16 9.3005
R63 VGND.n15 VGND.n2 9.3005
R64 VGND.n12 VGND.n11 9.3005
R65 VGND.n10 VGND.n3 9.3005
R66 VGND.n9 VGND.n8 9.3005
R67 VGND.n7 VGND.n4 9.3005
R68 VGND.n23 VGND.n21 8.28285
R69 VGND.n24 VGND.n23 7.65871
R70 VGND.n6 VGND.n5 7.46902
R71 VGND.n15 VGND.n14 5.31292
R72 VGND.n14 VGND.n12 3.01226
R73 VGND VGND.n24 0.16305
R74 VGND.n5 VGND.n4 0.152406
R75 VGND.n24 VGND.n0 0.144791
R76 VGND.n9 VGND.n4 0.122949
R77 VGND.n10 VGND.n9 0.122949
R78 VGND.n11 VGND.n10 0.122949
R79 VGND.n11 VGND.n2 0.122949
R80 VGND.n17 VGND.n2 0.122949
R81 VGND.n18 VGND.n17 0.122949
R82 VGND.n19 VGND.n18 0.122949
R83 VGND.n19 VGND.n0 0.122949
R84 A2.n0 A2.t1 231.629
R85 A2.n0 A2.t0 192.8
R86 A2 A2.n0 158.919
R87 a_768_74.t0 a_768_74.t1 45.0005
R88 A3.n0 A3.t0 293.514
R89 A3.n0 A3.t1 223.55
R90 A3 A3.n0 155.821
R91 a_979_74.t0 a_979_74.t1 45.0005
R92 S1.n1 S1.t0 1002.56
R93 S1.t0 S1.n0 448.901
R94 S1.n2 S1.t1 257.067
R95 S1.n2 S1.n1 187.981
R96 S1 S1.n2 154.522
R97 a_763_341.t0 a_763_341.t1 81.0265
R98 VPB.t9 VPB 2168.15
R99 VPB.t0 VPB.t2 1338.17
R100 VPB.n0 VPB 540.518
R101 VPB.t9 VPB.t5 509.342
R102 VPB.t1 VPB.t8 457.144
R103 VPB.t4 VPB.t3 295.238
R104 VPB VPB.t7 292.858
R105 VPB.n0 VPB.t1 247.619
R106 VPB.t6 VPB.t4 242.857
R107 VPB.t3 VPB.t9 240.476
R108 VPB.t5 VPB.t0 214.517
R109 VPB.t8 VPB.t6 214.286
R110 VPB.t7 VPB.n0 27.8008
R111 a_1396_99.t0 a_1396_99.n1 680.312
R112 a_1396_99.n1 a_1396_99.n0 263.762
R113 a_1396_99.n1 a_1396_99.t1 199.227
R114 VPWR.n7 VPWR.t0 833.578
R115 VPWR.n17 VPWR.n4 695.713
R116 VPWR.n8 VPWR.t2 418.995
R117 VPWR.n25 VPWR.n1 225.18
R118 VPWR.n1 VPWR.t1 52.7206
R119 VPWR.n4 VPWR.t3 46.2955
R120 VPWR.n4 VPWR.t4 46.2955
R121 VPWR.n1 VPWR.t5 37.1046
R122 VPWR.n19 VPWR.n18 36.1417
R123 VPWR.n19 VPWR.n2 36.1417
R124 VPWR.n23 VPWR.n2 36.1417
R125 VPWR.n24 VPWR.n23 36.1417
R126 VPWR.n11 VPWR.n10 36.1417
R127 VPWR.n12 VPWR.n11 36.1417
R128 VPWR.n12 VPWR.n5 36.1417
R129 VPWR.n16 VPWR.n5 36.1417
R130 VPWR.n10 VPWR.n7 15.8123
R131 VPWR.n18 VPWR.n17 10.9181
R132 VPWR.n25 VPWR.n24 10.9181
R133 VPWR.n10 VPWR.n9 9.3005
R134 VPWR.n11 VPWR.n6 9.3005
R135 VPWR.n13 VPWR.n12 9.3005
R136 VPWR.n14 VPWR.n5 9.3005
R137 VPWR.n16 VPWR.n15 9.3005
R138 VPWR.n18 VPWR.n3 9.3005
R139 VPWR.n20 VPWR.n19 9.3005
R140 VPWR.n21 VPWR.n2 9.3005
R141 VPWR.n23 VPWR.n22 9.3005
R142 VPWR.n24 VPWR.n0 9.3005
R143 VPWR.n26 VPWR.n25 8.08026
R144 VPWR.n8 VPWR.n7 7.49709
R145 VPWR.n17 VPWR.n16 0.376971
R146 VPWR VPWR.n26 0.163644
R147 VPWR.n9 VPWR.n8 0.152204
R148 VPWR.n26 VPWR.n0 0.144205
R149 VPWR.n9 VPWR.n6 0.122949
R150 VPWR.n13 VPWR.n6 0.122949
R151 VPWR.n14 VPWR.n13 0.122949
R152 VPWR.n15 VPWR.n14 0.122949
R153 VPWR.n15 VPWR.n3 0.122949
R154 VPWR.n20 VPWR.n3 0.122949
R155 VPWR.n21 VPWR.n20 0.122949
R156 VPWR.n22 VPWR.n21 0.122949
R157 VPWR.n22 VPWR.n0 0.122949
R158 X.n1 X.t0 279.738
R159 X.t0 X.n0 279.738
R160 X.n0 X 8.69186
R161 X X.n1 6.81532
R162 X.n1 X 5.53136
R163 X.n0 X 3.00297
R164 A0.n0 A0.t1 231.629
R165 A0.n0 A0.t0 192.8
R166 A0 A0.n0 159.758
R167 a_537_341.t0 a_537_341.t1 70.9205
R168 a_255_341.t0 a_255_341.t1 159.571
R169 a_1065_387.t0 a_1065_387.t1 53.1905
C0 A0 VPB 0.042012f
C1 S1 A1 5.8e-21
C2 A0 S0 0.106956f
C3 A3 VPB 0.06557f
C4 A0 VGND 0.013266f
C5 A3 X 4.21e-20
C6 S1 A2 8.96e-21
C7 A0 VPWR 0.026538f
C8 S1 VPB 0.091749f
C9 A3 S0 0.027815f
C10 A1 A2 0.123305f
C11 A3 VGND 0.025487f
C12 S1 X 0.001073f
C13 A3 a_846_74# 0.118929f
C14 A3 VPWR 0.017754f
C15 S1 S0 1.76e-19
C16 A1 VPB 0.03455f
C17 S1 VGND 0.07302f
C18 S1 a_846_74# 0.033075f
C19 A2 VPB 0.041275f
C20 S1 VPWR 0.018852f
C21 A1 S0 0.018342f
C22 A1 VGND 0.014902f
C23 A2 X 9.47e-21
C24 A3 a_1338_125# 7.88e-19
C25 A1 a_846_74# 4.53e-19
C26 X VPB 0.011892f
C27 A1 VPWR 0.013811f
C28 A2 S0 0.019282f
C29 A2 VGND 0.017187f
C30 S1 a_1338_125# 0.143989f
C31 A2 a_846_74# 0.013752f
C32 VPB S0 0.467071f
C33 VGND VPB 0.019906f
C34 X S0 2.44e-21
C35 A2 VPWR 0.015778f
C36 VPB a_846_74# 0.02072f
C37 X VGND 0.105718f
C38 VPB VPWR 0.244203f
C39 VGND S0 0.026515f
C40 X VPWR 0.078067f
C41 S0 a_846_74# 0.033896f
C42 VGND a_846_74# 0.417576f
C43 A2 a_1338_125# 4.47e-20
C44 S0 VPWR 0.14758f
C45 VGND VPWR 0.150907f
C46 VPB a_1338_125# 0.072686f
C47 VPWR a_846_74# 0.041141f
C48 X a_1338_125# 0.086414f
C49 A3 S1 0.028626f
C50 S0 a_1338_125# 2.67e-20
C51 VGND a_1338_125# 0.051206f
C52 a_846_74# a_1338_125# 0.173355f
C53 VPWR a_1338_125# 0.342765f
C54 VGND VNB 1.10767f
C55 X VNB 0.107907f
C56 A2 VNB 0.100559f
C57 A1 VNB 0.10039f
C58 S1 VNB 0.450779f
C59 A3 VNB 0.203717f
C60 A0 VNB 0.097384f
C61 VPWR VNB 0.882466f
C62 S0 VNB 0.500914f
C63 VPB VNB 2.28553f
C64 a_1338_125# VNB 0.146565f
C65 a_846_74# VNB 0.075485f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux2i_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2i_4 VNB VPB VPWR VGND S A0 A1 Y
X0 Y.t5 A0.t0 a_475_85.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 a_116_368.t3 A1.t0 Y.t14 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t2 S.t0 a_1030_268.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X3 a_1030_268.t0 S.t1 VPWR.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1862 ps=1.475 w=0.84 l=0.15
X4 a_1030_268.t2 S.t2 VGND.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 Y.t4 A0.t1 a_475_85.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 Y.t1 A0.t2 a_478_368.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1904 ps=1.46 w=1.12 l=0.15
X7 VPWR.t6 a_1030_268.t3 a_116_368.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2128 ps=1.5 w=1.12 l=0.15
X8 a_475_85.t7 a_1030_268.t4 VGND.t8 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.36 ps=2.83 w=0.74 l=0.15
X9 a_478_368.t5 S.t3 VPWR.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X10 a_475_85.t1 A0.t3 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_114_85.t3 A1.t1 Y.t15 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 VGND.t3 S.t4 a_114_85.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_475_85.t6 a_1030_268.t5 VGND.t7 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.20315 ps=1.49 w=0.74 l=0.15
X14 VGND.t4 S.t5 a_114_85.t6 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1887 pd=1.25 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VPWR.t5 a_1030_268.t6 a_116_368.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_116_368.t4 a_1030_268.t7 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.7504 ps=3.58 w=1.12 l=0.15
X17 Y.t8 A1.t2 a_116_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X18 Y.t9 A1.t3 a_114_85.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.13505 ps=1.105 w=0.74 l=0.15
X19 VGND.t6 a_1030_268.t8 a_475_85.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.19615 pd=1.41 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_116_368.t1 A1.t4 Y.t10 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 Y.t0 A0.t4 a_478_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X22 Y.t11 A1.t5 a_116_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_114_85.t5 S.t6 VGND.t2 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1887 ps=1.25 w=0.74 l=0.15
X24 a_114_85.t4 S.t7 VGND.t0 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19615 ps=1.41 w=0.74 l=0.15
X25 Y.t12 A1.t6 a_114_85.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 a_478_368.t1 A0.t5 Y.t6 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.1736 ps=1.43 w=1.12 l=0.15
X27 a_478_368.t0 A0.t6 Y.t7 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X28 a_478_368.t4 S.t8 VPWR.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X29 a_114_85.t0 A1.t7 Y.t13 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.13505 pd=1.105 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 a_475_85.t0 A0.t7 Y.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X31 VGND.t5 a_1030_268.t9 a_475_85.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.20315 pd=1.49 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A0.n0 A0.t4 307.142
R1 A0.n1 A0.t6 226.809
R2 A0.n4 A0.t2 226.809
R3 A0.n6 A0.t5 226.809
R4 A0.n6 A0.t3 180.531
R5 A0.n0 A0.t1 178.34
R6 A0.n5 A0.t0 178.34
R7 A0.n2 A0.t7 178.34
R8 A0.n7 A0 158.13
R9 A0 A0.n3 153.042
R10 A0.n9 A0.n8 152
R11 A0.n1 A0.n0 112.76
R12 A0.n8 A0.n7 49.6611
R13 A0.n4 A0.n3 38.7066
R14 A0.n3 A0.n2 29.9429
R15 A0.n7 A0.n6 10.955
R16 A0.n8 A0.n5 10.2247
R17 A0 A0.n9 9.07957
R18 A0.n9 A0 5.2098
R19 A0.n2 A0.n1 4.38232
R20 A0.n5 A0.n4 0.730803
R21 a_475_85.n2 a_475_85.n0 257.825
R22 a_475_85.n4 a_475_85.n3 253.142
R23 a_475_85.n2 a_475_85.n1 185
R24 a_475_85.n5 a_475_85.n4 185
R25 a_475_85.n4 a_475_85.n2 171.294
R26 a_475_85.n3 a_475_85.t1 34.0546
R27 a_475_85.n3 a_475_85.t3 22.7032
R28 a_475_85.n1 a_475_85.t5 22.7032
R29 a_475_85.n1 a_475_85.t7 22.7032
R30 a_475_85.n0 a_475_85.t4 22.7032
R31 a_475_85.n0 a_475_85.t6 22.7032
R32 a_475_85.n5 a_475_85.t2 22.7032
R33 a_475_85.t0 a_475_85.n5 22.7032
R34 Y.n13 Y.n12 585
R35 Y.n7 Y.t0 331.259
R36 Y.n9 Y.n8 300.733
R37 Y.n11 Y.n10 297.598
R38 Y.n9 Y.t14 293.408
R39 Y.n6 Y.t4 279.738
R40 Y.n1 Y.t15 207.595
R41 Y.n1 Y.n0 199.306
R42 Y.n5 Y.n4 185
R43 Y.n3 Y.n2 96.4473
R44 Y.n3 Y.n1 60.2814
R45 Y.n11 Y.n9 55.3417
R46 Y.n13 Y.n11 55.1936
R47 Y.n6 Y.n5 46.2372
R48 Y.n5 Y.n3 41.0127
R49 Y.n12 Y.t1 35.1791
R50 Y.n7 Y.n6 32.0389
R51 Y.n10 Y.t6 28.1434
R52 Y.n4 Y.t2 26.7573
R53 Y.n12 Y.t7 26.3844
R54 Y.n8 Y.t10 26.3844
R55 Y.n8 Y.t11 26.3844
R56 Y.n10 Y.t8 26.3844
R57 Y.n4 Y.t5 25.9464
R58 Y Y.n13 23.4908
R59 Y.n2 Y.t3 22.7032
R60 Y.n2 Y.t9 22.7032
R61 Y.n0 Y.t13 22.7032
R62 Y.n0 Y.t12 22.7032
R63 Y Y.n7 10.8917
R64 VNB.t2 VNB.t7 3718.64
R65 VNB.t13 VNB.t14 1524.41
R66 VNB.t4 VNB.t15 1362.73
R67 VNB.t5 VNB.t6 1362.73
R68 VNB.t10 VNB.t8 1189.5
R69 VNB.t12 VNB.t11 1154.86
R70 VNB.t1 VNB.t3 1154.86
R71 VNB VNB.t16 1143.31
R72 VNB.t3 VNB.t0 1097.11
R73 VNB.t14 VNB.t12 993.177
R74 VNB.t15 VNB.t13 993.177
R75 VNB.t6 VNB.t4 993.177
R76 VNB.t7 VNB.t5 993.177
R77 VNB.t0 VNB.t2 993.177
R78 VNB.t8 VNB.t1 993.177
R79 VNB.t9 VNB.t10 993.177
R80 VNB.t16 VNB.t9 993.177
R81 A1.n0 A1.t2 226.809
R82 A1.n2 A1.t4 226.809
R83 A1.n3 A1.t5 226.809
R84 A1.n5 A1.t0 226.809
R85 A1.n0 A1.t3 180.531
R86 A1.n5 A1.t1 179.802
R87 A1.n4 A1.t6 178.34
R88 A1.n10 A1.t7 178.34
R89 A1 A1.n1 155.721
R90 A1.n12 A1.n11 152
R91 A1.n9 A1.n8 152
R92 A1.n7 A1.n6 152
R93 A1.n2 A1.n1 46.0096
R94 A1.n10 A1.n9 46.0096
R95 A1.n6 A1.n4 32.8641
R96 A1.n6 A1.n5 28.4823
R97 A1.n1 A1.n0 19.7187
R98 A1.n9 A1.n3 12.4157
R99 A1.n8 A1.n7 10.1214
R100 A1.n12 A1 7.88887
R101 A1 A1.n12 6.4005
R102 A1.n4 A1.n3 4.38232
R103 A1.n11 A1.n2 3.65202
R104 A1.n11 A1.n10 3.65202
R105 A1.n8 A1 2.23306
R106 A1.n7 A1 1.93538
R107 a_116_368.n1 a_116_368.t6 834.093
R108 a_116_368.n1 a_116_368.n0 585
R109 a_116_368.n4 a_116_368.n3 346.034
R110 a_116_368.n3 a_116_368.n2 305.998
R111 a_116_368.n3 a_116_368.n1 276.051
R112 a_116_368.n0 a_116_368.t5 26.3844
R113 a_116_368.n0 a_116_368.t4 26.3844
R114 a_116_368.n2 a_116_368.t2 26.3844
R115 a_116_368.n2 a_116_368.t1 26.3844
R116 a_116_368.n4 a_116_368.t0 26.3844
R117 a_116_368.t3 a_116_368.n4 26.3844
R118 VPB.t6 VPB.t8 732.931
R119 VPB.t13 VPB.t12 510.753
R120 VPB.t9 VPB.t10 500.538
R121 VPB.t12 VPB.t11 487.769
R122 VPB VPB.t3 257.93
R123 VPB.t10 VPB.t13 255.376
R124 VPB.t4 VPB.t6 255.376
R125 VPB.t7 VPB.t4 255.376
R126 VPB.t5 VPB.t7 250.269
R127 VPB.t2 VPB.t5 234.946
R128 VPB.t11 VPB.t14 229.839
R129 VPB.t8 VPB.t9 229.839
R130 VPB.t1 VPB.t2 229.839
R131 VPB.t0 VPB.t1 229.839
R132 VPB.t3 VPB.t0 229.839
R133 S.n22 S.t8 261.863
R134 S.n4 S.n3 250.909
R135 S.n2 S.t3 250.909
R136 S.n19 S.n1 250.909
R137 S.n5 S.t0 248.207
R138 S.n7 S.t1 205.922
R139 S S.n22 155.911
R140 S.n21 S.t7 154.24
R141 S.n18 S.t5 154.24
R142 S.n13 S.t6 154.24
R143 S.n8 S.t4 154.24
R144 S.n5 S.t2 154.24
R145 S.n6 S 152.357
R146 S.n10 S.n9 152
R147 S.n12 S.n11 152
R148 S.n15 S.n14 152
R149 S.n17 S.n16 152
R150 S.n20 S.n0 152
R151 S.n8 S.n4 37.246
R152 S.n17 S.n2 35.7853
R153 S.n21 S.n20 33.5944
R154 S.n9 S.n7 26.2914
R155 S.n14 S.n13 26.2914
R156 S.n19 S.n18 24.1005
R157 S.n7 S.n6 23.3702
R158 S.n13 S.n12 23.3702
R159 S.n18 S.n17 20.449
R160 S.n22 S.n21 16.0672
R161 S.n14 S.n2 13.8763
R162 S.n6 S.n5 13.146
R163 S.n16 S.n15 12.0894
R164 S.n10 S 11.7338
R165 S.n11 S 10.3116
R166 S.n9 S.n8 10.2247
R167 S S.n0 8.88939
R168 S S.n0 8.17828
R169 S.n11 S 6.75606
R170 S S.n10 5.33383
R171 S.n20 S.n19 5.11262
R172 S.n16 S 3.2005
R173 S.n12 S.n4 2.19141
R174 S.n15 S 1.77828
R175 a_1030_268.n13 a_1030_268.n12 307.885
R176 a_1030_268.n5 a_1030_268.t7 240.44
R177 a_1030_268.n0 a_1030_268.t3 229.487
R178 a_1030_268.n9 a_1030_268.n2 229.487
R179 a_1030_268.n4 a_1030_268.t6 229.487
R180 a_1030_268.n12 a_1030_268.t2 207.471
R181 a_1030_268.n0 a_1030_268.t8 193.093
R182 a_1030_268.n12 a_1030_268.n11 189.079
R183 a_1030_268.n10 a_1030_268.t5 179.947
R184 a_1030_268.n5 a_1030_268.t4 154.24
R185 a_1030_268.n3 a_1030_268.t9 154.24
R186 a_1030_268.n8 a_1030_268.n7 152
R187 a_1030_268.n10 a_1030_268.n1 152
R188 a_1030_268.n11 a_1030_268.n0 152
R189 a_1030_268.n7 a_1030_268.n6 81.6328
R190 a_1030_268.n0 a_1030_268.n10 49.6611
R191 a_1030_268.n8 a_1030_268.n3 36.5157
R192 a_1030_268.n13 a_1030_268.t1 35.1791
R193 a_1030_268.t0 a_1030_268.n13 35.1791
R194 a_1030_268.n10 a_1030_268.n9 28.4823
R195 a_1030_268.n6 a_1030_268.n4 25.6895
R196 a_1030_268.n6 a_1030_268.n5 22.3626
R197 a_1030_268.n9 a_1030_268.n8 21.1793
R198 a_1030_268.n11 a_1030_268.n1 13.1884
R199 a_1030_268.n7 a_1030_268.n1 13.1884
R200 a_1030_268.n4 a_1030_268.n3 8.03383
R201 VPWR.n3 VPWR.t5 827.967
R202 VPWR.n9 VPWR.t3 809.364
R203 VPWR.n1 VPWR.n0 604.976
R204 VPWR.n3 VPWR.t4 442.084
R205 VPWR.n6 VPWR.t2 368.435
R206 VPWR.n4 VPWR.t1 335.3
R207 VPWR.n4 VPWR.n3 217.905
R208 VPWR.n5 VPWR.n4 50.2389
R209 VPWR.n0 VPWR.t0 35.1791
R210 VPWR.n10 VPWR.n1 28.6123
R211 VPWR.n8 VPWR.n5 27.1064
R212 VPWR.n0 VPWR.t6 26.3844
R213 VPWR.n9 VPWR.n8 25.6005
R214 VPWR.n10 VPWR.n9 21.8358
R215 VPWR.n8 VPWR.n7 9.3005
R216 VPWR.n9 VPWR.n2 9.3005
R217 VPWR.n11 VPWR.n10 9.3005
R218 VPWR.n12 VPWR.n1 6.85475
R219 VPWR.n6 VPWR.n5 6.77545
R220 VPWR VPWR.n12 1.74509
R221 VPWR.n7 VPWR.n6 0.632103
R222 VPWR.n12 VPWR.n11 0.162016
R223 VPWR.n7 VPWR.n2 0.122949
R224 VPWR.n11 VPWR.n2 0.122949
R225 VGND.n18 VGND.t8 391.56
R226 VGND.n2 VGND.n1 246.475
R227 VGND.n11 VGND.n10 220.173
R228 VGND.n5 VGND.n4 201.915
R229 VGND.n7 VGND.n6 123.767
R230 VGND.n1 VGND.t5 43.1743
R231 VGND.n4 VGND.t2 41.3519
R232 VGND.n4 VGND.t4 41.3519
R233 VGND.n10 VGND.t0 35.6762
R234 VGND.n10 VGND.t6 35.6762
R235 VGND.n9 VGND.n5 35.0123
R236 VGND.n6 VGND.t3 34.0546
R237 VGND.n13 VGND.n12 32.9284
R238 VGND.n17 VGND.n16 29.9622
R239 VGND.n18 VGND.n17 25.224
R240 VGND.n13 VGND.n2 24.973
R241 VGND.n1 VGND.t7 24.8648
R242 VGND.n6 VGND.t1 22.7032
R243 VGND.n11 VGND.n9 20.4554
R244 VGND.n17 VGND.n0 9.3005
R245 VGND.n16 VGND.n15 9.3005
R246 VGND.n14 VGND.n13 9.3005
R247 VGND.n12 VGND.n3 9.3005
R248 VGND.n9 VGND.n8 9.3005
R249 VGND.n19 VGND.n18 7.36261
R250 VGND.n7 VGND.n5 5.17976
R251 VGND.n12 VGND.n11 2.58636
R252 VGND VGND.n19 1.26109
R253 VGND.n16 VGND.n2 1.03484
R254 VGND.n8 VGND.n7 0.434826
R255 VGND.n19 VGND.n0 0.154009
R256 VGND.n8 VGND.n3 0.122949
R257 VGND.n14 VGND.n3 0.122949
R258 VGND.n15 VGND.n14 0.122949
R259 VGND.n15 VGND.n0 0.122949
R260 a_478_368.n3 a_478_368.n2 647.758
R261 a_478_368.n2 a_478_368.n1 585
R262 a_478_368.n0 a_478_368.t5 372.591
R263 a_478_368.n0 a_478_368.t4 322.144
R264 a_478_368.n2 a_478_368.n0 267.524
R265 a_478_368.n1 a_478_368.t0 35.1791
R266 a_478_368.n3 a_478_368.t1 33.4201
R267 a_478_368.n1 a_478_368.t2 26.3844
R268 a_478_368.t3 a_478_368.n3 26.3844
R269 a_114_85.n4 a_114_85.n2 445.483
R270 a_114_85.n5 a_114_85.n4 237.9
R271 a_114_85.n4 a_114_85.n3 197.994
R272 a_114_85.n2 a_114_85.n0 158.034
R273 a_114_85.n2 a_114_85.n1 91.1008
R274 a_114_85.n3 a_114_85.t2 36.487
R275 a_114_85.n1 a_114_85.t6 22.7032
R276 a_114_85.n1 a_114_85.t4 22.7032
R277 a_114_85.n0 a_114_85.t7 22.7032
R278 a_114_85.n0 a_114_85.t5 22.7032
R279 a_114_85.n3 a_114_85.t0 22.7032
R280 a_114_85.n5 a_114_85.t1 22.7032
R281 a_114_85.t3 a_114_85.n5 22.7032
C0 S VPWR 0.121198f
C1 A0 VGND 0.021141f
C2 VPWR VPB 0.247884f
C3 Y VPWR 0.102164f
C4 S VGND 0.115654f
C5 VGND VPB 0.012554f
C6 Y VGND 0.069242f
C7 VPWR VGND 0.167521f
C8 A1 A0 0.074829f
C9 A1 VPB 0.137796f
C10 A1 Y 0.341891f
C11 A0 VPB 0.146598f
C12 A1 VPWR 0.028059f
C13 A0 Y 0.318274f
C14 S VPB 0.218585f
C15 S Y 0.001454f
C16 A1 VGND 0.026668f
C17 A0 VPWR 0.02145f
C18 Y VPB 0.027863f
C19 VGND VNB 1.14104f
C20 VPWR VNB 0.935171f
C21 Y VNB 0.129862f
C22 S VNB 0.612437f
C23 A0 VNB 0.415032f
C24 A1 VNB 0.425136f
C25 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux2i_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2i_2 VNB VPB VPWR VGND A0 Y S A1
X0 a_922_72.t0 S.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2382 ps=1.555 w=1 l=0.15
X1 a_115_74.t1 A0.t0 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1369 pd=1.11 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 a_340_368.t3 a_922_72.t2 VPWR.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3021 ps=1.805 w=1.12 l=0.15
X3 a_118_368.t1 A0.t1 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.3416 ps=2.85 w=1.12 l=0.15
X4 Y.t4 A0.t2 a_118_368.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2632 pd=1.59 as=0.1904 ps=1.46 w=1.12 l=0.15
X5 VPWR.t1 a_922_72.t3 a_340_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t1 S.t1 a_337_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.215625 pd=1.505 as=0.1221 ps=1.07 w=0.74 l=0.15
X7 a_115_74.t2 a_922_72.t4 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.215625 ps=1.505 w=0.74 l=0.15
X8 a_340_368.t0 A1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.2632 ps=1.59 w=1.12 l=0.15
X9 a_337_74.t1 S.t2 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.36 ps=2.83 w=0.74 l=0.15
X10 Y.t1 A0.t3 a_115_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.188175 pd=1.355 as=0.1369 ps=1.11 w=0.74 l=0.15
X11 Y.t7 A1.t1 a_337_74.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.270675 ps=1.505 w=0.74 l=0.15
X12 a_922_72.t1 S.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X13 VPWR.t4 S.t4 a_118_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3021 pd=1.805 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y.t5 A1.t2 a_340_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3808 ps=1.8 w=1.12 l=0.15
X15 a_337_74.t0 A1.t3 Y.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.270675 pd=1.505 as=0.188175 ps=1.355 w=0.74 l=0.15
X16 VGND.t3 a_922_72.t5 a_115_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1221 ps=1.07 w=0.74 l=0.15
X17 a_118_368.t2 S.t5 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.581825 ps=3.6 w=1.12 l=0.15
R0 S S.n0 242.031
R1 S.n0 S.t0 230.581
R2 S.n2 S.t4 226.809
R3 S.n4 S.t5 226.809
R4 S.n0 S.t3 164.44
R5 S.n4 S.t2 159.644
R6 S.n2 S.t1 159.644
R7 S.n3 S.n1 152
R8 S.n6 S.n5 152
R9 S.n5 S.n3 49.6611
R10 S.n1 S 13.8932
R11 S.n5 S.n4 10.955
R12 S S.n6 9.52245
R13 S.n6 S 5.46391
R14 S.n3 S.n2 5.11262
R15 S S.n1 1.09318
R16 VPWR.n0 VPWR.t3 882.855
R17 VPWR.n5 VPWR.n4 607.607
R18 VPWR.n3 VPWR.n2 323.262
R19 VPWR.n2 VPWR.t2 46.2955
R20 VPWR.n4 VPWR.t0 43.0943
R21 VPWR.n4 VPWR.t4 42.2148
R22 VPWR.n7 VPWR.n6 36.1417
R23 VPWR.n2 VPWR.t1 35.4615
R24 VPWR.n7 VPWR.n0 15.4776
R25 VPWR.n6 VPWR.n5 13.6401
R26 VPWR.n9 VPWR.n0 11.8491
R27 VPWR.n5 VPWR.n3 11.5874
R28 VPWR.n6 VPWR.n1 9.3005
R29 VPWR.n8 VPWR.n7 9.3005
R30 VPWR VPWR.n9 0.772485
R31 VPWR.n3 VPWR.n1 0.523977
R32 VPWR.n9 VPWR.n8 0.150543
R33 VPWR.n8 VPWR.n1 0.122949
R34 a_922_72.t0 a_922_72.n3 407.3
R35 a_922_72.n0 a_922_72.t3 229.487
R36 a_922_72.n1 a_922_72.t2 229.487
R37 a_922_72.n3 a_922_72.n2 209.691
R38 a_922_72.n1 a_922_72.t4 156.431
R39 a_922_72.n0 a_922_72.t5 156.431
R40 a_922_72.n3 a_922_72.t1 131.947
R41 a_922_72.n2 a_922_72.n1 54.7732
R42 a_922_72.n2 a_922_72.n0 10.955
R43 VPB.t1 VPB.t2 592.473
R44 VPB.t0 VPB.t1 423.925
R45 VPB.t3 VPB.t6 324.329
R46 VPB.t8 VPB.t0 316.668
R47 VPB.t5 VPB.t4 298.791
R48 VPB VPB.t7 263.038
R49 VPB.t7 VPB.t8 250.269
R50 VPB.t6 VPB.t5 229.839
R51 VPB.t2 VPB.t3 229.839
R52 A0.n1 A0.t2 261.62
R53 A0.n3 A0.t1 261.62
R54 A0.n3 A0.t0 156.431
R55 A0.n1 A0.t3 156.431
R56 A0 A0.n4 153.558
R57 A0.n2 A0.n0 152
R58 A0.n4 A0.n2 49.6611
R59 A0.n2 A0.n1 10.955
R60 A0.n4 A0.n3 10.955
R61 A0 A0.n0 10.2059
R62 A0.n0 A0 6.4005
R63 Y.n2 Y.t5 934.861
R64 Y.n6 Y 589.444
R65 Y.n2 Y.n1 585
R66 Y.n6 Y.n0 585
R67 Y.n7 Y.n6 585
R68 Y.n4 Y.t7 371.964
R69 Y.n4 Y.n3 197.415
R70 Y.n5 Y.t2 132.03
R71 Y.n5 Y.n4 78.4882
R72 Y Y.n5 75.3784
R73 Y.n8 Y.n2 65.5064
R74 Y.n1 Y.t0 41.3353
R75 Y.n1 Y.t4 41.3353
R76 Y.n3 Y.t6 35.6762
R77 Y.n3 Y.t1 35.6762
R78 Y.n6 Y.t3 28.1434
R79 Y Y.n0 10.3116
R80 Y Y.n8 10.3116
R81 Y Y.n0 2.84494
R82 Y.n8 Y.n7 1.6005
R83 Y.n7 Y 1.24494
R84 a_115_74.n1 a_115_74.n0 655.407
R85 a_115_74.t1 a_115_74.n1 37.2978
R86 a_115_74.n0 a_115_74.t3 26.7573
R87 a_115_74.n0 a_115_74.t2 26.7573
R88 a_115_74.n1 a_115_74.t0 22.7032
R89 VNB.t8 VNB.t4 2609.97
R90 VNB.t2 VNB.t8 1986.35
R91 VNB.t5 VNB.t7 1397.38
R92 VNB.t0 VNB.t2 1362.73
R93 VNB.t6 VNB.t3 1339.63
R94 VNB.t1 VNB.t0 1201.05
R95 VNB VNB.t1 1154.86
R96 VNB.t7 VNB.t6 1108.66
R97 VNB.t4 VNB.t5 1108.66
R98 a_340_368.n1 a_340_368.n0 757.462
R99 a_340_368.n0 a_340_368.t0 58.4134
R100 a_340_368.n0 a_340_368.t1 57.6263
R101 a_340_368.t2 a_340_368.n1 26.3844
R102 a_340_368.n1 a_340_368.t3 26.3844
R103 a_118_368.n1 a_118_368.n0 1077.7
R104 a_118_368.t1 a_118_368.n1 33.4201
R105 a_118_368.n0 a_118_368.t3 26.3844
R106 a_118_368.n0 a_118_368.t2 26.3844
R107 a_118_368.n1 a_118_368.t0 26.3844
R108 a_337_74.n1 a_337_74.n0 504.817
R109 a_337_74.n1 a_337_74.t3 79.46
R110 a_337_74.t0 a_337_74.n1 35.6762
R111 a_337_74.n0 a_337_74.t2 26.7573
R112 a_337_74.n0 a_337_74.t1 26.7573
R113 VGND.n0 VGND.t0 374.921
R114 VGND.n5 VGND.n4 249.918
R115 VGND.n3 VGND.n2 216.04
R116 VGND.n2 VGND.t2 41.2505
R117 VGND.n4 VGND.t4 37.2978
R118 VGND.n4 VGND.t1 36.487
R119 VGND.n7 VGND.n6 36.1417
R120 VGND.n2 VGND.t3 30.6984
R121 VGND.n6 VGND.n5 13.5731
R122 VGND.n7 VGND.n0 13.4618
R123 VGND.n9 VGND.n0 12.8294
R124 VGND.n5 VGND.n3 11.5462
R125 VGND.n8 VGND.n7 9.3005
R126 VGND.n6 VGND.n1 9.3005
R127 VGND VGND.n9 0.773575
R128 VGND.n3 VGND.n1 0.500418
R129 VGND.n9 VGND.n8 0.14947
R130 VGND.n8 VGND.n1 0.122949
R131 A1.n0 A1.t2 226.809
R132 A1.n1 A1.t0 226.809
R133 A1.n1 A1.t3 198.204
R134 A1.n0 A1.t1 198.204
R135 A1.n7 A1.n6 152
R136 A1.n5 A1.n4 152
R137 A1.n3 A1.n2 152
R138 A1.n6 A1.n5 49.6611
R139 A1.n5 A1.n2 49.6611
R140 A1.n4 A1.n3 12.615
R141 A1.n7 A1 11.3164
R142 A1.n6 A1.n0 10.955
R143 A1.n2 A1.n1 10.955
R144 A1 A1.n7 6.49325
R145 A1.n3 A1 3.89615
R146 A1.n4 A1 1.29905
C0 S VGND 0.03731f
C1 Y VGND 0.337142f
C2 VPB VPWR 0.155214f
C3 VPB A0 0.066883f
C4 VPB A1 0.103882f
C5 VPWR A0 0.019908f
C6 VPWR A1 0.019427f
C7 VPB S 0.123919f
C8 A0 A1 0.050983f
C9 VPB Y 0.020567f
C10 VPWR S 0.095658f
C11 A0 S 3.01e-19
C12 VPWR Y 0.066025f
C13 VPB VGND 0.009744f
C14 A0 Y 0.144902f
C15 A1 S 0.038276f
C16 VPWR VGND 0.100142f
C17 A0 VGND 0.013548f
C18 A1 Y 0.145136f
C19 S Y 0.004125f
C20 A1 VGND 0.015901f
C21 VGND VNB 0.742867f
C22 Y VNB 0.142416f
C23 S VNB 0.334482f
C24 A1 VNB 0.271079f
C25 A0 VNB 0.24228f
C26 VPWR VNB 0.586404f
C27 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux2i_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2i_1 VNB VPB VPWR VGND S A1 A0 Y
X0 a_114_74.t1 S.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.231 pd=2.23 as=0.2394 ps=2.25 w=0.84 l=0.15
X1 a_399_368.t1 A1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_114_74.t0 S.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3 Y.t2 A0.t0 a_223_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4 a_426_74.t0 a_114_74.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 VGND.t1 S.t2 a_225_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_225_74.t1 A1.t1 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.26085 ps=1.445 w=0.74 l=0.15
X7 a_399_368.t0 a_114_74.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Y.t3 A0.t1 a_426_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.26085 pd=1.445 as=0.0888 ps=0.98 w=0.74 l=0.15
X9 VPWR.t1 S.t3 a_223_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
R0 S.n1 S.t3 339.274
R1 S.n2 S.n1 260.281
R2 S.n0 S.t0 232.661
R3 S.n2 S.t1 183.85
R4 S.n1 S.t2 163.077
R5 S S.n0 155.314
R6 S.n4 S.n3 152
R7 S.n3 S.n0 46.8234
R8 S.n3 S.n2 12.3948
R9 S S.n4 6.92756
R10 S.n4 S 4.21697
R11 VPWR.n1 VPWR.t0 428.098
R12 VPWR.n1 VPWR.n0 321.998
R13 VPWR.n0 VPWR.t2 26.3844
R14 VPWR.n0 VPWR.t1 26.3844
R15 VPWR VPWR.n1 0.152248
R16 a_114_74.t1 a_114_74.n1 446.161
R17 a_114_74.n1 a_114_74.t0 258.699
R18 a_114_74.n0 a_114_74.t3 250.909
R19 a_114_74.n1 a_114_74.n0 233.319
R20 a_114_74.n0 a_114_74.t2 220.113
R21 VPB.t3 VPB.t4 497.985
R22 VPB.t2 VPB.t1 497.985
R23 VPB VPB.t2 252.823
R24 VPB.t4 VPB.t0 229.839
R25 VPB.t1 VPB.t3 229.839
R26 A1.n0 A1.t0 277.526
R27 A1.n0 A1.t1 170.147
R28 A1 A1.n0 158.788
R29 Y.n1 Y.n0 367.779
R30 Y.n4 Y.n3 185
R31 Y.n2 Y.n1 185
R32 Y.n3 Y.n2 68.9194
R33 Y.n0 Y.t0 26.3844
R34 Y.n0 Y.t2 26.3844
R35 Y.n2 Y.t1 22.7032
R36 Y.n3 Y.t3 22.7032
R37 Y.n4 Y.n1 16.4853
R38 Y Y.n4 4.07323
R39 a_399_368.t0 a_399_368.t1 651.721
R40 VGND.n1 VGND.t0 255.815
R41 VGND.n1 VGND.n0 217.169
R42 VGND.n0 VGND.t2 34.0546
R43 VGND.n0 VGND.t1 34.0546
R44 VGND VGND.n1 0.143944
R45 VNB.t1 VNB.t0 2286.61
R46 VNB.t4 VNB.t3 1974.8
R47 VNB.t0 VNB.t2 1316.54
R48 VNB VNB.t1 1143.31
R49 VNB.t2 VNB.t4 900.788
R50 A0.n0 A0.t0 255.168
R51 A0.n0 A0.t1 249.034
R52 A0 A0.n0 156.316
R53 a_223_368.t0 a_223_368.t1 699.898
R54 a_426_74.t0 a_426_74.t1 38.9194
R55 a_225_74.t0 a_225_74.t1 455.281
C0 VPWR VGND 0.060801f
C1 A1 VPB 0.039933f
C2 A0 S 2.21e-19
C3 Y VGND 0.013114f
C4 VPWR VPB 0.114202f
C5 VPWR S 0.059726f
C6 Y VPB 0.004874f
C7 VGND VPB 0.010263f
C8 Y S 8.64e-19
C9 VGND S 0.055946f
C10 VPB S 0.124452f
C11 A0 A1 0.042888f
C12 A0 VPWR 0.007166f
C13 A0 Y 0.076012f
C14 A1 VPWR 0.006751f
C15 A1 Y 0.052541f
C16 A0 VGND 0.009062f
C17 VPWR Y 0.009109f
C18 A1 VGND 0.009993f
C19 A0 VPB 0.049505f
C20 VGND VNB 0.514799f
C21 Y VNB 0.027487f
C22 VPWR VNB 0.415927f
C23 A1 VNB 0.174945f
C24 A0 VNB 0.133946f
C25 S VNB 0.383772f
C26 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2_4 VNB VPB VPWR VGND A0 A1 X S
X0 VPWR.t8 S.t0 a_27_368.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2186 pd=1.52 as=0.295 ps=2.59 w=1 l=0.15
X1 VPWR.t3 a_193_241# X.t7 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.278 pd=1.775 as=0.275525 ps=1.675 w=1.12 l=0.15
X2 a_193_241# A0.t0 a_722_391.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.31 as=0.15 ps=1.3 w=1 l=0.15
X3 X.t6 a_193_241# VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.29075 pd=1.78 as=0.2186 ps=1.52 w=1.12 l=0.15
X4 X.t5 a_193_241# VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.275525 pd=1.675 as=0.290025 ps=1.775 w=1.12 l=0.15
X5 a_722_391.t2 A0.t1 a_193_241# VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.33 ps=2.66 w=1 l=0.15
X6 VGND.t6 S.t1 a_27_368.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1469 pd=1.16 as=0.1824 ps=1.85 w=0.64 l=0.15
X7 VPWR.t0 a_193_241# X.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.290025 pd=1.775 as=0.29075 ps=1.78 w=1.12 l=0.15
X8 a_709_119# S.t2 VGND.t8 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.232925 ps=1.455 w=0.64 l=0.15
X9 a_193_241# A1.t0 a_936_391.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.15 ps=1.3 w=1 l=0.15
X10 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2112 pd=1.94 as=0.0992 ps=0.95 w=0.64 l=0.15
X11 a_936_391.t0 A1.t1 a_193_241# VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.155 ps=1.31 w=1 l=0.15
X12 a_937_119.t2 A0.t2 a_193_241# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.096 pd=0.94 as=0.4992 ps=2.84 w=0.64 l=0.15
X13 VPWR.t4 a_27_368.t2 a_936_391.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4177 pd=3.02 as=0.15 ps=1.3 w=1 l=0.15
X14 VPWR.t7 S.t3 a_722_391.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.25385 pd=1.6 as=0.15 ps=1.3 w=1 l=0.15
X15 VGND.t3 a_193_241# X.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.1184 ps=1.06 w=0.74 l=0.15
X16 a_722_391.t0 S.t4 VPWR.t6 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.278 ps=1.775 w=1 l=0.15
X17 X.t2 a_193_241# VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1469 ps=1.16 w=0.74 l=0.15
X18 a_936_391.t2 a_27_368.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.25385 ps=1.6 w=1 l=0.15
X19 X.t1 a_193_241# VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1628 ps=1.18 w=0.74 l=0.15
X20 VGND.t5 a_27_368.t4 a_937_119.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.3692 pd=2.64 as=0.0896 ps=0.92 w=0.64 l=0.15
X21 a_937_119.t0 a_27_368.t5 VGND.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1568 ps=1.13 w=0.64 l=0.15
X22 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0992 pd=0.95 as=0.1056 ps=0.97 w=0.64 l=0.15
X23 VGND.t0 a_193_241# X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.232925 pd=1.455 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VGND.t7 S.t5 a_709_119# VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1568 pd=1.13 as=0.112 ps=0.99 w=0.64 l=0.15
R0 S S.n2 397.88
R1 S.n3 S.t0 230.919
R2 S.n0 S.t3 217.752
R3 S.n1 S.t4 215.561
R4 S.n3 S.t1 196.911
R5 S.n1 S.t2 176.588
R6 S.n0 S.t5 167.094
R7 S S.n3 154.03
R8 S.n2 S.n0 56.9641
R9 S.n2 S.n1 6.57323
R10 a_27_368.t1 a_27_368.n3 829.89
R11 a_27_368.t1 a_27_368.n4 735.255
R12 a_27_368.n2 a_27_368.t2 217.752
R13 a_27_368.n0 a_27_368.t3 215.561
R14 a_27_368.n4 a_27_368.t0 201.685
R15 a_27_368.n1 a_27_368.n0 14.5754
R16 a_27_368.n0 a_27_368.t5 167.094
R17 a_27_368.n2 a_27_368.t4 167.094
R18 a_27_368.n3 a_27_368.n1 400.233
R19 a_27_368.n1 a_27_368.n2 46.2748
R20 a_27_368.n4 a_27_368.n3 12.8005
R21 VPWR.n9 VPWR.t4 863.729
R22 VPWR.n6 VPWR.n5 614.765
R23 VPWR.n3 VPWR.n2 612.173
R24 VPWR.n22 VPWR.n1 604.107
R25 VPWR.n10 VPWR.n8 600.128
R26 VPWR.n5 VPWR.t6 55.1605
R27 VPWR.n1 VPWR.t8 47.2805
R28 VPWR.n8 VPWR.t5 46.2955
R29 VPWR.n8 VPWR.t7 46.2955
R30 VPWR.n2 VPWR.t1 41.3353
R31 VPWR.n2 VPWR.t0 41.3353
R32 VPWR.n21 VPWR.n20 36.1417
R33 VPWR.n17 VPWR.n16 36.1417
R34 VPWR.n12 VPWR.n11 36.1417
R35 VPWR.n16 VPWR.n15 32.9482
R36 VPWR.n5 VPWR.t3 31.6736
R37 VPWR.n1 VPWR.t2 28.5142
R38 VPWR.n12 VPWR.n6 19.4536
R39 VPWR.n22 VPWR.n21 15.4358
R40 VPWR.n10 VPWR.n9 14.5291
R41 VPWR.n20 VPWR.n3 14.1831
R42 VPWR.n11 VPWR.n7 9.3005
R43 VPWR.n13 VPWR.n12 9.3005
R44 VPWR.n15 VPWR.n14 9.3005
R45 VPWR.n16 VPWR.n4 9.3005
R46 VPWR.n18 VPWR.n17 9.3005
R47 VPWR.n20 VPWR.n19 9.3005
R48 VPWR.n21 VPWR.n0 9.3005
R49 VPWR.n23 VPWR.n22 7.53404
R50 VPWR.n17 VPWR.n3 4.39482
R51 VPWR.n11 VPWR.n10 3.76521
R52 VPWR.n15 VPWR.n6 2.31774
R53 VPWR.n9 VPWR.n7 0.772636
R54 VPWR VPWR.n23 0.161409
R55 VPWR.n23 VPWR.n0 0.146411
R56 VPWR.n13 VPWR.n7 0.122949
R57 VPWR.n14 VPWR.n13 0.122949
R58 VPWR.n14 VPWR.n4 0.122949
R59 VPWR.n18 VPWR.n4 0.122949
R60 VPWR.n19 VPWR.n18 0.122949
R61 VPWR.n19 VPWR.n0 0.122949
R62 VPB VPB.n1 415.168
R63 VPB.t1 VPB.t3 302.829
R64 VPB.t0 VPB.t1 302.829
R65 VPB.t2 VPB.t0 302.829
R66 VPB.t6 VPB 257.93
R67 VPB.n1 VPB.t6 176.21
R68 VPB.n1 VPB.t2 100.129
R69 VPB.n0 VPB 79.7039
R70 VPB.n0 VPB.t4 20.9327
R71 VPB.t3 VPB.t5 8.85643
R72 VPB.t3 VPB.n0 7.32698
R73 VPB.t4 VPB.t5 0.805585
R74 X.n6 X.n5 615.569
R75 X X.n2 587.213
R76 X.n4 X.n0 111.602
R77 X.n3 X.n1 107.365
R78 X.n5 X.t4 41.3353
R79 X.n5 X.t6 41.3353
R80 X.n2 X.t7 41.3353
R81 X.n2 X.t5 41.3353
R82 X.n0 X.t2 29.1897
R83 X.n0 X.t3 22.7032
R84 X.n1 X.t0 22.7032
R85 X.n1 X.t1 22.7032
R86 X X.n3 11.6711
R87 X X.n6 6.27501
R88 X.n4 X 3.01226
R89 X.n6 X.n4 2.76128
R90 X.n3 X 0.376971
R91 A0.n2 A0.t2 246.405
R92 A0.n1 A0.n0 244.214
R93 A0.n1 A0.t0 214.793
R94 A0.n2 A0.t1 212.883
R95 A0 A0.n3 154.715
R96 A0.n3 A0.n1 51.852
R97 A0.n3 A0.n2 11.6853
R98 a_722_391.n1 a_722_391.n0 1083.16
R99 a_722_391.n0 a_722_391.t3 29.5505
R100 a_722_391.n0 a_722_391.t2 29.5505
R101 a_722_391.t1 a_722_391.n1 29.5505
R102 a_722_391.n1 a_722_391.t0 29.5505
R103 VGND.n5 VGND.t5 324.594
R104 VGND.n7 VGND.n6 205.154
R105 VGND.n10 VGND.n9 125.681
R106 VGND.n1 VGND.n0 120.406
R107 VGND.n16 VGND.n15 117.419
R108 VGND.n9 VGND.t8 68.2541
R109 VGND.n6 VGND.t4 52.5005
R110 VGND.n9 VGND.t0 45.6041
R111 VGND.n6 VGND.t7 39.3755
R112 VGND.n0 VGND.t6 39.3755
R113 VGND.n15 VGND.t1 37.2978
R114 VGND.n14 VGND.n3 36.1417
R115 VGND.n18 VGND.n17 36.1417
R116 VGND.n0 VGND.t2 35.7861
R117 VGND.n15 VGND.t3 34.0546
R118 VGND.n8 VGND.n7 31.624
R119 VGND.n10 VGND.n8 25.977
R120 VGND.n10 VGND.n3 21.4593
R121 VGND.n20 VGND.n1 11.4685
R122 VGND.n17 VGND.n16 9.78874
R123 VGND.n19 VGND.n18 9.3005
R124 VGND.n17 VGND.n2 9.3005
R125 VGND.n14 VGND.n13 9.3005
R126 VGND.n12 VGND.n3 9.3005
R127 VGND.n11 VGND.n10 9.3005
R128 VGND.n8 VGND.n4 9.3005
R129 VGND.n18 VGND.n1 7.52991
R130 VGND.n7 VGND.n5 5.16544
R131 VGND.n16 VGND.n14 1.50638
R132 VGND.n5 VGND.n4 0.383817
R133 VGND VGND.n20 0.163644
R134 VGND.n20 VGND.n19 0.144205
R135 VGND.n11 VGND.n4 0.122949
R136 VGND.n12 VGND.n11 0.122949
R137 VGND.n13 VGND.n12 0.122949
R138 VGND.n13 VGND.n2 0.122949
R139 VGND.n19 VGND.n2 0.122949
R140 VNB.n0 VNB 6767.45
R141 VNB.t3 VNB.t7 3857.22
R142 VNB VNB.t0 2164.52
R143 VNB.t6 VNB 1667.64
R144 VNB.t4 VNB.t2 1478.22
R145 VNB.t1 VNB.t6 1462.39
R146 VNB.n0 VNB.t5 1247.24
R147 VNB.t0 VNB.t1 1205.83
R148 VNB.t5 VNB.t4 1154.86
R149 VNB.t2 VNB.t3 993.177
R150 VNB.t0 VNB.n0 123.603
R151 A1.n1 A1.n0 246.405
R152 A1.n4 A1.n3 244.214
R153 A1.n4 A1.t1 213.614
R154 A1.n1 A1.t0 212.883
R155 A1 A1.n2 158.788
R156 A1.n6 A1.n5 152
R157 A1.n5 A1.n2 49.6611
R158 A1.n6 A1 12.2187
R159 A1.n2 A1.n1 10.955
R160 A1 A1.n6 6.4005
R161 A1.n5 A1.n4 4.38232
R162 a_936_391.n1 a_936_391.n0 1093.07
R163 a_936_391.n0 a_936_391.t3 29.5505
R164 a_936_391.n0 a_936_391.t2 29.5505
R165 a_936_391.t1 a_936_391.n1 29.5505
R166 a_936_391.n1 a_936_391.t0 29.5505
R167 a_937_119.n0 a_937_119.t2 540.639
R168 a_937_119.t1 a_937_119.n0 26.2505
R169 a_937_119.n0 a_937_119.t0 26.2505
C0 a_709_119# A1 0.083213f
C1 S X 0.226064f
C2 VPB A0 0.078979f
C3 VGND a_193_241# 0.567789f
C4 a_709_119# VGND 0.171903f
C5 VPB a_193_241# 0.271741f
C6 S A0 7.61e-22
C7 VPWR X 0.037729f
C8 a_709_119# VPB 0.002762f
C9 S a_193_241# 0.153427f
C10 VPWR A0 0.014355f
C11 a_709_119# S 0.045412f
C12 VPWR a_193_241# 0.111404f
C13 X A0 4.72e-20
C14 a_709_119# VPWR 0.00548f
C15 X a_193_241# 0.160982f
C16 a_709_119# X 4.32e-19
C17 A1 VGND 0.012328f
C18 A0 a_193_241# 0.144887f
C19 VPB A1 0.081466f
C20 a_709_119# A0 0.062601f
C21 VPB VGND 0.015811f
C22 a_709_119# a_193_241# 0.272795f
C23 VPWR A1 0.018938f
C24 S VGND 0.090944f
C25 VPB S 0.131119f
C26 VPWR VGND 0.141394f
C27 X A1 3.1e-20
C28 VPB VPWR 0.217984f
C29 A0 A1 0.091601f
C30 X VGND 0.371736f
C31 VPB X 0.01255f
C32 S VPWR 0.078766f
C33 A1 a_193_241# 0.167779f
C34 A0 VGND 0.010801f
C35 VGND VNB 0.978512f
C36 A1 VNB 0.244746f
C37 A0 VNB 0.210289f
C38 X VNB 0.02879f
C39 VPWR VNB 0.78904f
C40 S VNB 0.315005f
C41 VPB VNB 2.04506f
C42 a_709_119# VNB 0.039253f
C43 a_193_241# VNB 1.20292f
.ends

* NGSPICE file created from sky130_fd_sc_hs__mux2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__mux2_2 VNB VPB VPWR VGND S A1 A0 X
X0 a_116_368.t1 A0.t0 a_27_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X1 VPWR.t4 a_116_368.t4 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.392 pd=2.94 as=0.168 ps=1.42 w=1.12 l=0.15
X2 X.t0 a_116_368.t5 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2086 ps=1.515 w=1.12 l=0.15
X3 a_38_74.t1 a_459_48.t2 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2183 pd=2.07 as=0.20535 ps=1.295 w=0.74 l=0.15
X4 X.t3 a_116_368.t6 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.137875 ps=1.155 w=0.74 l=0.15
X5 VPWR.t1 S.t0 a_27_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.295 ps=2.59 w=1 l=0.15
X6 a_116_368.t0 A0.t1 a_38_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.21275 pd=1.315 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 VGND.t2 a_116_368.t7 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_206_368.t1 A1.t0 a_116_368.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X9 VPWR.t2 S.t1 a_459_48.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2086 pd=1.515 as=0.2478 ps=2.27 w=0.84 l=0.15
X10 VGND.t0 S.t2 a_270_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.20535 pd=1.295 as=0.0888 ps=0.98 w=0.74 l=0.15
X11 a_206_368.t0 a_459_48.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2 ps=1.4 w=1 l=0.15
X12 a_270_74.t1 A1.t1 a_116_368.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.21275 ps=1.315 w=0.74 l=0.15
X13 VGND.t1 S.t3 a_459_48.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.137875 pd=1.155 as=0.15675 ps=1.67 w=0.55 l=0.15
R0 A0.n0 A0.t0 257.634
R1 A0.n0 A0.t1 169.535
R2 A0 A0.n0 158.788
R3 a_27_368.t0 a_27_368.t1 1157.21
R4 a_116_368.n3 a_116_368.n0 493.64
R5 a_116_368.n4 a_116_368.n3 327.286
R6 a_116_368.n3 a_116_368.n1 266.546
R7 a_116_368.n2 a_116_368.t5 253.202
R8 a_116_368.n0 a_116_368.t4 240.197
R9 a_116_368.n2 a_116_368.t6 179.947
R10 a_116_368.n0 a_116_368.t7 179.947
R11 a_116_368.n0 a_116_368.n2 70.4873
R12 a_116_368.n1 a_116_368.t0 47.8383
R13 a_116_368.n1 a_116_368.t2 45.4059
R14 a_116_368.n4 a_116_368.t3 29.5505
R15 a_116_368.t1 a_116_368.n4 29.5505
R16 VPB.t0 VPB.t3 618.011
R17 VPB.t6 VPB.t1 515.861
R18 VPB.t1 VPB.t0 280.914
R19 VPB.t3 VPB.t4 278.361
R20 VPB VPB.t2 257.93
R21 VPB.t4 VPB.t5 229.839
R22 VPB.t2 VPB.t6 229.839
R23 X X.n0 593.047
R24 X.n2 X.n1 185
R25 X.n0 X.t1 26.3844
R26 X.n0 X.t0 26.3844
R27 X.n1 X.t2 22.7032
R28 X.n1 X.t3 22.7032
R29 X X.n2 4.75479
R30 X.n2 X 2.01193
R31 VPWR.n5 VPWR.t4 842.01
R32 VPWR.n4 VPWR.n3 691.586
R33 VPWR.n1 VPWR.n0 604.976
R34 VPWR.n3 VPWR.t2 56.2862
R35 VPWR.n0 VPWR.t0 39.4005
R36 VPWR.n0 VPWR.t1 39.4005
R37 VPWR.n8 VPWR.n7 36.1417
R38 VPWR.n9 VPWR.n8 36.1417
R39 VPWR.n3 VPWR.t3 30.268
R40 VPWR.n7 VPWR.n4 20.3299
R41 VPWR.n9 VPWR.n1 17.6946
R42 VPWR.n7 VPWR.n6 9.3005
R43 VPWR.n8 VPWR.n2 9.3005
R44 VPWR.n10 VPWR.n9 9.3005
R45 VPWR.n11 VPWR.n1 7.42496
R46 VPWR.n5 VPWR.n4 6.70329
R47 VPWR.n6 VPWR.n5 0.692082
R48 VPWR VPWR.n11 0.52393
R49 VPWR.n11 VPWR.n10 0.152994
R50 VPWR.n6 VPWR.n2 0.122949
R51 VPWR.n10 VPWR.n2 0.122949
R52 a_459_48.t1 a_459_48.n1 753.759
R53 a_459_48.n0 a_459_48.t2 326.154
R54 a_459_48.n1 a_459_48.t0 290.147
R55 a_459_48.n0 a_459_48.t3 245.018
R56 a_459_48.n1 a_459_48.n0 209.689
R57 VGND.n1 VGND.n0 322.601
R58 VGND.n5 VGND.n4 201.904
R59 VGND.n3 VGND.t2 161.363
R60 VGND.n0 VGND.t4 67.2978
R61 VGND.n4 VGND.t1 52.3641
R62 VGND.n9 VGND.n1 41.1563
R63 VGND.n7 VGND.n6 36.1417
R64 VGND.n4 VGND.t3 31.639
R65 VGND.n0 VGND.t0 22.7032
R66 VGND.n6 VGND.n5 18.0711
R67 VGND.n6 VGND.n2 9.3005
R68 VGND.n8 VGND.n7 9.3005
R69 VGND.n5 VGND.n3 6.68354
R70 VGND.n7 VGND.n1 2.63579
R71 VGND.n3 VGND.n2 0.650615
R72 VGND VGND.n9 0.650547
R73 VGND.n9 VGND.n8 0.149466
R74 VGND.n8 VGND.n2 0.122949
R75 a_38_74.t0 a_38_74.t1 577.143
R76 VNB.t6 VNB.t3 3118.11
R77 VNB.t1 VNB.t2 1674.54
R78 VNB.t0 VNB.t6 1628.35
R79 VNB.t3 VNB.t5 1304.99
R80 VNB VNB.t1 1270.34
R81 VNB.t5 VNB.t4 993.177
R82 VNB.t2 VNB.t0 900.788
R83 S S.n0 303.346
R84 S.n1 S.t2 245.25
R85 S.n0 S.t1 241.464
R86 S.n1 S.t0 229.988
R87 S S.n1 159.565
R88 S.n0 S.t3 155.847
R89 A1.n0 A1.t0 258.738
R90 A1.n0 A1.t1 170.638
R91 A1 A1.n0 165.666
R92 a_206_368.t0 a_206_368.t1 1133.22
R93 a_270_74.t0 a_270_74.t1 38.9194
C0 S VPWR 0.02434f
C1 A0 VGND 0.009579f
C2 S X 0.00703f
C3 A1 VGND 0.007919f
C4 VPWR X 0.023888f
C5 S VGND 0.141054f
C6 VPWR VGND 0.085593f
C7 X VGND 0.094664f
C8 VPB A0 0.041613f
C9 VPB A1 0.042803f
C10 VPB S 0.113387f
C11 A0 A1 0.090561f
C12 VPB VPWR 0.153688f
C13 VPB X 0.003997f
C14 A1 S 0.046063f
C15 A0 VPWR 0.00648f
C16 A1 VPWR 0.006352f
C17 VPB VGND 0.012053f
C18 VGND VNB 0.688161f
C19 X VNB 0.017841f
C20 VPWR VNB 0.514098f
C21 S VNB 0.326481f
C22 A1 VNB 0.12558f
C23 A0 VNB 0.173043f
C24 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2b_4 VNB VPB VPWR VGND A_N Y B
X0 VGND.t2 A_N.t0 a_31_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 a_243_74.t7 B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2 a_243_74.t1 a_31_74.t3 Y.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t5 a_31_74.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.203 ps=1.505 w=1.12 l=0.15
X4 VPWR.t5 B.t1 Y.t7 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.1792 ps=1.44 w=1.12 l=0.15
X5 VGND.t3 B.t2 a_243_74.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.27935 pd=1.495 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_243_74.t5 B.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.27935 ps=1.495 w=0.74 l=0.15
X7 VPWR.t1 A_N.t1 a_31_74.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.126 ps=1.14 w=0.84 l=0.15
X8 a_31_74.t0 A_N.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.5376 ps=2.96 w=0.84 l=0.15
X9 VGND.t0 B.t4 a_243_74.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VPWR.t2 a_31_74.t5 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.896 pd=2.72 as=0.3808 ps=1.8 w=1.12 l=0.15
X11 Y.t6 B.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.896 ps=2.72 w=1.12 l=0.15
X12 a_243_74.t2 a_31_74.t6 Y.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15355 ps=1.155 w=0.74 l=0.15
X13 Y.t1 a_31_74.t7 a_243_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.15355 pd=1.155 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 Y.t0 a_31_74.t8 a_243_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
R0 A_N.n1 A_N.t1 286.822
R1 A_N.n4 A_N.t0 179.947
R2 A_N.n5 A_N.n4 179.786
R3 A_N.n1 A_N.t2 169.772
R4 A_N.n2 A_N 160.4
R5 A_N.n3 A_N.n0 152
R6 A_N.n3 A_N.n2 38.5605
R7 A_N.n2 A_N.n1 24.9511
R8 A_N.n4 A_N.n3 10.7746
R9 A_N.n5 A_N.n0 9.06717
R10 A_N A_N.n5 3.06717
R11 A_N A_N.n0 0.667167
R12 a_31_74.n8 a_31_74.n7 323.248
R13 a_31_74.n3 a_31_74.t8 279.933
R14 a_31_74.n7 a_31_74.t2 246.251
R15 a_31_74.n0 a_31_74.t5 226.809
R16 a_31_74.n4 a_31_74.t4 226.809
R17 a_31_74.n6 a_31_74.n5 152
R18 a_31_74.n0 a_31_74.t6 144.454
R19 a_31_74.n2 a_31_74.t7 142.994
R20 a_31_74.n3 a_31_74.t3 141.213
R21 a_31_74.n6 a_31_74.n1 90.0435
R22 a_31_74.n7 a_31_74.n6 44.0325
R23 a_31_74.n8 a_31_74.t1 35.1791
R24 a_31_74.t0 a_31_74.n8 35.1791
R25 a_31_74.n2 a_31_74.n1 27.3413
R26 a_31_74.n4 a_31_74.n3 26.0933
R27 a_31_74.n1 a_31_74.n0 23.1245
R28 a_31_74.n5 a_31_74.n2 19.9621
R29 a_31_74.n5 a_31_74.n4 7.30353
R30 VGND.n21 VGND.t2 278.688
R31 VGND.n13 VGND.n4 204.201
R32 VGND.n6 VGND.n5 185.119
R33 VGND.n8 VGND.n7 185
R34 VGND.n7 VGND.n6 77.0275
R35 VGND.n15 VGND.n14 36.1417
R36 VGND.n15 VGND.n1 36.1417
R37 VGND.n19 VGND.n1 36.1417
R38 VGND.n20 VGND.n19 36.1417
R39 VGND.n4 VGND.t0 34.0546
R40 VGND.n14 VGND.n13 32.377
R41 VGND.n9 VGND.n3 31.2884
R42 VGND.n21 VGND.n20 22.9652
R43 VGND.n6 VGND.t4 22.7032
R44 VGND.n7 VGND.t3 22.7032
R45 VGND.n4 VGND.t1 22.7032
R46 VGND.n13 VGND.n3 15.0593
R47 VGND.n10 VGND.n9 9.3005
R48 VGND.n11 VGND.n3 9.3005
R49 VGND.n13 VGND.n12 9.3005
R50 VGND.n14 VGND.n2 9.3005
R51 VGND.n16 VGND.n15 9.3005
R52 VGND.n17 VGND.n1 9.3005
R53 VGND.n19 VGND.n18 9.3005
R54 VGND.n20 VGND.n0 9.3005
R55 VGND.n10 VGND.n5 7.61187
R56 VGND.n22 VGND.n21 7.27223
R57 VGND.n8 VGND.n5 6.83134
R58 VGND.n9 VGND.n8 0.219929
R59 VGND VGND.n22 0.157962
R60 VGND.n22 VGND.n0 0.149814
R61 VGND.n11 VGND.n10 0.122949
R62 VGND.n12 VGND.n11 0.122949
R63 VGND.n12 VGND.n2 0.122949
R64 VGND.n16 VGND.n2 0.122949
R65 VGND.n17 VGND.n16 0.122949
R66 VGND.n18 VGND.n17 0.122949
R67 VGND.n18 VGND.n0 0.122949
R68 VNB.t2 VNB.t5 2448.29
R69 VNB.t3 VNB.t4 2090.29
R70 VNB.t6 VNB.t7 1304.99
R71 VNB VNB.t2 1189.5
R72 VNB.t0 VNB.t1 1154.86
R73 VNB.t1 VNB.t3 993.177
R74 VNB.t7 VNB.t0 993.177
R75 VNB.t8 VNB.t6 993.177
R76 VNB.t5 VNB.t8 993.177
R77 B.n1 B.t4 252.977
R78 B.n2 B.t1 240.197
R79 B.n7 B.t5 240.197
R80 B.n1 B.t0 179.947
R81 B.n9 B.t2 179.947
R82 B.n3 B.t3 179.947
R83 B.n4 B.n3 167.337
R84 B.n6 B.n5 152
R85 B.n8 B.n0 152
R86 B B.n10 72.9298
R87 B.n9 B.n8 48.2005
R88 B.n7 B.n6 43.0884
R89 B.n10 B.n1 34.0475
R90 B.n6 B.n2 25.5611
R91 B.n10 B.n9 22.038
R92 B.n5 B.n4 9.06717
R93 B.n3 B.n2 8.76414
R94 B B.n0 7.06717
R95 B.n8 B.n7 6.57323
R96 B B.n0 5.73383
R97 B.n5 B 2.0005
R98 B.n4 B 1.73383
R99 a_243_74.n1 a_243_74.t0 313.079
R100 a_243_74.n4 a_243_74.t5 227.862
R101 a_243_74.n1 a_243_74.n0 101.697
R102 a_243_74.n5 a_243_74.n4 95.243
R103 a_243_74.n3 a_243_74.n2 89.3175
R104 a_243_74.n3 a_243_74.n1 62.4507
R105 a_243_74.n4 a_243_74.n3 57.6712
R106 a_243_74.n2 a_243_74.t4 22.7032
R107 a_243_74.n2 a_243_74.t2 22.7032
R108 a_243_74.n0 a_243_74.t3 22.7032
R109 a_243_74.n0 a_243_74.t1 22.7032
R110 a_243_74.t6 a_243_74.n5 22.7032
R111 a_243_74.n5 a_243_74.t7 22.7032
R112 Y Y.n4 253.119
R113 Y.n3 Y.n1 252.924
R114 Y.n3 Y.n2 198.982
R115 Y.n5 Y.n0 105.587
R116 Y Y.n3 57.3054
R117 Y.n0 Y.t5 54.9164
R118 Y.n0 Y.t4 54.9163
R119 Y.n2 Y.t1 34.8654
R120 Y.n2 Y.t2 32.4329
R121 Y.n4 Y.t6 29.9023
R122 Y.n4 Y.t7 26.3844
R123 Y.n1 Y.t3 22.7032
R124 Y.n1 Y.t0 22.7032
R125 Y.n5 Y 14.5072
R126 Y Y.n5 5.97383
R127 Y.n5 Y 1.73023
R128 VPWR.n12 VPWR.n4 292.5
R129 VPWR.n14 VPWR.n13 292.5
R130 VPWR.n11 VPWR.n6 292.5
R131 VPWR.n10 VPWR.n9 292.5
R132 VPWR.n7 VPWR.t5 260.632
R133 VPWR.n2 VPWR.n1 233.293
R134 VPWR.n25 VPWR.t0 218.548
R135 VPWR.n13 VPWR.n11 75.6344
R136 VPWR.n11 VPWR.n10 73.8755
R137 VPWR.n13 VPWR.n12 73.8755
R138 VPWR.n1 VPWR.t1 55.1136
R139 VPWR.n24 VPWR.n23 36.1417
R140 VPWR.n20 VPWR.n19 36.1417
R141 VPWR.n10 VPWR.t4 31.6612
R142 VPWR.n19 VPWR.n18 31.3713
R143 VPWR.n1 VPWR.t3 29.6087
R144 VPWR.n12 VPWR.t2 26.3844
R145 VPWR.n25 VPWR.n24 10.5417
R146 VPWR.n8 VPWR.n5 9.3005
R147 VPWR.n16 VPWR.n15 9.3005
R148 VPWR.n18 VPWR.n17 9.3005
R149 VPWR.n19 VPWR.n3 9.3005
R150 VPWR.n21 VPWR.n20 9.3005
R151 VPWR.n23 VPWR.n22 9.3005
R152 VPWR.n24 VPWR.n0 9.3005
R153 VPWR.n9 VPWR.n7 7.94475
R154 VPWR.n26 VPWR.n25 6.67776
R155 VPWR.n23 VPWR.n2 6.4005
R156 VPWR.n14 VPWR.n6 5.02698
R157 VPWR.n20 VPWR.n2 4.89462
R158 VPWR.n9 VPWR.n8 4.6763
R159 VPWR.n15 VPWR.n4 4.5594
R160 VPWR.n18 VPWR.n4 1.05255
R161 VPWR.n7 VPWR.n5 0.584947
R162 VPWR.n15 VPWR.n14 0.351185
R163 VPWR.n8 VPWR.n6 0.23429
R164 VPWR.n26 VPWR.n0 0.157539
R165 VPWR VPWR.n26 0.150134
R166 VPWR.n16 VPWR.n5 0.122949
R167 VPWR.n17 VPWR.n16 0.122949
R168 VPWR.n17 VPWR.n3 0.122949
R169 VPWR.n21 VPWR.n3 0.122949
R170 VPWR.n22 VPWR.n21 0.122949
R171 VPWR.n22 VPWR.n0 0.122949
R172 VPB.t2 VPB.t4 893.817
R173 VPB VPB.t0 597.582
R174 VPB.t3 VPB.t2 423.925
R175 VPB.t1 VPB.t3 273.253
R176 VPB.t4 VPB.t5 240.054
R177 VPB.t0 VPB.t1 229.839
C0 VPB B 0.149731f
C1 VPB VPWR 0.198333f
C2 VPB A_N 0.133012f
C3 B VPWR 0.087891f
C4 VPB Y 0.021593f
C5 B Y 0.195853f
C6 VPWR A_N 0.101808f
C7 VPB VGND 0.011868f
C8 VPWR Y 0.588731f
C9 B VGND 0.064642f
C10 VPWR VGND 0.099362f
C11 A_N Y 0.001188f
C12 A_N VGND 0.025671f
C13 Y VGND 0.029585f
C14 VGND VNB 0.681592f
C15 Y VNB 0.023717f
C16 A_N VNB 0.290898f
C17 VPWR VNB 0.596758f
C18 B VNB 0.481854f
C19 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2b_2 VNB VPB VPWR VGND B Y A_N
X0 Y.t3 B.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t4 A_N.t0 a_27_74.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.4613 pd=1.97 as=0.295 ps=2.59 w=1 l=0.15
X2 VPWR.t0 a_27_74.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t1 a_27_74.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4613 ps=1.97 w=1.12 l=0.15
X4 a_242_74.t3 B.t1 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10545 ps=1.025 w=0.74 l=0.15
X5 a_242_74.t1 a_27_74.t4 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VGND.t0 A_N.t1 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.16675 pd=1.81 as=0.1824 ps=1.85 w=0.64 l=0.15
X7 Y.t5 a_27_74.t5 a_242_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.20635 ps=2.05 w=0.74 l=0.15
X8 VGND.t1 B.t2 a_242_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t2 B.t3 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B.n1 B.t0 230.459
R1 B.n0 B.t3 226.809
R2 B.n0 B.t1 197.475
R3 B.n1 B.t2 196.013
R4 B B.n2 154.522
R5 B.n2 B.n0 35.7853
R6 B.n2 B.n1 26.2914
R7 VPWR.n4 VPWR.t2 882.412
R8 VPWR.n3 VPWR.n2 605.365
R9 VPWR.n8 VPWR.n1 313.414
R10 VPWR.n1 VPWR.t1 80.1994
R11 VPWR.n1 VPWR.t4 69.4596
R12 VPWR.n7 VPWR.n6 36.1417
R13 VPWR.n2 VPWR.t3 26.3844
R14 VPWR.n2 VPWR.t0 26.3844
R15 VPWR.n6 VPWR.n3 25.224
R16 VPWR.n6 VPWR.n5 9.3005
R17 VPWR.n7 VPWR.n0 9.3005
R18 VPWR.n9 VPWR.n8 8.08026
R19 VPWR.n8 VPWR.n7 7.90638
R20 VPWR.n4 VPWR.n3 6.50549
R21 VPWR.n5 VPWR.n4 0.686474
R22 VPWR VPWR.n9 0.163644
R23 VPWR.n9 VPWR.n0 0.144205
R24 VPWR.n5 VPWR.n0 0.122949
R25 Y.n2 Y.n0 607.051
R26 Y Y.n3 596.621
R27 Y Y.n1 249.623
R28 Y.n3 Y.t0 26.3844
R29 Y.n3 Y.t1 26.3844
R30 Y.n0 Y.t2 26.3844
R31 Y.n0 Y.t3 26.3844
R32 Y.n1 Y.t4 22.7032
R33 Y.n1 Y.t5 22.7032
R34 Y.n2 Y 13.357
R35 Y Y.n2 2.86366
R36 VPB.t4 VPB.t1 510.753
R37 VPB VPB.t4 257.93
R38 VPB.t3 VPB.t2 229.839
R39 VPB.t0 VPB.t3 229.839
R40 VPB.t1 VPB.t0 229.839
R41 A_N.n0 A_N.t1 236.18
R42 A_N.n0 A_N.t0 234.738
R43 A_N A_N.n0 159.442
R44 a_27_74.t0 a_27_74.n3 478.24
R45 a_27_74.n0 a_27_74.t2 300.255
R46 a_27_74.n3 a_27_74.n2 294.993
R47 a_27_74.n2 a_27_74.t3 283.041
R48 a_27_74.n0 a_27_74.t4 203.589
R49 a_27_74.n1 a_27_74.t5 186.374
R50 a_27_74.n3 a_27_74.t1 184.489
R51 a_27_74.n1 a_27_74.n0 94.7938
R52 a_27_74.n2 a_27_74.n1 20.8872
R53 VGND.n1 VGND.t0 249.962
R54 VGND.n1 VGND.n0 139.904
R55 VGND.n0 VGND.t2 23.514
R56 VGND.n0 VGND.t1 22.7032
R57 VGND VGND.n1 0.200718
R58 a_242_74.n0 a_242_74.t3 493.377
R59 a_242_74.n1 a_242_74.n0 156.517
R60 a_242_74.n0 a_242_74.t0 112.532
R61 a_242_74.n1 a_242_74.t2 22.7032
R62 a_242_74.t1 a_242_74.n1 22.7032
R63 VNB.t2 VNB.t0 2482.94
R64 VNB VNB.t2 1143.31
R65 VNB.t3 VNB.t4 1004.72
R66 VNB.t1 VNB.t3 993.177
R67 VNB.t0 VNB.t1 993.177
C0 VPWR Y 0.034395f
C1 VGND VPB 0.006753f
C2 VGND A_N 0.015538f
C3 VGND B 0.050305f
C4 VGND VPWR 0.057776f
C5 VGND Y 0.014644f
C6 VPB A_N 0.044549f
C7 VPB B 0.063274f
C8 VPB VPWR 0.100871f
C9 A_N VPWR 0.015137f
C10 VPB Y 0.004886f
C11 A_N Y 8.24e-20
C12 B VPWR 0.031614f
C13 B Y 0.090004f
C14 VGND VNB 0.444863f
C15 Y VNB 0.01378f
C16 VPWR VNB 0.363767f
C17 B VNB 0.219263f
C18 A_N VNB 0.17134f
C19 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2b_1 VNB VPB VPWR VGND A_N B Y
X0 VPWR.t0 A_N.t0 a_27_112.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2786 pd=1.64 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VPWR.t1 a_27_112.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_269_74.t0 B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.224125 ps=1.365 w=0.74 l=0.15
X3 Y.t2 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2786 ps=1.64 w=1.12 l=0.15
X4 Y.t0 a_27_112.t3 a_269_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3182 pd=2.34 as=0.0888 ps=0.98 w=0.74 l=0.15
X5 VGND.t0 A_N.t1 a_27_112.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.224125 pd=1.365 as=0.15675 ps=1.67 w=0.55 l=0.15
R0 A_N.n1 A_N.t0 195.21
R1 A_N.n3 A_N.n2 184.864
R2 A_N.n1 A_N.n0 167.337
R3 A_N.n2 A_N.t1 149.421
R4 A_N.n3 A_N.n0 9.06717
R5 A_N A_N.n3 3.06717
R6 A_N.n2 A_N.n1 1.46111
R7 A_N.n0 A_N 0.667167
R8 a_27_112.t1 a_27_112.n1 451.139
R9 a_27_112.n1 a_27_112.t0 335.628
R10 a_27_112.n0 a_27_112.t2 264.298
R11 a_27_112.n0 a_27_112.t3 204.048
R12 a_27_112.n1 a_27_112.n0 152
R13 VPWR.n1 VPWR.t1 884.038
R14 VPWR.n1 VPWR.n0 337.363
R15 VPWR.n0 VPWR.t0 63.5958
R16 VPWR.n0 VPWR.t2 43.9461
R17 VPWR VPWR.n1 0.382628
R18 VPB.t0 VPB.t2 342.204
R19 VPB VPB.t0 257.93
R20 VPB.t2 VPB.t1 255.376
R21 Y Y.n0 588.333
R22 Y.n2 Y.n0 585
R23 Y.n1 Y.t0 265.57
R24 Y.n0 Y.t1 35.1791
R25 Y.n0 Y.t2 26.3844
R26 Y Y.n2 6.26717
R27 Y.n2 Y.n1 2.13383
R28 Y.n1 Y 1.46717
R29 B.n0 B.t1 250.909
R30 B.n0 B.t0 220.113
R31 B B.n0 153.935
R32 VGND VGND.n0 96.6906
R33 VGND.n0 VGND.t0 59.618
R34 VGND.n0 VGND.t1 51.2672
R35 a_269_74.t0 a_269_74.t1 38.9194
R36 VNB.t0 VNB.t1 1790.03
R37 VNB VNB.t0 1143.31
R38 VNB.t1 VNB.t2 900.788
C0 B VPWR 0.006625f
C1 VPB B 0.03685f
C2 B A_N 0.068354f
C3 VPB VPWR 0.084627f
C4 B Y 0.015151f
C5 VPWR A_N 0.015521f
C6 VPB A_N 0.059327f
C7 VPWR Y 0.197241f
C8 B VGND 0.015884f
C9 VPB Y 0.020621f
C10 VPWR VGND 0.041756f
C11 A_N Y 0.001095f
C12 VPB VGND 0.007503f
C13 A_N VGND 0.016873f
C14 Y VGND 0.064137f
C15 VGND VNB 0.340772f
C16 Y VNB 0.103376f
C17 A_N VNB 0.197616f
C18 VPWR VNB 0.286967f
C19 B VNB 0.109889f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand2_8 VNB VPB VPWR VGND B A Y
X0 Y.t8 A.t0 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X2 Y.t7 A.t1 a_27_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_27_74.t8 B.t0 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 Y.t0 A.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3808 ps=1.8 w=1.12 l=0.15
X6 Y.t6 A.t3 a_27_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t1 B.t1 Y.t9 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.8904 pd=2.71 as=0.196 ps=1.47 w=1.12 l=0.15
X8 VGND.t6 B.t2 a_27_74.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2035 ps=2.03 w=0.74 l=0.15
X9 VGND.t5 B.t3 a_27_74.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1184 ps=1.06 w=0.74 l=0.15
X10 a_27_74.t11 B.t4 VGND.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.222 ps=1.34 w=0.74 l=0.15
X11 a_27_74.t4 A.t4 Y.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 Y.t4 A.t5 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2368 ps=1.38 w=0.74 l=0.15
X13 Y.t10 B.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=1.4952 ps=4.91 w=1.12 l=0.15
X14 a_27_74.t12 B.t6 VGND.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_27_74.t13 B.t7 VGND.t2 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_27_74.t2 A.t6 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2368 pd=1.38 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_27_74.t1 A.t7 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.19805 pd=2.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VPWR.t3 B.t8 Y.t11 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.196 ps=1.47 w=1.12 l=0.15
X20 a_27_74.t0 A.t8 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 Y.t12 B.t9 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.8904 ps=2.71 w=1.12 l=0.15
X22 VGND.t1 B.t10 a_27_74.t14 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=1.34 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 VGND.t0 B.t11 a_27_74.t15 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n15 A.t3 281.168
R1 A.n5 A.n4 262.349
R2 A.n3 A.t2 261.62
R3 A.n12 A.n2 261.62
R4 A.n20 A.n13 261.62
R5 A.n18 A.n17 165.189
R6 A.n11 A.t6 154.24
R7 A.n6 A.t5 154.24
R8 A.n5 A.t7 154.24
R9 A A.n7 152.8
R10 A.n19 A.n18 152
R11 A.n9 A.n8 152
R12 A.n10 A.n0 152
R13 A.n24 A.n23 152
R14 A.n22 A.n1 152
R15 A.n15 A.t4 142.994
R16 A.n14 A.t8 142.994
R17 A.n21 A.t0 142.994
R18 A.n16 A.t1 140.06
R19 A.n16 A.n15 135.576
R20 A.n10 A.n9 49.6611
R21 A.n23 A.n22 48.9608
R22 A.n11 A.n10 40.1672
R23 A.n7 A.n5 38.7066
R24 A.n17 A.n16 32.3873
R25 A.n17 A.n14 29.7128
R26 A.n20 A.n19 25.0909
R27 A.n7 A.n6 24.1005
R28 A.n9 A.n3 23.3702
R29 A.n21 A.n20 16.5073
R30 A.n19 A.n14 15.1868
R31 A.n18 A.n1 12.1529
R32 A.n12 A.n11 8.03383
R33 A.n24 A.n1 7.77193
R34 A A.n0 7.2005
R35 A.n8 A 6.97193
R36 A.n8 A 4.0005
R37 A A.n0 3.77193
R38 A.n22 A.n21 3.30187
R39 A.n6 A.n3 2.19141
R40 A.n23 A.n12 1.46111
R41 A A.n24 0.571929
R42 a_27_74.n0 a_27_74.t1 257.834
R43 a_27_74.n5 a_27_74.t9 211.566
R44 a_27_74.n3 a_27_74.n2 185
R45 a_27_74.n1 a_27_74.n0 185
R46 a_27_74.n13 a_27_74.n12 185
R47 a_27_74.n15 a_27_74.n14 185
R48 a_27_74.n9 a_27_74.n8 105.6
R49 a_27_74.n7 a_27_74.n6 104.127
R50 a_27_74.n5 a_27_74.n4 102.538
R51 a_27_74.n11 a_27_74.n10 86.1054
R52 a_27_74.n11 a_27_74.n9 73.7803
R53 a_27_74.n9 a_27_74.n7 69.2711
R54 a_27_74.n2 a_27_74.n1 58.3789
R55 a_27_74.n13 a_27_74.n11 56.8241
R56 a_27_74.n14 a_27_74.n3 44.0325
R57 a_27_74.n14 a_27_74.n13 44.0325
R58 a_27_74.n7 a_27_74.n5 29.7199
R59 a_27_74.n8 a_27_74.t10 25.9464
R60 a_27_74.n8 a_27_74.t11 25.9464
R61 a_27_74.n10 a_27_74.t5 22.7032
R62 a_27_74.n10 a_27_74.t12 22.7032
R63 a_27_74.n4 a_27_74.t15 22.7032
R64 a_27_74.n4 a_27_74.t8 22.7032
R65 a_27_74.n6 a_27_74.t14 22.7032
R66 a_27_74.n6 a_27_74.t13 22.7032
R67 a_27_74.n12 a_27_74.t6 22.7032
R68 a_27_74.n12 a_27_74.t4 22.7032
R69 a_27_74.n1 a_27_74.t3 22.7032
R70 a_27_74.n2 a_27_74.t2 22.7032
R71 a_27_74.n15 a_27_74.t7 22.7032
R72 a_27_74.t0 a_27_74.n15 22.7032
R73 a_27_74.n3 a_27_74.n0 18.4325
R74 Y.n2 Y.n0 349.971
R75 Y.n4 Y.t0 337.296
R76 Y.n2 Y.n1 202.457
R77 Y.n4 Y.n3 185
R78 Y.n6 Y.n5 185
R79 Y.n8 Y.n7 185
R80 Y.n10 Y.n9 185
R81 Y.n6 Y.n4 55.7719
R82 Y.n8 Y.n6 39.3148
R83 Y.n0 Y.t9 35.1791
R84 Y Y.n2 31.3256
R85 Y.n10 Y.n8 31.0801
R86 Y.n1 Y.t11 26.3844
R87 Y.n1 Y.t12 26.3844
R88 Y.n0 Y.t10 26.3844
R89 Y.n9 Y.t5 22.7032
R90 Y.n9 Y.t6 22.7032
R91 Y.n7 Y.t1 22.7032
R92 Y.n7 Y.t7 22.7032
R93 Y.n5 Y.t3 22.7032
R94 Y.n5 Y.t8 22.7032
R95 Y.n3 Y.t2 22.7032
R96 Y.n3 Y.t4 22.7032
R97 Y Y.n10 9.24753
R98 VNB.t2 VNB.t3 1824.67
R99 VNB.t14 VNB.t11 1732.28
R100 VNB VNB.t9 1120.21
R101 VNB.t11 VNB.t10 1085.56
R102 VNB.t3 VNB.t1 993.177
R103 VNB.t7 VNB.t2 993.177
R104 VNB.t0 VNB.t7 993.177
R105 VNB.t6 VNB.t0 993.177
R106 VNB.t4 VNB.t6 993.177
R107 VNB.t5 VNB.t4 993.177
R108 VNB.t12 VNB.t5 993.177
R109 VNB.t10 VNB.t12 993.177
R110 VNB.t13 VNB.t14 993.177
R111 VNB.t15 VNB.t13 993.177
R112 VNB.t8 VNB.t15 993.177
R113 VNB.t9 VNB.t8 993.177
R114 VPWR.n22 VPWR.n21 292.5
R115 VPWR.n20 VPWR.n19 292.5
R116 VPWR.n7 VPWR.n6 292.5
R117 VPWR.n13 VPWR.n12 292.5
R118 VPWR.n10 VPWR.t3 258.875
R119 VPWR.n9 VPWR.t0 202.784
R120 VPWR.n3 VPWR.n2 195
R121 VPWR.n28 VPWR.n1 195
R122 VPWR.n30 VPWR.n1 170.423
R123 VPWR.n20 VPWR.n6 80.0317
R124 VPWR.n21 VPWR.n20 74.755
R125 VPWR.n12 VPWR.n6 71.2371
R126 VPWR.n2 VPWR.n1 59.8041
R127 VPWR.n24 VPWR.n23 36.1417
R128 VPWR.n13 VPWR.n11 27.7188
R129 VPWR.n2 VPWR.t2 27.2639
R130 VPWR.n12 VPWR.t4 27.2639
R131 VPWR.n21 VPWR.t1 26.3844
R132 VPWR.n11 VPWR.n10 24.0946
R133 VPWR.n24 VPWR.n3 15.3548
R134 VPWR.n31 VPWR.n30 10.1681
R135 VPWR.n11 VPWR.n8 9.3005
R136 VPWR.n15 VPWR.n14 9.3005
R137 VPWR.n18 VPWR.n17 9.3005
R138 VPWR.n16 VPWR.n5 9.3005
R139 VPWR.n23 VPWR.n4 9.3005
R140 VPWR.n25 VPWR.n24 9.3005
R141 VPWR.n27 VPWR.n26 9.3005
R142 VPWR.n29 VPWR.n0 9.3005
R143 VPWR.n10 VPWR.n9 6.61379
R144 VPWR.n14 VPWR.n7 4.49472
R145 VPWR.n19 VPWR.n18 4.21028
R146 VPWR.n22 VPWR.n5 3.5845
R147 VPWR.n29 VPWR.n28 2.70903
R148 VPWR.n23 VPWR.n22 1.87783
R149 VPWR.n30 VPWR.n29 1.5862
R150 VPWR.n27 VPWR.n3 1.48582
R151 VPWR.n28 VPWR.n27 1.48582
R152 VPWR.n19 VPWR.n5 1.25206
R153 VPWR.n18 VPWR.n7 0.967611
R154 VPWR.n9 VPWR.n8 0.229721
R155 VPWR VPWR.n31 0.161993
R156 VPWR.n31 VPWR.n0 0.145835
R157 VPWR.n15 VPWR.n8 0.122949
R158 VPWR.n17 VPWR.n15 0.122949
R159 VPWR.n17 VPWR.n16 0.122949
R160 VPWR.n16 VPWR.n4 0.122949
R161 VPWR.n25 VPWR.n4 0.122949
R162 VPWR.n26 VPWR.n25 0.122949
R163 VPWR.n26 VPWR.n0 0.122949
R164 VPWR.n14 VPWR.n13 0.114278
R165 VPB.t3 VPB.t0 1246.24
R166 VPB VPB.t2 1062.37
R167 VPB.t1 VPB.t4 888.711
R168 VPB.t2 VPB.t1 255.376
R169 VPB.t4 VPB.t3 229.839
R170 B.n0 B.t8 344.433
R171 B.n4 B.t2 281.168
R172 B.n7 B.t5 221.827
R173 B.n10 B.t1 214.758
R174 B.n0 B.t9 204.048
R175 B.n3 B.t4 196.013
R176 B.n16 B.t3 196.013
R177 B.n1 B.t6 196.013
R178 B.n7 B.t10 163.442
R179 B.n18 B.n17 152
R180 B.n15 B.n14 152
R181 B.n13 B.n2 152
R182 B.n12 B.n11 152
R183 B.n9 B.n8 152
R184 B.n4 B.t0 142.994
R185 B.n5 B.t11 142.994
R186 B.n6 B.t7 142.994
R187 B.n6 B.n5 138.173
R188 B.n5 B.n4 138.173
R189 B.n1 B.n0 128.873
R190 B.n7 B.n6 111.445
R191 B.n15 B.n2 50.1285
R192 B.n10 B.n9 47.5578
R193 B.n11 B.n3 46.2725
R194 B.n17 B.n16 43.7018
R195 B.n13 B.n12 11.6098
R196 B.n17 B.n1 11.5685
R197 B.n8 B 10.2703
R198 B.n14 B 10.1214
R199 B.n9 B.n7 9.6405
R200 B.n18 B 7.44236
R201 B B.n18 6.84701
R202 B.n16 B.n15 6.42717
R203 B.n14 B 4.16794
R204 B.n8 B 4.0191
R205 B.n3 B.n2 3.8565
R206 B.n11 B.n10 1.9285
R207 B B.n13 1.48887
R208 B.n12 B 1.1912
R209 VGND.n6 VGND.n3 215.157
R210 VGND.n9 VGND.n2 211.183
R211 VGND.n12 VGND.n11 116.156
R212 VGND.n5 VGND.n4 93.4416
R213 VGND.n4 VGND.t4 45.8493
R214 VGND.n4 VGND.t1 45.153
R215 VGND.n9 VGND.n1 32.7534
R216 VGND.n12 VGND.n10 25.224
R217 VGND.n3 VGND.t3 22.7032
R218 VGND.n3 VGND.t5 22.7032
R219 VGND.n2 VGND.t2 22.7032
R220 VGND.n2 VGND.t0 22.7032
R221 VGND.n11 VGND.t7 22.7032
R222 VGND.n11 VGND.t6 22.7032
R223 VGND.n10 VGND.n9 14.6829
R224 VGND.n5 VGND.n1 12.424
R225 VGND.n7 VGND.n1 9.3005
R226 VGND.n9 VGND.n8 9.3005
R227 VGND.n10 VGND.n0 9.3005
R228 VGND.n13 VGND.n12 7.16028
R229 VGND.n6 VGND.n5 6.20359
R230 VGND.n7 VGND.n6 0.592618
R231 VGND VGND.n13 0.156488
R232 VGND.n13 VGND.n0 0.151269
R233 VGND.n8 VGND.n7 0.122949
R234 VGND.n8 VGND.n0 0.122949
C0 VPB B 0.277183f
C1 VPB A 0.206318f
C2 VPB VPWR 0.26631f
C3 B A 0.073893f
C4 B VPWR 0.117729f
C5 VPB Y 0.025485f
C6 B Y 0.297417f
C7 A VPWR 0.132374f
C8 VPB VGND 0.016116f
C9 A Y 0.578857f
C10 B VGND 0.144875f
C11 VPWR Y 1.00552f
C12 A VGND 0.050161f
C13 VPWR VGND 0.14287f
C14 Y VGND 0.043823f
C15 VGND VNB 0.924687f
C16 Y VNB 0.082666f
C17 VPWR VNB 0.773233f
C18 A VNB 0.767358f
C19 B VNB 0.805489f
C20 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand3b_2 VNB VPB VPWR VGND Y A_N C B
X0 VGND.t1 C.t0 a_206_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.19445 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 Y.t5 a_27_94.t2 a_403_54.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.24845 ps=2.6 w=0.74 l=0.15
X2 a_206_74.t3 B.t0 a_403_54.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1816 ps=1.38 w=0.74 l=0.15
X3 Y.t2 C.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.1934 ps=1.475 w=1.12 l=0.15
X4 a_206_74.t0 C.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1165 ps=1.065 w=0.74 l=0.15
X5 VPWR.t0 A_N.t0 a_27_94.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.295 ps=2.59 w=1 l=0.15
X6 VPWR.t4 a_27_94.t3 Y.t7 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2856 pd=1.63 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_403_54.t2 a_27_94.t4 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1816 pd=1.38 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 Y.t6 a_27_94.t5 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X9 a_403_54.t0 B.t1 a_206_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VGND.t2 A_N.t1 a_27_94.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.1728 ps=1.82 w=0.64 l=0.15
X11 Y.t3 B.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.2856 ps=1.63 w=1.12 l=0.15
X12 VPWR.t1 C.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1932 ps=1.465 w=1.12 l=0.15
X13 VPWR.t5 B.t3 Y.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2016 ps=1.48 w=1.12 l=0.15
R0 C.n0 C.t3 234.599
R1 C.n2 C.t1 226.809
R2 C.n2 C.t2 201.565
R3 C C.n0 152.732
R4 C.n4 C.n3 152
R5 C.n1 C.t0 142.994
R6 C.n1 C.n0 22.3965
R7 C C.n4 11.7034
R8 C.n3 C.n1 10.7116
R9 C.n3 C.n2 7.30353
R10 C.n4 C 5.85193
R11 a_206_74.n1 a_206_74.n0 330.63
R12 a_206_74.n0 a_206_74.t2 22.7032
R13 a_206_74.n0 a_206_74.t3 22.7032
R14 a_206_74.n1 a_206_74.t1 22.7032
R15 a_206_74.t0 a_206_74.n1 22.7032
R16 VGND.n1 VGND.t1 236.727
R17 VGND.n1 VGND.n0 222.581
R18 VGND.n0 VGND.t0 31.0986
R19 VGND.n0 VGND.t2 26.2505
R20 VGND VGND.n1 0.522834
R21 VNB.t1 VNB.t3 2390.55
R22 VNB.t4 VNB.t6 1293.44
R23 VNB VNB.t5 1108.66
R24 VNB.t5 VNB.t0 1097.11
R25 VNB.t6 VNB.t2 993.177
R26 VNB.t3 VNB.t4 993.177
R27 VNB.t0 VNB.t1 993.177
R28 a_27_94.t0 a_27_94.n3 299.791
R29 a_27_94.n3 a_27_94.n2 263.435
R30 a_27_94.n1 a_27_94.t5 241.166
R31 a_27_94.n0 a_27_94.t3 226.809
R32 a_27_94.n0 a_27_94.t4 205.596
R33 a_27_94.n3 a_27_94.t1 180.733
R34 a_27_94.n2 a_27_94.t2 171.161
R35 a_27_94.n1 a_27_94.n0 25.8219
R36 a_27_94.n2 a_27_94.n1 2.56433
R37 a_403_54.n1 a_403_54.t3 385.498
R38 a_403_54.n1 a_403_54.n0 224.232
R39 a_403_54.t0 a_403_54.n1 211.847
R40 a_403_54.n0 a_403_54.t1 33.2437
R41 a_403_54.n0 a_403_54.t2 33.2437
R42 Y.n3 Y.n1 263.36
R43 Y.n4 Y.n0 256.353
R44 Y Y.n5 207.576
R45 Y.n3 Y.n2 203.315
R46 Y.n0 Y.t0 36.938
R47 Y.n1 Y.t1 30.7817
R48 Y.n1 Y.t2 29.9023
R49 Y.n0 Y.t3 26.3844
R50 Y.n2 Y.t7 26.3844
R51 Y.n2 Y.t6 26.3844
R52 Y.n5 Y.t4 22.7032
R53 Y.n5 Y.t5 22.7032
R54 Y Y.n4 17.2223
R55 Y.n4 Y.n3 16.1065
R56 B.n2 B.t2 242.023
R57 B.n0 B.t3 226.809
R58 B.n0 B.t1 157.893
R59 B.n2 B.t0 154.24
R60 B.n4 B.n3 152
R61 B.n2 B.n1 152
R62 B.n3 B.n2 49.6611
R63 B.n1 B 11.1633
R64 B.n3 B.n0 9.49444
R65 B B.n4 7.29352
R66 B.n4 B 6.99585
R67 B.n1 B 3.12608
R68 VPWR.n14 VPWR.n1 324.034
R69 VPWR.n3 VPWR.n2 316.353
R70 VPWR.n7 VPWR.n5 316.353
R71 VPWR.n6 VPWR.t5 256.281
R72 VPWR.n5 VPWR.t6 48.371
R73 VPWR.n5 VPWR.t4 41.3353
R74 VPWR.n13 VPWR.n12 36.1417
R75 VPWR.n9 VPWR.n8 36.1417
R76 VPWR.n1 VPWR.t0 35.4605
R77 VPWR.n2 VPWR.t1 35.1791
R78 VPWR.n1 VPWR.t2 32.4757
R79 VPWR.n2 VPWR.t3 26.3844
R80 VPWR.n15 VPWR.n14 15.9861
R81 VPWR.n8 VPWR.n7 11.2946
R82 VPWR.n12 VPWR.n3 9.41227
R83 VPWR.n14 VPWR.n13 9.41227
R84 VPWR.n8 VPWR.n4 9.3005
R85 VPWR.n10 VPWR.n9 9.3005
R86 VPWR.n12 VPWR.n11 9.3005
R87 VPWR.n13 VPWR.n0 9.3005
R88 VPWR.n7 VPWR.n6 7.24479
R89 VPWR.n9 VPWR.n3 1.88285
R90 VPWR.n6 VPWR.n4 0.537576
R91 VPWR VPWR.n15 0.163644
R92 VPWR.n15 VPWR.n0 0.144205
R93 VPWR.n10 VPWR.n4 0.122949
R94 VPWR.n11 VPWR.n10 0.122949
R95 VPWR.n11 VPWR.n0 0.122949
R96 VPB VPB.t0 354.974
R97 VPB.t4 VPB.t6 337.098
R98 VPB.t6 VPB.t5 260.485
R99 VPB.t0 VPB.t2 257.93
R100 VPB.t1 VPB.t3 255.376
R101 VPB.t2 VPB.t1 252.823
R102 VPB.t3 VPB.t4 229.839
R103 A_N.n0 A_N.t0 261.983
R104 A_N.n0 A_N.t1 235.821
R105 A_N A_N.n0 160.922
C0 Y VGND 0.011428f
C1 VGND VPB 0.008322f
C2 Y A_N 9.01e-19
C3 VPB A_N 0.068523f
C4 Y C 0.081528f
C5 VGND A_N 0.017291f
C6 VPWR Y 0.565569f
C7 VPB C 0.072358f
C8 VPWR VPB 0.128633f
C9 VGND C 0.032763f
C10 Y B 0.122856f
C11 VPWR VGND 0.072136f
C12 VPB B 0.074647f
C13 A_N C 0.037256f
C14 VPWR A_N 0.017253f
C15 VGND B 0.012329f
C16 VPWR C 0.034278f
C17 VPWR B 0.073578f
C18 Y VPB 0.014639f
C19 VGND VNB 0.533593f
C20 Y VNB 0.018574f
C21 VPWR VNB 0.465812f
C22 B VNB 0.230291f
C23 C VNB 0.233805f
C24 A_N VNB 0.170546f
C25 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand3b_1 VNB VPB VPWR VGND A_N C Y B
X0 Y.t1 C.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.231 ps=1.555 w=1.12 l=0.15
X1 VGND.t0 A_N.t0 a_27_116.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.224125 pd=1.365 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 a_347_78.t0 B.t0 a_269_78.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0888 ps=0.98 w=0.74 l=0.15
X3 Y.t2 a_27_116.t2 a_347_78.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.3404 pd=2.4 as=0.1443 ps=1.13 w=0.74 l=0.15
X4 VPWR.t2 A_N.t1 a_27_116.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 Y.t0 a_27_116.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6 a_269_78.t0 C.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.224125 ps=1.365 w=0.74 l=0.15
X7 VPWR.t3 B.t1 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
R0 C.n0 C.t0 250.909
R1 C.n0 C.t1 213.688
R2 C C.n0 153.935
R3 VPWR.n2 VPWR.n1 321.978
R4 VPWR.n2 VPWR.n0 236.361
R5 VPWR.n0 VPWR.t2 56.9746
R6 VPWR.n0 VPWR.t1 36.6268
R7 VPWR.n1 VPWR.t0 35.1791
R8 VPWR.n1 VPWR.t3 35.1791
R9 VPWR VPWR.n2 0.552453
R10 Y.n3 Y.n2 585
R11 Y.n2 Y.n0 291.433
R12 Y.n4 Y.n1 255.935
R13 Y Y.t2 184.504
R14 Y.n2 Y.t0 26.3844
R15 Y.n1 Y.t3 26.3844
R16 Y.n1 Y.t1 26.3844
R17 Y Y.n4 7.4454
R18 Y Y.n0 5.84378
R19 Y.n0 Y 3.77493
R20 Y.n4 Y.n3 1.30662
R21 Y.n3 Y 0.914786
R22 VPB VPB.t2 337.098
R23 VPB.t2 VPB.t1 298.791
R24 VPB.t3 VPB.t0 280.914
R25 VPB.t1 VPB.t3 229.839
R26 A_N.n0 A_N.t1 204.225
R27 A_N.n0 A_N.t0 181.464
R28 A_N A_N.n0 154.133
R29 a_27_116.t0 a_27_116.n1 398.901
R30 a_27_116.n1 a_27_116.n0 305.661
R31 a_27_116.n0 a_27_116.t3 258.942
R32 a_27_116.n1 a_27_116.t1 225.501
R33 a_27_116.n0 a_27_116.t2 204.048
R34 VGND VGND.n0 96.7685
R35 VGND.n0 VGND.t0 58.915
R36 VGND.n0 VGND.t1 51.6632
R37 VNB.t0 VNB.t2 1790.03
R38 VNB.t1 VNB.t3 1247.24
R39 VNB VNB.t0 1143.31
R40 VNB.t2 VNB.t1 900.788
R41 B.n0 B.t1 250.909
R42 B.n0 B.t0 213.688
R43 B B.n0 156.614
R44 a_269_78.t0 a_269_78.t1 38.9194
R45 a_347_78.t0 a_347_78.t1 63.2437
C0 B VPWR 0.015707f
C1 VPB A_N 0.045064f
C2 VPB Y 0.026528f
C3 C A_N 0.069013f
C4 C Y 0.015379f
C5 VPB VGND 0.006692f
C6 C VGND 0.016392f
C7 B Y 0.054653f
C8 VPWR A_N 0.02157f
C9 VPWR Y 0.340682f
C10 B VGND 0.009854f
C11 VPWR VGND 0.048058f
C12 VPB C 0.035886f
C13 A_N Y 0.001006f
C14 VPB B 0.033732f
C15 A_N VGND 0.014507f
C16 VPB VPWR 0.088332f
C17 C B 0.092062f
C18 Y VGND 0.06861f
C19 C VPWR 0.033493f
C20 VGND VNB 0.392955f
C21 Y VNB 0.117287f
C22 A_N VNB 0.141498f
C23 VPWR VNB 0.319113f
C24 B VNB 0.101216f
C25 C VNB 0.108811f
C26 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand3_4 VNB VPB VPWR VGND C B A Y
X0 VPWR.t1 A.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.4592 ps=1.94 w=1.12 l=0.15
X1 Y.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.4592 pd=1.94 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VGND.t3 C.t0 a_456_82.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_27_82.t4 A.t2 Y.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 Y.t4 A.t3 a_27_82.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19525 ps=2.03 w=0.74 l=0.15
X5 VGND.t2 C.t1 a_456_82.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_27_82.t0 B.t0 a_456_82.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.19525 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_27_82.t7 B.t1 a_456_82.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t3 B.t2 Y.t7 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.742 pd=2.445 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_456_82.t2 C.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2035 ps=2.03 w=0.74 l=0.15
X10 Y.t6 B.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X11 a_27_82.t2 A.t4 Y.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_456_82.t6 B.t4 a_27_82.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t4 C.t3 Y.t8 VPB.t4 sky130_fd_pr__pfet_01v8 ad=1.484 pd=4.89 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_456_82.t5 B.t5 a_27_82.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 Y.t9 C.t4 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.742 ps=2.445 w=1.12 l=0.15
X16 Y.t2 A.t5 a_27_82.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_456_82.t1 C.t5 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t0 226.809
R1 A.n4 A.t1 226.809
R2 A.n0 A.t4 220.007
R3 A A.n1 159.591
R4 A.n8 A.n7 152
R5 A.n5 A.n2 152
R6 A.n4 A.t3 145.113
R7 A.n6 A.t2 142.994
R8 A.n3 A.t5 142.994
R9 A.n7 A.n3 33.3697
R10 A.n6 A.n5 23.8357
R11 A.n5 A.n4 19.5983
R12 A.n7 A.n6 12.1829
R13 A.n1 A.n0 11.1236
R14 A.n8 A.n2 10.1214
R15 A.n3 A.n1 2.64885
R16 A A.n8 2.53073
R17 A.n2 A 1.63771
R18 Y.n2 Y.n0 323.221
R19 Y.n2 Y.n1 203.127
R20 Y.n7 Y.n5 138.5
R21 Y.n7 Y.n6 98.5941
R22 Y.n4 Y.n3 83.8909
R23 Y.n3 Y.t0 63.7309
R24 Y.n3 Y.t1 63.7308
R25 Y.n4 Y.n2 50.4476
R26 Y Y.n4 44.8987
R27 Y.n0 Y.t8 26.3844
R28 Y.n0 Y.t9 26.3844
R29 Y.n1 Y.t7 26.3844
R30 Y.n1 Y.t6 26.3844
R31 Y.n5 Y.t3 22.7032
R32 Y.n5 Y.t2 22.7032
R33 Y.n6 Y.t5 22.7032
R34 Y.n6 Y.t4 22.7032
R35 Y Y.n7 19.9534
R36 VPWR.n22 VPWR.t0 342.877
R37 VPWR.n2 VPWR.n1 315.928
R38 VPWR.n14 VPWR.n13 292.5
R39 VPWR.n12 VPWR.n11 292.5
R40 VPWR.n6 VPWR.n5 292.5
R41 VPWR.n7 VPWR.t4 141.335
R42 VPWR.n12 VPWR.n5 89.7059
R43 VPWR.n13 VPWR.n12 88.8264
R44 VPWR.n21 VPWR.n20 36.1417
R45 VPWR.n1 VPWR.t2 35.1791
R46 VPWR.n7 VPWR.n6 29.8731
R47 VPWR.n16 VPWR.n15 29.4305
R48 VPWR.n5 VPWR.t5 27.2639
R49 VPWR.n13 VPWR.t3 27.2639
R50 VPWR.n1 VPWR.t1 26.3844
R51 VPWR.n20 VPWR.n2 25.224
R52 VPWR.n16 VPWR.n2 22.2123
R53 VPWR.n22 VPWR.n21 20.7064
R54 VPWR.n10 VPWR.n9 9.3005
R55 VPWR.n8 VPWR.n4 9.3005
R56 VPWR.n15 VPWR.n3 9.3005
R57 VPWR.n17 VPWR.n16 9.3005
R58 VPWR.n18 VPWR.n2 9.3005
R59 VPWR.n20 VPWR.n19 9.3005
R60 VPWR.n21 VPWR.n0 9.3005
R61 VPWR.n23 VPWR.n22 9.3005
R62 VPWR.n14 VPWR.n4 5.29117
R63 VPWR.n11 VPWR.n10 5.00672
R64 VPWR.n10 VPWR.n6 0.796944
R65 VPWR.n9 VPWR.n7 0.767524
R66 VPWR.n11 VPWR.n4 0.455611
R67 VPWR.n15 VPWR.n14 0.171167
R68 VPWR.n9 VPWR.n8 0.122949
R69 VPWR.n8 VPWR.n3 0.122949
R70 VPWR.n17 VPWR.n3 0.122949
R71 VPWR.n18 VPWR.n17 0.122949
R72 VPWR.n19 VPWR.n18 0.122949
R73 VPWR.n19 VPWR.n0 0.122949
R74 VPWR.n23 VPWR.n0 0.122949
R75 VPWR VPWR.n23 0.0617245
R76 VPB.t3 VPB.t5 753.361
R77 VPB.t0 VPB.t1 495.43
R78 VPB VPB.t0 257.93
R79 VPB.t1 VPB.t2 255.376
R80 VPB.t5 VPB.t4 229.839
R81 VPB.t2 VPB.t3 229.839
R82 C.n1 C.t4 288.64
R83 C.n3 C.t3 229.487
R84 C.n10 C.t0 193.093
R85 C.n9 C.t5 179.947
R86 C.n4 C.t2 179.947
R87 C.n2 C.t1 179.947
R88 C.n6 C.n1 164.75
R89 C.n11 C.n10 152
R90 C.n9 C.n8 152
R91 C.n7 C.n0 152
R92 C.n6 C.n5 152
R93 C.n10 C.n9 49.6611
R94 C.n9 C.n0 49.6611
R95 C.n5 C.n2 36.5157
R96 C.n5 C.n4 26.2914
R97 C.n4 C.n3 16.7975
R98 C.n2 C.n0 13.146
R99 C.n8 C.n7 9.89141
R100 C C.n6 9.01868
R101 C C.n11 7.27323
R102 C.n11 C 6.69141
R103 C.n3 C.n1 6.57323
R104 C.n8 C 3.2005
R105 C.n7 C 0.873227
R106 a_456_82.n3 a_456_82.n2 142.929
R107 a_456_82.n4 a_456_82.n0 123.79
R108 a_456_82.n3 a_456_82.n1 98.2648
R109 a_456_82.n5 a_456_82.n4 96.6547
R110 a_456_82.n4 a_456_82.n3 63.2325
R111 a_456_82.n1 a_456_82.t3 22.7032
R112 a_456_82.n1 a_456_82.t2 22.7032
R113 a_456_82.n2 a_456_82.t4 22.7032
R114 a_456_82.n2 a_456_82.t1 22.7032
R115 a_456_82.n0 a_456_82.t7 22.7032
R116 a_456_82.n0 a_456_82.t5 22.7032
R117 a_456_82.t0 a_456_82.n5 22.7032
R118 a_456_82.n5 a_456_82.t6 22.7032
R119 VGND.n0 VGND.t1 292.783
R120 VGND.n3 VGND.n2 207.691
R121 VGND.n1 VGND.t3 173.927
R122 VGND.n4 VGND.n3 28.9887
R123 VGND.n2 VGND.t0 22.7032
R124 VGND.n2 VGND.t2 22.7032
R125 VGND.n4 VGND.n0 10.9181
R126 VGND.n5 VGND.n4 9.3005
R127 VGND.n6 VGND.n0 8.02692
R128 VGND.n3 VGND.n1 6.21929
R129 VGND VGND.n6 1.01964
R130 VGND.n5 VGND.n1 0.735283
R131 VGND.n6 VGND.n5 0.149471
R132 VNB.t0 VNB.t2 2240.42
R133 VNB VNB.t7 1120.21
R134 VNB.t1 VNB.t4 993.177
R135 VNB.t3 VNB.t1 993.177
R136 VNB.t2 VNB.t3 993.177
R137 VNB.t10 VNB.t0 993.177
R138 VNB.t11 VNB.t10 993.177
R139 VNB.t9 VNB.t11 993.177
R140 VNB.t6 VNB.t9 993.177
R141 VNB.t5 VNB.t6 993.177
R142 VNB.t8 VNB.t5 993.177
R143 VNB.t7 VNB.t8 993.177
R144 a_27_82.n4 a_27_82.t3 282.094
R145 a_27_82.n2 a_27_82.t0 271.432
R146 a_27_82.n2 a_27_82.n1 200.495
R147 a_27_82.n5 a_27_82.n4 199.306
R148 a_27_82.n3 a_27_82.n0 110.049
R149 a_27_82.n4 a_27_82.n3 64.7534
R150 a_27_82.n3 a_27_82.n2 57.6005
R151 a_27_82.n1 a_27_82.t6 22.7032
R152 a_27_82.n1 a_27_82.t7 22.7032
R153 a_27_82.n0 a_27_82.t5 22.7032
R154 a_27_82.n0 a_27_82.t2 22.7032
R155 a_27_82.n5 a_27_82.t1 22.7032
R156 a_27_82.t4 a_27_82.n5 22.7032
R157 B.n3 B.t3 262.565
R158 B.n2 B.t2 204.048
R159 B.n8 B.t0 193.613
R160 B.n7 B.t4 183.161
R161 B.n3 B.t5 183.161
R162 B.n1 B.t1 183.161
R163 B.n5 B.n4 169.026
R164 B.n9 B.n8 152
R165 B.n7 B.n0 152
R166 B.n6 B.n5 152
R167 B.n8 B.n7 39.4897
R168 B.n7 B.n6 39.4897
R169 B.n2 B.n1 24.3909
R170 B.n4 B.n2 15.0993
R171 B.n6 B.n1 10.4535
R172 B.n4 B.n3 10.4535
R173 B.n9 B.n0 10.1214
R174 B.n5 B 9.22841
R175 B B.n9 3.27492
R176 B B.n0 0.893523
C0 VPB A 0.110809f
C1 VPWR VGND 0.107719f
C2 VPB B 0.126803f
C3 Y VGND 0.026507f
C4 VPB C 0.15481f
C5 A B 0.060041f
C6 A C 2.85e-20
C7 VPB VPWR 0.187428f
C8 A VPWR 0.044169f
C9 B C 0.063015f
C10 VPB Y 0.025107f
C11 B VPWR 0.054135f
C12 A Y 0.329871f
C13 B Y 0.177432f
C14 C VPWR 0.185625f
C15 C Y 0.052845f
C16 VPB VGND 0.010567f
C17 VPWR Y 0.772794f
C18 A VGND 0.022637f
C19 B VGND 0.02304f
C20 C VGND 0.100196f
C21 VGND VNB 0.757715f
C22 Y VNB 0.073255f
C23 VPWR VNB 0.610374f
C24 C VNB 0.441582f
C25 B VNB 0.361662f
C26 A VNB 0.358432f
C27 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand3_2 VNB VPB VPWR VGND Y C B A
X0 Y.t6 A.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1932 ps=1.465 w=1.12 l=0.15
X1 a_283_74.t1 B.t0 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.176975 pd=1.375 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t7 C.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_27_74.t2 C.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 Y.t2 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.196 ps=1.47 w=1.12 l=0.15
X5 VGND.t0 C.t2 a_27_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1998 ps=2.02 w=0.74 l=0.15
X6 VPWR.t3 A.t1 Y.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.1708 ps=1.425 w=1.12 l=0.15
X7 a_27_74.t1 B.t2 a_283_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.179175 ps=1.375 w=0.74 l=0.15
X8 VPWR.t0 C.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_283_74.t3 A.t2 Y.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.179175 pd=1.375 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 Y.t4 A.t3 a_283_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.176975 ps=1.375 w=0.74 l=0.15
X11 VPWR.t1 B.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n0 A.t0 238.494
R1 A.n1 A.t1 226.809
R2 A.n1 A.t3 180.531
R3 A.n0 A.t2 178.34
R4 A A.n2 154.522
R5 A.n2 A.n1 32.1338
R6 A.n2 A.n0 28.4823
R7 VPWR.n8 VPWR.n2 612.393
R8 VPWR.n4 VPWR.n3 605.753
R9 VPWR.n5 VPWR.t1 266.168
R10 VPWR.n10 VPWR.t5 259.171
R11 VPWR.n2 VPWR.t0 35.1791
R12 VPWR.n3 VPWR.t3 34.2996
R13 VPWR.n8 VPWR.n7 27.4829
R14 VPWR.n10 VPWR.n9 26.7299
R15 VPWR.n2 VPWR.t2 26.3844
R16 VPWR.n3 VPWR.t4 26.3844
R17 VPWR.n9 VPWR.n8 25.977
R18 VPWR.n7 VPWR.n4 25.224
R19 VPWR.n7 VPWR.n6 9.3005
R20 VPWR.n8 VPWR.n1 9.3005
R21 VPWR.n9 VPWR.n0 9.3005
R22 VPWR.n11 VPWR.n10 9.3005
R23 VPWR.n5 VPWR.n4 6.59649
R24 VPWR.n6 VPWR.n5 0.612104
R25 VPWR.n6 VPWR.n1 0.122949
R26 VPWR.n1 VPWR.n0 0.122949
R27 VPWR.n11 VPWR.n0 0.122949
R28 VPWR VPWR.n11 0.0617245
R29 Y.n6 Y.n3 348.824
R30 Y.n2 Y.n0 314.231
R31 Y.n5 Y.n4 291.017
R32 Y.n2 Y.n1 194.847
R33 Y.n6 Y.n2 34.7617
R34 Y.n4 Y.t5 27.2639
R35 Y.n4 Y.t2 26.3844
R36 Y.n3 Y.t1 26.3844
R37 Y.n3 Y.t6 26.3844
R38 Y.n1 Y.t0 26.3844
R39 Y.n1 Y.t7 26.3844
R40 Y.n0 Y.t3 22.7032
R41 Y.n0 Y.t4 22.7032
R42 Y.n6 Y.n5 6.71693
R43 Y.n5 Y 5.40377
R44 Y Y.n6 2.13383
R45 VPB VPB.t5 257.93
R46 VPB.t0 VPB.t2 255.376
R47 VPB.t3 VPB.t4 252.823
R48 VPB.t2 VPB.t3 232.393
R49 VPB.t4 VPB.t1 229.839
R50 VPB.t5 VPB.t0 229.839
R51 B.n2 B.n0 266.022
R52 B.n0 B.t3 258.942
R53 B.n1 B.t1 250.909
R54 B.n1 B.t0 220.113
R55 B.n0 B.t2 192.8
R56 B.n2 B.n1 156.731
R57 B B.n2 0.544688
R58 a_27_74.n0 a_27_74.t1 273.952
R59 a_27_74.n0 a_27_74.t3 194.704
R60 a_27_74.n1 a_27_74.n0 94.3463
R61 a_27_74.t0 a_27_74.n1 22.7032
R62 a_27_74.n1 a_27_74.t2 22.7032
R63 a_283_74.n1 a_283_74.n0 517.907
R64 a_283_74.n1 a_283_74.t2 39.2741
R65 a_283_74.n0 a_283_74.t0 33.2437
R66 a_283_74.n0 a_283_74.t3 32.4329
R67 a_283_74.t1 a_283_74.n1 23.0813
R68 VNB.t5 VNB.t0 1281.89
R69 VNB.t1 VNB.t4 1281.89
R70 VNB VNB.t3 1108.66
R71 VNB.t4 VNB.t5 993.177
R72 VNB.t2 VNB.t1 993.177
R73 VNB.t3 VNB.t2 993.177
R74 C.n0 C.t3 266.002
R75 C.n1 C.t0 261.62
R76 C C.n2 166.357
R77 C.n1 C.t2 157.893
R78 C.n0 C.t1 154.24
R79 C.n2 C.n0 49.6611
R80 C.n2 C.n1 9.49444
R81 VGND VGND.n0 210.24
R82 VGND.n0 VGND.t1 22.7032
R83 VGND.n0 VGND.t0 22.7032
C0 VPB C 0.062405f
C1 VPB B 0.07289f
C2 VPB Y 0.013319f
C3 C B 0.05791f
C4 VPB A 0.06302f
C5 VPB VGND 0.006254f
C6 C Y 0.096018f
C7 VPB VPWR 0.113649f
C8 B Y 0.261487f
C9 C VGND 0.029513f
C10 B A 0.204938f
C11 C VPWR 0.051036f
C12 A Y 0.07557f
C13 B VGND 0.018352f
C14 B VPWR 0.083949f
C15 Y VGND 0.012977f
C16 VPWR Y 0.467737f
C17 A VGND 0.011063f
C18 A VPWR 0.032705f
C19 VPWR VGND 0.056542f
C20 VGND VNB 0.418374f
C21 Y VNB 0.031208f
C22 VPWR VNB 0.429105f
C23 A VNB 0.189149f
C24 B VNB 0.259338f
C25 C VNB 0.239262f
C26 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand3_1 VNB VPB VPWR VGND C Y B A
X0 a_233_74.t0 B.t0 a_155_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 VPWR.t2 B.t1 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t0 C.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.42 ps=2.99 w=1.12 l=0.15
X3 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.54 w=1.12 l=0.15
X4 a_155_74.t1 C.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 Y.t3 A.t1 a_233_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
R0 B.n0 B.t1 285.719
R1 B.n0 B.t0 178.34
R2 B B.n0 158.788
R3 a_155_74.t0 a_155_74.t1 38.9194
R4 a_233_74.t0 a_233_74.t1 68.1086
R5 VNB VNB.t2 1616.8
R6 VNB.t0 VNB.t1 1316.54
R7 VNB.t2 VNB.t0 900.788
R8 Y.n2 Y 588.636
R9 Y.n2 Y.n0 585
R10 Y.n3 Y.n2 585
R11 Y.n1 Y.t1 231.4
R12 Y.n1 Y.t3 201.327
R13 Y Y.n1 56.1716
R14 Y.n2 Y.t2 26.3844
R15 Y.n2 Y.t0 26.3844
R16 Y Y.n3 9.74595
R17 Y Y.n0 8.43686
R18 Y Y.n0 2.32777
R19 Y.n3 Y 1.01868
R20 VPWR.n1 VPWR.t0 280.007
R21 VPWR.n1 VPWR.n0 227.593
R22 VPWR.n0 VPWR.t1 38.6969
R23 VPWR.n0 VPWR.t2 35.1791
R24 VPWR VPWR.n1 0.352459
R25 VPB VPB.t0 334.543
R26 VPB.t2 VPB.t1 291.13
R27 VPB.t0 VPB.t2 229.839
R28 C.n0 C.t0 261.62
R29 C.n0 C.t1 160.814
R30 C.n1 C.n0 90.4558
R31 C C.n1 10.4704
R32 C.n1 C 5.75841
R33 A.n0 A.t0 285.719
R34 A.n0 A.t1 178.34
R35 A A.n0 158.4
R36 VGND VGND.t0 162.57
C0 VPWR Y 0.399091f
C1 VGND A 0.010836f
C2 VGND VPWR 0.041234f
C3 VGND Y 0.056053f
C4 VPB C 0.050137f
C5 VPB B 0.030385f
C6 C B 0.096253f
C7 VPB A 0.035925f
C8 VPB VPWR 0.082994f
C9 C VPWR 0.034399f
C10 B A 0.079111f
C11 VPB Y 0.032409f
C12 B VPWR 0.019601f
C13 C Y 0.040305f
C14 VGND VPB 0.006613f
C15 A VPWR 0.015659f
C16 B Y 0.086353f
C17 VGND C 0.058007f
C18 A Y 0.116279f
C19 VGND B 0.064331f
C20 VGND VNB 0.368479f
C21 Y VNB 0.128369f
C22 VPWR VNB 0.311409f
C23 A VNB 0.137698f
C24 B VNB 0.113343f
C25 C VNB 0.191167f
C26 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand3b_4 VNB VPB VPWR VGND A_N C B Y
X0 a_744_74.t7 a_89_172.t3 Y.t8 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_297_82.t7 C.t0 VGND.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.203425 ps=1.425 w=0.74 l=0.15
X2 VGND.t3 C.t1 a_297_82.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.19935 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 VPWR.t2 B.t0 Y.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=1.7472 pd=5.36 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4424 ps=1.91 w=1.12 l=0.15
X5 a_744_74.t6 a_89_172.t4 Y.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11285 ps=1.045 w=0.74 l=0.15
X6 a_744_74.t0 B.t1 a_297_82.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1976 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_297_82.t5 C.t2 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2715 ps=1.56 w=0.74 l=0.15
X8 Y.t6 a_89_172.t5 a_744_74.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_744_74.t1 B.t2 a_297_82.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VPWR.t0 A_N.t0 a_89_172.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.6202 pd=2.25 as=0.126 ps=1.14 w=0.84 l=0.15
X11 a_89_172.t2 A_N.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.5754 ps=3.05 w=0.84 l=0.15
X12 Y.t4 a_89_172.t6 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3808 pd=1.8 as=0.2604 ps=1.585 w=1.12 l=0.15
X13 a_297_82.t2 B.t3 a_744_74.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 Y.t5 a_89_172.t7 a_744_74.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1962 ps=2.05 w=0.74 l=0.15
X15 VGND.t1 C.t3 a_297_82.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2715 pd=1.56 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_297_82.t3 B.t4 a_744_74.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 VPWR.t3 a_89_172.t8 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.4424 pd=1.91 as=0.3808 ps=1.8 w=1.12 l=0.15
X18 VPWR.t6 C.t4 Y.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2604 pd=1.585 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t2 C.t5 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.6202 ps=2.25 w=1.12 l=0.15
X20 VGND.t0 A_N.t2 a_89_172.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.203425 pd=1.425 as=0.19515 ps=2.05 w=0.74 l=0.15
R0 a_89_172.n7 a_89_172.n6 658.471
R1 a_89_172.n1 a_89_172.t3 281.168
R2 a_89_172.n6 a_89_172.t0 264.401
R3 a_89_172.n4 a_89_172.t6 248.321
R4 a_89_172.n0 a_89_172.t8 240.197
R5 a_89_172.n6 a_89_172.n5 187.951
R6 a_89_172.n5 a_89_172.n4 152
R7 a_89_172.n1 a_89_172.t5 142.994
R8 a_89_172.n3 a_89_172.t7 142.994
R9 a_89_172.n0 a_89_172.t4 142.994
R10 a_89_172.n0 a_89_172.n1 122.198
R11 a_89_172.n5 a_89_172.n2 84.114
R12 a_89_172.t1 a_89_172.n7 35.1791
R13 a_89_172.n7 a_89_172.t2 35.1791
R14 a_89_172.n4 a_89_172.n3 34.1196
R15 a_89_172.n2 a_89_172.n0 26.9332
R16 a_89_172.n3 a_89_172.n2 18.5209
R17 Y.n5 Y.t0 860.333
R18 Y.n1 Y.n0 652.232
R19 Y.n2 Y.n1 585
R20 Y.n4 Y.n3 585
R21 Y.n9 Y.n6 209.048
R22 Y.n8 Y.n7 185
R23 Y.n3 Y.n2 66.8398
R24 Y.n5 Y.n4 29.8005
R25 Y.n3 Y.t3 26.3844
R26 Y.n2 Y.t4 26.3844
R27 Y.n0 Y.t1 26.3844
R28 Y.n0 Y.t2 26.3844
R29 Y.n6 Y.t7 25.1356
R30 Y.n6 Y.t5 24.3248
R31 Y.n7 Y.t8 22.7032
R32 Y.n7 Y.t6 22.7032
R33 Y.n4 Y.n1 15.2005
R34 Y Y.n5 13.357
R35 Y Y.n9 9.48125
R36 Y.n8 Y 2.13383
R37 Y.n9 Y.n8 1.67669
R38 a_744_74.n4 a_744_74.t4 255.303
R39 a_744_74.n1 a_744_74.t0 244.671
R40 a_744_74.n1 a_744_74.n0 185
R41 a_744_74.n3 a_744_74.n2 185
R42 a_744_74.n5 a_744_74.n4 185
R43 a_744_74.n4 a_744_74.n3 45.7685
R44 a_744_74.n3 a_744_74.n1 34.4005
R45 a_744_74.n2 a_744_74.t7 34.0546
R46 a_744_74.n2 a_744_74.t3 22.7032
R47 a_744_74.n0 a_744_74.t2 22.7032
R48 a_744_74.n0 a_744_74.t1 22.7032
R49 a_744_74.n5 a_744_74.t5 22.7032
R50 a_744_74.t6 a_744_74.n5 22.7032
R51 VNB.t2 VNB.t9 2286.61
R52 VNB VNB.t0 1859.32
R53 VNB.t5 VNB.t4 1732.28
R54 VNB.t0 VNB.t1 1397.38
R55 VNB.t12 VNB.t8 1154.86
R56 VNB.t4 VNB.t2 1154.86
R57 VNB.t9 VNB.t11 1050.92
R58 VNB.t7 VNB.t3 993.177
R59 VNB.t6 VNB.t7 993.177
R60 VNB.t8 VNB.t6 993.177
R61 VNB.t10 VNB.t12 993.177
R62 VNB.t11 VNB.t10 993.177
R63 VNB.t1 VNB.t5 993.177
R64 C.n2 C.t0 265.012
R65 C.n1 C.t4 226.809
R66 C.n8 C.t5 226.809
R67 C C.n3 156.316
R68 C.n10 C.n9 152
R69 C.n7 C.n0 152
R70 C.n5 C.n4 152
R71 C.n1 C.t1 144.583
R72 C.n2 C.t3 142.994
R73 C.n6 C.t2 142.994
R74 C.n5 C.n3 36.0181
R75 C.n9 C.n8 34.4291
R76 C.n6 C.n5 33.8994
R77 C.n9 C.n1 13.2423
R78 C.n10 C.n0 10.1214
R79 C.n3 C.n2 9.53457
R80 C.n4 C 8.48422
R81 C.n4 C 5.80515
R82 C C.n10 2.53073
R83 C.n7 C.n6 2.11918
R84 C C.n0 1.63771
R85 C.n8 C.n7 1.58951
R86 VGND.n5 VGND.t3 238.608
R87 VGND.n1 VGND.n0 218.444
R88 VGND.n4 VGND.n3 205
R89 VGND.n3 VGND.t2 48.6491
R90 VGND.n3 VGND.t1 48.6491
R91 VGND.n0 VGND.t4 37.2978
R92 VGND.n0 VGND.t0 36.487
R93 VGND.n9 VGND.n8 32.1868
R94 VGND.n11 VGND.n1 28.288
R95 VGND.n8 VGND.n7 25.9931
R96 VGND.n5 VGND.n4 25.4896
R97 VGND.n10 VGND.n9 9.3005
R98 VGND.n8 VGND.n2 9.3005
R99 VGND.n7 VGND.n6 9.3005
R100 VGND.n9 VGND.n1 2.45707
R101 VGND.n7 VGND.n4 1.20392
R102 VGND.n6 VGND.n5 1.17936
R103 VGND VGND.n11 0.163644
R104 VGND.n11 VGND.n10 0.144205
R105 VGND.n6 VGND.n2 0.122949
R106 VGND.n10 VGND.n2 0.122949
R107 a_297_82.n4 a_297_82.n2 857.777
R108 a_297_82.n5 a_297_82.n4 258.387
R109 a_297_82.n2 a_297_82.n0 249.754
R110 a_297_82.n2 a_297_82.n1 185
R111 a_297_82.n4 a_297_82.n3 185
R112 a_297_82.t6 a_297_82.n5 34.0546
R113 a_297_82.n3 a_297_82.t4 22.7032
R114 a_297_82.n3 a_297_82.t7 22.7032
R115 a_297_82.n0 a_297_82.t1 22.7032
R116 a_297_82.n0 a_297_82.t3 22.7032
R117 a_297_82.n1 a_297_82.t0 22.7032
R118 a_297_82.n1 a_297_82.t2 22.7032
R119 a_297_82.n5 a_297_82.t5 22.7032
R120 B.n8 B.n7 314.341
R121 B.n2 B.t1 220.879
R122 B.n9 B.t0 214.758
R123 B.n8 B.t4 186.374
R124 B.n5 B.t2 186.374
R125 B.n1 B.t3 186.374
R126 B B.n2 154.452
R127 B.n4 B.n3 152
R128 B.n6 B.n0 152
R129 B.n11 B.n10 152
R130 B.n10 B.n6 40.4647
R131 B.n5 B.n4 35.7042
R132 B.n2 B.n1 24.9931
R133 B.n4 B.n1 15.4721
R134 B.n11 B.n0 9.26007
R135 B.n3 B 6.80901
R136 B.n3 B 6.26433
R137 B.n6 B.n5 4.76099
R138 B.n10 B.n9 4.16593
R139 B B.n0 2.99624
R140 B.n9 B.n8 1.78569
R141 B B.n11 0.817521
R142 VPWR.n29 VPWR.t1 744.032
R143 VPWR.n16 VPWR.n6 598.317
R144 VPWR.n22 VPWR.n21 585
R145 VPWR.n23 VPWR.n22 585
R146 VPWR.n22 VPWR.n1 585
R147 VPWR.n9 VPWR.n7 585
R148 VPWR.n10 VPWR.n9 585
R149 VPWR.n8 VPWR.t2 181.263
R150 VPWR.n9 VPWR.t3 103.487
R151 VPWR.n22 VPWR.t5 78.6111
R152 VPWR.t5 VPWR.t0 47.6269
R153 VPWR.n6 VPWR.t4 41.3353
R154 VPWR.n6 VPWR.t6 40.4559
R155 VPWR.n28 VPWR.n27 36.1417
R156 VPWR.n20 VPWR.n4 36.1417
R157 VPWR.n15 VPWR.n14 36.1417
R158 VPWR.n16 VPWR.n15 33.8829
R159 VPWR.n27 VPWR.n1 24.5966
R160 VPWR.n29 VPWR.n28 20.7064
R161 VPWR.n10 VPWR.n8 19.0108
R162 VPWR.n12 VPWR.n11 9.3005
R163 VPWR.n14 VPWR.n13 9.3005
R164 VPWR.n15 VPWR.n5 9.3005
R165 VPWR.n17 VPWR.n16 9.3005
R166 VPWR.n18 VPWR.n4 9.3005
R167 VPWR.n20 VPWR.n19 9.3005
R168 VPWR.n3 VPWR.n2 9.3005
R169 VPWR.n25 VPWR.n24 9.3005
R170 VPWR.n27 VPWR.n26 9.3005
R171 VPWR.n28 VPWR.n0 9.3005
R172 VPWR.n30 VPWR.n29 9.3005
R173 VPWR.n21 VPWR.n20 8.40834
R174 VPWR.n24 VPWR.n23 5.77305
R175 VPWR.n11 VPWR.n7 4.93645
R176 VPWR.n14 VPWR.n7 4.26717
R177 VPWR.n21 VPWR.n3 4.01619
R178 VPWR.n11 VPWR.n10 3.26325
R179 VPWR.n23 VPWR.n3 2.25932
R180 VPWR.n16 VPWR.n4 1.12991
R181 VPWR.n12 VPWR.n8 0.445341
R182 VPWR.n24 VPWR.n1 0.418801
R183 VPWR.n13 VPWR.n12 0.122949
R184 VPWR.n13 VPWR.n5 0.122949
R185 VPWR.n17 VPWR.n5 0.122949
R186 VPWR.n18 VPWR.n17 0.122949
R187 VPWR.n19 VPWR.n18 0.122949
R188 VPWR.n19 VPWR.n2 0.122949
R189 VPWR.n25 VPWR.n2 0.122949
R190 VPWR.n26 VPWR.n25 0.122949
R191 VPWR.n26 VPWR.n0 0.122949
R192 VPWR.n30 VPWR.n0 0.122949
R193 VPWR VPWR.n30 0.0617245
R194 VPB.t3 VPB.t2 709.947
R195 VPB.t0 VPB.t5 653.764
R196 VPB VPB.t1 457.125
R197 VPB.t4 VPB.t3 423.925
R198 VPB.t6 VPB.t4 314.113
R199 VPB.t5 VPB.t6 229.839
R200 VPB.t1 VPB.t0 229.839
R201 A_N.n0 A_N.t0 258.558
R202 A_N.n2 A_N.t2 183.161
R203 A_N A_N.n2 178.311
R204 A_N A_N.n0 160.781
R205 A_N.n1 A_N.t1 159.06
R206 A_N.n2 A_N.n1 10.4535
R207 A_N.n1 A_N.n0 4.06556
C0 VPB C 0.122616f
C1 VPB B 0.136917f
C2 VPB VPWR 0.227984f
C3 C VPWR 0.048138f
C4 VPB A_N 0.095813f
C5 C A_N 0.032021f
C6 VPB Y 0.015718f
C7 B VPWR 0.047618f
C8 C Y 0.058855f
C9 VPB VGND 0.011374f
C10 B Y 0.045151f
C11 VPWR A_N 0.021318f
C12 C VGND 0.048871f
C13 VPWR Y 0.095052f
C14 B VGND 0.027056f
C15 A_N Y 3.61e-20
C16 VPWR VGND 0.133528f
C17 A_N VGND 0.012223f
C18 Y VGND 0.027129f
C19 VGND VNB 0.887022f
C20 Y VNB 0.027275f
C21 A_N VNB 0.206562f
C22 VPWR VNB 0.738828f
C23 B VNB 0.412047f
C24 C VNB 0.388728f
C25 VPB VNB 1.79899f
.ends

* NGSPICE file created from sky130_fd_sc_hs__nand4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4_1 VNB VPB VPWR VGND C Y D B A
X0 Y.t2 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2576 ps=1.58 w=1.12 l=0.15
X1 a_259_74.t0 C.t0 a_181_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X2 a_181_74.t0 D.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2923 ps=2.72 w=0.74 l=0.15
X3 Y.t0 A.t0 a_373_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2085 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X4 a_373_74.t1 B.t1 a_259_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 VPWR.t3 C.t1 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2576 pd=1.58 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t3 D.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X7 VPWR.t0 A.t1 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
R0 B.n0 B.t0 285.719
R1 B.n0 B.t1 178.34
R2 B B.n0 158.746
R3 VPWR.n2 VPWR.n1 315.812
R4 VPWR.n7 VPWR.t2 256.943
R5 VPWR.n3 VPWR.t0 256.817
R6 VPWR.n1 VPWR.t1 41.3353
R7 VPWR.n1 VPWR.t3 39.5764
R8 VPWR.n6 VPWR.n5 36.1417
R9 VPWR.n8 VPWR.n7 19.4652
R10 VPWR.n5 VPWR.n2 15.0593
R11 VPWR.n5 VPWR.n4 9.3005
R12 VPWR.n6 VPWR.n0 9.3005
R13 VPWR.n3 VPWR.n2 7.08651
R14 VPWR.n7 VPWR.n6 1.12991
R15 VPWR.n4 VPWR.n3 0.569455
R16 VPWR.n4 VPWR.n0 0.122949
R17 VPWR.n8 VPWR.n0 0.122949
R18 VPWR VPWR.n8 0.0617245
R19 Y.n2 Y.t0 378.428
R20 Y Y.n0 220.571
R21 Y.n2 Y.n1 203.72
R22 Y.n0 Y.t1 35.1791
R23 Y.n0 Y.t2 26.3844
R24 Y.n1 Y.t4 26.3844
R25 Y.n1 Y.t3 26.3844
R26 Y Y.n2 15.1278
R27 VPB VPB.t2 416.264
R28 VPB.t3 VPB.t1 311.56
R29 VPB.t1 VPB.t0 255.376
R30 VPB.t2 VPB.t3 229.839
R31 C.n0 C.t1 285.719
R32 C.n0 C.t0 178.34
R33 C C.n0 158.746
R34 a_181_74.t0 a_181_74.t1 38.9194
R35 a_259_74.t0 a_259_74.t1 68.1086
R36 VNB VNB.t1 1917.06
R37 VNB.t3 VNB.t0 1316.54
R38 VNB.t2 VNB.t3 1316.54
R39 VNB.t1 VNB.t2 900.788
R40 D.n0 D.t1 285.719
R41 D.n0 D.t0 178.34
R42 D D.n0 158.788
R43 VGND VGND.t0 149.5
R44 A.n0 A.t1 277.849
R45 A.n0 A.t0 170.471
R46 A A.n0 158.788
R47 a_373_74.t0 a_373_74.t1 68.1086
C0 A Y 0.055971f
C1 A VGND 0.011866f
C2 VPWR Y 0.446211f
C3 VPB A 0.040569f
C4 VPWR VGND 0.049838f
C5 VPB VPWR 0.106914f
C6 Y VGND 0.147261f
C7 D VPWR 0.019305f
C8 VPB Y 0.022978f
C9 D Y 0.12162f
C10 B A 0.08779f
C11 C VPWR 0.015559f
C12 VPB VGND 0.008813f
C13 D VGND 0.015901f
C14 C Y 0.093919f
C15 B VPWR 0.018034f
C16 VPB D 0.034573f
C17 C VGND 0.009144f
C18 B Y 0.115095f
C19 VPB C 0.031198f
C20 B VGND 0.010631f
C21 D C 0.091737f
C22 VPB B 0.03272f
C23 C B 0.071259f
C24 A VPWR 0.050274f
C25 VGND VNB 0.397535f
C26 Y VNB 0.117345f
C27 VPWR VNB 0.378137f
C28 A VNB 0.169063f
C29 B VNB 0.11093f
C30 C VNB 0.106744f
C31 D VNB 0.133471f
C32 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtn_2 VNB VPB VPWR VGND D GATE_N RESET_B Q
X0 a_232_98.t0 GATE_N.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.168 ps=1.24 w=0.84 l=0.15
X1 Q.t1 a_913_406.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4984 ps=2.01 w=1.12 l=0.15
X2 a_697_74.t1 a_27_136.t2 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.4209 ps=1.98 w=0.64 l=0.15
X3 Q.t3 a_913_406.t4 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.34225 ps=1.665 w=0.74 l=0.15
X4 VGND.t4 a_232_98.t2 a_373_82.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.4209 pd=1.98 as=0.2294 ps=2.1 w=0.74 l=0.15
X5 a_1153_74.t0 a_670_392.t4 a_913_406.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VPWR.t7 a_232_98.t3 a_373_82.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.25825 pd=1.68 as=0.2478 ps=2.27 w=0.84 l=0.15
X7 VPWR.t6 RESET_B.t0 a_913_406.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.4984 pd=2.01 as=0.1736 ps=1.43 w=1.12 l=0.15
X8 a_870_74.t1 a_373_82.t2 a_670_392.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.05775 pd=0.695 as=0.09575 ps=0.965 w=0.42 l=0.15
X9 a_670_392.t0 a_232_98.t4 a_697_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.09575 pd=0.965 as=0.0768 ps=0.88 w=0.64 l=0.15
X10 VPWR.t0 D.t0 a_27_136.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X11 VGND.t2 a_913_406.t5 a_870_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05775 ps=0.695 w=0.42 l=0.15
X12 VPWR.t3 a_913_406.t6 a_778_504.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.26915 pd=1.96 as=0.1449 ps=1.11 w=0.42 l=0.15
X13 VGND.t6 D.t1 a_27_136.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.200625 pd=1.49 as=0.15675 ps=1.67 w=0.55 l=0.15
X14 VGND.t0 a_913_406.t7 Q.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_778_504.t1 a_232_98.t5 a_670_392.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1449 pd=1.11 as=0.16855 ps=1.39 w=0.42 l=0.15
X16 a_670_392.t3 a_373_82.t3 a_586_392.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.16855 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X17 a_232_98.t1 GATE_N.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=2.09 as=0.200625 ps=1.49 w=0.74 l=0.15
X18 a_913_406.t2 a_670_392.t5 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.26915 ps=1.96 w=1.12 l=0.15
X19 a_586_392.t1 a_27_136.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.25825 ps=1.68 w=1 l=0.15
X20 VPWR.t4 a_913_406.t8 Q.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3976 pd=2.95 as=0.168 ps=1.42 w=1.12 l=0.15
R0 GATE_N.n0 GATE_N.t0 213.954
R1 GATE_N.n0 GATE_N.t1 213.688
R2 GATE_N GATE_N.n0 154.133
R3 VPWR.n25 VPWR.n24 712.104
R4 VPWR.n17 VPWR.n16 585
R5 VPWR.n15 VPWR.n14 585
R6 VPWR.n32 VPWR.n1 323.534
R7 VPWR.n9 VPWR.n8 318.089
R8 VPWR.n10 VPWR.t4 266.05
R9 VPWR.n16 VPWR.n15 234.524
R10 VPWR.n8 VPWR.t2 102.897
R11 VPWR.n16 VPWR.t3 70.3576
R12 VPWR.n24 VPWR.t7 65.6672
R13 VPWR.n8 VPWR.t6 53.6478
R14 VPWR.n15 VPWR.t8 48.602
R15 VPWR.n1 VPWR.t5 46.9053
R16 VPWR.n1 VPWR.t0 46.9053
R17 VPWR.n30 VPWR.n2 36.1417
R18 VPWR.n31 VPWR.n30 36.1417
R19 VPWR.n18 VPWR.n4 36.1417
R20 VPWR.n22 VPWR.n4 36.1417
R21 VPWR.n23 VPWR.n22 36.1417
R22 VPWR.n24 VPWR.t1 35.5684
R23 VPWR.n13 VPWR.n7 34.667
R24 VPWR.n26 VPWR.n23 32.4855
R25 VPWR.n9 VPWR.n7 24.0946
R26 VPWR.n25 VPWR.n2 20.3706
R27 VPWR.n18 VPWR.n17 14.3615
R28 VPWR.n33 VPWR.n32 12.5979
R29 VPWR.n11 VPWR.n7 9.3005
R30 VPWR.n13 VPWR.n12 9.3005
R31 VPWR.n6 VPWR.n5 9.3005
R32 VPWR.n19 VPWR.n18 9.3005
R33 VPWR.n20 VPWR.n4 9.3005
R34 VPWR.n22 VPWR.n21 9.3005
R35 VPWR.n23 VPWR.n3 9.3005
R36 VPWR.n27 VPWR.n26 9.3005
R37 VPWR.n28 VPWR.n2 9.3005
R38 VPWR.n30 VPWR.n29 9.3005
R39 VPWR.n31 VPWR.n0 9.3005
R40 VPWR.n10 VPWR.n9 7.03588
R41 VPWR.n32 VPWR.n31 6.4005
R42 VPWR.n14 VPWR.n6 5.54445
R43 VPWR.n17 VPWR.n6 2.60942
R44 VPWR.n14 VPWR.n13 2.2833
R45 VPWR.n26 VPWR.n25 2.19149
R46 VPWR.n11 VPWR.n10 0.248854
R47 VPWR VPWR.n33 0.163644
R48 VPWR.n33 VPWR.n0 0.144205
R49 VPWR.n12 VPWR.n11 0.122949
R50 VPWR.n12 VPWR.n5 0.122949
R51 VPWR.n19 VPWR.n5 0.122949
R52 VPWR.n20 VPWR.n19 0.122949
R53 VPWR.n21 VPWR.n20 0.122949
R54 VPWR.n21 VPWR.n3 0.122949
R55 VPWR.n27 VPWR.n3 0.122949
R56 VPWR.n28 VPWR.n27 0.122949
R57 VPWR.n29 VPWR.n28 0.122949
R58 VPWR.n29 VPWR.n0 0.122949
R59 a_232_98.t0 a_232_98.n1 770.614
R60 a_232_98.t0 a_232_98.n4 768.644
R61 a_232_98.n0 a_232_98.t4 432.779
R62 a_232_98.n1 a_232_98.n0 392.976
R63 a_232_98.n2 a_232_98.t3 284.916
R64 a_232_98.n3 a_232_98.t1 279.125
R65 a_232_98.n3 a_232_98.n2 253.22
R66 a_232_98.n2 a_232_98.t2 200.03
R67 a_232_98.n0 a_232_98.t5 114.341
R68 a_232_98.n4 a_232_98.n3 31.7782
R69 a_232_98.n4 a_232_98.n1 16.0826
R70 VPB.t9 VPB.t2 531.183
R71 VPB.t5 VPB.t8 515.861
R72 VPB.t3 VPB.t10 505.646
R73 VPB.t7 VPB.t3 429.033
R74 VPB VPB.t0 344.759
R75 VPB.t8 VPB.t1 316.668
R76 VPB.t0 VPB.t5 280.914
R77 VPB.t6 VPB.t7 275.807
R78 VPB.t10 VPB.t9 234.946
R79 VPB.t2 VPB.t4 229.839
R80 VPB.t1 VPB.t6 214.517
R81 a_913_406.n3 a_913_406.t5 471.289
R82 a_913_406.n0 a_913_406.t8 303.125
R83 a_913_406.n1 a_913_406.t3 303.125
R84 a_913_406.n2 a_913_406.n1 296.099
R85 a_913_406.n0 a_913_406.t7 206.458
R86 a_913_406.n1 a_913_406.t4 206.458
R87 a_913_406.n5 a_913_406.n4 198.084
R88 a_913_406.n2 a_913_406.t0 195.151
R89 a_913_406.n4 a_913_406.n3 185.434
R90 a_913_406.n3 a_913_406.t6 138.441
R91 a_913_406.n1 a_913_406.n0 86.7605
R92 a_913_406.n5 a_913_406.t2 28.1434
R93 a_913_406.t1 a_913_406.n5 26.3844
R94 a_913_406.n4 a_913_406.n2 8.13229
R95 Q.n2 Q 587.319
R96 Q.n2 Q.n0 585
R97 Q.n3 Q.n2 585
R98 Q Q.n1 145.02
R99 Q.n2 Q.t0 26.3844
R100 Q.n2 Q.t1 26.3844
R101 Q.n1 Q.t2 22.7032
R102 Q.n1 Q.t3 22.7032
R103 Q Q.n3 6.21499
R104 Q Q.n0 5.38021
R105 Q Q.n0 1.48456
R106 Q.n3 Q 0.649775
R107 a_27_136.t0 a_27_136.n1 455.235
R108 a_27_136.n1 a_27_136.n0 355.474
R109 a_27_136.n0 a_27_136.t2 332.58
R110 a_27_136.n0 a_27_136.t3 287.861
R111 a_27_136.n1 a_27_136.t1 215.546
R112 VGND.n1 VGND.n0 275.382
R113 VGND.n17 VGND.t2 244.976
R114 VGND.n11 VGND.n10 185.744
R115 VGND.n26 VGND.n25 185
R116 VGND.n24 VGND.n3 185
R117 VGND.n8 VGND.t0 161.395
R118 VGND.n10 VGND.n9 92.5005
R119 VGND.n25 VGND.n24 82.4101
R120 VGND.n0 VGND.t6 55.6369
R121 VGND.n16 VGND.n7 36.1417
R122 VGND.n18 VGND.n5 36.1417
R123 VGND.n22 VGND.n5 36.1417
R124 VGND.n31 VGND.n30 36.1417
R125 VGND.n32 VGND.n31 36.1417
R126 VGND.n25 VGND.t5 35.0269
R127 VGND.n10 VGND.t1 34.0546
R128 VGND.n17 VGND.n16 33.1299
R129 VGND.n24 VGND.t4 31.3528
R130 VGND.n0 VGND.t3 30.0005
R131 VGND.n23 VGND.n22 28.232
R132 VGND.n32 VGND.n1 22.7142
R133 VGND.n30 VGND.n3 20.8319
R134 VGND.n18 VGND.n17 14.3064
R135 VGND.n27 VGND.n26 12.2833
R136 VGND.n11 VGND.n7 11.7175
R137 VGND.n34 VGND.n1 9.36437
R138 VGND.n33 VGND.n32 9.3005
R139 VGND.n31 VGND.n2 9.3005
R140 VGND.n30 VGND.n29 9.3005
R141 VGND.n28 VGND.n27 9.3005
R142 VGND.n23 VGND.n4 9.3005
R143 VGND.n22 VGND.n21 9.3005
R144 VGND.n20 VGND.n5 9.3005
R145 VGND.n19 VGND.n18 9.3005
R146 VGND.n17 VGND.n6 9.3005
R147 VGND.n16 VGND.n15 9.3005
R148 VGND.n14 VGND.n7 9.3005
R149 VGND.n13 VGND.n12 9.3005
R150 VGND.n9 VGND.n8 8.08165
R151 VGND.n12 VGND.n9 4.5594
R152 VGND.n27 VGND.n3 2.45707
R153 VGND.n12 VGND.n11 2.16306
R154 VGND.n13 VGND.n8 0.587633
R155 VGND VGND.n34 0.161675
R156 VGND.n34 VGND.n33 0.146149
R157 VGND.n26 VGND.n23 0.129793
R158 VGND.n14 VGND.n13 0.122949
R159 VGND.n15 VGND.n14 0.122949
R160 VGND.n15 VGND.n6 0.122949
R161 VGND.n19 VGND.n6 0.122949
R162 VGND.n20 VGND.n19 0.122949
R163 VGND.n21 VGND.n20 0.122949
R164 VGND.n21 VGND.n4 0.122949
R165 VGND.n28 VGND.n4 0.122949
R166 VGND.n29 VGND.n28 0.122949
R167 VGND.n29 VGND.n2 0.122949
R168 VGND.n33 VGND.n2 0.122949
R169 a_697_74.t0 a_697_74.t1 45.0005
R170 VNB.t7 VNB.t3 3383.73
R171 VNB.t4 VNB.t6 2690.81
R172 VNB.t6 VNB.t8 2679.26
R173 VNB.t2 VNB.t7 2286.61
R174 VNB.t9 VNB.t4 1362.73
R175 VNB VNB.t9 1143.31
R176 VNB.t5 VNB.t0 1097.11
R177 VNB.t3 VNB.t1 993.177
R178 VNB.t0 VNB.t2 981.628
R179 VNB.t8 VNB.t5 900.788
R180 a_373_82.t0 a_373_82.n1 748.972
R181 a_373_82.n0 a_373_82.t2 412.647
R182 a_373_82.n0 a_373_82.t3 383.628
R183 a_373_82.n1 a_373_82.t1 330.545
R184 a_373_82.n1 a_373_82.n0 79.7666
R185 a_670_392.n3 a_670_392.n2 727.995
R186 a_670_392.n2 a_670_392.n0 291.327
R187 a_670_392.n1 a_670_392.t5 226.809
R188 a_670_392.n2 a_670_392.n1 215.536
R189 a_670_392.n1 a_670_392.t4 203.762
R190 a_670_392.n3 a_670_392.t1 112.572
R191 a_670_392.n0 a_670_392.t0 40.5809
R192 a_670_392.n0 a_670_392.t2 40.0005
R193 a_670_392.n4 a_670_392.t3 24.0586
R194 a_670_392.n5 a_670_392.n4 11.7119
R195 a_670_392.n4 a_670_392.n3 4.33463
R196 RESET_B.n1 RESET_B.t0 285.719
R197 RESET_B.n1 RESET_B.n0 178.34
R198 RESET_B RESET_B.n1 159.785
R199 a_870_74.t0 a_870_74.t1 78.5719
R200 D.n0 D.t0 212.907
R201 D.n0 D.t1 182.113
R202 D D.n0 153.358
R203 a_778_504.t0 a_778_504.t1 323.644
R204 a_586_392.t0 a_586_392.t1 53.1905
C0 VPB RESET_B 0.034618f
C1 RESET_B VGND 0.04071f
C2 VPB VGND 0.018591f
C3 VPWR RESET_B 0.01832f
C4 VPB VPWR 0.250713f
C5 RESET_B Q 0.004302f
C6 VPWR VGND 0.150774f
C7 VPB Q 0.00964f
C8 VPB D 0.051079f
C9 VGND Q 0.169496f
C10 D VGND 0.008351f
C11 VPWR Q 0.265373f
C12 VPWR D 0.023358f
C13 VPB GATE_N 0.050695f
C14 D Q 7.84e-21
C15 GATE_N VGND 0.007592f
C16 VPWR GATE_N 0.029433f
C17 GATE_N Q 7.46e-21
C18 D GATE_N 0.070924f
C19 Q VNB 0.036266f
C20 VGND VNB 1.01149f
C21 RESET_B VNB 0.112449f
C22 GATE_N VNB 0.10527f
C23 D VNB 0.130177f
C24 VPWR VNB 0.798574f
C25 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtn_4 VNB VPB VPWR VGND D GATE_N RESET_B Q
X0 VPWR.t9 a_888_406# a_747_504.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.21315 pd=1.59 as=0.1512 ps=1.14 w=0.42 l=0.15
X1 a_888_406# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1554 pd=1.21 as=0.147 ps=1.19 w=0.84 l=0.15
X2 a_232_98.t0 GATE_N.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.168 ps=1.24 w=0.84 l=0.15
X3 VGND.t10 a_888_406# a_839_74.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05775 ps=0.695 w=0.42 l=0.15
X4 a_1035_74.t2 RESET_B.t0 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 Q.t7 a_888_406# VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_888_406# a_639_392.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21315 ps=1.59 w=0.84 l=0.15
X7 a_839_74.t0 a_348_392.t2 a_639_392.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.05775 pd=0.695 as=0.09575 ps=0.965 w=0.42 l=0.15
X8 a_747_504.t0 a_232_98.t2 a_639_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.14 as=0.16855 ps=1.39 w=0.42 l=0.15
X9 VPWR RESET_B a_888_406# VPB sky130_fd_pr__pfet_01v8 ad=0.2206 pd=1.555 as=0.1554 ps=1.21 w=0.84 l=0.15
X10 VGND.t3 RESET_B.t1 a_1035_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X11 a_639_392.t3 a_348_392.t3 a_561_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.16855 pd=1.39 as=0.12 ps=1.24 w=1 l=0.15
X12 a_666_74.t1 a_27_136.t2 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.392625 ps=1.975 w=0.64 l=0.15
X13 Q.t3 a_888_406# VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.196 ps=1.47 w=1.12 l=0.15
X14 a_561_392.t1 a_27_136.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.25825 ps=1.68 w=1 l=0.15
X15 a_888_406# a_639_392.t5 a_1035_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X16 Q.t6 a_888_406# VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t1 D.t0 a_27_136.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.200625 pd=1.49 as=0.15675 ps=1.67 w=0.55 l=0.15
X18 VPWR.t0 a_232_98.t3 a_348_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.25825 pd=1.68 as=0.2478 ps=2.27 w=0.84 l=0.15
X19 VPWR.t4 D.t1 a_27_136.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X20 VGND.t2 a_232_98.t4 a_348_392.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.392625 pd=1.975 as=0.2109 ps=2.05 w=0.74 l=0.15
X21 a_1035_74.t0 a_639_392.t6 a_888_406# VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X22 VPWR.t7 a_888_406# Q.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X23 VGND.t6 a_888_406# Q.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 Q.t1 a_888_406# VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2206 ps=1.555 w=1.12 l=0.15
X25 a_232_98.t1 GATE_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2886 pd=2.26 as=0.200625 ps=1.49 w=0.74 l=0.15
X26 VGND.t9 a_888_406# Q.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 a_639_392.t0 a_232_98.t5 a_666_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.09575 pd=0.965 as=0.0768 ps=0.88 w=0.64 l=0.15
X28 VPWR.t5 a_888_406# Q.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
R0 a_747_504.t0 a_747_504.t1 337.714
R1 VPWR.n34 VPWR.n33 712.104
R2 VPWR.n26 VPWR.n25 585
R3 VPWR.n24 VPWR.n23 585
R4 VPWR.n16 VPWR.t6 357.474
R5 VPWR.n12 VPWR.t5 349.731
R6 VPWR.n41 VPWR.n1 323.534
R7 VPWR.n11 VPWR.n10 315.832
R8 VPWR.n25 VPWR.n24 187.619
R9 VPWR.n25 VPWR.t9 70.3576
R10 VPWR.n33 VPWR.t0 65.6672
R11 VPWR.n24 VPWR.t3 62.1493
R12 VPWR.n1 VPWR.t2 46.9053
R13 VPWR.n1 VPWR.t4 46.9053
R14 VPWR.n39 VPWR.n2 36.1417
R15 VPWR.n40 VPWR.n39 36.1417
R16 VPWR.n27 VPWR.n4 36.1417
R17 VPWR.n31 VPWR.n4 36.1417
R18 VPWR.n32 VPWR.n31 36.1417
R19 VPWR.n35 VPWR.n32 36.1417
R20 VPWR.n18 VPWR.n17 36.1417
R21 VPWR.n15 VPWR.n9 36.1417
R22 VPWR.n33 VPWR.t1 35.5684
R23 VPWR.n22 VPWR.n7 35.3887
R24 VPWR.n10 VPWR.t7 35.1791
R25 VPWR.n10 VPWR.t8 26.3844
R26 VPWR.n23 VPWR.n22 17.7498
R27 VPWR.n41 VPWR.n40 16.9417
R28 VPWR.n18 VPWR.n7 12.0476
R29 VPWR.n34 VPWR.n2 11.5998
R30 VPWR.n11 VPWR.n9 9.41227
R31 VPWR.n13 VPWR.n9 9.3005
R32 VPWR.n15 VPWR.n14 9.3005
R33 VPWR.n17 VPWR.n8 9.3005
R34 VPWR.n19 VPWR.n18 9.3005
R35 VPWR.n20 VPWR.n7 9.3005
R36 VPWR.n22 VPWR.n21 9.3005
R37 VPWR.n6 VPWR.n5 9.3005
R38 VPWR.n28 VPWR.n27 9.3005
R39 VPWR.n29 VPWR.n4 9.3005
R40 VPWR.n31 VPWR.n30 9.3005
R41 VPWR.n32 VPWR.n3 9.3005
R42 VPWR.n36 VPWR.n35 9.3005
R43 VPWR.n37 VPWR.n2 9.3005
R44 VPWR.n39 VPWR.n38 9.3005
R45 VPWR.n40 VPWR.n0 9.3005
R46 VPWR.n12 VPWR.n11 8.9986
R47 VPWR.n35 VPWR.n34 8.58799
R48 VPWR.n42 VPWR.n41 7.52053
R49 VPWR.n17 VPWR.n16 6.4005
R50 VPWR.n27 VPWR.n26 4.94977
R51 VPWR.n16 VPWR.n15 4.89462
R52 VPWR.n26 VPWR.n6 4.64763
R53 VPWR.n23 VPWR.n6 1.87566
R54 VPWR.n13 VPWR.n12 0.647735
R55 VPWR VPWR.n42 0.161231
R56 VPWR.n42 VPWR.n0 0.146587
R57 VPWR.n14 VPWR.n13 0.122949
R58 VPWR.n14 VPWR.n8 0.122949
R59 VPWR.n19 VPWR.n8 0.122949
R60 VPWR.n20 VPWR.n19 0.122949
R61 VPWR.n21 VPWR.n20 0.122949
R62 VPWR.n21 VPWR.n5 0.122949
R63 VPWR.n28 VPWR.n5 0.122949
R64 VPWR.n29 VPWR.n28 0.122949
R65 VPWR.n30 VPWR.n29 0.122949
R66 VPWR.n30 VPWR.n3 0.122949
R67 VPWR.n36 VPWR.n3 0.122949
R68 VPWR.n37 VPWR.n36 0.122949
R69 VPWR.n38 VPWR.n37 0.122949
R70 VPWR.n38 VPWR.n0 0.122949
R71 VPB.t3 VPB.t8 1049.6
R72 VPB.t2 VPB.t0 523.521
R73 VPB.t11 VPB.t3 459.678
R74 VPB.t6 VPB.t11 444.356
R75 VPB.t0 VPB.t1 316.668
R76 VPB.t10 VPB.t7 280.914
R77 VPB.t5 VPB.t2 280.914
R78 VPB.t4 VPB.t6 275.807
R79 VPB VPB.t5 273.253
R80 VPB.t9 VPB.t10 255.376
R81 VPB.t8 VPB.t9 229.839
R82 VPB.t1 VPB.t4 199.195
R83 RESET_B.n5 RESET_B.n1 283.236
R84 RESET_B.n3 RESET_B.n2 278.562
R85 RESET_B.n6 RESET_B.n5 152
R86 RESET_B.n4 RESET_B.n0 152
R87 RESET_B.n5 RESET_B.t0 138.173
R88 RESET_B.n3 RESET_B.t1 138.173
R89 RESET_B.n5 RESET_B.n4 34.8686
R90 RESET_B.n6 RESET_B.n0 13.1884
R91 RESET_B.n4 RESET_B.n3 9.23029
R92 RESET_B.n0 RESET_B 3.49141
R93 RESET_B RESET_B.n6 1.93989
R94 GATE_N.n0 GATE_N.t0 213.954
R95 GATE_N.n0 GATE_N.t1 213.688
R96 GATE_N GATE_N.n0 153.423
R97 a_232_98.t0 a_232_98.n1 768.644
R98 a_232_98.t0 a_232_98.n4 768.644
R99 a_232_98.n0 a_232_98.t5 432.779
R100 a_232_98.n1 a_232_98.n0 394.966
R101 a_232_98.n3 a_232_98.t1 282.231
R102 a_232_98.n3 a_232_98.n2 211.886
R103 a_232_98.n2 a_232_98.t3 195.21
R104 a_232_98.n2 a_232_98.t4 192.102
R105 a_232_98.n0 a_232_98.t2 114.341
R106 a_232_98.n4 a_232_98.n3 24.6288
R107 a_232_98.n4 a_232_98.n1 14.516
R108 a_839_74.t0 a_839_74.t1 78.5719
R109 VGND.n12 VGND.t6 300.51
R110 VGND.n1 VGND.n0 275.382
R111 VGND.n24 VGND.t10 244.976
R112 VGND.n11 VGND.n10 209.243
R113 VGND.n18 VGND.n17 204.976
R114 VGND.n31 VGND.n3 185
R115 VGND.n33 VGND.n32 185
R116 VGND.n31 VGND.t2 144.808
R117 VGND.n15 VGND.t8 138.75
R118 VGND.n32 VGND.n31 70.121
R119 VGND.n0 VGND.t1 55.6369
R120 VGND.n22 VGND.n7 36.1417
R121 VGND.n23 VGND.n22 36.1417
R122 VGND.n25 VGND.n5 36.1417
R123 VGND.n29 VGND.n5 36.1417
R124 VGND.n38 VGND.n37 36.1417
R125 VGND.n39 VGND.n38 36.1417
R126 VGND.n30 VGND.n29 35.8765
R127 VGND.n16 VGND.n15 35.7652
R128 VGND.n32 VGND.t5 35.0269
R129 VGND.n18 VGND.n7 33.5064
R130 VGND.n0 VGND.t0 30.0005
R131 VGND.n11 VGND.n9 28.2358
R132 VGND.n17 VGND.t4 26.2505
R133 VGND.n17 VGND.t3 26.2505
R134 VGND.n10 VGND.t7 22.7032
R135 VGND.n10 VGND.t9 22.7032
R136 VGND.n39 VGND.n1 22.1206
R137 VGND.n37 VGND.n3 14.9677
R138 VGND.n18 VGND.n16 13.9299
R139 VGND.n15 VGND.n9 11.6711
R140 VGND.n40 VGND.n39 9.3005
R141 VGND.n38 VGND.n2 9.3005
R142 VGND.n37 VGND.n36 9.3005
R143 VGND.n35 VGND.n34 9.3005
R144 VGND.n30 VGND.n4 9.3005
R145 VGND.n29 VGND.n28 9.3005
R146 VGND.n27 VGND.n5 9.3005
R147 VGND.n26 VGND.n25 9.3005
R148 VGND.n23 VGND.n6 9.3005
R149 VGND.n22 VGND.n21 9.3005
R150 VGND.n20 VGND.n7 9.3005
R151 VGND.n19 VGND.n18 9.3005
R152 VGND.n16 VGND.n8 9.3005
R153 VGND.n15 VGND.n14 9.3005
R154 VGND.n13 VGND.n9 9.3005
R155 VGND.n41 VGND.n1 9.10055
R156 VGND.n24 VGND.n23 8.65932
R157 VGND.n34 VGND.n33 7.12398
R158 VGND.n12 VGND.n11 6.26985
R159 VGND.n34 VGND.n3 3.67354
R160 VGND.n33 VGND.n30 3.56224
R161 VGND.n25 VGND.n24 2.63579
R162 VGND.n13 VGND.n12 0.733933
R163 VGND VGND.n41 0.161517
R164 VGND.n41 VGND.n40 0.146304
R165 VGND.n14 VGND.n13 0.122949
R166 VGND.n14 VGND.n8 0.122949
R167 VGND.n19 VGND.n8 0.122949
R168 VGND.n20 VGND.n19 0.122949
R169 VGND.n21 VGND.n20 0.122949
R170 VGND.n21 VGND.n6 0.122949
R171 VGND.n26 VGND.n6 0.122949
R172 VGND.n27 VGND.n26 0.122949
R173 VGND.n28 VGND.n27 0.122949
R174 VGND.n28 VGND.n4 0.122949
R175 VGND.n35 VGND.n4 0.122949
R176 VGND.n36 VGND.n35 0.122949
R177 VGND.n36 VGND.n2 0.122949
R178 VGND.n40 VGND.n2 0.122949
R179 VNB.t0 VNB.t4 2529.13
R180 VNB.t4 VNB.t9 2482.94
R181 VNB.t6 VNB.t13 2286.61
R182 VNB.t14 VNB.t7 2286.61
R183 VNB.t2 VNB.t0 1362.73
R184 VNB VNB.t2 1143.31
R185 VNB.t3 VNB.t8 1097.11
R186 VNB.t12 VNB.t11 993.177
R187 VNB.t10 VNB.t12 993.177
R188 VNB.t13 VNB.t10 993.177
R189 VNB.t5 VNB.t6 993.177
R190 VNB.t1 VNB.t5 993.177
R191 VNB.t7 VNB.t1 993.177
R192 VNB.t8 VNB.t14 981.628
R193 VNB.t9 VNB.t3 900.788
R194 a_1035_74.n1 a_1035_74.t3 196.63
R195 a_1035_74.t2 a_1035_74.n1 189.601
R196 a_1035_74.n1 a_1035_74.n0 88.1174
R197 a_1035_74.n0 a_1035_74.t1 26.2505
R198 a_1035_74.n0 a_1035_74.t0 26.2505
R199 Q.n2 Q.n0 256.635
R200 Q.n2 Q.n1 202.203
R201 Q.n5 Q.n4 158.883
R202 Q.n5 Q.n3 96.9112
R203 Q Q.n2 50.2294
R204 Q.n1 Q.t0 35.1791
R205 Q.n1 Q.t3 35.1791
R206 Q.n0 Q.t2 26.3844
R207 Q.n0 Q.t1 26.3844
R208 Q.n3 Q.t5 22.7032
R209 Q.n3 Q.t6 22.7032
R210 Q.n4 Q.t4 22.7032
R211 Q.n4 Q.t7 22.7032
R212 Q Q.n5 14.9338
R213 a_639_392.n6 a_639_392.n5 735.731
R214 a_639_392.n5 a_639_392.n0 279.781
R215 a_639_392.n2 a_639_392.n1 221.988
R216 a_639_392.n4 a_639_392.t4 221.988
R217 a_639_392.n2 a_639_392.t6 148.488
R218 a_639_392.n3 a_639_392.t5 138.173
R219 a_639_392.n6 a_639_392.t1 112.572
R220 a_639_392.n5 a_639_392.n4 100.383
R221 a_639_392.n0 a_639_392.t0 40.5809
R222 a_639_392.n0 a_639_392.t2 40.0005
R223 a_639_392.n3 a_639_392.n2 24.8199
R224 a_639_392.n7 a_639_392.t3 24.0586
R225 a_639_392.n8 a_639_392.n7 11.7119
R226 a_639_392.n4 a_639_392.n3 7.55423
R227 a_639_392.n7 a_639_392.n6 4.33463
R228 a_348_392.t0 a_348_392.n1 721.119
R229 a_348_392.n0 a_348_392.t2 410.514
R230 a_348_392.n0 a_348_392.t3 390.322
R231 a_348_392.n1 a_348_392.t1 335.399
R232 a_348_392.n1 a_348_392.n0 79.5727
R233 a_561_392.t0 a_561_392.t1 47.2805
R234 a_27_136.t1 a_27_136.n1 457.394
R235 a_27_136.n0 a_27_136.t2 348.647
R236 a_27_136.n1 a_27_136.n0 342.923
R237 a_27_136.n0 a_27_136.t3 266.44
R238 a_27_136.n1 a_27_136.t0 215.546
R239 a_666_74.t0 a_666_74.t1 45.0005
R240 D.n0 D.t1 213.595
R241 D.n0 D.t0 182.8
R242 D D.n0 153.745
C0 RESET_B Q 0.005819f
C1 a_888_406# D 4.53e-21
C2 a_888_406# RESET_B 0.234205f
C3 VGND Q 0.281251f
C4 a_888_406# VGND 0.107418f
C5 a_888_406# Q 0.385895f
C6 VPB VPWR 0.288962f
C7 VPB GATE_N 0.048809f
C8 VPB D 0.049102f
C9 VPB RESET_B 0.104552f
C10 VPWR GATE_N 0.021394f
C11 VPWR D 0.036534f
C12 VPB VGND 0.019057f
C13 VPWR RESET_B 0.039877f
C14 D GATE_N 0.074091f
C15 VPB Q 0.019083f
C16 VPWR VGND 0.157916f
C17 GATE_N VGND 0.009685f
C18 a_888_406# VPB 0.301743f
C19 D VGND 0.007993f
C20 VPWR Q 0.421202f
C21 RESET_B VGND 0.048193f
C22 GATE_N Q 1.14e-21
C23 a_888_406# VPWR 0.525097f
C24 a_888_406# GATE_N 2.29e-21
C25 D Q 3.75e-21
C26 Q VNB 0.075008f
C27 VGND VNB 1.15003f
C28 RESET_B VNB 0.239445f
C29 GATE_N VNB 0.104353f
C30 D VNB 0.129662f
C31 VPWR VNB 0.906433f
C32 VPB VNB 2.22754f
C33 a_888_406# VNB 0.59258f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtp_1 VNB VPB VPWR VGND Q GATE RESET_B D
X0 Q.t1 a_817_48.t3 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2309 ps=1.55 w=1.12 l=0.15
X1 a_1045_74# a_643_74.t4 a_817_48.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VGND.t2 a_216_424.t2 a_363_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1277 pd=1.1 as=0.32225 ps=2.64 w=0.74 l=0.15
X3 a_769_74.t0 a_216_424.t3 a_643_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.14535 ps=1.12 w=0.42 l=0.15
X4 a_643_74.t3 a_363_74.t2 a_565_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.14535 pd=1.12 as=0.0768 ps=0.88 w=0.64 l=0.15
X5 Q.t0 a_817_48.t4 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1332 ps=1.1 w=0.74 l=0.15
X6 VPWR.t2 a_216_424.t4 a_363_74.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2078 pd=1.43 as=0.2478 ps=2.27 w=0.84 l=0.15
X7 VGND.t0 D.t0 a_27_424.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1467 pd=1.175 as=0.15675 ps=1.67 w=0.55 l=0.15
X8 a_216_424.t1 GATE.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1467 ps=1.175 w=0.74 l=0.15
X9 VGND RESET_B a_1045_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X10 VPWR.t3 D.t1 a_27_424.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X11 VPWR.t1 RESET_B.t0 a_817_48.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2309 pd=1.55 as=0.175 ps=1.35 w=1 l=0.15
X12 VGND.t4 a_817_48.t5 a_769_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 a_643_74.t0 a_216_424.t5 a_568_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X14 a_565_74.t1 a_27_424.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1277 ps=1.1 w=0.64 l=0.15
X15 a_568_392.t0 a_27_424.t3 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2078 ps=1.43 w=1 l=0.15
X16 a_759_508.t0 a_363_74.t3 a_643_74.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.10605 pd=0.925 as=0.1664 ps=1.385 w=0.42 l=0.15
X17 a_817_48.t2 a_643_74.t5 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.20495 ps=1.61 w=1 l=0.15
X18 a_216_424.t0 GATE.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.43935 pd=2.87 as=0.147 ps=1.19 w=0.84 l=0.15
X19 VPWR.t5 a_817_48.t6 a_759_508.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.20495 pd=1.61 as=0.10605 ps=0.925 w=0.42 l=0.15
R0 a_817_48.n2 a_817_48.t5 518.953
R1 a_817_48.n0 a_817_48.t3 285.719
R2 a_817_48.n1 a_817_48.n0 223.459
R3 a_817_48.n4 a_817_48.n3 199.167
R4 a_817_48.n3 a_817_48.n2 178.351
R5 a_817_48.n0 a_817_48.t4 178.34
R6 a_817_48.n1 a_817_48.t1 164.294
R7 a_817_48.n2 a_817_48.t6 138.565
R8 a_817_48.n3 a_817_48.n1 64.2154
R9 a_817_48.n4 a_817_48.t2 39.4005
R10 a_817_48.t0 a_817_48.n4 29.5505
R11 VPWR.n16 VPWR.n4 611.27
R12 VPWR.n22 VPWR.n1 604.976
R13 VPWR.n9 VPWR.n8 585
R14 VPWR.n7 VPWR.n6 227.905
R15 VPWR.n8 VPWR.t5 143.06
R16 VPWR.n8 VPWR.t7 106.334
R17 VPWR.n4 VPWR.t2 60.9767
R18 VPWR.n1 VPWR.t3 46.9053
R19 VPWR.n6 VPWR.t4 43.3107
R20 VPWR.n6 VPWR.t1 39.4005
R21 VPWR.n20 VPWR.n2 36.1417
R22 VPWR.n21 VPWR.n20 36.1417
R23 VPWR.n14 VPWR.n5 36.1417
R24 VPWR.n15 VPWR.n14 36.1417
R25 VPWR.n1 VPWR.t0 35.1791
R26 VPWR.n4 VPWR.t6 33.1589
R27 VPWR.n16 VPWR.n15 31.2476
R28 VPWR.n10 VPWR.n5 28.8214
R29 VPWR.n22 VPWR.n21 19.2005
R30 VPWR.n16 VPWR.n2 12.8005
R31 VPWR.n9 VPWR.n7 11.9372
R32 VPWR.n11 VPWR.n10 9.3005
R33 VPWR.n12 VPWR.n5 9.3005
R34 VPWR.n14 VPWR.n13 9.3005
R35 VPWR.n15 VPWR.n3 9.3005
R36 VPWR.n17 VPWR.n16 9.3005
R37 VPWR.n18 VPWR.n2 9.3005
R38 VPWR.n20 VPWR.n19 9.3005
R39 VPWR.n21 VPWR.n0 9.3005
R40 VPWR.n23 VPWR.n22 7.43488
R41 VPWR.n10 VPWR.n9 3.26325
R42 VPWR.n11 VPWR.n7 0.535194
R43 VPWR VPWR.n23 0.160103
R44 VPWR.n23 VPWR.n0 0.1477
R45 VPWR.n12 VPWR.n11 0.122949
R46 VPWR.n13 VPWR.n12 0.122949
R47 VPWR.n13 VPWR.n3 0.122949
R48 VPWR.n17 VPWR.n3 0.122949
R49 VPWR.n18 VPWR.n17 0.122949
R50 VPWR.n19 VPWR.n18 0.122949
R51 VPWR.n19 VPWR.n0 0.122949
R52 Q.n0 Q.t1 312.998
R53 Q.n0 Q.t0 207.703
R54 Q Q.n0 4.90517
R55 VPB VPB.n0 1483.74
R56 VPB.t5 VPB.t8 388.173
R57 VPB.t4 VPB.t5 334.543
R58 VPB.t1 VPB.t6 296.238
R59 VPB.t3 VPB.t4 273.253
R60 VPB.t8 VPB.t1 255.376
R61 VPB.n0 VPB.t3 143.012
R62 VPB.n0 VPB 133.523
R63 VPB.n0 VPB.t0 33.7646
R64 VPB.t0 VPB.t7 24.5562
R65 VPB.t7 VPB.t2 24.5562
R66 a_643_74.n3 a_643_74.n2 640.471
R67 a_643_74.n2 a_643_74.n0 251.636
R68 a_643_74.n1 a_643_74.t4 248.775
R69 a_643_74.n2 a_643_74.n1 242.31
R70 a_643_74.n1 a_643_74.t5 221.731
R71 a_643_74.n3 a_643_74.t1 110.227
R72 a_643_74.n0 a_643_74.t2 80.0005
R73 a_643_74.n0 a_643_74.t3 37.5005
R74 a_643_74.t0 a_643_74.n3 30.9107
R75 VNB.t1 VNB.t2 2436.75
R76 VNB.t6 VNB.t5 2286.61
R77 VNB.t5 VNB.t7 2078.74
R78 VNB.t8 VNB.t3 1455.12
R79 VNB VNB.t0 1385.83
R80 VNB.t0 VNB.t1 1351.18
R81 VNB.t2 VNB.t4 1177.95
R82 VNB.t3 VNB.t6 900.788
R83 VNB.t4 VNB.t8 900.788
R84 a_216_424.t0 a_216_424.n3 785.99
R85 a_216_424.n0 a_216_424.t5 439.224
R86 a_216_424.n1 a_216_424.n0 420.964
R87 a_216_424.n3 a_216_424.n2 261.253
R88 a_216_424.n2 a_216_424.t4 251.809
R89 a_216_424.n2 a_216_424.t2 244.579
R90 a_216_424.n0 a_216_424.t3 227.143
R91 a_216_424.n1 a_216_424.t1 141.708
R92 a_216_424.n3 a_216_424.n1 36.9012
R93 a_363_74.t1 a_363_74.n1 822.346
R94 a_363_74.n0 a_363_74.t3 481.45
R95 a_363_74.n1 a_363_74.t0 358.361
R96 a_363_74.n0 a_363_74.t2 314.274
R97 a_363_74.n1 a_363_74.n0 74.617
R98 VGND.n7 VGND.t5 253.607
R99 VGND.n6 VGND.t4 247.498
R100 VGND.n4 VGND.n3 202.123
R101 VGND.n1 VGND.n0 137.833
R102 VGND.n0 VGND.t0 63.6442
R103 VGND.n10 VGND.n9 36.1417
R104 VGND.n11 VGND.n10 36.1417
R105 VGND.n16 VGND.n15 36.1417
R106 VGND.n17 VGND.n16 36.1417
R107 VGND.n3 VGND.t3 35.6255
R108 VGND.n11 VGND.n4 33.1299
R109 VGND.n3 VGND.t2 28.2861
R110 VGND.n19 VGND.n1 26.5273
R111 VGND.n0 VGND.t1 21.9497
R112 VGND.n17 VGND.n1 17.3181
R113 VGND.n15 VGND.n4 10.1652
R114 VGND.n9 VGND.n6 9.78874
R115 VGND.n18 VGND.n17 9.3005
R116 VGND.n16 VGND.n2 9.3005
R117 VGND.n15 VGND.n14 9.3005
R118 VGND.n13 VGND.n4 9.3005
R119 VGND.n12 VGND.n11 9.3005
R120 VGND.n10 VGND.n5 9.3005
R121 VGND.n9 VGND.n8 9.3005
R122 VGND.n7 VGND.n6 9.01336
R123 VGND.n8 VGND.n7 0.291092
R124 VGND VGND.n19 0.163644
R125 VGND.n19 VGND.n18 0.144205
R126 VGND.n8 VGND.n5 0.122949
R127 VGND.n12 VGND.n5 0.122949
R128 VGND.n13 VGND.n12 0.122949
R129 VGND.n14 VGND.n13 0.122949
R130 VGND.n14 VGND.n2 0.122949
R131 VGND.n18 VGND.n2 0.122949
R132 a_769_74.t0 a_769_74.t1 68.5719
R133 a_565_74.t0 a_565_74.t1 45.0005
R134 D.n0 D.t1 290.69
R135 D.n0 D.t0 174.624
R136 D D.n0 155.067
R137 a_27_424.t1 a_27_424.n1 780.348
R138 a_27_424.t1 a_27_424.n2 768.644
R139 a_27_424.n1 a_27_424.n0 345.507
R140 a_27_424.n2 a_27_424.t0 299.729
R141 a_27_424.n0 a_27_424.t2 274.74
R142 a_27_424.n0 a_27_424.t3 231.629
R143 a_27_424.n2 a_27_424.n1 4.4805
R144 GATE.n0 GATE.t1 253.073
R145 GATE.n0 GATE.t0 251.2
R146 GATE GATE.n0 153.262
R147 RESET_B.n1 RESET_B.t0 263.762
R148 RESET_B.n1 RESET_B.n0 220.113
R149 RESET_B RESET_B.n1 156.912
R150 a_568_392.t0 a_568_392.t1 53.1905
R151 a_759_508.t0 a_759_508.t1 236.869
C0 RESET_B VPWR 0.026217f
C1 GATE VGND 0.024621f
C2 D Q 1.81e-20
C3 a_1045_74# Q 5.03e-19
C4 RESET_B VGND 0.014929f
C5 VPWR VGND 0.107097f
C6 RESET_B Q 0.008506f
C7 VPWR Q 0.120803f
C8 VGND Q 0.097381f
C9 VPB D 0.0677f
C10 VPB GATE 0.059308f
C11 VPB RESET_B 0.045109f
C12 D GATE 0.050599f
C13 VPB VPWR 0.191313f
C14 VPB VGND 0.014989f
C15 D VPWR 0.012861f
C16 a_1045_74# VPWR 7.95e-19
C17 GATE VPWR 0.014758f
C18 VPB Q 0.015692f
C19 D VGND 0.008396f
C20 a_1045_74# VGND 0.008746f
C21 Q VNB 0.1184f
C22 VGND VNB 0.834558f
C23 VPWR VNB 0.632804f
C24 RESET_B VNB 0.103826f
C25 GATE VNB 0.123045f
C26 D VNB 0.192787f
C27 VPB VNB 1.55959f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtp_2 VNB VPB VPWR VGND D GATE RESET_B Q
X0 a_235_74.t1 GATE.t0 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X1 VPWR.t3 D.t0 a_27_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.23945 pd=1.6 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 a_646_74.t0 a_347_98.t2 a_568_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.160775 pd=1.18 as=0.0768 ps=0.88 w=0.64 l=0.15
X3 a_646_74.t2 a_235_74.t2 a_565_392.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X4 a_565_392.t0 a_27_392.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.243825 ps=1.595 w=1 l=0.15
X5 a_756_508.t1 a_347_98.t3 a_646_74.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.11235 pd=0.955 as=0.1664 ps=1.385 w=0.42 l=0.15
X6 Q.t0 a_832_55.t3 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.224 ps=1.52 w=1.12 l=0.15
X7 a_784_81.t1 a_235_74.t3 a_646_74.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.160775 ps=1.18 w=0.42 l=0.15
X8 VGND.t3 a_832_55.t4 Q.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1073 ps=1.03 w=0.74 l=0.15
X9 VPWR.t4 a_832_55.t5 a_756_508.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2303 pd=1.775 as=0.11235 ps=0.955 w=0.42 l=0.15
X10 VGND.t4 RESET_B.t0 a_1060_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.0888 ps=0.98 w=0.74 l=0.15
X11 VPWR.t7 a_235_74.t4 a_347_98.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.243825 pd=1.595 as=0.2478 ps=2.27 w=0.84 l=0.15
X12 a_1060_74.t1 a_646_74.t4 a_832_55.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 a_568_74.t0 a_27_392.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.19135 ps=1.49 w=0.64 l=0.15
X14 Q.t1 a_832_55.t6 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1628 ps=1.18 w=0.74 l=0.15
X15 VGND.t0 D.t1 a_27_392.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X16 VGND.t1 a_235_74.t5 a_347_98.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.19135 pd=1.49 as=0.2701 ps=2.21 w=0.74 l=0.15
X17 VGND.t7 a_832_55.t7 a_784_81.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X18 a_235_74.t0 GATE.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.23945 ps=1.6 w=0.84 l=0.15
X19 VPWR.t5 RESET_B.t1 a_832_55.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_832_55.t0 a_646_74.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2303 ps=1.775 w=1.12 l=0.15
R0 GATE.n0 GATE.t1 272.866
R1 GATE.n0 GATE.t0 178.34
R2 GATE GATE.n0 160.615
R3 VGND.n11 VGND.t7 248.856
R4 VGND.n7 VGND.t3 248.38
R5 VGND.n18 VGND.n17 243.073
R6 VGND.n26 VGND.n25 118.88
R7 VGND.n6 VGND.n5 116.109
R8 VGND.n25 VGND.t0 51.1752
R9 VGND.n17 VGND.t1 50.5955
R10 VGND.n5 VGND.t4 37.2978
R11 VGND.n10 VGND.n9 36.1417
R12 VGND.n15 VGND.n3 36.1417
R13 VGND.n16 VGND.n15 36.1417
R14 VGND.n19 VGND.n16 36.1417
R15 VGND.n23 VGND.n1 36.1417
R16 VGND.n24 VGND.n23 36.1417
R17 VGND.n5 VGND.t6 34.0546
R18 VGND.n25 VGND.t2 32.4566
R19 VGND.n11 VGND.n10 32.0005
R20 VGND.n17 VGND.t5 25.8859
R21 VGND.n9 VGND.n6 17.6946
R22 VGND.n26 VGND.n24 16.5652
R23 VGND.n11 VGND.n3 15.4358
R24 VGND.n18 VGND.n1 15.1848
R25 VGND.n24 VGND.n0 9.3005
R26 VGND.n23 VGND.n22 9.3005
R27 VGND.n21 VGND.n1 9.3005
R28 VGND.n20 VGND.n19 9.3005
R29 VGND.n16 VGND.n2 9.3005
R30 VGND.n15 VGND.n14 9.3005
R31 VGND.n13 VGND.n3 9.3005
R32 VGND.n12 VGND.n11 9.3005
R33 VGND.n10 VGND.n4 9.3005
R34 VGND.n9 VGND.n8 9.3005
R35 VGND.n27 VGND.n26 7.53404
R36 VGND.n7 VGND.n6 6.96039
R37 VGND.n19 VGND.n18 4.64364
R38 VGND.n8 VGND.n7 0.594857
R39 VGND VGND.n27 0.161409
R40 VGND.n27 VGND.n0 0.146411
R41 VGND.n8 VGND.n4 0.122949
R42 VGND.n12 VGND.n4 0.122949
R43 VGND.n13 VGND.n12 0.122949
R44 VGND.n14 VGND.n13 0.122949
R45 VGND.n14 VGND.n2 0.122949
R46 VGND.n20 VGND.n2 0.122949
R47 VGND.n21 VGND.n20 0.122949
R48 VGND.n22 VGND.n21 0.122949
R49 VGND.n22 VGND.n0 0.122949
R50 a_235_74.t0 a_235_74.n3 795.176
R51 a_235_74.n0 a_235_74.t2 456.293
R52 a_235_74.n1 a_235_74.n0 416.967
R53 a_235_74.n0 a_235_74.t3 231.361
R54 a_235_74.n3 a_235_74.n2 211.886
R55 a_235_74.n2 a_235_74.t4 195.21
R56 a_235_74.n2 a_235_74.t5 186.115
R57 a_235_74.n1 a_235_74.t1 131.46
R58 a_235_74.n3 a_235_74.n1 41.6969
R59 VNB.t1 VNB.t7 2482.94
R60 VNB.t10 VNB.t2 2286.61
R61 VNB.t6 VNB.t8 1593.7
R62 VNB.t4 VNB.t9 1362.73
R63 VNB.t7 VNB.t5 1362.73
R64 VNB.t0 VNB.t1 1339.63
R65 VNB VNB.t0 1201.05
R66 VNB.t9 VNB.t3 1016.27
R67 VNB.t2 VNB.t4 900.788
R68 VNB.t8 VNB.t10 900.788
R69 VNB.t5 VNB.t6 900.788
R70 D.n0 D.t1 218.828
R71 D.n0 D.t0 208.386
R72 D D.n0 160.922
R73 a_27_392.t1 a_27_392.n1 771.861
R74 a_27_392.t1 a_27_392.n2 761.966
R75 a_27_392.n1 a_27_392.n0 339.86
R76 a_27_392.n2 a_27_392.t0 305.399
R77 a_27_392.n0 a_27_392.t3 265.101
R78 a_27_392.n0 a_27_392.t2 239.661
R79 a_27_392.n2 a_27_392.n1 7.09239
R80 VPWR.n23 VPWR.n1 698.433
R81 VPWR.n16 VPWR.n15 676.107
R82 VPWR.n8 VPWR.n7 585
R83 VPWR.n6 VPWR.n5 227.294
R84 VPWR.n7 VPWR.t2 142.56
R85 VPWR.n7 VPWR.t4 140.714
R86 VPWR.n15 VPWR.t7 64.4945
R87 VPWR.n1 VPWR.t1 55.1136
R88 VPWR.n1 VPWR.t3 55.1136
R89 VPWR.n21 VPWR.n2 36.1417
R90 VPWR.n22 VPWR.n21 36.1417
R91 VPWR.n13 VPWR.n4 36.1417
R92 VPWR.n14 VPWR.n13 36.1417
R93 VPWR.n17 VPWR.n14 36.1417
R94 VPWR.n15 VPWR.t0 35.6631
R95 VPWR.n5 VPWR.t6 35.1791
R96 VPWR.n5 VPWR.t5 35.1791
R97 VPWR.n9 VPWR.n4 29.6998
R98 VPWR.n23 VPWR.n22 16.5652
R99 VPWR.n8 VPWR.n6 11.7597
R100 VPWR.n10 VPWR.n9 9.3005
R101 VPWR.n11 VPWR.n4 9.3005
R102 VPWR.n13 VPWR.n12 9.3005
R103 VPWR.n14 VPWR.n3 9.3005
R104 VPWR.n18 VPWR.n17 9.3005
R105 VPWR.n19 VPWR.n2 9.3005
R106 VPWR.n21 VPWR.n20 9.3005
R107 VPWR.n22 VPWR.n0 9.3005
R108 VPWR.n16 VPWR.n2 9.03579
R109 VPWR.n24 VPWR.n23 7.53404
R110 VPWR.n9 VPWR.n8 3.43057
R111 VPWR.n17 VPWR.n16 2.25932
R112 VPWR.n10 VPWR.n6 0.526721
R113 VPWR VPWR.n24 0.161409
R114 VPWR.n24 VPWR.n0 0.146411
R115 VPWR.n11 VPWR.n10 0.122949
R116 VPWR.n12 VPWR.n11 0.122949
R117 VPWR.n12 VPWR.n3 0.122949
R118 VPWR.n18 VPWR.n3 0.122949
R119 VPWR.n19 VPWR.n18 0.122949
R120 VPWR.n20 VPWR.n19 0.122949
R121 VPWR.n20 VPWR.n0 0.122949
R122 VPB.t1 VPB.t8 515.861
R123 VPB.t4 VPB.t2 411.156
R124 VPB.t7 VPB.t4 349.866
R125 VPB.t3 VPB.t1 316.668
R126 VPB.t8 VPB.t0 314.113
R127 VPB.t5 VPB.t6 280.914
R128 VPB.t9 VPB.t7 273.253
R129 VPB VPB.t3 257.93
R130 VPB.t2 VPB.t5 229.839
R131 VPB.t0 VPB.t9 214.517
R132 a_347_98.t0 a_347_98.n1 829.712
R133 a_347_98.n0 a_347_98.t3 492.317
R134 a_347_98.n0 a_347_98.t2 314.274
R135 a_347_98.n1 a_347_98.t1 269.252
R136 a_347_98.n1 a_347_98.n0 70.8349
R137 a_568_74.t0 a_568_74.t1 45.0005
R138 a_646_74.n3 a_646_74.n2 634.318
R139 a_646_74.n2 a_646_74.n1 304.053
R140 a_646_74.n2 a_646_74.n0 258.036
R141 a_646_74.n1 a_646_74.t5 226.809
R142 a_646_74.n1 a_646_74.t4 200.519
R143 a_646_74.n3 a_646_74.t1 110.227
R144 a_646_74.n0 a_646_74.t3 68.0406
R145 a_646_74.n0 a_646_74.t0 41.8163
R146 a_646_74.t2 a_646_74.n3 30.9107
R147 a_565_392.t0 a_565_392.t1 53.1905
R148 a_756_508.t0 a_756_508.t1 250.94
R149 a_832_55.n5 a_832_55.t7 461.945
R150 a_832_55.n1 a_832_55.n0 242.268
R151 a_832_55.n2 a_832_55.t3 241.657
R152 a_832_55.n7 a_832_55.n6 197.218
R153 a_832_55.n4 a_832_55.t1 194.888
R154 a_832_55.n6 a_832_55.n5 183.047
R155 a_832_55.n1 a_832_55.t4 179.947
R156 a_832_55.n2 a_832_55.t6 179.947
R157 a_832_55.n5 a_832_55.t5 138.441
R158 a_832_55.n4 a_832_55.n3 119.737
R159 a_832_55.n3 a_832_55.n1 35.5081
R160 a_832_55.n7 a_832_55.t2 26.3844
R161 a_832_55.t0 a_832_55.n7 26.3844
R162 a_832_55.n3 a_832_55.n2 22.038
R163 a_832_55.n6 a_832_55.n4 9.06891
R164 Q Q.t0 302.176
R165 Q Q.n0 128.53
R166 Q.n0 Q.t2 24.3248
R167 Q.n0 Q.t1 22.7032
R168 a_784_81.t0 a_784_81.t1 68.5719
R169 RESET_B.n0 RESET_B.t1 285.719
R170 RESET_B.n0 RESET_B.t0 178.34
R171 RESET_B RESET_B.n0 160.304
R172 a_1060_74.t0 a_1060_74.t1 38.9194
C0 VGND Q 0.169803f
C1 VPWR GATE 0.009115f
C2 D GATE 0.036621f
C3 RESET_B VPB 0.030201f
C4 RESET_B VPWR 0.020576f
C5 VGND VPB 0.016057f
C6 VGND VPWR 0.118297f
C7 Q VPB 0.009104f
C8 VGND D 0.01281f
C9 Q VPWR 0.221829f
C10 Q D 5.74e-21
C11 VGND GATE 0.01918f
C12 VPB VPWR 0.213682f
C13 RESET_B VGND 0.034341f
C14 VPB D 0.052031f
C15 RESET_B Q 0.003671f
C16 VPWR D 0.008441f
C17 VPB GATE 0.04628f
C18 Q VNB 0.063704f
C19 VGND VNB 0.899701f
C20 RESET_B VNB 0.10724f
C21 GATE VNB 0.121477f
C22 D VNB 0.159248f
C23 VPWR VNB 0.699893f
C24 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtp_4 VNB VPB VPWR VGND D GATE RESET_B Q
X0 VPWR RESET_B a_797_48# VPB sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X1 VGND.t9 a_797_48# Q.t7 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_755_74.t1 a_240_394.t2 a_640_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.12775 ps=1.065 w=0.42 l=0.15
X3 VGND.t0 a_240_394.t3 a_364_120.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.149425 pd=1.335 as=0.2294 ps=2.1 w=0.74 l=0.15
X4 a_797_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.147 ps=1.19 w=0.84 l=0.15
X5 VGND.t10 a_797_48# a_755_74.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_938_74.t1 RESET_B.t0 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X7 a_640_74.t0 a_364_120.t2 a_559_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12775 pd=1.065 as=0.0816 ps=0.895 w=0.64 l=0.15
X8 a_938_74.t3 a_640_74.t4 a_797_48# VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0912 ps=0.925 w=0.64 l=0.15
X9 VGND.t8 a_797_48# Q.t6 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_559_74.t0 a_27_126.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0816 pd=0.895 as=0.149425 ps=1.335 w=0.64 l=0.15
X11 a_240_394.t0 GATE.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.294 pd=2.38 as=0.22785 ps=1.52 w=0.84 l=0.15
X12 VPWR.t0 a_240_394.t4 a_364_120.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1903 pd=1.395 as=0.2478 ps=2.27 w=0.84 l=0.15
X13 a_240_394.t1 GATE.t1 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.194525 ps=1.285 w=0.74 l=0.15
X14 a_797_48# a_640_74.t5 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2093 ps=1.735 w=0.84 l=0.15
X15 Q.t3 a_797_48# VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2072 pd=1.49 as=0.196 ps=1.47 w=1.12 l=0.15
X16 VGND.t4 RESET_B.t1 a_938_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X17 a_640_74.t2 a_240_394.t5 a_562_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.12 ps=1.24 w=1 l=0.15
X18 VPWR.t4 D.t0 a_27_126.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.22785 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X19 Q.t5 a_797_48# VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_562_392.t0 a_27_126.t3 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.1903 ps=1.395 w=1 l=0.15
X21 a_747_508.t0 a_364_120.t3 a_640_74.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1664 ps=1.385 w=0.42 l=0.15
X22 VPWR.t5 a_797_48# a_747_508.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2093 pd=1.735 as=0.09975 ps=0.895 w=0.42 l=0.15
X23 VPWR.t7 a_797_48# Q.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_797_48# a_640_74.t6 a_938_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0912 pd=0.925 as=0.1824 ps=1.85 w=0.64 l=0.15
X25 Q.t4 a_797_48# VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X26 Q.t1 a_797_48# VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.203 ps=1.505 w=1.12 l=0.15
X27 VGND.t3 D.t1 a_27_126.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.194525 pd=1.285 as=0.15675 ps=1.67 w=0.55 l=0.15
X28 VPWR.t9 a_797_48# Q.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.364 pd=2.89 as=0.2072 ps=1.49 w=1.12 l=0.15
R0 RESET_B.n6 RESET_B.n1 259.478
R1 RESET_B.n3 RESET_B.n2 243.411
R2 RESET_B.n7 RESET_B.n6 152
R3 RESET_B.n4 RESET_B.n0 152
R4 RESET_B.n3 RESET_B.t1 150.589
R5 RESET_B.n5 RESET_B.t0 138.173
R6 RESET_B.n5 RESET_B.n4 43.0884
R7 RESET_B.n7 RESET_B.n0 13.1884
R8 RESET_B.n4 RESET_B.n3 7.30353
R9 RESET_B.n6 RESET_B.n5 6.57323
R10 RESET_B.n0 RESET_B 5.23686
R11 RESET_B RESET_B.n7 0.194439
R12 VPWR.n35 VPWR.n1 646.804
R13 VPWR.n29 VPWR.n4 608.593
R14 VPWR.n22 VPWR.n21 588.519
R15 VPWR.n21 VPWR.t1 408.894
R16 VPWR.n11 VPWR.t9 356
R17 VPWR.n10 VPWR.n9 318.089
R18 VPWR.n14 VPWR.t6 262.769
R19 VPWR.n21 VPWR.t5 121.953
R20 VPWR.n4 VPWR.t0 56.2862
R21 VPWR.n1 VPWR.t2 55.1136
R22 VPWR.n1 VPWR.t4 55.1136
R23 VPWR.n33 VPWR.n2 36.1417
R24 VPWR.n34 VPWR.n33 36.1417
R25 VPWR.n27 VPWR.n5 36.1417
R26 VPWR.n28 VPWR.n27 36.1417
R27 VPWR.n20 VPWR.n19 36.1417
R28 VPWR.n15 VPWR.n7 36.1417
R29 VPWR.n9 VPWR.t7 35.1791
R30 VPWR.n14 VPWR.n13 35.0123
R31 VPWR.n29 VPWR.n28 34.2593
R32 VPWR.n4 VPWR.t3 31.1891
R33 VPWR.n9 VPWR.t8 26.3844
R34 VPWR.n23 VPWR.n5 23.5508
R35 VPWR.n35 VPWR.n34 16.5652
R36 VPWR.n22 VPWR.n20 14.8502
R37 VPWR.n29 VPWR.n2 13.177
R38 VPWR.n15 VPWR.n14 12.424
R39 VPWR.n13 VPWR.n10 11.6711
R40 VPWR.n19 VPWR.n7 11.2946
R41 VPWR.n13 VPWR.n12 9.3005
R42 VPWR.n14 VPWR.n8 9.3005
R43 VPWR.n16 VPWR.n15 9.3005
R44 VPWR.n17 VPWR.n7 9.3005
R45 VPWR.n19 VPWR.n18 9.3005
R46 VPWR.n20 VPWR.n6 9.3005
R47 VPWR.n24 VPWR.n23 9.3005
R48 VPWR.n25 VPWR.n5 9.3005
R49 VPWR.n27 VPWR.n26 9.3005
R50 VPWR.n28 VPWR.n3 9.3005
R51 VPWR.n30 VPWR.n29 9.3005
R52 VPWR.n31 VPWR.n2 9.3005
R53 VPWR.n33 VPWR.n32 9.3005
R54 VPWR.n34 VPWR.n0 9.3005
R55 VPWR.n36 VPWR.n35 7.53404
R56 VPWR.n11 VPWR.n10 7.14239
R57 VPWR.n23 VPWR.n22 1.08808
R58 VPWR.n12 VPWR.n11 0.61555
R59 VPWR VPWR.n36 0.161409
R60 VPWR.n36 VPWR.n0 0.146411
R61 VPWR.n12 VPWR.n8 0.122949
R62 VPWR.n16 VPWR.n8 0.122949
R63 VPWR.n17 VPWR.n16 0.122949
R64 VPWR.n18 VPWR.n17 0.122949
R65 VPWR.n18 VPWR.n6 0.122949
R66 VPWR.n24 VPWR.n6 0.122949
R67 VPWR.n25 VPWR.n24 0.122949
R68 VPWR.n26 VPWR.n25 0.122949
R69 VPWR.n26 VPWR.n3 0.122949
R70 VPWR.n30 VPWR.n3 0.122949
R71 VPWR.n31 VPWR.n30 0.122949
R72 VPWR.n32 VPWR.n31 0.122949
R73 VPWR.n32 VPWR.n0 0.122949
R74 VPB VPB.n0 1465.86
R75 VPB.t2 VPB.t7 1013.84
R76 VPB.t0 VPB.t3 581.466
R77 VPB.t9 VPB.t2 390.726
R78 VPB.t3 VPB.t5 338.507
R79 VPB.t11 VPB.t9 319.221
R80 VPB.t4 VPB.t0 297.558
R81 VPB.t5 VPB 275.719
R82 VPB.t1 VPB.t11 273.253
R83 VPB.t10 VPB.t6 265.591
R84 VPB.t8 VPB.t10 255.376
R85 VPB.t7 VPB.t8 229.839
R86 VPB.n0 VPB.t1 130.243
R87 VPB.n0 VPB.t4 73.7074
R88 Q.n2 Q.n0 261.986
R89 Q.n2 Q.n1 207.6
R90 Q.n5 Q.n4 138.7
R91 Q.n5 Q.n3 98.0421
R92 Q Q.n2 42.5744
R93 Q.n1 Q.t3 35.1791
R94 Q.n1 Q.t0 29.9023
R95 Q Q.n5 28.5167
R96 Q.n0 Q.t2 26.3844
R97 Q.n0 Q.t1 26.3844
R98 Q.n3 Q.t6 22.7032
R99 Q.n3 Q.t5 22.7032
R100 Q.n4 Q.t7 22.7032
R101 Q.n4 Q.t4 22.7032
R102 VGND.n10 VGND.t8 300.51
R103 VGND.n20 VGND.t10 254.696
R104 VGND.n28 VGND.n27 240.149
R105 VGND.n35 VGND.n34 215.061
R106 VGND.n9 VGND.n8 205.559
R107 VGND.n6 VGND.n5 204.976
R108 VGND.n13 VGND.t6 169.403
R109 VGND.n34 VGND.t3 60.0005
R110 VGND.n27 VGND.t0 48.0756
R111 VGND.n34 VGND.t2 45.745
R112 VGND.n19 VGND.n18 36.1417
R113 VGND.n21 VGND.n19 36.1417
R114 VGND.n25 VGND.n3 36.1417
R115 VGND.n26 VGND.n25 36.1417
R116 VGND.n32 VGND.n1 36.1417
R117 VGND.n33 VGND.n32 36.1417
R118 VGND.n14 VGND.n13 35.7652
R119 VGND.n28 VGND.n26 34.2593
R120 VGND.n18 VGND.n6 33.5064
R121 VGND.n12 VGND.n9 28.2358
R122 VGND.n5 VGND.t5 26.2505
R123 VGND.n5 VGND.t4 26.2505
R124 VGND.n8 VGND.t7 22.7032
R125 VGND.n8 VGND.t9 22.7032
R126 VGND.n27 VGND.t1 19.8358
R127 VGND.n13 VGND.n12 16.9417
R128 VGND.n35 VGND.n33 14.3064
R129 VGND.n14 VGND.n6 13.9299
R130 VGND.n28 VGND.n1 13.177
R131 VGND.n33 VGND.n0 9.3005
R132 VGND.n32 VGND.n31 9.3005
R133 VGND.n30 VGND.n1 9.3005
R134 VGND.n29 VGND.n28 9.3005
R135 VGND.n26 VGND.n2 9.3005
R136 VGND.n25 VGND.n24 9.3005
R137 VGND.n23 VGND.n3 9.3005
R138 VGND.n22 VGND.n21 9.3005
R139 VGND.n19 VGND.n4 9.3005
R140 VGND.n18 VGND.n17 9.3005
R141 VGND.n16 VGND.n6 9.3005
R142 VGND.n15 VGND.n14 9.3005
R143 VGND.n13 VGND.n7 9.3005
R144 VGND.n12 VGND.n11 9.3005
R145 VGND.n21 VGND.n20 9.03579
R146 VGND.n20 VGND.n3 8.28285
R147 VGND.n36 VGND.n35 7.61102
R148 VGND.n10 VGND.n9 6.26985
R149 VGND.n11 VGND.n10 0.733933
R150 VGND VGND.n36 0.162422
R151 VGND.n36 VGND.n0 0.145411
R152 VGND.n11 VGND.n7 0.122949
R153 VGND.n15 VGND.n7 0.122949
R154 VGND.n16 VGND.n15 0.122949
R155 VGND.n17 VGND.n16 0.122949
R156 VGND.n17 VGND.n4 0.122949
R157 VGND.n22 VGND.n4 0.122949
R158 VGND.n23 VGND.n22 0.122949
R159 VGND.n24 VGND.n23 0.122949
R160 VGND.n24 VGND.n2 0.122949
R161 VGND.n29 VGND.n2 0.122949
R162 VGND.n30 VGND.n29 0.122949
R163 VGND.n31 VGND.n30 0.122949
R164 VGND.n31 VGND.n0 0.122949
R165 VNB.t5 VNB.t1 2344.36
R166 VNB.t9 VNB.t10 2286.61
R167 VNB.t13 VNB.t4 2286.61
R168 VNB.t6 VNB.t5 1605.25
R169 VNB.t7 VNB.t0 1328.08
R170 VNB.t1 VNB.t2 1189.5
R171 VNB VNB.t6 1143.31
R172 VNB.t4 VNB.t3 1004.72
R173 VNB.t11 VNB.t12 993.177
R174 VNB.t14 VNB.t11 993.177
R175 VNB.t10 VNB.t14 993.177
R176 VNB.t8 VNB.t9 993.177
R177 VNB.t3 VNB.t8 993.177
R178 VNB.t2 VNB.t7 935.433
R179 VNB.t0 VNB.t13 831.496
R180 a_240_394.t0 a_240_394.n3 766.091
R181 a_240_394.n0 a_240_394.t5 431.276
R182 a_240_394.n1 a_240_394.n0 421.774
R183 a_240_394.n0 a_240_394.t2 222.41
R184 a_240_394.n3 a_240_394.n2 218.458
R185 a_240_394.n2 a_240_394.t4 187.178
R186 a_240_394.n2 a_240_394.t3 156.431
R187 a_240_394.n1 a_240_394.t1 140.589
R188 a_240_394.n3 a_240_394.n1 31.9178
R189 a_640_74.n6 a_640_74.n5 647.131
R190 a_640_74.n5 a_640_74.n0 254.44
R191 a_640_74.n2 a_640_74.n1 250.105
R192 a_640_74.n5 a_640_74.n4 249.293
R193 a_640_74.n2 a_640_74.t4 224.131
R194 a_640_74.n3 a_640_74.t6 220.688
R195 a_640_74.n4 a_640_74.t5 200.757
R196 a_640_74.n6 a_640_74.t3 110.227
R197 a_640_74.n3 a_640_74.n2 86.7605
R198 a_640_74.n0 a_640_74.t1 72.3671
R199 a_640_74.n0 a_640_74.t0 31.876
R200 a_640_74.t2 a_640_74.n6 30.9107
R201 a_640_74.n4 a_640_74.n3 10.3291
R202 a_755_74.t0 a_755_74.t1 60.0005
R203 a_364_120.t0 a_364_120.n1 834.534
R204 a_364_120.n0 a_364_120.t3 480.164
R205 a_364_120.n0 a_364_120.t2 314.274
R206 a_364_120.n1 a_364_120.t1 285.651
R207 a_364_120.n1 a_364_120.n0 63.228
R208 a_938_74.n1 a_938_74.t2 194.186
R209 a_938_74.t1 a_938_74.n1 190.827
R210 a_938_74.n1 a_938_74.n0 88.1117
R211 a_938_74.n0 a_938_74.t0 26.2505
R212 a_938_74.n0 a_938_74.t3 26.2505
R213 a_559_74.t0 a_559_74.t1 47.813
R214 a_27_126.t0 a_27_126.n1 774.963
R215 a_27_126.t0 a_27_126.n2 768.644
R216 a_27_126.n1 a_27_126.n0 332.084
R217 a_27_126.n2 a_27_126.t1 304.567
R218 a_27_126.n0 a_27_126.t2 274.74
R219 a_27_126.n0 a_27_126.t3 231.629
R220 a_27_126.n2 a_27_126.n1 5.88158
R221 GATE.n0 GATE.t1 229.754
R222 GATE.n0 GATE.t0 213.954
R223 GATE GATE.n0 153.94
R224 a_562_392.t0 a_562_392.t1 47.2805
R225 D.n0 D.t0 211.062
R226 D.n0 D.t1 196.335
R227 D D.n0 160.922
R228 a_747_508.t0 a_747_508.t1 222.798
C0 VPB GATE 0.049089f
C1 VPWR D 0.009582f
C2 a_797_48# VPB 0.29693f
C3 VPB RESET_B 0.067465f
C4 VPWR GATE 0.010191f
C5 D GATE 0.032124f
C6 a_797_48# VPWR 0.476535f
C7 a_797_48# D 6.84e-22
C8 VPWR RESET_B 0.029339f
C9 VPB VGND 0.018514f
C10 a_797_48# GATE 5.06e-20
C11 VPWR VGND 0.149098f
C12 VPB Q 0.018087f
C13 D VGND 0.011143f
C14 a_797_48# RESET_B 0.170952f
C15 VPWR Q 0.439694f
C16 GATE VGND 0.017585f
C17 D Q 2.15e-21
C18 a_797_48# VGND 0.135312f
C19 GATE Q 7.26e-21
C20 RESET_B VGND 0.03138f
C21 a_797_48# Q 0.397207f
C22 RESET_B Q 0.00315f
C23 VGND Q 0.29289f
C24 VPB VPWR 0.291255f
C25 VPB D 0.052584f
C26 Q VNB 0.073652f
C27 VGND VNB 1.12092f
C28 RESET_B VNB 0.231609f
C29 GATE VNB 0.115136f
C30 D VNB 0.153338f
C31 VPWR VNB 0.868612f
C32 VPB VNB 2.10038f
C33 a_797_48# VNB 0.643964f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxbn_1 VNB VPB VPWR VGND D Q_N Q GATE_N
X0 a_863_294.t0 a_653_79.t4 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.2225 ps=1.695 w=1.12 l=0.15
X1 Q_N.t0 a_1347_424# VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3136 ps=2.8 w=1.12 l=0.15
X2 VGND.t7 a_232_82.t2 a_343_80.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.180625 pd=1.39 as=0.3182 ps=2.34 w=0.74 l=0.15
X3 a_232_82.t0 GATE_N.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.147 ps=1.19 w=0.84 l=0.15
X4 VPWR.t0 a_232_82.t3 a_343_80.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1903 pd=1.395 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_863_294.t1 a_653_79.t5 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2183 pd=2.07 as=0.139825 ps=1.16 w=0.74 l=0.15
X6 a_653_79.t0 a_232_82.t4 a_575_79.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.20495 pd=1.485 as=0.0768 ps=0.88 w=0.64 l=0.15
X7 a_232_82.t1 GATE_N.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.189025 ps=1.41 w=0.74 l=0.15
X8 VGND.t4 a_863_294.t2 a_852_123.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.139825 pd=1.16 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 a_653_79.t3 a_343_80.t2 a_571_392.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.20285 pd=1.6 as=0.135 ps=1.27 w=1 l=0.15
X10 a_571_392.t0 a_27_120.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.1903 ps=1.395 w=1 l=0.15
X11 a_852_123.t1 a_343_80.t3 a_653_79.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.20495 ps=1.485 w=0.42 l=0.15
X12 VPWR.t4 D.t0 a_27_120.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.294 ps=2.38 w=0.84 l=0.15
X13 VGND.t3 a_863_294.t3 Q.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.12275 pd=1.1 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 Q_N.t1 a_1347_424# VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 a_805_392.t1 a_232_82.t5 a_653_79.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.07035 pd=0.755 as=0.20285 ps=1.6 w=0.42 l=0.15
X16 a_575_79.t0 a_27_120.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.180625 ps=1.39 w=0.64 l=0.15
X17 VPWR.t6 a_863_294.t4 a_805_392.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2225 pd=1.695 as=0.07035 ps=0.755 w=0.42 l=0.15
X18 VGND.t2 D.t1 a_27_120.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.189025 pd=1.41 as=0.15675 ps=1.67 w=0.55 l=0.15
X19 VPWR.t7 a_863_294.t5 Q.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.3136 ps=2.8 w=1.12 l=0.15
R0 a_653_79.n5 a_653_79.n4 643.467
R1 a_653_79.n0 a_653_79.t4 262.288
R2 a_653_79.n1 a_653_79.n0 219.114
R3 a_653_79.n4 a_653_79.n3 187.087
R4 a_653_79.n2 a_653_79.n1 185
R5 a_653_79.n0 a_653_79.t5 176.333
R6 a_653_79.n5 a_653_79.t1 161.821
R7 a_653_79.n6 a_653_79.t3 156.113
R8 a_653_79.n3 a_653_79.n2 132.857
R9 a_653_79.t3 a_653_79.n5 88.7387
R10 a_653_79.n3 a_653_79.t0 56.2951
R11 a_653_79.n2 a_653_79.t2 40.0005
R12 a_653_79.n4 a_653_79.n1 8.34833
R13 VPWR.n21 VPWR.n4 614.664
R14 VPWR.n9 VPWR.t7 358.2
R15 VPWR.n27 VPWR.n1 316.399
R16 VPWR.n15 VPWR.n7 289.678
R17 VPWR.n10 VPWR.t5 265.038
R18 VPWR.n7 VPWR.t6 153.448
R19 VPWR.n7 VPWR.t3 68.9444
R20 VPWR.n4 VPWR.t0 56.2862
R21 VPWR.n1 VPWR.t1 46.9053
R22 VPWR.n25 VPWR.n2 36.1417
R23 VPWR.n26 VPWR.n25 36.1417
R24 VPWR.n19 VPWR.n5 36.1417
R25 VPWR.n20 VPWR.n19 36.1417
R26 VPWR.n13 VPWR.n8 36.1417
R27 VPWR.n14 VPWR.n13 36.1417
R28 VPWR.n1 VPWR.t4 35.1791
R29 VPWR.n4 VPWR.t2 31.1891
R30 VPWR.n21 VPWR.n20 30.8711
R31 VPWR.n15 VPWR.n5 30.1181
R32 VPWR.n9 VPWR.n8 22.5887
R33 VPWR.n21 VPWR.n2 16.5652
R34 VPWR.n27 VPWR.n26 10.1652
R35 VPWR.n11 VPWR.n8 9.3005
R36 VPWR.n13 VPWR.n12 9.3005
R37 VPWR.n14 VPWR.n6 9.3005
R38 VPWR.n16 VPWR.n15 9.3005
R39 VPWR.n17 VPWR.n5 9.3005
R40 VPWR.n19 VPWR.n18 9.3005
R41 VPWR.n20 VPWR.n3 9.3005
R42 VPWR.n22 VPWR.n21 9.3005
R43 VPWR.n23 VPWR.n2 9.3005
R44 VPWR.n25 VPWR.n24 9.3005
R45 VPWR.n26 VPWR.n0 9.3005
R46 VPWR.n28 VPWR.n27 8.8332
R47 VPWR.n10 VPWR.n9 7.10322
R48 VPWR.n15 VPWR.n14 1.50638
R49 VPWR.n11 VPWR.n10 0.497626
R50 VPWR VPWR.n28 0.163644
R51 VPWR.n28 VPWR.n0 0.144205
R52 VPWR.n12 VPWR.n11 0.122949
R53 VPWR.n12 VPWR.n6 0.122949
R54 VPWR.n16 VPWR.n6 0.122949
R55 VPWR.n17 VPWR.n16 0.122949
R56 VPWR.n18 VPWR.n17 0.122949
R57 VPWR.n18 VPWR.n3 0.122949
R58 VPWR.n22 VPWR.n3 0.122949
R59 VPWR.n23 VPWR.n22 0.122949
R60 VPWR.n24 VPWR.n23 0.122949
R61 VPWR.n24 VPWR.n0 0.122949
R62 a_863_294.n3 a_863_294.n1 278.221
R63 a_863_294.n5 a_863_294.t5 247.131
R64 a_863_294.t0 a_863_294.n7 233.619
R65 a_863_294.n0 a_863_294.t2 231
R66 a_863_294.n6 a_863_294.n5 226.944
R67 a_863_294.n7 a_863_294.n0 201.888
R68 a_863_294.n6 a_863_294.t1 151.478
R69 a_863_294.n4 a_863_294.t3 142.994
R70 a_863_294.n0 a_863_294.t4 138.082
R71 a_863_294.n3 a_863_294.n2 90.1093
R72 a_863_294.n4 a_863_294.n3 56.9113
R73 a_863_294.n7 a_863_294.n6 17.5158
R74 a_863_294.n5 a_863_294.n4 1.69801
R75 VPB.t4 VPB.t8 766.13
R76 VPB.t2 VPB.t0 541.399
R77 VPB.t6 VPB.t4 508.2
R78 VPB.t9 VPB.t1 383.065
R79 VPB.t5 VPB.t6 370.296
R80 VPB VPB.t7 344.759
R81 VPB.t0 VPB.t3 278.361
R82 VPB.t7 VPB.t2 255.376
R83 VPB.t1 VPB.t5 247.715
R84 VPB.t3 VPB.t9 214.517
R85 Q_N.n3 Q_N 589.777
R86 Q_N.n3 Q_N.n0 585
R87 Q_N.n4 Q_N.n3 585
R88 Q_N.n2 Q_N.t1 281.43
R89 Q_N.t1 Q_N.n1 281.43
R90 Q_N.n3 Q_N.t0 26.3844
R91 Q_N Q_N.n4 12.8005
R92 Q_N.n1 Q_N 12.4184
R93 Q_N Q_N.n0 11.0811
R94 Q_N Q_N.n2 9.36169
R95 Q_N.n2 Q_N 4.77662
R96 Q_N Q_N.n0 3.05722
R97 Q_N.n1 Q_N 1.7199
R98 Q_N.n4 Q_N 1.33781
R99 a_232_82.n2 a_232_82.t4 409.471
R100 a_232_82.n3 a_232_82.n2 387.693
R101 a_232_82.t0 a_232_82.n3 340.265
R102 a_232_82.n0 a_232_82.t3 309.017
R103 a_232_82.n1 a_232_82.t1 300.825
R104 a_232_82.n1 a_232_82.n0 260.606
R105 a_232_82.n0 a_232_82.t2 174.323
R106 a_232_82.n2 a_232_82.t5 134.999
R107 a_232_82.n3 a_232_82.n1 60.2358
R108 a_343_80.t0 a_343_80.n1 764.657
R109 a_343_80.n0 a_343_80.t3 408.43
R110 a_343_80.n0 a_343_80.t2 383.628
R111 a_343_80.n1 a_343_80.t1 314.582
R112 a_343_80.n1 a_343_80.n0 34.9505
R113 VGND.n9 VGND.t3 264.389
R114 VGND.n1 VGND.n0 242.279
R115 VGND.n4 VGND.n3 216.69
R116 VGND.n10 VGND.t6 177.683
R117 VGND.n16 VGND.n15 117.856
R118 VGND.n15 VGND.t4 66.3746
R119 VGND.n0 VGND.t2 55.6369
R120 VGND.n3 VGND.t7 43.5449
R121 VGND.n13 VGND.n8 36.1417
R122 VGND.n14 VGND.n13 36.1417
R123 VGND.n17 VGND.n6 36.1417
R124 VGND.n21 VGND.n6 36.1417
R125 VGND.n22 VGND.n21 36.1417
R126 VGND.n27 VGND.n26 36.1417
R127 VGND.n28 VGND.n27 36.1417
R128 VGND.n23 VGND.n22 34.4114
R129 VGND.n15 VGND.t5 32.0505
R130 VGND.n0 VGND.t1 30.0005
R131 VGND.n3 VGND.t0 25.7805
R132 VGND.n28 VGND.n1 22.7142
R133 VGND.n9 VGND.n8 22.5887
R134 VGND.n26 VGND.n4 17.8201
R135 VGND.n17 VGND.n16 10.9181
R136 VGND.n30 VGND.n1 9.36437
R137 VGND.n29 VGND.n28 9.3005
R138 VGND.n27 VGND.n2 9.3005
R139 VGND.n26 VGND.n25 9.3005
R140 VGND.n24 VGND.n23 9.3005
R141 VGND.n22 VGND.n5 9.3005
R142 VGND.n21 VGND.n20 9.3005
R143 VGND.n19 VGND.n6 9.3005
R144 VGND.n18 VGND.n17 9.3005
R145 VGND.n14 VGND.n7 9.3005
R146 VGND.n13 VGND.n12 9.3005
R147 VGND.n11 VGND.n8 9.3005
R148 VGND.n10 VGND.n9 7.12578
R149 VGND.n23 VGND.n4 3.49141
R150 VGND.n11 VGND.n10 0.478668
R151 VGND.n16 VGND.n14 0.376971
R152 VGND VGND.n30 0.161675
R153 VGND.n30 VGND.n29 0.146149
R154 VGND.n12 VGND.n11 0.122949
R155 VGND.n12 VGND.n7 0.122949
R156 VGND.n18 VGND.n7 0.122949
R157 VGND.n19 VGND.n18 0.122949
R158 VGND.n20 VGND.n19 0.122949
R159 VGND.n20 VGND.n5 0.122949
R160 VGND.n24 VGND.n5 0.122949
R161 VGND.n25 VGND.n24 0.122949
R162 VGND.n25 VGND.n2 0.122949
R163 VGND.n29 VGND.n2 0.122949
R164 VNB.n1 VNB 13153.8
R165 VNB.t3 VNB.t7 3464.57
R166 VNB VNB.n1 2734.58
R167 VNB.t9 VNB.t1 2621.52
R168 VNB.t6 VNB.t8 2298.16
R169 VNB.t1 VNB.t2 1362.73
R170 VNB.t0 VNB.t9 1339.63
R171 VNB.t2 VNB 1143.31
R172 VNB.n1 VNB.t3 1097.11
R173 VNB.t4 VNB.t6 900.788
R174 VNB.t8 VNB.t0 900.788
R175 VNB.n0 VNB.t5 139.38
R176 VNB.n0 VNB.t4 52.1919
R177 VNB.n1 VNB.n0 46.0518
R178 GATE_N.n0 GATE_N.t1 297.233
R179 GATE_N.n0 GATE_N.t0 205.922
R180 GATE_N GATE_N.n0 158.012
R181 a_575_79.t0 a_575_79.t1 45.0005
R182 a_852_123.t0 a_852_123.t1 68.5719
R183 a_571_392.t0 a_571_392.t1 53.1905
R184 a_27_120.t1 a_27_120.n1 463.83
R185 a_27_120.n1 a_27_120.n0 344.673
R186 a_27_120.n0 a_27_120.t2 289.83
R187 a_27_120.n1 a_27_120.t0 215.546
R188 a_27_120.n0 a_27_120.t3 195.305
R189 D.n0 D.t0 233.607
R190 D.n0 D.t1 167.341
R191 D D.n0 68.4016
R192 Q.n0 Q.t0 295.498
R193 Q.n1 Q.t1 279.738
R194 Q.t1 Q.n0 267.106
R195 Q.n1 Q 12.2358
R196 Q.n0 Q 3.57697
R197 Q Q.n1 1.69462
R198 a_805_392.t0 a_805_392.t1 157.131
C0 VPB VGND 0.021259f
C1 GATE_N VPWR 0.02601f
C2 D VGND 0.009951f
C3 a_1347_424# VPB 0.070564f
C4 GATE_N Q 2.23e-20
C5 GATE_N VGND 0.009856f
C6 VPWR Q_N 0.127503f
C7 VPWR Q 0.119368f
C8 VPWR VGND 0.144503f
C9 Q_N VGND 0.102688f
C10 Q VGND 0.103106f
C11 a_1347_424# VPWR 0.246097f
C12 a_1347_424# Q_N 0.070412f
C13 a_1347_424# Q 0.033884f
C14 a_1347_424# VGND 0.160932f
C15 VPB D 0.063309f
C16 VPB GATE_N 0.069203f
C17 D GATE_N 0.090112f
C18 VPB VPWR 0.278958f
C19 VPB Q_N 0.013928f
C20 VPB Q 0.013195f
C21 D VPWR 0.026313f
C22 VGND VNB 0.989302f
C23 Q_N VNB 0.110205f
C24 Q VNB 0.010347f
C25 VPWR VNB 0.760219f
C26 GATE_N VNB 0.10633f
C27 D VNB 0.145839f
C28 VPB VNB 1.9164f
C29 a_1347_424# VNB 0.188284f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxbn_2 VNB VPB VPWR VGND D GATE_N Q Q_N
X0 VPWR.t7 a_887_270.t2 a_814_392.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2473 pd=1.635 as=0.0798 ps=0.8 w=0.42 l=0.15
X1 VPWR.t0 a_1442_94.t2 Q_N.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Q_N.t2 a_1442_94.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_839_123.t1 a_343_74.t2 a_647_79.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0651 pd=0.73 as=0.1976 ps=1.45 w=0.42 l=0.15
X4 a_232_98.t1 GATE_N.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.147 ps=1.19 w=0.84 l=0.15
X5 a_887_270.t0 a_647_79.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.12505 ps=1.145 w=0.74 l=0.15
X6 a_647_79.t2 a_343_74.t3 a_565_392.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2186 pd=1.675 as=0.135 ps=1.27 w=1 l=0.15
X7 a_814_392.t0 a_232_98.t2 a_647_79.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0798 pd=0.8 as=0.2186 ps=1.675 w=0.42 l=0.15
X8 a_565_392.t0 a_27_136.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.1853 ps=1.385 w=1 l=0.15
X9 a_569_79.t0 a_27_136.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.192975 ps=1.395 w=0.64 l=0.15
X10 VGND.t7 a_887_270.t3 a_839_123.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.12505 pd=1.145 as=0.0651 ps=0.73 w=0.42 l=0.15
X11 VPWR.t8 a_232_98.t3 a_343_74.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2478 ps=2.27 w=0.84 l=0.15
X12 a_1442_94.t1 a_887_270.t4 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.1934 ps=1.475 w=1 l=0.15
X13 VPWR.t3 D.t0 a_27_136.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.3192 ps=2.44 w=0.84 l=0.15
X14 VGND.t4 a_1442_94.t4 Q_N.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VPWR.t6 a_887_270.t5 Q.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_1442_94.t0 a_887_270.t6 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X17 VGND.t1 D.t1 a_27_136.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.200625 pd=1.49 as=0.15675 ps=1.67 w=0.55 l=0.15
X18 VGND.t10 a_232_98.t4 a_343_74.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.192975 pd=1.395 as=0.2817 ps=2.29 w=0.74 l=0.15
X19 Q.t1 a_887_270.t7 VGND.t9 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X20 a_887_270.t1 a_647_79.t5 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2473 ps=1.635 w=1.12 l=0.15
X21 Q_N.t0 a_1442_94.t5 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X22 a_647_79.t1 a_232_98.t5 a_569_79.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1976 pd=1.45 as=0.0768 ps=0.88 w=0.64 l=0.15
X23 a_232_98.t0 GATE_N.t1 VGND.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.200625 ps=1.49 w=0.74 l=0.15
X24 VGND.t8 a_887_270.t8 Q.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_887_270.n9 a_887_270.t0 321.43
R1 a_887_270.n3 a_887_270.t4 255.971
R2 a_887_270.n5 a_887_270.t5 240.197
R3 a_887_270.n1 a_887_270.n0 240.197
R4 a_887_270.t1 a_887_270.n10 221.49
R5 a_887_270.n9 a_887_270.n8 199.013
R6 a_887_270.n1 a_887_270.t7 193.53
R7 a_887_270.n8 a_887_270.t3 192.091
R8 a_887_270.n4 a_887_270.t8 179.947
R9 a_887_270.n8 a_887_270.t2 169.867
R10 a_887_270.n7 a_887_270.n2 165.189
R11 a_887_270.n3 a_887_270.t6 163.881
R12 a_887_270.n7 a_887_270.n6 152
R13 a_887_270.n10 a_887_270.n7 144.1
R14 a_887_270.n6 a_887_270.n3 50.3914
R15 a_887_270.n2 a_887_270.n1 36.5157
R16 a_887_270.n6 a_887_270.n5 20.449
R17 a_887_270.n4 a_887_270.n2 15.3369
R18 a_887_270.n5 a_887_270.n4 13.8763
R19 a_887_270.n10 a_887_270.n9 12.7226
R20 a_814_392.t0 a_814_392.t1 178.238
R21 VPWR.n28 VPWR.n4 614.994
R22 VPWR.n15 VPWR.n10 606.333
R23 VPWR.n34 VPWR.n1 316.399
R24 VPWR.n12 VPWR.t0 266.248
R25 VPWR.n11 VPWR.t1 259.171
R26 VPWR.n21 VPWR.n7 216.255
R27 VPWR.n7 VPWR.t7 78.6598
R28 VPWR.n4 VPWR.t8 55.1136
R29 VPWR.n1 VPWR.t4 46.9053
R30 VPWR.n7 VPWR.t9 45.2807
R31 VPWR.n10 VPWR.t5 40.3855
R32 VPWR.n32 VPWR.n2 36.1417
R33 VPWR.n33 VPWR.n32 36.1417
R34 VPWR.n22 VPWR.n5 36.1417
R35 VPWR.n26 VPWR.n5 36.1417
R36 VPWR.n27 VPWR.n26 36.1417
R37 VPWR.n1 VPWR.t3 35.1791
R38 VPWR.n21 VPWR.n20 33.1299
R39 VPWR.n28 VPWR.n27 32.377
R40 VPWR.n4 VPWR.t2 30.4598
R41 VPWR.n15 VPWR.n14 30.1181
R42 VPWR.n20 VPWR.n8 27.8593
R43 VPWR.n10 VPWR.t6 27.6909
R44 VPWR.n16 VPWR.n8 25.6005
R45 VPWR.n14 VPWR.n11 25.224
R46 VPWR.n16 VPWR.n15 17.3181
R47 VPWR.n34 VPWR.n33 16.5652
R48 VPWR.n28 VPWR.n2 15.0593
R49 VPWR.n14 VPWR.n13 9.3005
R50 VPWR.n15 VPWR.n9 9.3005
R51 VPWR.n17 VPWR.n16 9.3005
R52 VPWR.n18 VPWR.n8 9.3005
R53 VPWR.n20 VPWR.n19 9.3005
R54 VPWR.n21 VPWR.n6 9.3005
R55 VPWR.n23 VPWR.n22 9.3005
R56 VPWR.n24 VPWR.n5 9.3005
R57 VPWR.n26 VPWR.n25 9.3005
R58 VPWR.n27 VPWR.n3 9.3005
R59 VPWR.n29 VPWR.n28 9.3005
R60 VPWR.n30 VPWR.n2 9.3005
R61 VPWR.n32 VPWR.n31 9.3005
R62 VPWR.n33 VPWR.n0 9.3005
R63 VPWR.n22 VPWR.n21 8.28285
R64 VPWR.n35 VPWR.n34 7.53404
R65 VPWR.n12 VPWR.n11 6.95806
R66 VPWR.n13 VPWR.n12 0.546775
R67 VPWR VPWR.n35 0.161409
R68 VPWR.n35 VPWR.n0 0.146411
R69 VPWR.n13 VPWR.n9 0.122949
R70 VPWR.n17 VPWR.n9 0.122949
R71 VPWR.n18 VPWR.n17 0.122949
R72 VPWR.n19 VPWR.n18 0.122949
R73 VPWR.n19 VPWR.n6 0.122949
R74 VPWR.n23 VPWR.n6 0.122949
R75 VPWR.n24 VPWR.n23 0.122949
R76 VPWR.n25 VPWR.n24 0.122949
R77 VPWR.n25 VPWR.n3 0.122949
R78 VPWR.n29 VPWR.n3 0.122949
R79 VPWR.n30 VPWR.n29 0.122949
R80 VPWR.n31 VPWR.n30 0.122949
R81 VPWR.n31 VPWR.n0 0.122949
R82 VPB.t11 VPB.t6 745.699
R83 VPB.t5 VPB.t9 574.597
R84 VPB.t7 VPB.t1 515.861
R85 VPB.t10 VPB.t2 421.372
R86 VPB.t8 VPB.t11 339.651
R87 VPB VPB.t4 301.344
R88 VPB.t9 VPB.t3 273.253
R89 VPB.t2 VPB.t8 270.7
R90 VPB.t6 VPB.t7 257.93
R91 VPB.t4 VPB.t5 255.376
R92 VPB.t1 VPB.t0 229.839
R93 VPB.t3 VPB.t10 214.517
R94 a_1442_94.t1 a_1442_94.n3 249.685
R95 a_1442_94.n0 a_1442_94.t2 236.889
R96 a_1442_94.n2 a_1442_94.t3 234.841
R97 a_1442_94.n0 a_1442_94.t4 188.571
R98 a_1442_94.n1 a_1442_94.t5 186.374
R99 a_1442_94.n3 a_1442_94.t0 147.739
R100 a_1442_94.n3 a_1442_94.n2 126.84
R101 a_1442_94.n1 a_1442_94.n0 61.4051
R102 a_1442_94.n2 a_1442_94.n1 4.38232
R103 Q_N.n2 Q_N 589.85
R104 Q_N.n2 Q_N.n0 585
R105 Q_N.n3 Q_N.n2 585
R106 Q_N Q_N.n1 163.368
R107 Q_N.n2 Q_N.t3 26.3844
R108 Q_N.n2 Q_N.t2 26.3844
R109 Q_N.n1 Q_N.t1 22.7032
R110 Q_N.n1 Q_N.t0 22.7032
R111 Q_N Q_N.n3 12.9944
R112 Q_N Q_N.n0 11.249
R113 Q_N Q_N.n0 3.10353
R114 Q_N.n3 Q_N 1.35808
R115 a_343_74.t0 a_343_74.n1 779.231
R116 a_343_74.n0 a_343_74.t3 383.628
R117 a_343_74.n1 a_343_74.t1 339.889
R118 a_343_74.n0 a_343_74.t2 309.974
R119 a_343_74.n1 a_343_74.n0 71.418
R120 a_647_79.n5 a_647_79.n4 326.332
R121 a_647_79.n0 a_647_79.t5 285.719
R122 a_647_79.n1 a_647_79.n0 236.541
R123 a_647_79.n4 a_647_79.n3 188.724
R124 a_647_79.n2 a_647_79.n1 185
R125 a_647_79.n0 a_647_79.t4 178.34
R126 a_647_79.n6 a_647_79.t2 156.113
R127 a_647_79.n5 a_647_79.t0 146.493
R128 a_647_79.t2 a_647_79.n5 116.733
R129 a_647_79.n3 a_647_79.n2 110.001
R130 a_647_79.n3 a_647_79.t1 69.1523
R131 a_647_79.n2 a_647_79.t3 40.0005
R132 a_647_79.n4 a_647_79.n1 7.37441
R133 a_839_123.t0 a_839_123.t1 88.5719
R134 VNB.t2 VNB.t12 2471.39
R135 VNB.t8 VNB.t4 2448.29
R136 VNB.t0 VNB.t7 2286.61
R137 VNB.t10 VNB.t11 2217.32
R138 VNB.t12 VNB.t3 1420.47
R139 VNB.t1 VNB.t2 1362.73
R140 VNB.t6 VNB.t8 1339.63
R141 VNB.t9 VNB.t0 1281.89
R142 VNB VNB.t1 1143.31
R143 VNB.t11 VNB.t9 1062.47
R144 VNB.t4 VNB.t5 993.177
R145 VNB.t7 VNB.t6 993.177
R146 VNB.t3 VNB.t10 900.788
R147 GATE_N.n0 GATE_N.t1 271.527
R148 GATE_N.n0 GATE_N.t0 205.922
R149 GATE_N GATE_N.n0 158.012
R150 a_232_98.n3 a_232_98.n0 408.747
R151 a_232_98.n0 a_232_98.t5 400.207
R152 a_232_98.t1 a_232_98.n3 331.56
R153 a_232_98.n1 a_232_98.t3 323.378
R154 a_232_98.n2 a_232_98.t0 296.639
R155 a_232_98.n2 a_232_98.n1 270.106
R156 a_232_98.n1 a_232_98.t4 167.094
R157 a_232_98.n0 a_232_98.t2 127.731
R158 a_232_98.n3 a_232_98.n2 68.8946
R159 VGND.n8 VGND.t9 306.106
R160 VGND.n1 VGND.n0 275.382
R161 VGND.n23 VGND.n22 210.268
R162 VGND.n4 VGND.n3 209.835
R163 VGND.n11 VGND.t4 170.706
R164 VGND.n10 VGND.t3 154.727
R165 VGND.n15 VGND.n14 116.644
R166 VGND.n0 VGND.t1 55.6369
R167 VGND.n22 VGND.t0 52.3146
R168 VGND.n3 VGND.t2 50.6255
R169 VGND.n22 VGND.t7 47.1434
R170 VGND.n14 VGND.t6 41.2505
R171 VGND.n21 VGND.n20 36.1417
R172 VGND.n24 VGND.n6 36.1417
R173 VGND.n28 VGND.n6 36.1417
R174 VGND.n29 VGND.n28 36.1417
R175 VGND.n30 VGND.n29 36.1417
R176 VGND.n34 VGND.n33 36.1417
R177 VGND.n35 VGND.n34 36.1417
R178 VGND.n15 VGND.n13 32.7534
R179 VGND.n14 VGND.t8 30.6984
R180 VGND.n16 VGND.n8 30.4946
R181 VGND.n0 VGND.t5 30.0005
R182 VGND.n3 VGND.t10 25.3115
R183 VGND.n13 VGND.n10 22.9652
R184 VGND.n20 VGND.n8 22.9652
R185 VGND.n35 VGND.n1 22.7142
R186 VGND.n16 VGND.n15 14.6829
R187 VGND.n33 VGND.n4 13.9375
R188 VGND.n37 VGND.n1 9.36437
R189 VGND.n36 VGND.n35 9.3005
R190 VGND.n34 VGND.n2 9.3005
R191 VGND.n33 VGND.n32 9.3005
R192 VGND.n31 VGND.n30 9.3005
R193 VGND.n29 VGND.n5 9.3005
R194 VGND.n28 VGND.n27 9.3005
R195 VGND.n26 VGND.n6 9.3005
R196 VGND.n25 VGND.n24 9.3005
R197 VGND.n21 VGND.n7 9.3005
R198 VGND.n20 VGND.n19 9.3005
R199 VGND.n18 VGND.n8 9.3005
R200 VGND.n17 VGND.n16 9.3005
R201 VGND.n13 VGND.n12 9.3005
R202 VGND.n15 VGND.n9 9.3005
R203 VGND.n11 VGND.n10 6.6595
R204 VGND.n24 VGND.n23 5.27109
R205 VGND.n30 VGND.n4 4.65505
R206 VGND.n23 VGND.n21 1.88285
R207 VGND.n12 VGND.n11 0.655456
R208 VGND VGND.n37 0.161675
R209 VGND.n37 VGND.n36 0.146149
R210 VGND.n12 VGND.n9 0.122949
R211 VGND.n17 VGND.n9 0.122949
R212 VGND.n18 VGND.n17 0.122949
R213 VGND.n19 VGND.n18 0.122949
R214 VGND.n19 VGND.n7 0.122949
R215 VGND.n25 VGND.n7 0.122949
R216 VGND.n26 VGND.n25 0.122949
R217 VGND.n27 VGND.n26 0.122949
R218 VGND.n27 VGND.n5 0.122949
R219 VGND.n31 VGND.n5 0.122949
R220 VGND.n32 VGND.n31 0.122949
R221 VGND.n32 VGND.n2 0.122949
R222 VGND.n36 VGND.n2 0.122949
R223 a_565_392.t0 a_565_392.t1 53.1905
R224 a_27_136.t1 a_27_136.n1 449.882
R225 a_27_136.n1 a_27_136.n0 346.546
R226 a_27_136.n0 a_27_136.t2 298.572
R227 a_27_136.n1 a_27_136.t0 215.546
R228 a_27_136.n0 a_27_136.t3 186.374
R229 a_569_79.t0 a_569_79.t1 45.0005
R230 D.n0 D.t0 252.744
R231 D.n0 D.t1 181.784
R232 D D.n0 153.196
R233 Q Q.t2 889.909
R234 Q Q.n0 116.751
R235 Q.n0 Q.t0 22.7032
R236 Q.n0 Q.t1 22.7032
C0 VPB GATE_N 0.070761f
C1 D GATE_N 0.066434f
C2 VPB VPWR 0.308141f
C3 D VPWR 0.030649f
C4 VPB VGND 0.022727f
C5 VPB Q 0.005143f
C6 GATE_N VPWR 0.022249f
C7 D VGND 0.00819f
C8 GATE_N VGND 0.007781f
C9 D Q 4.23e-21
C10 VPB Q_N 0.007055f
C11 D Q_N 2.26e-21
C12 GATE_N Q 2.56e-20
C13 VPWR VGND 0.164918f
C14 GATE_N Q_N 8.57e-21
C15 VPWR Q 0.020778f
C16 VGND Q 0.151706f
C17 VPWR Q_N 0.215471f
C18 VGND Q_N 0.15956f
C19 VPB D 0.060373f
C20 Q_N VNB 0.030997f
C21 Q VNB 0.013217f
C22 VGND VNB 1.12468f
C23 VPWR VNB 0.881865f
C24 GATE_N VNB 0.102461f
C25 D VNB 0.135259f
C26 VPB VNB 2.1204f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxbp_1 VNB VPB VPWR VGND Q_N Q GATE D
X0 a_815_124.t1 a_231_74.t2 a_664_392.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1514 ps=1.23 w=0.42 l=0.15
X1 VGND.t0 D.t0 a_27_413.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 a_231_74.t0 GATE.t0 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X3 a_863_98.t0 a_664_392.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2114 ps=1.685 w=1.12 l=0.15
X4 VPWR.t4 a_231_74.t3 a_373_82.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.243825 pd=1.595 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 VGND.t4 a_231_74.t4 a_373_82.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.209725 pd=1.465 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 Q_N a_1347_424# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.3248 ps=2.82 w=1.12 l=0.15
X7 VGND.t2 a_863_98.t2 Q.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.12 pd=1.09 as=0.2072 ps=2.04 w=0.74 l=0.15
X8 a_589_80.t1 a_27_413.t2 VGND.t7 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.209725 ps=1.465 w=0.64 l=0.15
X9 a_863_98.t1 a_664_392.t5 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1471 ps=1.17 w=0.74 l=0.15
X10 VPWR.t0 D.t1 a_27_413.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2338 pd=1.59 as=0.2436 ps=2.26 w=0.84 l=0.15
X11 Q_N.t0 a_1347_424# VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 a_770_508.t0 a_373_82.t2 a_664_392.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.10605 pd=0.925 as=0.1639 ps=1.38 w=0.42 l=0.15
X13 a_231_74.t1 GATE.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2338 ps=1.59 w=0.84 l=0.15
X14 a_664_392.t1 a_373_82.t3 a_589_80.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1514 pd=1.23 as=0.0768 ps=0.88 w=0.64 l=0.15
X15 a_664_392.t2 a_231_74.t5 a_586_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1639 pd=1.38 as=0.12 ps=1.24 w=1 l=0.15
X16 VGND.t3 a_863_98.t3 a_815_124.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1471 pd=1.17 as=0.0504 ps=0.66 w=0.42 l=0.15
X17 VPWR.t2 a_863_98.t4 a_770_508.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2114 pd=1.685 as=0.10605 ps=0.925 w=0.42 l=0.15
X18 a_1347_424# a_863_98.t5 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.12 ps=1.09 w=0.55 l=0.15
X19 a_586_392.t1 a_27_413.t3 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.243825 ps=1.595 w=1 l=0.15
X20 VPWR.t5 a_863_98.t6 Q.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 a_231_74.t1 a_231_74.n2 798.371
R1 a_231_74.t2 a_231_74.t5 706.933
R2 a_231_74.n0 a_231_74.t2 432.635
R3 a_231_74.n1 a_231_74.t4 221.72
R4 a_231_74.n1 a_231_74.t3 184.012
R5 a_231_74.n0 a_231_74.t0 134.325
R6 a_231_74.n2 a_231_74.n1 105.871
R7 a_231_74.n2 a_231_74.n0 39.5512
R8 a_664_392.t2 a_664_392.n2 877.356
R9 a_664_392.n1 a_664_392.t4 292.32
R10 a_664_392.n2 a_664_392.n0 262.93
R11 a_664_392.n2 a_664_392.n1 228.048
R12 a_664_392.n1 a_664_392.t5 184.059
R13 a_664_392.t2 a_664_392.t0 140.435
R14 a_664_392.n0 a_664_392.t3 84.2862
R15 a_664_392.n0 a_664_392.t1 72.0094
R16 a_815_124.t0 a_815_124.t1 68.5719
R17 VNB.t0 VNB.t1 2783.2
R18 VNB.t10 VNB.t6 2644.62
R19 VNB.t9 VNB.t8 2286.61
R20 VNB.t4 VNB.t7 1709.19
R21 VNB.t6 VNB.t5 1489.76
R22 VNB.t2 VNB.t0 1339.63
R23 VNB.t3 VNB.t10 1339.63
R24 VNB.t1 VNB.t9 1154.86
R25 VNB VNB.t3 1154.86
R26 VNB.t7 VNB.t2 900.788
R27 VNB.t5 VNB.t4 900.788
R28 D.n0 D.t1 228.269
R29 D.n0 D.t0 166.35
R30 D D.n0 68.654
R31 a_27_413.t1 a_27_413.n1 776.634
R32 a_27_413.t1 a_27_413.n2 761.621
R33 a_27_413.n1 a_27_413.n0 353.995
R34 a_27_413.n2 a_27_413.t0 306.909
R35 a_27_413.n0 a_27_413.t2 260.884
R36 a_27_413.n0 a_27_413.t3 227.411
R37 a_27_413.n2 a_27_413.n1 15.0266
R38 VGND.n7 VGND.n6 228.776
R39 VGND.n21 VGND.n20 213.945
R40 VGND.n8 VGND.t5 177.679
R41 VGND.n29 VGND.n28 119.719
R42 VGND.n14 VGND.n13 117.663
R43 VGND.n13 VGND.t3 67.0573
R44 VGND.n28 VGND.t0 51.1959
R45 VGND.n20 VGND.t4 50.4716
R46 VGND.n6 VGND.t6 38.1823
R47 VGND.n11 VGND.n5 36.1417
R48 VGND.n12 VGND.n11 36.1417
R49 VGND.n18 VGND.n3 36.1417
R50 VGND.n19 VGND.n18 36.1417
R51 VGND.n26 VGND.n1 36.1417
R52 VGND.n27 VGND.n26 36.1417
R53 VGND.n14 VGND.n3 33.1299
R54 VGND.n28 VGND.t8 32.4366
R55 VGND.n6 VGND.t2 31.639
R56 VGND.n22 VGND.n19 31.1981
R57 VGND.n13 VGND.t1 28.6551
R58 VGND.n20 VGND.t7 27.5561
R59 VGND.n7 VGND.n5 22.2123
R60 VGND.n21 VGND.n1 19.596
R61 VGND.n29 VGND.n27 18.0711
R62 VGND.n14 VGND.n12 14.3064
R63 VGND.n9 VGND.n5 9.3005
R64 VGND.n11 VGND.n10 9.3005
R65 VGND.n12 VGND.n4 9.3005
R66 VGND.n15 VGND.n14 9.3005
R67 VGND.n16 VGND.n3 9.3005
R68 VGND.n18 VGND.n17 9.3005
R69 VGND.n19 VGND.n2 9.3005
R70 VGND.n23 VGND.n22 9.3005
R71 VGND.n24 VGND.n1 9.3005
R72 VGND.n26 VGND.n25 9.3005
R73 VGND.n27 VGND.n0 9.3005
R74 VGND.n30 VGND.n29 7.47871
R75 VGND.n8 VGND.n7 7.13856
R76 VGND.n22 VGND.n21 2.45707
R77 VGND.n9 VGND.n8 0.479515
R78 VGND VGND.n30 0.16068
R79 VGND.n30 VGND.n0 0.14713
R80 VGND.n10 VGND.n9 0.122949
R81 VGND.n10 VGND.n4 0.122949
R82 VGND.n15 VGND.n4 0.122949
R83 VGND.n16 VGND.n15 0.122949
R84 VGND.n17 VGND.n16 0.122949
R85 VGND.n17 VGND.n2 0.122949
R86 VGND.n23 VGND.n2 0.122949
R87 VGND.n24 VGND.n23 0.122949
R88 VGND.n25 VGND.n24 0.122949
R89 VGND.n25 VGND.n0 0.122949
R90 GATE.n0 GATE.t1 300.983
R91 GATE.n0 GATE.t0 178.34
R92 GATE GATE.n0 158.788
R93 VPWR.n19 VPWR.n18 687.019
R94 VPWR.n12 VPWR.n3 676.107
R95 VPWR.n6 VPWR.n5 599.562
R96 VPWR.n7 VPWR.t5 363.344
R97 VPWR.n5 VPWR.t1 121.453
R98 VPWR.n5 VPWR.t2 119.608
R99 VPWR.n3 VPWR.t4 64.4945
R100 VPWR.n18 VPWR.t3 53.941
R101 VPWR.n18 VPWR.t0 53.941
R102 VPWR.n16 VPWR.n1 36.1417
R103 VPWR.n17 VPWR.n16 36.1417
R104 VPWR.n10 VPWR.n4 36.1417
R105 VPWR.n11 VPWR.n10 36.1417
R106 VPWR.n3 VPWR.t6 35.6631
R107 VPWR.n6 VPWR.n4 30.8711
R108 VPWR.n12 VPWR.n11 30.8711
R109 VPWR.n19 VPWR.n17 21.3031
R110 VPWR.n12 VPWR.n1 16.5652
R111 VPWR.n20 VPWR.n19 9.62791
R112 VPWR.n8 VPWR.n4 9.3005
R113 VPWR.n10 VPWR.n9 9.3005
R114 VPWR.n11 VPWR.n2 9.3005
R115 VPWR.n13 VPWR.n12 9.3005
R116 VPWR.n14 VPWR.n1 9.3005
R117 VPWR.n16 VPWR.n15 9.3005
R118 VPWR.n17 VPWR.n0 9.3005
R119 VPWR.n7 VPWR.n6 4.24299
R120 VPWR.n8 VPWR.n7 0.232061
R121 VPWR VPWR.n20 0.161949
R122 VPWR.n20 VPWR.n0 0.145878
R123 VPWR.n9 VPWR.n8 0.122949
R124 VPWR.n9 VPWR.n2 0.122949
R125 VPWR.n13 VPWR.n2 0.122949
R126 VPWR.n14 VPWR.n13 0.122949
R127 VPWR.n15 VPWR.n14 0.122949
R128 VPWR.n15 VPWR.n0 0.122949
R129 a_863_98.n5 a_863_98.t3 365.298
R130 a_863_98.n1 a_863_98.n0 264.832
R131 a_863_98.n3 a_863_98.t6 234.841
R132 a_863_98.n4 a_863_98.n3 231.603
R133 a_863_98.t0 a_863_98.n6 224.459
R134 a_863_98.n6 a_863_98.n5 186.588
R135 a_863_98.n2 a_863_98.t2 179.947
R136 a_863_98.n4 a_863_98.t1 164.843
R137 a_863_98.n5 a_863_98.t4 154.508
R138 a_863_98.n1 a_863_98.t5 151.612
R139 a_863_98.n2 a_863_98.n1 70.8399
R140 a_863_98.n6 a_863_98.n4 16.8284
R141 a_863_98.n3 a_863_98.n2 2.92171
R142 VPB.t3 VPB.t5 577.152
R143 VPB.t1 VPB.t7 515.861
R144 VPB.t8 VPB.t1 365.188
R145 VPB.t2 VPB.t8 334.543
R146 VPB.t5 VPB.t6 314.113
R147 VPB.t0 VPB.t3 311.56
R148 VPB.t4 VPB.t2 270.7
R149 VPB VPB.t0 255.376
R150 VPB.t6 VPB.t4 199.195
R151 a_373_82.t0 a_373_82.n1 815.152
R152 a_373_82.n0 a_373_82.t1 358.784
R153 a_373_82.n1 a_373_82.t2 345.717
R154 a_373_82.n0 a_373_82.t3 314.274
R155 a_373_82.n1 a_373_82.n0 76.7765
R156 Q_N.n3 Q_N.n0 1214.34
R157 Q_N.n2 Q_N.t0 279.738
R158 Q_N.t0 Q_N.n1 279.738
R159 Q_N Q_N.n3 12.8005
R160 Q_N.n1 Q_N 12.4184
R161 Q_N Q_N.n2 9.36169
R162 Q_N Q_N.n0 7.47404
R163 Q_N.n0 Q_N 6.58162
R164 Q_N.n2 Q_N 4.77662
R165 Q_N.n1 Q_N 1.7199
R166 Q_N.n3 Q_N 1.33781
R167 Q.n0 Q.t0 292.108
R168 Q.t1 Q.n0 281.43
R169 Q.n1 Q.t1 281.43
R170 Q.n1 Q 11.8308
R171 Q.n0 Q 5.62474
R172 Q Q.n1 2.52171
R173 a_589_80.t0 a_589_80.t1 45.0005
R174 a_770_508.t0 a_770_508.t1 236.869
R175 a_586_392.t0 a_586_392.t1 47.2805
C0 GATE Q 4.01e-21
C1 VPWR a_1347_424# 0.227776f
C2 GATE Q_N 1.89e-21
C3 VGND Q 0.100648f
C4 VGND Q_N 0.101699f
C5 GATE a_1347_424# 2.57e-21
C6 VGND a_1347_424# 0.145898f
C7 VPB VPWR 0.253345f
C8 Q a_1347_424# 0.032978f
C9 VPB D 0.05985f
C10 Q_N a_1347_424# 0.065392f
C11 VPB GATE 0.054724f
C12 VPWR D 0.01426f
C13 VPB VGND 0.02099f
C14 VPWR GATE 0.010078f
C15 VPB Q 0.012467f
C16 VPWR VGND 0.150558f
C17 D GATE 0.089612f
C18 VPB Q_N 0.013933f
C19 D VGND 0.036579f
C20 VPWR Q 0.116373f
C21 VPWR Q_N 0.128805f
C22 GATE VGND 0.020051f
C23 VPB a_1347_424# 0.07935f
C24 Q_N VNB 0.110208f
C25 Q VNB 0.014248f
C26 VGND VNB 1.00303f
C27 GATE VNB 0.120964f
C28 D VNB 0.15192f
C29 VPWR VNB 0.756881f
C30 VPB VNB 1.90613f
C31 a_1347_424# VNB 0.200829f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlygate4sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlygate4sd1_1 VNB VPB VPWR VGND A X
X0 VPWR.t1 A.t0 a_28_74.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.31125 pd=1.695 as=0.1176 ps=1.4 w=0.42 l=0.15
X1 a_288_74.t0 a_28_74.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.31125 ps=1.695 w=1 l=0.18
X2 X.t1 a_405_138.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.11485 ps=1.085 w=0.74 l=0.15
X3 VGND.t1 A.t1 a_28_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15435 pd=1.155 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VGND.t0 a_288_74.t2 a_405_138.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.11485 pd=1.085 as=0.2562 ps=2.06 w=0.42 l=0.15
X5 X.t0 a_405_138.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.194 ps=1.475 w=1.12 l=0.15
X6 VPWR.t0 a_288_74.t3 a_405_138.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.475 as=0.58 ps=3.16 w=1 l=0.18
X7 a_288_74.t1 a_28_74.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.15435 ps=1.155 w=0.42 l=0.15
R0 A.n0 A.t0 313.837
R1 A.n0 A.t1 220.113
R2 A A.n0 159.929
R3 a_28_74.n0 a_28_74.t0 737.053
R4 a_28_74.t1 a_28_74.n3 289.522
R5 a_28_74.n1 a_28_74.t2 192.639
R6 a_28_74.n2 a_28_74.t3 192.639
R7 a_28_74.n1 a_28_74.n0 152
R8 a_28_74.n3 a_28_74.n2 152
R9 a_28_74.n2 a_28_74.n1 32.7765
R10 a_28_74.n3 a_28_74.n0 13.1884
R11 VPWR.n2 VPWR.n1 621.289
R12 VPWR.n2 VPWR.n0 323.997
R13 VPWR.n1 VPWR.t2 103.425
R14 VPWR.n1 VPWR.t1 67.4965
R15 VPWR.n0 VPWR.t0 40.3855
R16 VPWR.n0 VPWR.t3 27.3314
R17 VPWR VPWR.n2 0.195508
R18 VPB.t2 VPB.t0 684.409
R19 VPB.t1 VPB.t2 439.248
R20 VPB.t0 VPB.t3 265.591
R21 VPB VPB.t1 252.823
R22 a_288_74.t0 a_288_74.n1 665.54
R23 a_288_74.n1 a_288_74.t1 272.24
R24 a_288_74.n0 a_288_74.t3 190.123
R25 a_288_74.n1 a_288_74.n0 138.701
R26 a_288_74.n0 a_288_74.t2 130.725
R27 a_405_138.t1 a_405_138.n1 744.612
R28 a_405_138.n1 a_405_138.t0 389.591
R29 a_405_138.n0 a_405_138.t3 265.637
R30 a_405_138.n0 a_405_138.t2 202.44
R31 a_405_138.n1 a_405_138.n0 152
R32 VGND.n2 VGND.n0 217.103
R33 VGND.n2 VGND.n1 212.748
R34 VGND.n1 VGND.t2 154.286
R35 VGND.n0 VGND.t0 60.0005
R36 VGND.n1 VGND.t1 55.7148
R37 VGND.n0 VGND.t3 21.8924
R38 VGND VGND.n2 0.196947
R39 X.n1 X 588.702
R40 X.n1 X.n0 585
R41 X.n2 X.n1 585
R42 X.t1 X.n3 284.623
R43 X.n4 X.t1 282.358
R44 X.n1 X.t0 27.2639
R45 X.n2 X 10.333
R46 X.n3 X 9.87038
R47 X X.n4 9.06207
R48 X.n0 X 8.01978
R49 X.n4 X 3.54749
R50 X.n0 X 3.39327
R51 X.n3 X 1.54267
R52 X X.n2 1.08002
R53 VNB.t2 VNB.t0 3106.56
R54 VNB.t1 VNB.t2 2044.09
R55 VNB.t0 VNB.t3 1143.31
R56 VNB VNB.t1 1108.66
C0 VPB A 0.092768f
C1 VPWR X 0.134114f
C2 VPWR VGND 0.063785f
C3 X VGND 0.092359f
C4 VPB VPWR 0.128753f
C5 VPB X 0.020957f
C6 A VPWR 0.01616f
C7 VPB VGND 0.010293f
C8 A X 1.81e-19
C9 A VGND 0.017399f
C10 VGND VNB 0.506354f
C11 X VNB 0.119844f
C12 VPWR VNB 0.396994f
C13 A VNB 0.218678f
C14 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxtp_1 VNB VPB VPWR VGND D Q GATE
X0 VGND.t4 a_592_149.t4 a_386_326.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.19615 pd=1.41 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 a_592_149.t0 a_562_123.t1 a_229_392.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.295 ps=2.59 w=1 l=0.15
X2 a_685_59.t0 a_562_123.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.19615 ps=1.41 w=0.74 l=0.15
X3 a_116_424.t0 D.t0 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1815 pd=1.76 as=0.1705 ps=1.72 w=0.55 l=0.15
X4 a_419_392.t1 a_685_59.t2 a_592_149.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.19295 pd=1.83 as=0.1664 ps=1.385 w=0.42 l=0.15
X5 VPWR.t4 GATE.t0 a_562_123.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 a_419_392.t0 a_386_326.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.193575 ps=1.7 w=0.42 l=0.15
X7 Q.t0 a_386_326.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.261625 ps=1.545 w=0.74 l=0.15
X8 VPWR.t6 a_116_424.t2 a_229_392.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.193575 pd=1.7 as=0.295 ps=2.59 w=1 l=0.15
X9 a_239_85.t0 a_685_59.t3 a_592_149.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=2.08 as=0.13765 ps=1.205 w=0.74 l=0.15
X10 a_116_424.t1 D.t1 VPWR.t5 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2478 ps=2.27 w=0.84 l=0.15
X11 a_592_149.t1 a_562_123.t3 a_514_149.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.13765 pd=1.205 as=0.0504 ps=0.66 w=0.42 l=0.15
X12 a_685_59.t1 a_562_123.t4 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.30135 ps=1.94 w=0.84 l=0.15
X13 VPWR.t3 a_592_149.t5 a_386_326.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.30135 pd=1.94 as=0.3696 ps=2.9 w=1.12 l=0.15
X14 VGND.t3 a_116_424.t3 a_239_85.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.19645 pd=1.485 as=0.2238 ps=2.14 w=0.74 l=0.15
X15 a_514_149.t0 a_386_326.t4 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.19645 ps=1.485 w=0.42 l=0.15
X16 Q.t1 a_386_326.t5 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.231 ps=1.555 w=1.12 l=0.15
R0 a_592_149.t0 a_592_149.n2 931.005
R1 a_592_149.n2 a_592_149.n0 338.515
R2 a_592_149.n0 a_592_149.t5 287.058
R3 a_592_149.n2 a_592_149.n1 185
R4 a_592_149.n0 a_592_149.t4 168.701
R5 a_592_149.t0 a_592_149.t2 142.493
R6 a_592_149.n1 a_592_149.t1 64.2862
R7 a_592_149.n1 a_592_149.t3 53.1279
R8 a_386_326.t1 a_386_326.n3 875.845
R9 a_386_326.t4 a_386_326.t2 480.394
R10 a_386_326.n2 a_386_326.t4 463.541
R11 a_386_326.n1 a_386_326.n0 363.796
R12 a_386_326.n3 a_386_326.t0 279.738
R13 a_386_326.t0 a_386_326.n2 279.738
R14 a_386_326.n0 a_386_326.t5 258.582
R15 a_386_326.n0 a_386_326.t3 197.261
R16 a_386_326.n3 a_386_326.n1 17.4085
R17 a_386_326.n2 a_386_326.n1 5.6325
R18 VGND.n8 VGND.t0 293.791
R19 VGND.n24 VGND.t5 248.733
R20 VGND.n2 VGND.n1 222.042
R21 VGND.n7 VGND.n6 220.173
R22 VGND.n1 VGND.t1 165.714
R23 VGND.n12 VGND.n11 36.1417
R24 VGND.n12 VGND.n4 36.1417
R25 VGND.n16 VGND.n4 36.1417
R26 VGND.n17 VGND.n16 36.1417
R27 VGND.n18 VGND.n17 36.1417
R28 VGND.n23 VGND.n22 36.1417
R29 VGND.n22 VGND.n2 35.7652
R30 VGND.n6 VGND.t2 35.6762
R31 VGND.n6 VGND.t4 35.6762
R32 VGND.n11 VGND.n10 33.9171
R33 VGND.n1 VGND.t3 31.6993
R34 VGND.n8 VGND.n7 26.5057
R35 VGND.n24 VGND.n23 20.7064
R36 VGND.n18 VGND.n2 11.6711
R37 VGND.n25 VGND.n24 9.3005
R38 VGND.n23 VGND.n0 9.3005
R39 VGND.n22 VGND.n21 9.3005
R40 VGND.n20 VGND.n2 9.3005
R41 VGND.n10 VGND.n9 9.3005
R42 VGND.n11 VGND.n5 9.3005
R43 VGND.n13 VGND.n12 9.3005
R44 VGND.n14 VGND.n4 9.3005
R45 VGND.n16 VGND.n15 9.3005
R46 VGND.n17 VGND.n3 9.3005
R47 VGND.n19 VGND.n18 9.3005
R48 VGND.n10 VGND.n7 3.10353
R49 VGND.n9 VGND.n8 0.242475
R50 VGND.n9 VGND.n5 0.122949
R51 VGND.n13 VGND.n5 0.122949
R52 VGND.n14 VGND.n13 0.122949
R53 VGND.n15 VGND.n14 0.122949
R54 VGND.n15 VGND.n3 0.122949
R55 VGND.n19 VGND.n3 0.122949
R56 VGND.n20 VGND.n19 0.122949
R57 VGND.n21 VGND.n20 0.122949
R58 VGND.n21 VGND.n0 0.122949
R59 VGND.n25 VGND.n0 0.122949
R60 VGND VGND.n25 0.0617245
R61 VNB.n0 VNB 13546.5
R62 VNB VNB.n1 10333.7
R63 VNB.n0 VNB.t1 3048.82
R64 VNB.t4 VNB.t7 2494.49
R65 VNB.t0 VNB.t4 2067.19
R66 VNB.n1 VNB.t6 1898.29
R67 VNB.t6 VNB.t2 1483.43
R68 VNB.t5 VNB.t3 1420.47
R69 VNB.n1 VNB.t5 1408.92
R70 VNB.t7 VNB 1201.05
R71 VNB.t2 VNB.n0 1030.86
R72 VNB.t3 VNB.t0 900.788
R73 a_562_123.n2 a_562_123.n1 407.899
R74 a_562_123.t0 a_562_123.n2 325.716
R75 a_562_123.n2 a_562_123.n0 325.327
R76 a_562_123.n1 a_562_123.t1 238.108
R77 a_562_123.n0 a_562_123.t4 233.502
R78 a_562_123.n0 a_562_123.t2 183.161
R79 a_562_123.n1 a_562_123.t3 175.448
R80 a_229_392.t0 a_229_392.t1 1139.45
R81 VPB.t6 VPB.t5 648.657
R82 VPB.t4 VPB.t8 577.152
R83 VPB.t1 VPB.t7 515.861
R84 VPB.t2 VPB.t3 515.861
R85 VPB.t8 VPB.t6 316.668
R86 VPB.t5 VPB.t0 298.791
R87 VPB.t7 VPB.t4 273.253
R88 VPB.t3 VPB.t1 257.93
R89 VPB VPB.t2 257.93
R90 a_685_59.n1 a_685_59.t0 330.81
R91 a_685_59.n1 a_685_59.n0 329.163
R92 a_685_59.t1 a_685_59.n1 323.392
R93 a_685_59.n0 a_685_59.t2 320.2
R94 a_685_59.n0 a_685_59.t3 171.841
R95 D.n0 D.t1 235.377
R96 D.n1 D.t0 173.52
R97 D D.n0 154.861
R98 D.n2 D.n1 152
R99 D.n1 D.n0 49.6611
R100 D D.n2 6.4005
R101 D.n2 D 3.6771
R102 a_116_424.t1 a_116_424.n1 433.349
R103 a_116_424.n0 a_116_424.t2 317.317
R104 a_116_424.n1 a_116_424.t0 253.871
R105 a_116_424.n1 a_116_424.n0 197.337
R106 a_116_424.n0 a_116_424.t3 170.308
R107 a_419_392.t0 a_419_392.t1 1492.43
R108 GATE.n1 GATE.n0 207.261
R109 GATE.n1 GATE.t0 205.922
R110 GATE GATE.n1 156.614
R111 VPWR.n8 VPWR.n7 869.418
R112 VPWR.n17 VPWR.n16 715.178
R113 VPWR.n24 VPWR.t5 409.56
R114 VPWR.n6 VPWR.n5 333.574
R115 VPWR.n16 VPWR.t0 105.537
R116 VPWR.n7 VPWR.t2 65.6672
R117 VPWR.n5 VPWR.t4 55.1136
R118 VPWR.n5 VPWR.t1 38.522
R119 VPWR.n23 VPWR.n22 36.1417
R120 VPWR.n10 VPWR.n9 36.1417
R121 VPWR.n10 VPWR.n3 36.1417
R122 VPWR.n14 VPWR.n3 36.1417
R123 VPWR.n15 VPWR.n14 36.1417
R124 VPWR.n18 VPWR.n15 36.1417
R125 VPWR.n22 VPWR.n1 35.1923
R126 VPWR.n7 VPWR.t3 34.0942
R127 VPWR.n16 VPWR.t6 25.791
R128 VPWR.n9 VPWR.n8 24.7881
R129 VPWR.n24 VPWR.n23 20.7064
R130 VPWR.n18 VPWR.n17 17.1545
R131 VPWR.n9 VPWR.n4 9.3005
R132 VPWR.n11 VPWR.n10 9.3005
R133 VPWR.n12 VPWR.n3 9.3005
R134 VPWR.n14 VPWR.n13 9.3005
R135 VPWR.n15 VPWR.n2 9.3005
R136 VPWR.n19 VPWR.n18 9.3005
R137 VPWR.n20 VPWR.n1 9.3005
R138 VPWR.n22 VPWR.n21 9.3005
R139 VPWR.n23 VPWR.n0 9.3005
R140 VPWR.n25 VPWR.n24 9.3005
R141 VPWR.n8 VPWR.n6 8.17974
R142 VPWR.n17 VPWR.n1 4.03528
R143 VPWR.n6 VPWR.n4 0.165473
R144 VPWR.n11 VPWR.n4 0.122949
R145 VPWR.n12 VPWR.n11 0.122949
R146 VPWR.n13 VPWR.n12 0.122949
R147 VPWR.n13 VPWR.n2 0.122949
R148 VPWR.n19 VPWR.n2 0.122949
R149 VPWR.n20 VPWR.n19 0.122949
R150 VPWR.n21 VPWR.n20 0.122949
R151 VPWR.n21 VPWR.n0 0.122949
R152 VPWR.n25 VPWR.n0 0.122949
R153 VPWR VPWR.n25 0.0617245
R154 Q.n1 Q 589.385
R155 Q.n1 Q.n0 585
R156 Q.n2 Q.n1 585
R157 Q Q.t0 202.212
R158 Q.n1 Q.t1 26.3844
R159 Q Q.n2 11.7484
R160 Q Q.n0 10.1704
R161 Q Q.n0 2.80598
R162 Q.n2 Q 1.2279
R163 a_239_85.t0 a_239_85.t1 670.255
R164 a_514_149.t0 a_514_149.t1 68.5719
C0 VPB GATE 0.047552f
C1 VPWR D 0.048707f
C2 VPWR GATE 0.019175f
C3 VPB Q 0.015418f
C4 VPB VGND 0.02138f
C5 VPWR Q 0.12796f
C6 VPWR VGND 0.12516f
C7 GATE Q 0.005492f
C8 D VGND 0.051723f
C9 GATE VGND 0.011131f
C10 Q VGND 0.041794f
C11 VPB VPWR 0.246565f
C12 VPB D 0.069875f
C13 VGND VNB 0.945089f
C14 Q VNB 0.110683f
C15 GATE VNB 0.109127f
C16 D VNB 0.189991f
C17 VPWR VNB 0.745493f
C18 VPB VNB 1.83163f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxtn_4 VNB VPB VPWR VGND D GATE_N Q
X0 VPWR.t1 a_840_395.t3 a_789_508.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.21945 pd=1.62 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR.t5 a_840_395.t4 Q.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_789_508.t1 a_230_424.t2 a_675_392.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.17375 ps=1.42 w=0.42 l=0.15
X3 Q.t2 a_840_395.t5 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t3 a_840_395.t6 Q.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.21 ps=1.495 w=1.12 l=0.15
X5 VPWR.t9 a_675_392.t4 a_840_395.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.1491 ps=1.195 w=0.84 l=0.15
X6 VPWR.t0 D.t0 a_27_115.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X7 a_230_424.t0 GATE_N.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.201575 ps=1.57 w=0.74 l=0.15
X8 VGND.t8 a_230_424.t3 a_369_392.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2397 pd=1.45 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 VPWR.t6 a_230_424.t4 a_369_392.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2503 pd=1.515 as=0.2478 ps=2.27 w=0.84 l=0.15
X10 a_840_395.t1 a_675_392.t5 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1491 pd=1.195 as=0.21945 ps=1.62 w=0.84 l=0.15
X11 a_675_392.t1 a_230_424.t5 a_658_79.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.16295 pd=1.285 as=0.0768 ps=0.88 w=0.64 l=0.15
X12 Q.t0 a_840_395.t7 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.495 as=0.1862 ps=1.475 w=1.12 l=0.15
X13 a_230_424.t1 GATE_N.t1 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.168 ps=1.24 w=0.84 l=0.15
X14 Q.t6 a_840_395.t8 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1369 pd=1.11 as=0.1293 ps=1.105 w=0.74 l=0.15
X15 VGND.t4 a_840_395.t9 a_895_123.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1031 pd=1 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_675_392.t0 a_369_392.t2 a_591_392.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.17375 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t2 a_840_395.t10 Q.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1369 ps=1.11 w=0.74 l=0.15
X18 a_591_392.t1 a_27_115.t2 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2503 ps=1.515 w=1 l=0.15
X19 a_895_123.t0 a_369_392.t3 a_675_392.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.16295 ps=1.285 w=0.42 l=0.15
X20 VGND.t7 D.t1 a_27_115.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.201575 pd=1.57 as=0.15675 ps=1.67 w=0.55 l=0.15
X21 Q.t4 a_840_395.t11 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_658_79.t0 a_27_115.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2397 ps=1.45 w=0.64 l=0.15
X23 a_840_395.t2 a_675_392.t6 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1031 ps=1 w=0.64 l=0.15
R0 a_840_395.n0 a_840_395.t9 375.411
R1 a_840_395.n17 a_840_395.n16 302.587
R2 a_840_395.n4 a_840_395.t4 236.862
R3 a_840_395.n5 a_840_395.t5 234.841
R4 a_840_395.n9 a_840_395.t6 234.841
R5 a_840_395.n12 a_840_395.t7 234.841
R6 a_840_395.n12 a_840_395.t8 188.565
R7 a_840_395.n4 a_840_395.n3 186.374
R8 a_840_395.n10 a_840_395.t10 186.374
R9 a_840_395.n2 a_840_395.t11 186.374
R10 a_840_395.n16 a_840_395.n0 181.48
R11 a_840_395.n0 a_840_395.t3 173.131
R12 a_840_395.n15 a_840_395.t2 169.268
R13 a_840_395.n7 a_840_395.n6 165.189
R14 a_840_395.n14 a_840_395.n13 152
R15 a_840_395.n11 a_840_395.n1 152
R16 a_840_395.n8 a_840_395.n7 152
R17 a_840_395.n13 a_840_395.n11 49.6611
R18 a_840_395.n6 a_840_395.n4 46.0096
R19 a_840_395.n17 a_840_395.t1 43.3874
R20 a_840_395.t0 a_840_395.n17 39.8695
R21 a_840_395.n9 a_840_395.n8 33.5944
R22 a_840_395.n16 a_840_395.n15 29.4451
R23 a_840_395.n8 a_840_395.n2 26.2914
R24 a_840_395.n15 a_840_395.n14 21.7217
R25 a_840_395.n6 a_840_395.n5 17.5278
R26 a_840_395.n7 a_840_395.n1 13.1884
R27 a_840_395.n14 a_840_395.n1 13.1884
R28 a_840_395.n11 a_840_395.n10 13.146
R29 a_840_395.n13 a_840_395.n12 10.955
R30 a_840_395.n5 a_840_395.n2 5.84292
R31 a_840_395.n10 a_840_395.n9 2.92171
R32 a_789_508.t0 a_789_508.t1 126.644
R33 VPWR.n28 VPWR.n4 606.284
R34 VPWR.n21 VPWR.n20 585
R35 VPWR.n19 VPWR.n18 585
R36 VPWR.n9 VPWR.t5 349.373
R37 VPWR.n11 VPWR.n10 317.716
R38 VPWR.n8 VPWR.n7 317.152
R39 VPWR.n34 VPWR.n1 315.926
R40 VPWR.n20 VPWR.n19 215.762
R41 VPWR.n20 VPWR.t1 72.7029
R42 VPWR.n4 VPWR.t6 70.3576
R43 VPWR.n1 VPWR.t7 46.9053
R44 VPWR.n1 VPWR.t0 46.9053
R45 VPWR.n19 VPWR.t10 45.7326
R46 VPWR.n7 VPWR.t9 42.2148
R47 VPWR.n4 VPWR.t8 38.2012
R48 VPWR.n7 VPWR.t2 36.8622
R49 VPWR.n32 VPWR.n2 36.1417
R50 VPWR.n33 VPWR.n32 36.1417
R51 VPWR.n26 VPWR.n5 36.1417
R52 VPWR.n27 VPWR.n26 36.1417
R53 VPWR.n17 VPWR.n16 29.8649
R54 VPWR.n10 VPWR.t4 26.3844
R55 VPWR.n10 VPWR.t3 26.3844
R56 VPWR.n21 VPWR.n5 25.3586
R57 VPWR.n12 VPWR.n11 25.224
R58 VPWR.n12 VPWR.n8 25.224
R59 VPWR.n28 VPWR.n27 22.5887
R60 VPWR.n16 VPWR.n8 22.2123
R61 VPWR.n34 VPWR.n33 17.6946
R62 VPWR.n28 VPWR.n2 15.0593
R63 VPWR.n13 VPWR.n12 9.3005
R64 VPWR.n14 VPWR.n8 9.3005
R65 VPWR.n16 VPWR.n15 9.3005
R66 VPWR.n17 VPWR.n6 9.3005
R67 VPWR.n23 VPWR.n22 9.3005
R68 VPWR.n24 VPWR.n5 9.3005
R69 VPWR.n26 VPWR.n25 9.3005
R70 VPWR.n27 VPWR.n3 9.3005
R71 VPWR.n29 VPWR.n28 9.3005
R72 VPWR.n30 VPWR.n2 9.3005
R73 VPWR.n32 VPWR.n31 9.3005
R74 VPWR.n33 VPWR.n0 9.3005
R75 VPWR.n35 VPWR.n34 7.49287
R76 VPWR.n22 VPWR.n18 6.51686
R77 VPWR.n11 VPWR.n9 6.50549
R78 VPWR.n18 VPWR.n17 0.931409
R79 VPWR.n13 VPWR.n9 0.686474
R80 VPWR.n22 VPWR.n21 0.621106
R81 VPWR VPWR.n35 0.160867
R82 VPWR.n35 VPWR.n0 0.146947
R83 VPWR.n14 VPWR.n13 0.122949
R84 VPWR.n15 VPWR.n14 0.122949
R85 VPWR.n15 VPWR.n6 0.122949
R86 VPWR.n23 VPWR.n6 0.122949
R87 VPWR.n24 VPWR.n23 0.122949
R88 VPWR.n25 VPWR.n24 0.122949
R89 VPWR.n25 VPWR.n3 0.122949
R90 VPWR.n29 VPWR.n3 0.122949
R91 VPWR.n30 VPWR.n29 0.122949
R92 VPWR.n31 VPWR.n30 0.122949
R93 VPWR.n31 VPWR.n0 0.122949
R94 VPB.t8 VPB.t7 582.259
R95 VPB.t5 VPB.t12 475
R96 VPB.t7 VPB.t9 339.651
R97 VPB.t6 VPB.t10 291.13
R98 VPB.t0 VPB.t8 280.914
R99 VPB.t1 VPB.t2 268.146
R100 VPB VPB.t0 268.146
R101 VPB.t11 VPB.t1 257.93
R102 VPB.t12 VPB.t11 257.93
R103 VPB.t3 VPB.t4 229.839
R104 VPB.t2 VPB.t3 229.839
R105 VPB.t10 VPB.t5 214.517
R106 VPB.t9 VPB.t6 214.517
R107 Q.n2 Q.n1 261.731
R108 Q.n2 Q.n0 203.512
R109 Q.n4 Q.n3 151.298
R110 Q.n4 Q.t4 144.683
R111 Q.n3 Q.t5 35.6762
R112 Q.n1 Q.t1 35.1791
R113 Q.n1 Q.t0 30.7817
R114 Q Q.n4 27.6465
R115 Q.n0 Q.t3 26.3844
R116 Q.n0 Q.t2 26.3844
R117 Q.n3 Q.t6 24.3248
R118 Q Q.n2 15.7096
R119 a_230_424.t1 a_230_424.n1 777.014
R120 a_230_424.t1 a_230_424.n4 768.644
R121 a_230_424.n1 a_230_424.n0 509.591
R122 a_230_424.n3 a_230_424.t0 292.892
R123 a_230_424.n0 a_230_424.t2 287.058
R124 a_230_424.n0 a_230_424.t5 256.045
R125 a_230_424.n2 a_230_424.t4 189.855
R126 a_230_424.n2 a_230_424.t3 164.97
R127 a_230_424.n3 a_230_424.n2 92.6775
R128 a_230_424.n4 a_230_424.n3 41.6612
R129 a_230_424.n4 a_230_424.n1 5.16973
R130 a_675_392.n8 a_675_392.n7 402.656
R131 a_675_392.n2 a_675_392.t5 269.945
R132 a_675_392.n1 a_675_392.t4 266.293
R133 a_675_392.n4 a_675_392.n3 216.172
R134 a_675_392.n2 a_675_392.t6 194.407
R135 a_675_392.n1 a_675_392.n0 194.407
R136 a_675_392.n7 a_675_392.n6 185
R137 a_675_392.n5 a_675_392.n4 185
R138 a_675_392.n8 a_675_392.t2 140.645
R139 a_675_392.n6 a_675_392.n5 104.287
R140 a_675_392.n3 a_675_392.n1 54.7732
R141 a_675_392.n5 a_675_392.t3 40.0005
R142 a_675_392.n6 a_675_392.t1 27.7237
R143 a_675_392.t0 a_675_392.n8 17.5044
R144 a_675_392.n7 a_675_392.n4 14.1581
R145 a_675_392.n3 a_675_392.n2 8.03383
R146 D.n0 D.t0 286.418
R147 D.n0 D.t1 160.832
R148 D D.n0 155.601
R149 a_27_115.t0 a_27_115.n1 478.693
R150 a_27_115.n1 a_27_115.n0 375.43
R151 a_27_115.n0 a_27_115.t2 298.572
R152 a_27_115.n1 a_27_115.t1 227.256
R153 a_27_115.n0 a_27_115.t3 217.192
R154 GATE_N.n0 GATE_N.t1 240.732
R155 GATE_N.n0 GATE_N.t0 204.048
R156 GATE_N GATE_N.n0 155.298
R157 VGND.n1 VGND.n0 288.024
R158 VGND.n9 VGND.t3 244.566
R159 VGND.n12 VGND.n11 227.24
R160 VGND.n8 VGND.n7 214.695
R161 VGND.n19 VGND.n18 116.674
R162 VGND.n18 VGND.t8 97.6196
R163 VGND.n0 VGND.t7 55.6369
R164 VGND.n11 VGND.t5 50.5809
R165 VGND.n11 VGND.t4 40.0005
R166 VGND.n16 VGND.n5 36.1417
R167 VGND.n17 VGND.n16 36.1417
R168 VGND.n23 VGND.n3 36.1417
R169 VGND.n24 VGND.n23 36.1417
R170 VGND.n25 VGND.n24 36.1417
R171 VGND.n19 VGND.n17 34.2593
R172 VGND.n18 VGND.t0 30.0005
R173 VGND.n12 VGND.n10 28.6123
R174 VGND.n0 VGND.t6 26.4679
R175 VGND.n12 VGND.n5 24.8476
R176 VGND.n7 VGND.t1 22.7032
R177 VGND.n7 VGND.t2 22.7032
R178 VGND.n25 VGND.n1 22.1206
R179 VGND.n10 VGND.n9 17.3181
R180 VGND.n19 VGND.n3 13.177
R181 VGND.n26 VGND.n25 9.3005
R182 VGND.n24 VGND.n2 9.3005
R183 VGND.n23 VGND.n22 9.3005
R184 VGND.n21 VGND.n3 9.3005
R185 VGND.n10 VGND.n6 9.3005
R186 VGND.n13 VGND.n12 9.3005
R187 VGND.n14 VGND.n5 9.3005
R188 VGND.n16 VGND.n15 9.3005
R189 VGND.n17 VGND.n4 9.3005
R190 VGND.n20 VGND.n19 9.3005
R191 VGND.n27 VGND.n1 9.10055
R192 VGND.n9 VGND.n8 7.08017
R193 VGND.n8 VGND.n6 0.490489
R194 VGND VGND.n27 0.161517
R195 VGND.n27 VGND.n26 0.146304
R196 VGND.n13 VGND.n6 0.122949
R197 VGND.n14 VGND.n13 0.122949
R198 VGND.n15 VGND.n14 0.122949
R199 VGND.n15 VGND.n4 0.122949
R200 VGND.n20 VGND.n4 0.122949
R201 VGND.n21 VGND.n20 0.122949
R202 VGND.n22 VGND.n21 0.122949
R203 VGND.n22 VGND.n2 0.122949
R204 VGND.n26 VGND.n2 0.122949
R205 VNB.t6 VNB.t9 2933.33
R206 VNB.t5 VNB.t4 2182.68
R207 VNB.t9 VNB.t0 1986.35
R208 VNB.t8 VNB.t10 1836.22
R209 VNB.t7 VNB.t6 1362.73
R210 VNB.t4 VNB.t2 1201.05
R211 VNB.t3 VNB.t5 1177.95
R212 VNB VNB.t7 1143.31
R213 VNB.t2 VNB.t1 993.177
R214 VNB.t0 VNB.t8 900.788
R215 VNB.t10 VNB.t3 831.496
R216 a_369_392.t0 a_369_392.n1 772.505
R217 a_369_392.n0 a_369_392.t3 401.034
R218 a_369_392.n0 a_369_392.t2 383.628
R219 a_369_392.n1 a_369_392.t1 256.087
R220 a_369_392.n1 a_369_392.n0 74.7356
R221 a_658_79.t0 a_658_79.t1 45.0005
R222 a_895_123.t0 a_895_123.t1 60.0005
R223 a_591_392.t0 a_591_392.t1 53.1905
C0 D GATE_N 0.041736f
C1 VPB VPWR 0.230753f
C2 D VPWR 0.018614f
C3 VPB VGND 0.016034f
C4 GATE_N VPWR 0.020999f
C5 D VGND 0.007731f
C6 VPB Q 0.016914f
C7 GATE_N VGND 0.007281f
C8 VPWR VGND 0.134687f
C9 VPWR Q 0.411291f
C10 VGND Q 0.306113f
C11 VPB D 0.066304f
C12 VPB GATE_N 0.064627f
C13 Q VNB 0.076423f
C14 VGND VNB 0.978057f
C15 VPWR VNB 0.761013f
C16 GATE_N VNB 0.099337f
C17 D VNB 0.180465f
C18 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxtn_2 VNB VPB VPWR VGND D GATE_N Q
X0 VPWR.t6 a_842_405.t2 Q.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1932 ps=1.465 w=1.12 l=0.15
X1 a_842_405.t0 a_669_392.t4 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.24815 ps=1.86 w=1.12 l=0.15
X2 a_875_139.t0 a_369_392.t2 a_669_392.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.14015 ps=1.265 w=0.42 l=0.15
X3 a_232_82.t0 GATE_N.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.168 ps=1.24 w=0.84 l=0.15
X4 a_232_82.t1 GATE_N.t1 VGND.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.189025 ps=1.41 w=0.74 l=0.15
X5 VGND.t4 a_232_82.t2 a_369_392.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2397 pd=1.45 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VPWR.t2 a_232_82.t3 a_369_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.255125 pd=1.615 as=0.2478 ps=2.27 w=0.84 l=0.15
X7 a_669_392.t3 a_232_82.t4 a_658_79.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.14015 pd=1.265 as=0.0768 ps=0.88 w=0.64 l=0.15
X8 a_842_405.t1 a_669_392.t5 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1212 ps=1.1 w=0.74 l=0.15
X9 VPWR.t5 a_842_405.t3 a_791_503.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.24815 pd=1.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR.t3 D.t0 a_27_120.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X11 a_669_392.t2 a_369_392.t3 a_585_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.202575 pd=1.46 as=0.135 ps=1.27 w=1 l=0.15
X12 a_791_503.t0 a_232_82.t5 a_669_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.202575 ps=1.46 w=0.42 l=0.15
X13 a_585_392.t1 a_27_120.t2 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.255125 ps=1.615 w=1 l=0.15
X14 Q.t1 a_842_405.t4 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 VGND.t0 D.t1 a_27_120.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.189025 pd=1.41 as=0.15675 ps=1.67 w=0.55 l=0.15
X16 a_658_79.t0 a_27_120.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2397 ps=1.45 w=0.64 l=0.15
X17 VGND.t5 a_842_405.t5 a_875_139.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_842_405.n6 a_842_405.t5 383.993
R1 a_842_405.n2 a_842_405.t2 243.833
R2 a_842_405.n3 a_842_405.n0 241.536
R3 a_842_405.t0 a_842_405.n7 222.964
R4 a_842_405.n7 a_842_405.n6 187.304
R5 a_842_405.n2 a_842_405.n1 178.34
R6 a_842_405.n4 a_842_405.t4 178.34
R7 a_842_405.n5 a_842_405.t1 167.865
R8 a_842_405.n6 a_842_405.t3 147.206
R9 a_842_405.n5 a_842_405.n4 112.691
R10 a_842_405.n3 a_842_405.n2 70.1096
R11 a_842_405.n7 a_842_405.n5 27.5166
R12 a_842_405.n4 a_842_405.n3 1.46111
R13 Q.n0 Q.t0 764.87
R14 Q Q.t1 205.745
R15 Q Q.n0 8.02183
R16 Q.n0 Q 4.6085
R17 VPWR.n17 VPWR.n4 671.601
R18 VPWR.n10 VPWR.n9 585
R19 VPWR.n8 VPWR.n7 585
R20 VPWR.n23 VPWR.n1 316.493
R21 VPWR.n6 VPWR.t6 266.873
R22 VPWR.n9 VPWR.n8 204.036
R23 VPWR.n9 VPWR.t5 70.3576
R24 VPWR.n4 VPWR.t2 66.8398
R25 VPWR.n8 VPWR.t4 48.7502
R26 VPWR.n1 VPWR.t0 46.9053
R27 VPWR.n1 VPWR.t3 46.9053
R28 VPWR.n4 VPWR.t1 36.7421
R29 VPWR.n21 VPWR.n2 36.1417
R30 VPWR.n22 VPWR.n21 36.1417
R31 VPWR.n15 VPWR.n5 36.1417
R32 VPWR.n16 VPWR.n15 36.1417
R33 VPWR.n17 VPWR.n16 31.2476
R34 VPWR.n10 VPWR.n5 23.7563
R35 VPWR.n17 VPWR.n2 15.0593
R36 VPWR.n24 VPWR.n23 11.092
R37 VPWR.n12 VPWR.n11 9.3005
R38 VPWR.n13 VPWR.n5 9.3005
R39 VPWR.n15 VPWR.n14 9.3005
R40 VPWR.n16 VPWR.n3 9.3005
R41 VPWR.n18 VPWR.n17 9.3005
R42 VPWR.n19 VPWR.n2 9.3005
R43 VPWR.n21 VPWR.n20 9.3005
R44 VPWR.n22 VPWR.n0 9.3005
R45 VPWR.n7 VPWR.n6 8.83746
R46 VPWR.n23 VPWR.n22 7.90638
R47 VPWR.n11 VPWR.n7 6.48151
R48 VPWR.n11 VPWR.n10 0.567589
R49 VPWR.n12 VPWR.n6 0.167537
R50 VPWR VPWR.n24 0.163644
R51 VPWR.n24 VPWR.n0 0.144205
R52 VPWR.n13 VPWR.n12 0.122949
R53 VPWR.n14 VPWR.n13 0.122949
R54 VPWR.n14 VPWR.n3 0.122949
R55 VPWR.n18 VPWR.n3 0.122949
R56 VPWR.n19 VPWR.n18 0.122949
R57 VPWR.n20 VPWR.n19 0.122949
R58 VPWR.n20 VPWR.n0 0.122949
R59 VPB.t6 VPB.t8 768.683
R60 VPB.t2 VPB.t4 515.861
R61 VPB.t7 VPB.t6 454.57
R62 VPB VPB.t5 334.543
R63 VPB.t4 VPB.t3 324.329
R64 VPB.t1 VPB.t0 311.56
R65 VPB.t5 VPB.t2 280.914
R66 VPB.t0 VPB.t7 214.517
R67 VPB.t3 VPB.t1 214.517
R68 a_669_392.n3 a_669_392.n2 388.351
R69 a_669_392.n0 a_669_392.t4 258.942
R70 a_669_392.n2 a_669_392.n0 249.608
R71 a_669_392.n0 a_669_392.t5 200.833
R72 a_669_392.n2 a_669_392.n1 185
R73 a_669_392.n3 a_669_392.t0 128.988
R74 a_669_392.n1 a_669_392.t1 78.7866
R75 a_669_392.n1 a_669_392.t3 74.6145
R76 a_669_392.n4 a_669_392.t2 23.8017
R77 a_669_392.n5 a_669_392.n4 16.7852
R78 a_669_392.n4 a_669_392.n3 11.8093
R79 a_369_392.t0 a_369_392.n1 777.297
R80 a_369_392.n0 a_369_392.t3 383.628
R81 a_369_392.n0 a_369_392.t2 383.38
R82 a_369_392.n1 a_369_392.t1 260.183
R83 a_369_392.n1 a_369_392.n0 75.5798
R84 a_875_139.t0 a_875_139.t1 68.5719
R85 VNB VNB.n0 10929.8
R86 VNB.t2 VNB.t8 2933.33
R87 VNB.t3 VNB.t7 2317.02
R88 VNB.t4 VNB.t2 1986.35
R89 VNB.t1 VNB.t5 1605.25
R90 VNB.t8 VNB.t0 1362.73
R91 VNB.t6 VNB.t3 1193.62
R92 VNB.t0 VNB 1143.31
R93 VNB.t5 VNB.t4 900.788
R94 VNB.n0 VNB.t1 854.593
R95 VNB.n0 VNB.t6 23.2502
R96 GATE_N.n0 GATE_N.t0 254.121
R97 GATE_N.n0 GATE_N.t1 239.393
R98 GATE_N GATE_N.n0 153.358
R99 a_232_82.t0 a_232_82.n1 778.163
R100 a_232_82.t0 a_232_82.n4 768.644
R101 a_232_82.n1 a_232_82.n0 491.702
R102 a_232_82.n2 a_232_82.t3 306.339
R103 a_232_82.n3 a_232_82.t1 297.082
R104 a_232_82.n0 a_232_82.t4 277.954
R105 a_232_82.n0 a_232_82.t5 258.942
R106 a_232_82.n2 a_232_82.t2 187.981
R107 a_232_82.n3 a_232_82.n2 163.709
R108 a_232_82.n4 a_232_82.n3 44.8231
R109 a_232_82.n4 a_232_82.n1 8.53383
R110 VGND.n1 VGND.n0 242.279
R111 VGND.n9 VGND.n6 199.546
R112 VGND.n9 VGND.n8 185
R113 VGND.n11 VGND.t6 172.115
R114 VGND.n17 VGND.n16 116.719
R115 VGND.n16 VGND.t4 97.6196
R116 VGND.n7 VGND.t5 61.4291
R117 VGND.n0 VGND.t0 55.6369
R118 VGND.n8 VGND.t2 52.5005
R119 VGND.t2 VGND.n6 40.0005
R120 VGND.n14 VGND.n5 36.1417
R121 VGND.n15 VGND.n14 36.1417
R122 VGND.n21 VGND.n3 36.1417
R123 VGND.n22 VGND.n21 36.1417
R124 VGND.n23 VGND.n22 36.1417
R125 VGND.n17 VGND.n15 34.2593
R126 VGND.n0 VGND.t1 30.0005
R127 VGND.n16 VGND.t3 30.0005
R128 VGND.n23 VGND.n1 22.7142
R129 VGND.n10 VGND.n9 19.9763
R130 VGND.n10 VGND.n5 19.577
R131 VGND.n17 VGND.n3 13.177
R132 VGND.n25 VGND.n1 9.36437
R133 VGND.n24 VGND.n23 9.3005
R134 VGND.n22 VGND.n2 9.3005
R135 VGND.n21 VGND.n20 9.3005
R136 VGND.n19 VGND.n3 9.3005
R137 VGND.n12 VGND.n5 9.3005
R138 VGND.n14 VGND.n13 9.3005
R139 VGND.n15 VGND.n4 9.3005
R140 VGND.n18 VGND.n17 9.3005
R141 VGND.n11 VGND.n10 6.98251
R142 VGND.n8 VGND.n7 1.8755
R143 VGND.n7 VGND.n6 1.42907
R144 VGND.n12 VGND.n11 0.497471
R145 VGND VGND.n25 0.161675
R146 VGND.n25 VGND.n24 0.146149
R147 VGND.n13 VGND.n12 0.122949
R148 VGND.n13 VGND.n4 0.122949
R149 VGND.n18 VGND.n4 0.122949
R150 VGND.n19 VGND.n18 0.122949
R151 VGND.n20 VGND.n19 0.122949
R152 VGND.n20 VGND.n2 0.122949
R153 VGND.n24 VGND.n2 0.122949
R154 a_658_79.t0 a_658_79.t1 45.0005
R155 a_791_503.t0 a_791_503.t1 126.644
R156 D.n0 D.t0 293.558
R157 D D.n0 185.542
R158 D.n0 D.t1 136.567
R159 a_27_120.t1 a_27_120.n1 468.906
R160 a_27_120.n1 a_27_120.n0 373.928
R161 a_27_120.n0 a_27_120.t2 277.151
R162 a_27_120.n0 a_27_120.t3 259.697
R163 a_27_120.n1 a_27_120.t0 225.554
R164 a_585_392.t0 a_585_392.t1 53.1905
C0 VPB D 0.075811f
C1 VPB Q 0.007274f
C2 VPB GATE_N 0.06251f
C3 VPB VPWR 0.22747f
C4 D GATE_N 0.056171f
C5 VPB VGND 0.018883f
C6 D VPWR 0.017872f
C7 VPWR Q 0.19816f
C8 GATE_N VPWR 0.023641f
C9 D VGND 0.006362f
C10 VGND Q 0.161284f
C11 GATE_N VGND 0.00984f
C12 VPWR VGND 0.129507f
C13 Q VNB 0.030256f
C14 VGND VNB 0.901164f
C15 VPWR VNB 0.718043f
C16 GATE_N VNB 0.107927f
C17 D VNB 0.18737f
C18 VPB VNB 1.69507f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlymetal6s4s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlymetal6s4s_1 VNB VPB VPWR VGND X A
X0 VPWR.t4 X.t2 a_604_138.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1757 pd=1.49 as=0.1155 ps=1.39 w=0.42 l=0.15
X1 a_209_74.t0 a_28_138.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1729 ps=1.485 w=1.12 l=0.15
X2 a_209_74.t1 a_28_138.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X3 VGND.t2 a_209_74.t2 a_316_138.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VGND.t4 X.t3 a_604_138.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VPWR.t2 A.t0 a_28_138.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.1155 ps=1.39 w=0.42 l=0.15
X6 X.t0 a_316_138.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X7 a_785_74.t0 a_604_138.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X8 VPWR.t0 a_209_74.t3 a_316_138.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.1155 ps=1.39 w=0.42 l=0.15
X9 a_785_74.t1 a_604_138.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1757 ps=1.49 w=1.12 l=0.15
X10 VGND.t1 A.t1 a_28_138.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 X.t1 a_316_138.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1729 ps=1.485 w=1.12 l=0.15
R0 X.n2 X.t1 230.347
R1 X.n1 X.n0 173.629
R2 X.n1 X.t0 158.536
R3 X.n0 X.t2 152.297
R4 X.n0 X.t3 138.373
R5 X.n2 X.n1 23.9942
R6 X.n3 X.n2 9.73488
R7 X.n3 X 1.37053
R8 X.n4 X 1.05932
R9 X X.n4 0.316289
R10 X.n4 X.n3 0.0520351
R11 a_604_138.n1 a_604_138.t0 701.467
R12 a_604_138.t1 a_604_138.n1 282.86
R13 a_604_138.n0 a_604_138.t3 270.991
R14 a_604_138.n0 a_604_138.t2 193.385
R15 a_604_138.n1 a_604_138.n0 152
R16 VPWR.n5 VPWR.n4 328.675
R17 VPWR.n3 VPWR.n2 321.303
R18 VPWR.n9 VPWR.n1 321.303
R19 VPWR.n4 VPWR.t4 107.882
R20 VPWR.n1 VPWR.t2 105.537
R21 VPWR.n2 VPWR.t0 105.537
R22 VPWR.n8 VPWR.n7 36.1417
R23 VPWR.n7 VPWR.n3 31.624
R24 VPWR.n1 VPWR.t3 24.6255
R25 VPWR.n2 VPWR.t1 24.6255
R26 VPWR.n4 VPWR.t5 24.6255
R27 VPWR.n9 VPWR.n8 23.7181
R28 VPWR.n7 VPWR.n6 9.3005
R29 VPWR.n8 VPWR.n0 9.3005
R30 VPWR.n10 VPWR.n9 7.35695
R31 VPWR.n5 VPWR.n3 6.7737
R32 VPWR.n6 VPWR.n5 0.217413
R33 VPWR VPWR.n10 0.159077
R34 VPWR.n10 VPWR.n0 0.148713
R35 VPWR.n6 VPWR.n0 0.122949
R36 VPB.t1 VPB.t4 495.43
R37 VPB.t3 VPB.t0 495.43
R38 VPB.t4 VPB.t5 265.591
R39 VPB.t0 VPB.t1 263.038
R40 VPB.t2 VPB.t3 263.038
R41 VPB VPB.t2 250.269
R42 a_28_138.n1 a_28_138.t1 717.919
R43 a_28_138.t0 a_28_138.n1 281.202
R44 a_28_138.n0 a_28_138.t2 270.991
R45 a_28_138.n0 a_28_138.t3 193.385
R46 a_28_138.n1 a_28_138.n0 152
R47 a_209_74.t0 a_209_74.n1 255.185
R48 a_209_74.n1 a_209_74.n0 175.614
R49 a_209_74.n1 a_209_74.t1 159.993
R50 a_209_74.n0 a_209_74.t3 154.308
R51 a_209_74.n0 a_209_74.t2 140.383
R52 VGND.n4 VGND.n3 218.977
R53 VGND.n2 VGND.n1 212.928
R54 VGND.n9 VGND.n8 212.928
R55 VGND.n3 VGND.t4 57.1434
R56 VGND.n1 VGND.t2 57.1434
R57 VGND.n8 VGND.t1 57.1434
R58 VGND.n7 VGND.n6 36.1417
R59 VGND.n6 VGND.n2 26.3534
R60 VGND.n3 VGND.t5 23.321
R61 VGND.n1 VGND.t0 23.321
R62 VGND.n8 VGND.t3 23.321
R63 VGND.n9 VGND.n7 21.0829
R64 VGND.n6 VGND.n5 9.3005
R65 VGND.n7 VGND.n0 9.3005
R66 VGND.n10 VGND.n9 7.35695
R67 VGND.n4 VGND.n2 6.93311
R68 VGND.n5 VGND.n4 0.22537
R69 VGND VGND.n10 0.159077
R70 VGND.n10 VGND.n0 0.148713
R71 VGND.n5 VGND.n0 0.122949
R72 VNB.t0 VNB.t4 2194.23
R73 VNB.t3 VNB.t2 2194.23
R74 VNB.t4 VNB.t5 1131.76
R75 VNB.t2 VNB.t0 1131.76
R76 VNB.t1 VNB.t3 1131.76
R77 VNB VNB.t1 1108.66
R78 a_316_138.n1 a_316_138.t1 707.567
R79 a_316_138.t0 a_316_138.n1 280.661
R80 a_316_138.n0 a_316_138.t3 270.991
R81 a_316_138.n0 a_316_138.t2 193.385
R82 a_316_138.n1 a_316_138.n0 152
R83 A A.n0 159.18
R84 A.n0 A.t0 156.827
R85 A.n0 A.t1 142.904
R86 a_785_74.t1 a_785_74.t0 433.267
C0 VPB A 0.042383f
C1 VPWR A 0.005539f
C2 VPB X 0.101527f
C3 VPB VGND 0.014614f
C4 VPWR X 0.359489f
C5 A X 6.41e-19
C6 VPWR VGND 0.029794f
C7 A VGND 0.01019f
C8 X VGND 0.176468f
C9 VPB VPWR 0.190004f
C10 VGND VNB 0.63349f
C11 X VNB 0.17277f
C12 A VNB 0.155573f
C13 VPWR VNB 0.488651f
C14 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlymetal6s2s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlymetal6s2s_1 VNB VPB VPWR VGND X A
X0 VPWR.t2 a_497_74.t2 a_604_138.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1757 pd=1.49 as=0.1155 ps=1.39 w=0.42 l=0.15
X1 X.t0 a_28_138.t2 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1729 ps=1.485 w=1.12 l=0.15
X2 X.t1 a_28_138.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X3 VGND.t5 X.t2 a_316_138.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VGND.t1 a_497_74.t3 a_604_138.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VPWR.t0 A.t0 a_28_138.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.1155 ps=1.39 w=0.42 l=0.15
X6 a_497_74.t1 a_316_138.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X7 a_785_74.t1 a_604_138.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X8 VPWR.t1 X.t3 a_316_138.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.1155 ps=1.39 w=0.42 l=0.15
X9 a_785_74.t0 a_604_138.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1757 ps=1.49 w=1.12 l=0.15
X10 VGND.t4 A.t1 a_28_138.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 a_497_74.t0 a_316_138.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1729 ps=1.485 w=1.12 l=0.15
R0 a_497_74.t0 a_497_74.n1 254.341
R1 a_497_74.n1 a_497_74.n0 173.629
R2 a_497_74.n1 a_497_74.t1 158.536
R3 a_497_74.n0 a_497_74.t2 152.297
R4 a_497_74.n0 a_497_74.t3 138.373
R5 a_604_138.n1 a_604_138.t1 701.467
R6 a_604_138.t0 a_604_138.n1 282.86
R7 a_604_138.n0 a_604_138.t3 270.991
R8 a_604_138.n0 a_604_138.t2 193.385
R9 a_604_138.n1 a_604_138.n0 152
R10 VPWR.n5 VPWR.n4 328.675
R11 VPWR.n3 VPWR.n2 321.303
R12 VPWR.n9 VPWR.n1 321.303
R13 VPWR.n4 VPWR.t2 107.882
R14 VPWR.n1 VPWR.t0 105.537
R15 VPWR.n2 VPWR.t1 105.537
R16 VPWR.n8 VPWR.n7 36.1417
R17 VPWR.n7 VPWR.n3 31.624
R18 VPWR.n1 VPWR.t5 24.6255
R19 VPWR.n2 VPWR.t3 24.6255
R20 VPWR.n4 VPWR.t4 24.6255
R21 VPWR.n9 VPWR.n8 23.7181
R22 VPWR.n7 VPWR.n6 9.3005
R23 VPWR.n8 VPWR.n0 9.3005
R24 VPWR.n10 VPWR.n9 7.35695
R25 VPWR.n5 VPWR.n3 6.7737
R26 VPWR.n6 VPWR.n5 0.217413
R27 VPWR VPWR.n10 0.159077
R28 VPWR.n10 VPWR.n0 0.148713
R29 VPWR.n6 VPWR.n0 0.122949
R30 VPB.t3 VPB.t2 495.43
R31 VPB.t5 VPB.t1 495.43
R32 VPB.t2 VPB.t4 265.591
R33 VPB.t1 VPB.t3 263.038
R34 VPB.t0 VPB.t5 263.038
R35 VPB VPB.t0 250.269
R36 a_28_138.n1 a_28_138.t0 717.919
R37 a_28_138.t1 a_28_138.n1 281.202
R38 a_28_138.n0 a_28_138.t2 270.991
R39 a_28_138.n0 a_28_138.t3 193.385
R40 a_28_138.n1 a_28_138.n0 152
R41 X.n2 X.t0 230.238
R42 X.n1 X.n0 175.614
R43 X.n1 X.t1 159.993
R44 X.n0 X.t3 154.308
R45 X.n0 X.t2 140.383
R46 X.n2 X.n1 24.9478
R47 X.n3 X.n2 9.79659
R48 X X.n3 0.31171
R49 X.n3 X 0.0520351
R50 VGND.n4 VGND.n3 218.977
R51 VGND.n2 VGND.n1 212.928
R52 VGND.n9 VGND.n8 212.928
R53 VGND.n3 VGND.t1 57.1434
R54 VGND.n1 VGND.t5 57.1434
R55 VGND.n8 VGND.t4 57.1434
R56 VGND.n7 VGND.n6 36.1417
R57 VGND.n6 VGND.n2 26.3534
R58 VGND.n3 VGND.t2 23.321
R59 VGND.n1 VGND.t3 23.321
R60 VGND.n8 VGND.t0 23.321
R61 VGND.n9 VGND.n7 21.0829
R62 VGND.n6 VGND.n5 9.3005
R63 VGND.n7 VGND.n0 9.3005
R64 VGND.n10 VGND.n9 7.35695
R65 VGND.n4 VGND.n2 6.93311
R66 VGND.n5 VGND.n4 0.22537
R67 VGND VGND.n10 0.159077
R68 VGND.n10 VGND.n0 0.148713
R69 VGND.n5 VGND.n0 0.122949
R70 VNB.t3 VNB.t1 2194.23
R71 VNB.t0 VNB.t5 2194.23
R72 VNB.t1 VNB.t2 1131.76
R73 VNB.t5 VNB.t3 1131.76
R74 VNB.t4 VNB.t0 1131.76
R75 VNB VNB.t4 1108.66
R76 a_316_138.n1 a_316_138.t0 707.567
R77 a_316_138.t1 a_316_138.n1 280.661
R78 a_316_138.n0 a_316_138.t3 270.991
R79 a_316_138.n0 a_316_138.t2 193.385
R80 a_316_138.n1 a_316_138.n0 152
R81 A A.n0 159.18
R82 A.n0 A.t0 156.827
R83 A.n0 A.t1 142.904
R84 a_785_74.t0 a_785_74.t1 433.267
C0 VPB VPWR 0.190004f
C1 VPB A 0.042383f
C2 VPWR A 0.005539f
C3 VPB X 0.098601f
C4 VPWR X 0.357365f
C5 VPB VGND 0.014614f
C6 A X 0.006645f
C7 VPWR VGND 0.029794f
C8 A VGND 0.01019f
C9 X VGND 0.169016f
C10 VGND VNB 0.63349f
C11 X VNB 0.17413f
C12 A VNB 0.155573f
C13 VPWR VNB 0.488651f
C14 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlygate4sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlygate4sd3_1 VNB VPB VPWR VGND A X
X0 a_289_74.t0 a_28_74.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1092 pd=1.36 as=0.1491 ps=1.13 w=0.42 l=0.18
X1 VPWR.t2 A.t0 a_28_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15125 pd=1.375 as=0.1176 ps=1.4 w=0.42 l=0.15
X2 X.t0 a_405_138.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.11485 ps=1.085 w=0.74 l=0.15
X3 VPWR.t3 a_289_74.t2 a_405_138.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.475 as=0.26 ps=2.52 w=1 l=0.5
X4 VGND.t3 A.t1 a_28_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.13 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VGND.t2 a_289_74.t3 a_405_138.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.11485 pd=1.085 as=0.2436 ps=2 w=0.42 l=0.18
X6 X.t1 a_405_138.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.194 ps=1.475 w=1.12 l=0.15
X7 a_289_74.t1 a_28_74.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.15125 ps=1.375 w=1 l=0.5
R0 a_28_74.n0 a_28_74.t0 737.053
R1 a_28_74.t1 a_28_74.n3 289.522
R2 a_28_74.n2 a_28_74.t2 163.185
R3 a_28_74.n1 a_28_74.n0 152
R4 a_28_74.n3 a_28_74.n2 152
R5 a_28_74.n1 a_28_74.t3 79.5305
R6 a_28_74.n2 a_28_74.n1 32.7765
R7 a_28_74.n3 a_28_74.n0 13.1884
R8 VGND.n2 VGND.n0 217.103
R9 VGND.n2 VGND.n1 212.748
R10 VGND.n1 VGND.t0 147.143
R11 VGND.n0 VGND.t2 60.0005
R12 VGND.n1 VGND.t3 55.7148
R13 VGND.n0 VGND.t1 21.8924
R14 VGND VGND.n2 0.196947
R15 a_289_74.n1 a_289_74.t1 665.54
R16 a_289_74.t0 a_289_74.n1 270.81
R17 a_289_74.n0 a_289_74.t3 123.017
R18 a_289_74.n1 a_289_74.n0 111.117
R19 a_289_74.n0 a_289_74.t2 84.3505
R20 VNB.t0 VNB.t2 3095.01
R21 VNB.t3 VNB.t0 2021
R22 VNB.t2 VNB.t1 1177.95
R23 VNB VNB.t3 1108.66
R24 A.n0 A.t0 313.837
R25 A.n0 A.t1 220.113
R26 A A.n0 159.929
R27 VPWR.n2 VPWR.n1 621.289
R28 VPWR.n2 VPWR.n0 323.997
R29 VPWR.n1 VPWR.t2 79.7386
R30 VPWR.n1 VPWR.t1 64.8571
R31 VPWR.n0 VPWR.t3 40.3855
R32 VPWR.n0 VPWR.t0 27.3314
R33 VPWR VPWR.n2 0.195508
R34 VPB.t1 VPB.t3 684.409
R35 VPB.t2 VPB.t1 357.527
R36 VPB.t3 VPB.t0 347.312
R37 VPB VPB.t2 252.823
R38 a_405_138.n1 a_405_138.t1 893.652
R39 a_405_138.t0 a_405_138.n1 381.021
R40 a_405_138.n0 a_405_138.t3 265.637
R41 a_405_138.n0 a_405_138.t2 202.44
R42 a_405_138.n1 a_405_138.n0 152
R43 X.n1 X 588.702
R44 X.n1 X.n0 585
R45 X.n2 X.n1 585
R46 X.t0 X.n3 284.623
R47 X.n4 X.t0 282.358
R48 X.n1 X.t1 27.2639
R49 X.n2 X 10.333
R50 X.n3 X 9.87038
R51 X X.n4 9.06207
R52 X.n0 X 8.01978
R53 X.n4 X 3.54749
R54 X.n0 X 3.39327
R55 X.n3 X 1.54267
R56 X X.n2 1.08002
C0 VPB A 0.090912f
C1 VPB VPWR 0.123898f
C2 VPB VGND 0.009448f
C3 VPB X 0.020957f
C4 A VPWR 0.01616f
C5 A VGND 0.017398f
C6 A X 1.81e-19
C7 VPWR VGND 0.062419f
C8 VPWR X 0.134114f
C9 X VGND 0.092359f
C10 VGND VNB 0.50594f
C11 X VNB 0.119844f
C12 VPWR VNB 0.397646f
C13 A VNB 0.218416f
C14 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlygate4sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlygate4sd2_1 VNB VPB VPWR VGND A X
X0 VPWR.t2 A.t0 a_28_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.27625 pd=1.625 as=0.1176 ps=1.4 w=0.42 l=0.15
X1 a_288_74.t0 a_28_74.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X2 X.t0 a_405_138.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.11485 ps=1.085 w=0.74 l=0.15
X3 VPWR.t1 a_288_74.t2 a_405_138.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.475 as=0.51 ps=3.02 w=1 l=0.25
X4 VGND.t2 A.t1 a_28_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VGND.t1 a_288_74.t3 a_405_138.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.11485 pd=1.085 as=0.2436 ps=2 w=0.42 l=0.18
X6 X.t1 a_405_138.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.194 ps=1.475 w=1.12 l=0.15
X7 a_288_74.t1 a_28_74.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.27625 ps=1.625 w=1 l=0.25
R0 A.n0 A.t0 313.837
R1 A.n0 A.t1 220.113
R2 A A.n0 159.929
R3 a_28_74.n0 a_28_74.t0 737.053
R4 a_28_74.t1 a_28_74.n3 289.522
R5 a_28_74.n2 a_28_74.t2 163.185
R6 a_28_74.n1 a_28_74.n0 152
R7 a_28_74.n3 a_28_74.n2 152
R8 a_28_74.n1 a_28_74.t3 143.155
R9 a_28_74.n2 a_28_74.n1 32.7765
R10 a_28_74.n3 a_28_74.n0 13.1884
R11 VPWR.n2 VPWR.n1 621.289
R12 VPWR.n2 VPWR.n0 323.997
R13 VPWR.n1 VPWR.t3 89.6355
R14 VPWR.n1 VPWR.t2 67.4965
R15 VPWR.n0 VPWR.t1 40.3855
R16 VPWR.n0 VPWR.t0 27.3314
R17 VPWR VPWR.n2 0.195508
R18 VPB.t3 VPB.t1 684.409
R19 VPB.t2 VPB.t3 421.372
R20 VPB.t1 VPB.t0 283.469
R21 VPB VPB.t2 252.823
R22 VGND.n2 VGND.n0 217.103
R23 VGND.n2 VGND.n1 212.748
R24 VGND.n1 VGND.t3 145.714
R25 VGND.n0 VGND.t1 60.0005
R26 VGND.n1 VGND.t2 55.7148
R27 VGND.n0 VGND.t0 21.8924
R28 VGND VGND.n2 0.196947
R29 a_288_74.t1 a_288_74.n1 665.54
R30 a_288_74.n1 a_288_74.t0 272.24
R31 a_288_74.n0 a_288_74.t2 136.888
R32 a_288_74.n1 a_288_74.n0 133.589
R33 a_288_74.n0 a_288_74.t3 112.224
R34 VNB.t3 VNB.t0 3106.56
R35 VNB.t2 VNB.t3 2009.45
R36 VNB.t0 VNB.t1 1177.95
R37 VNB VNB.t2 1108.66
R38 a_405_138.t1 a_405_138.n1 730.823
R39 a_405_138.n1 a_405_138.t0 381.021
R40 a_405_138.n0 a_405_138.t3 265.637
R41 a_405_138.n0 a_405_138.t2 202.44
R42 a_405_138.n1 a_405_138.n0 152
R43 X.n1 X 588.702
R44 X.n1 X.n0 585
R45 X.n2 X.n1 585
R46 X.t0 X.n3 284.623
R47 X.n4 X.t0 282.358
R48 X.n1 X.t1 27.2639
R49 X.n2 X 10.333
R50 X.n3 X 9.87038
R51 X X.n4 9.06207
R52 X.n0 X 8.01978
R53 X.n4 X 3.54749
R54 X.n0 X 3.39327
R55 X.n3 X 1.54267
R56 X X.n2 1.08002
C0 VPB VGND 0.010116f
C1 A X 1.81e-19
C2 A VGND 0.017398f
C3 VPWR X 0.134114f
C4 VPWR VGND 0.06344f
C5 X VGND 0.092359f
C6 VPB A 0.092465f
C7 VPB VPWR 0.127881f
C8 A VPWR 0.01616f
C9 VPB X 0.020957f
C10 VGND VNB 0.506019f
C11 X VNB 0.119844f
C12 VPWR VNB 0.397096f
C13 A VNB 0.218363f
C14 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlymetal6s6s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlymetal6s6s_1 VNB VPB VPWR VGND X A
X0 VPWR.t3 a_497_74.t2 a_604_138.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1757 pd=1.49 as=0.1155 ps=1.39 w=0.42 l=0.15
X1 a_209_74.t1 a_28_138.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1729 ps=1.485 w=1.12 l=0.15
X2 a_209_74.t0 a_28_138.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X3 VGND.t3 a_209_74.t2 a_316_138.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VGND.t2 a_497_74.t3 a_604_138.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VPWR.t1 A.t0 a_28_138.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.1155 ps=1.39 w=0.42 l=0.15
X6 a_497_74.t1 a_316_138.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X7 X.t0 a_604_138.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1138 ps=1.08 w=0.74 l=0.15
X8 VPWR.t4 a_209_74.t3 a_316_138.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.1155 ps=1.39 w=0.42 l=0.15
X9 X.t1 a_604_138.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1757 ps=1.49 w=1.12 l=0.15
X10 VGND.t0 A.t1 a_28_138.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 a_497_74.t0 a_316_138.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1729 ps=1.485 w=1.12 l=0.15
R0 a_497_74.t0 a_497_74.n1 254.341
R1 a_497_74.n1 a_497_74.n0 173.629
R2 a_497_74.n1 a_497_74.t1 158.536
R3 a_497_74.n0 a_497_74.t2 152.297
R4 a_497_74.n0 a_497_74.t3 138.373
R5 a_604_138.n1 a_604_138.t1 701.467
R6 a_604_138.t0 a_604_138.n1 282.86
R7 a_604_138.n0 a_604_138.t3 270.991
R8 a_604_138.n0 a_604_138.t2 193.385
R9 a_604_138.n1 a_604_138.n0 152
R10 VPWR.n5 VPWR.n4 328.675
R11 VPWR.n3 VPWR.n2 321.303
R12 VPWR.n9 VPWR.n1 321.303
R13 VPWR.n4 VPWR.t3 107.882
R14 VPWR.n1 VPWR.t1 105.537
R15 VPWR.n2 VPWR.t4 105.537
R16 VPWR.n8 VPWR.n7 36.1417
R17 VPWR.n7 VPWR.n3 31.624
R18 VPWR.n1 VPWR.t2 24.6255
R19 VPWR.n2 VPWR.t0 24.6255
R20 VPWR.n4 VPWR.t5 24.6255
R21 VPWR.n9 VPWR.n8 23.7181
R22 VPWR.n7 VPWR.n6 9.3005
R23 VPWR.n8 VPWR.n0 9.3005
R24 VPWR.n10 VPWR.n9 7.35695
R25 VPWR.n5 VPWR.n3 6.7737
R26 VPWR.n6 VPWR.n5 0.217413
R27 VPWR VPWR.n10 0.159077
R28 VPWR.n10 VPWR.n0 0.148713
R29 VPWR.n6 VPWR.n0 0.122949
R30 VPB.t0 VPB.t3 495.43
R31 VPB.t2 VPB.t4 495.43
R32 VPB.t3 VPB.t5 265.591
R33 VPB.t4 VPB.t0 263.038
R34 VPB.t1 VPB.t2 263.038
R35 VPB VPB.t1 250.269
R36 a_28_138.n1 a_28_138.t0 717.919
R37 a_28_138.t1 a_28_138.n1 281.202
R38 a_28_138.n0 a_28_138.t2 270.991
R39 a_28_138.n0 a_28_138.t3 193.385
R40 a_28_138.n1 a_28_138.n0 152
R41 a_209_74.t1 a_209_74.n1 255.185
R42 a_209_74.n1 a_209_74.n0 175.614
R43 a_209_74.n1 a_209_74.t0 159.993
R44 a_209_74.n0 a_209_74.t3 154.308
R45 a_209_74.n0 a_209_74.t2 140.383
R46 VGND.n4 VGND.n3 218.977
R47 VGND.n2 VGND.n1 212.928
R48 VGND.n9 VGND.n8 212.928
R49 VGND.n3 VGND.t2 57.1434
R50 VGND.n1 VGND.t3 57.1434
R51 VGND.n8 VGND.t0 57.1434
R52 VGND.n7 VGND.n6 36.1417
R53 VGND.n6 VGND.n2 26.3534
R54 VGND.n3 VGND.t5 23.321
R55 VGND.n1 VGND.t4 23.321
R56 VGND.n8 VGND.t1 23.321
R57 VGND.n9 VGND.n7 21.0829
R58 VGND.n6 VGND.n5 9.3005
R59 VGND.n7 VGND.n0 9.3005
R60 VGND.n10 VGND.n9 7.35695
R61 VGND.n4 VGND.n2 6.93311
R62 VGND.n5 VGND.n4 0.22537
R63 VGND VGND.n10 0.159077
R64 VGND.n10 VGND.n0 0.148713
R65 VGND.n5 VGND.n0 0.122949
R66 VNB.t4 VNB.t2 2194.23
R67 VNB.t1 VNB.t3 2194.23
R68 VNB.t2 VNB.t5 1131.76
R69 VNB.t3 VNB.t4 1131.76
R70 VNB.t0 VNB.t1 1131.76
R71 VNB VNB.t0 1108.66
R72 a_316_138.n1 a_316_138.t1 707.567
R73 a_316_138.t0 a_316_138.n1 280.661
R74 a_316_138.n0 a_316_138.t3 270.991
R75 a_316_138.n0 a_316_138.t2 193.385
R76 a_316_138.n1 a_316_138.n0 152
R77 A A.n0 159.18
R78 A.n0 A.t0 156.827
R79 A.n0 A.t1 142.904
R80 X.n0 X.t1 230.284
R81 X.n0 X.t0 202.984
R82 X.n1 X.n0 9.76893
R83 X.n1 X 2.11815
R84 X X.n1 0.632079
C0 VPB VPWR 0.190004f
C1 VPB A 0.042383f
C2 VPB X 0.053653f
C3 VPWR A 0.005539f
C4 VPB VGND 0.014614f
C5 VPWR X 0.334303f
C6 A X 5.4e-19
C7 VPWR VGND 0.029794f
C8 A VGND 0.01019f
C9 X VGND 0.152076f
C10 VGND VNB 0.63349f
C11 X VNB 0.142888f
C12 A VNB 0.155573f
C13 VPWR VNB 0.488651f
C14 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlxtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxtn_1 VNB VPB VPWR VGND Q GATE_N D
X0 VPWR.t4 a_863_441.t2 a_812_508.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.22205 pd=1.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 Q.t0 a_863_441.t3 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_655_79.t1 a_27_115.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2349 ps=1.435 w=0.64 l=0.15
X3 a_812_508.t0 a_217_419.t2 a_669_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.2564 ps=1.565 w=0.42 l=0.15
X4 a_217_419.t0 GATE_N.t0 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.44 as=0.147 ps=1.19 w=0.84 l=0.15
X5 VGND.t3 a_863_441.t4 a_871_139.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.11745 pd=1.05 as=0.0504 ps=0.66 w=0.42 l=0.15
X6 a_863_441.t0 a_669_392.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.11745 ps=1.05 w=0.64 l=0.15
X7 a_217_419.t1 GATE_N.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.201575 ps=1.57 w=0.74 l=0.15
X8 a_863_441.t1 a_669_392.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.22205 ps=1.65 w=1 l=0.15
X9 VGND.t1 a_217_419.t3 a_369_392.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2349 pd=1.435 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 VPWR.t2 a_217_419.t4 a_369_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.255125 pd=1.615 as=0.2478 ps=2.27 w=0.84 l=0.15
X11 a_871_139.t1 a_369_392.t2 a_669_392.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1393 ps=1.26 w=0.42 l=0.15
X12 a_669_392.t0 a_217_419.t5 a_655_79.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1393 pd=1.26 as=0.0768 ps=0.88 w=0.64 l=0.15
X13 a_669_392.t2 a_369_392.t3 a_585_392.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2564 pd=1.565 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t5 D.t0 a_27_115.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X15 a_585_392.t0 a_27_115.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.255125 ps=1.615 w=1 l=0.15
X16 VGND.t5 D.t1 a_27_115.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.201575 pd=1.57 as=0.15675 ps=1.67 w=0.55 l=0.15
R0 a_863_441.n3 a_863_441.t4 379.776
R1 a_863_441.n1 a_863_441.t3 241.804
R2 a_863_441.t1 a_863_441.n4 229.077
R3 a_863_441.n2 a_863_441.n1 223.608
R4 a_863_441.n4 a_863_441.n3 182.238
R5 a_863_441.n1 a_863_441.n0 181.368
R6 a_863_441.n2 a_863_441.t0 155.599
R7 a_863_441.n3 a_863_441.t2 141.09
R8 a_863_441.n4 a_863_441.n2 35.8671
R9 a_812_508.t0 a_812_508.t1 126.644
R10 VPWR.n17 VPWR.n4 671.601
R11 VPWR.n10 VPWR.n9 585
R12 VPWR.n8 VPWR.n7 585
R13 VPWR.n23 VPWR.n1 318.683
R14 VPWR.n6 VPWR.t3 265.072
R15 VPWR.n9 VPWR.n8 161.821
R16 VPWR.n9 VPWR.t4 72.7029
R17 VPWR.n4 VPWR.t2 66.8398
R18 VPWR.n1 VPWR.t5 46.9053
R19 VPWR.n4 VPWR.t0 36.7421
R20 VPWR.n21 VPWR.n2 36.1417
R21 VPWR.n22 VPWR.n21 36.1417
R22 VPWR.n15 VPWR.n5 36.1417
R23 VPWR.n16 VPWR.n15 36.1417
R24 VPWR.n1 VPWR.t6 35.1791
R25 VPWR.n17 VPWR.n16 31.2476
R26 VPWR.n11 VPWR.n5 30.6596
R27 VPWR.n8 VPWR.t1 29.5505
R28 VPWR.n23 VPWR.n22 18.824
R29 VPWR.n17 VPWR.n2 15.0593
R30 VPWR.n12 VPWR.n11 9.3005
R31 VPWR.n13 VPWR.n5 9.3005
R32 VPWR.n15 VPWR.n14 9.3005
R33 VPWR.n16 VPWR.n3 9.3005
R34 VPWR.n18 VPWR.n17 9.3005
R35 VPWR.n19 VPWR.n2 9.3005
R36 VPWR.n21 VPWR.n20 9.3005
R37 VPWR.n22 VPWR.n0 9.3005
R38 VPWR.n7 VPWR.n6 8.12709
R39 VPWR.n24 VPWR.n23 7.44972
R40 VPWR.n10 VPWR.n7 4.9623
R41 VPWR.n11 VPWR.n10 1.07915
R42 VPWR.n12 VPWR.n6 0.470223
R43 VPWR VPWR.n24 0.160299
R44 VPWR.n24 VPWR.n0 0.147507
R45 VPWR.n13 VPWR.n12 0.122949
R46 VPWR.n14 VPWR.n13 0.122949
R47 VPWR.n14 VPWR.n3 0.122949
R48 VPWR.n18 VPWR.n3 0.122949
R49 VPWR.n19 VPWR.n18 0.122949
R50 VPWR.n20 VPWR.n19 0.122949
R51 VPWR.n20 VPWR.n0 0.122949
R52 VPB.t7 VPB.t3 615.457
R53 VPB.t1 VPB.t4 515.861
R54 VPB.t5 VPB.t1 408.603
R55 VPB.t8 VPB.t2 365.188
R56 VPB.t3 VPB.t0 324.329
R57 VPB VPB.t6 260.485
R58 VPB.t6 VPB.t7 255.376
R59 VPB.t2 VPB.t5 214.517
R60 VPB.t0 VPB.t8 214.517
R61 Q.n1 Q 589.777
R62 Q.n1 Q.n0 585
R63 Q.n2 Q.n1 585
R64 Q.n1 Q.t0 26.3844
R65 Q Q.n2 12.8005
R66 Q Q.n0 11.0811
R67 Q Q.n0 3.05722
R68 Q.n2 Q 1.33781
R69 a_27_115.t0 a_27_115.n1 478.534
R70 a_27_115.n1 a_27_115.n0 376.942
R71 a_27_115.n0 a_27_115.t3 297.233
R72 a_27_115.n1 a_27_115.t1 230.541
R73 a_27_115.n0 a_27_115.t2 222.743
R74 VGND.n1 VGND.n0 288.024
R75 VGND.n7 VGND.n4 142.895
R76 VGND.n6 VGND.n5 116.719
R77 VGND.n5 VGND.t1 97.6196
R78 VGND.n4 VGND.t3 76.0861
R79 VGND.n0 VGND.t5 55.6369
R80 VGND.n10 VGND.n3 36.1417
R81 VGND.n11 VGND.n10 36.1417
R82 VGND.n12 VGND.n11 36.1417
R83 VGND.n5 VGND.t2 27.188
R84 VGND.n0 VGND.t4 26.4679
R85 VGND.n12 VGND.n1 22.1206
R86 VGND.n4 VGND.t0 20.5121
R87 VGND.n6 VGND.n3 13.177
R88 VGND.n13 VGND.n12 9.3005
R89 VGND.n11 VGND.n2 9.3005
R90 VGND.n10 VGND.n9 9.3005
R91 VGND.n8 VGND.n3 9.3005
R92 VGND.n14 VGND.n1 9.10055
R93 VGND.n7 VGND.n6 7.57984
R94 VGND VGND.n14 0.161517
R95 VGND.n8 VGND.n7 0.160525
R96 VGND.n14 VGND.n13 0.146304
R97 VGND.n9 VGND.n8 0.122949
R98 VGND.n9 VGND.n2 0.122949
R99 VGND.n13 VGND.n2 0.122949
R100 a_655_79.t0 a_655_79.t1 45.0005
R101 VNB.t5 VNB.t1 2933.33
R102 VNB.t1 VNB.t3 1951.71
R103 VNB.t2 VNB.t6 1593.7
R104 VNB.t7 VNB.t5 1362.73
R105 VNB.t4 VNB.t0 1293.44
R106 VNB VNB.t7 1143.31
R107 VNB.t6 VNB.t4 900.788
R108 VNB.t3 VNB.t2 900.788
R109 a_217_419.t0 a_217_419.n1 734.351
R110 a_217_419.t0 a_217_419.n4 727.567
R111 a_217_419.n1 a_217_419.n0 476.411
R112 a_217_419.n3 a_217_419.t1 292.892
R113 a_217_419.n0 a_217_419.t5 284.964
R114 a_217_419.n0 a_217_419.t2 273.67
R115 a_217_419.n2 a_217_419.t4 213.954
R116 a_217_419.n2 a_217_419.t3 166.181
R117 a_217_419.n3 a_217_419.n2 100.093
R118 a_217_419.n4 a_217_419.n3 39.9413
R119 a_217_419.n4 a_217_419.n1 7.2965
R120 a_669_392.n3 a_669_392.n2 383.012
R121 a_669_392.n0 a_669_392.t5 275.812
R122 a_669_392.n2 a_669_392.n0 225.887
R123 a_669_392.n0 a_669_392.t4 187.981
R124 a_669_392.n2 a_669_392.n1 185
R125 a_669_392.n3 a_669_392.t1 88.5098
R126 a_669_392.n1 a_669_392.t0 76.3792
R127 a_669_392.n1 a_669_392.t3 75.2572
R128 a_669_392.t2 a_669_392.n3 47.2805
R129 GATE_N.n0 GATE_N.t0 232.341
R130 GATE_N.n0 GATE_N.t1 202.35
R131 GATE_N GATE_N.n0 154.941
R132 a_871_139.t0 a_871_139.t1 68.5719
R133 a_369_392.t1 a_369_392.n1 781.664
R134 a_369_392.n0 a_369_392.t3 383.628
R135 a_369_392.n0 a_369_392.t2 382.805
R136 a_369_392.n1 a_369_392.t0 256.344
R137 a_369_392.n1 a_369_392.n0 72.8829
R138 a_585_392.t0 a_585_392.t1 53.1905
R139 D.n0 D.t0 337.132
R140 D D.n0 176.775
R141 D.n0 D.t1 166.559
C0 VPB D 0.059265f
C1 VPB GATE_N 0.063957f
C2 VPB VPWR 0.202103f
C3 D GATE_N 0.044779f
C4 VPB VGND 0.016621f
C5 D VPWR 0.019996f
C6 GATE_N VPWR 0.026542f
C7 VPB Q 0.013721f
C8 D VGND 0.00821f
C9 GATE_N VGND 0.008017f
C10 VPWR VGND 0.117798f
C11 GATE_N Q 2.46e-21
C12 VPWR Q 0.128805f
C13 VGND Q 0.101699f
C14 Q VNB 0.109861f
C15 VGND VNB 0.824058f
C16 VPWR VNB 0.628123f
C17 GATE_N VNB 0.101728f
C18 D VNB 0.178797f
C19 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvn_8 VNB VPB VPWR VGND A TE_B Z
X0 a_293_74.t7 a_126_74.t2 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_239_368.t11 A.t0 Z.t7 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Z.t6 A.t1 a_239_368.t10 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VPWR.t7 TE_B.t0 a_239_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_239_368.t9 A.t2 Z.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VGND.t4 a_126_74.t3 a_293_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VPWR.t6 TE_B.t1 a_239_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 a_239_368.t12 TE_B.t2 VPWR.t5 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8 Z.t4 A.t3 a_239_368.t8 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Z.t15 A.t4 a_293_74.t8 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_239_368.t7 A.t5 Z.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X11 Z.t14 A.t6 a_293_74.t9 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X12 a_126_74.t1 TE_B.t3 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 a_293_74.t5 a_126_74.t4 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X14 a_293_74.t10 A.t7 Z.t13 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X15 a_293_74.t4 a_126_74.t5 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 VPWR.t4 TE_B.t4 a_239_368.t15 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_293_74.t11 A.t8 Z.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_239_368.t2 TE_B.t5 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X19 Z.t2 A.t9 a_239_368.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_239_368.t3 TE_B.t6 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X21 a_239_368.t5 A.t10 Z.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X22 Z.t0 A.t11 a_239_368.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_293_74.t12 A.t12 Z.t11 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VGND.t1 a_126_74.t6 a_293_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 VGND.t0 a_126_74.t7 a_293_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 a_126_74.t0 TE_B.t7 VPWR.t8 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X27 Z.t10 A.t13 a_293_74.t13 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VPWR.t1 TE_B.t8 a_239_368.t13 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X29 VGND.t7 a_126_74.t8 a_293_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X30 a_293_74.t0 a_126_74.t9 VGND.t6 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 a_239_368.t14 TE_B.t9 VPWR.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X32 Z.t9 A.t14 a_293_74.t14 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 a_293_74.t15 A.t15 Z.t8 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_126_74.n0 a_126_74.t9 281.168
R1 a_126_74.t0 a_126_74.n7 273.32
R2 a_126_74.n7 a_126_74.n6 237.3
R3 a_126_74.n2 a_126_74.n1 160.667
R4 a_126_74.n4 a_126_74.n3 160.667
R5 a_126_74.n6 a_126_74.t8 142.994
R6 a_126_74.n5 a_126_74.t2 142.994
R7 a_126_74.n4 a_126_74.t7 142.994
R8 a_126_74.n3 a_126_74.t5 142.994
R9 a_126_74.n2 a_126_74.t6 142.994
R10 a_126_74.n1 a_126_74.t4 142.994
R11 a_126_74.n0 a_126_74.t3 142.994
R12 a_126_74.n7 a_126_74.t1 141.993
R13 a_126_74.n1 a_126_74.n0 138.173
R14 a_126_74.n3 a_126_74.n2 138.173
R15 a_126_74.n5 a_126_74.n4 138.173
R16 a_126_74.n6 a_126_74.n5 138.173
R17 VGND.n22 VGND.t8 156.062
R18 VGND.n15 VGND.n14 124.29
R19 VGND.n7 VGND.n6 121.306
R20 VGND.n5 VGND.n4 116.644
R21 VGND.n12 VGND.n11 116.644
R22 VGND.n10 VGND.n3 36.1417
R23 VGND.n16 VGND.n13 36.1417
R24 VGND.n20 VGND.n1 36.1417
R25 VGND.n21 VGND.n20 36.1417
R26 VGND.n4 VGND.t3 34.0546
R27 VGND.n11 VGND.t2 34.0546
R28 VGND.n6 VGND.t6 22.7032
R29 VGND.n6 VGND.t4 22.7032
R30 VGND.n4 VGND.t1 22.7032
R31 VGND.n11 VGND.t0 22.7032
R32 VGND.n14 VGND.t5 22.7032
R33 VGND.n14 VGND.t7 22.7032
R34 VGND.n22 VGND.n21 16.1887
R35 VGND.n15 VGND.n1 14.6829
R36 VGND.n7 VGND.n5 13.0424
R37 VGND.n23 VGND.n22 9.3005
R38 VGND.n21 VGND.n0 9.3005
R39 VGND.n20 VGND.n19 9.3005
R40 VGND.n18 VGND.n1 9.3005
R41 VGND.n8 VGND.n3 9.3005
R42 VGND.n10 VGND.n9 9.3005
R43 VGND.n13 VGND.n2 9.3005
R44 VGND.n17 VGND.n16 9.3005
R45 VGND.n13 VGND.n12 7.15344
R46 VGND.n5 VGND.n3 4.89462
R47 VGND.n12 VGND.n10 4.14168
R48 VGND.n16 VGND.n15 2.63579
R49 VGND.n8 VGND.n7 1.11297
R50 VGND.n9 VGND.n8 0.122949
R51 VGND.n9 VGND.n2 0.122949
R52 VGND.n17 VGND.n2 0.122949
R53 VGND.n18 VGND.n17 0.122949
R54 VGND.n19 VGND.n18 0.122949
R55 VGND.n19 VGND.n0 0.122949
R56 VGND.n23 VGND.n0 0.122949
R57 VGND VGND.n23 0.0617245
R58 a_293_74.n12 a_293_74.t1 225.41
R59 a_293_74.n2 a_293_74.t10 205.042
R60 a_293_74.n3 a_293_74.n0 187.327
R61 a_293_74.n2 a_293_74.n1 185
R62 a_293_74.n5 a_293_74.n4 185
R63 a_293_74.n11 a_293_74.n10 119.427
R64 a_293_74.n13 a_293_74.n12 119.427
R65 a_293_74.n9 a_293_74.n8 114.82
R66 a_293_74.n9 a_293_74.n7 89.5921
R67 a_293_74.n7 a_293_74.n6 86.1054
R68 a_293_74.n11 a_293_74.n9 55.8085
R69 a_293_74.n12 a_293_74.n11 51.2005
R70 a_293_74.n3 a_293_74.n2 49.7334
R71 a_293_74.n7 a_293_74.n5 44.6993
R72 a_293_74.n5 a_293_74.n3 34.5048
R73 a_293_74.n0 a_293_74.t11 34.0546
R74 a_293_74.n8 a_293_74.t6 22.7032
R75 a_293_74.n8 a_293_74.t5 22.7032
R76 a_293_74.n6 a_293_74.t14 22.7032
R77 a_293_74.n6 a_293_74.t0 22.7032
R78 a_293_74.n4 a_293_74.t13 22.7032
R79 a_293_74.n4 a_293_74.t12 22.7032
R80 a_293_74.n1 a_293_74.t8 22.7032
R81 a_293_74.n1 a_293_74.t15 22.7032
R82 a_293_74.n0 a_293_74.t9 22.7032
R83 a_293_74.n10 a_293_74.t3 22.7032
R84 a_293_74.n10 a_293_74.t4 22.7032
R85 a_293_74.n13 a_293_74.t2 22.7032
R86 a_293_74.t7 a_293_74.n13 22.7032
R87 VNB.t8 VNB.t1 2933.33
R88 VNB.t9 VNB.t11 1316.54
R89 VNB VNB.t8 1281.89
R90 VNB.t12 VNB.t10 1154.86
R91 VNB.t3 VNB.t5 1154.86
R92 VNB.t2 VNB.t4 1154.86
R93 VNB.t16 VNB.t9 993.177
R94 VNB.t10 VNB.t16 993.177
R95 VNB.t14 VNB.t12 993.177
R96 VNB.t13 VNB.t14 993.177
R97 VNB.t15 VNB.t13 993.177
R98 VNB.t0 VNB.t15 993.177
R99 VNB.t6 VNB.t0 993.177
R100 VNB.t5 VNB.t6 993.177
R101 VNB.t4 VNB.t3 993.177
R102 VNB.t7 VNB.t2 993.177
R103 VNB.t1 VNB.t7 993.177
R104 A.n0 A.t0 226.809
R105 A.n1 A.t1 226.809
R106 A.n22 A.t2 226.809
R107 A.n3 A.t3 226.809
R108 A.n5 A.t5 226.809
R109 A.n12 A.t9 226.809
R110 A.n8 A.t10 226.809
R111 A.n6 A.t11 226.809
R112 A.n6 A.t14 197.475
R113 A.n0 A.t7 197.475
R114 A.n7 A.t12 196.013
R115 A.n11 A.t13 196.013
R116 A.n10 A.t8 196.013
R117 A.n4 A.t6 196.013
R118 A.n21 A.t15 196.013
R119 A.n2 A.t4 196.013
R120 A.n14 A.n9 162.121
R121 A.n28 A.n27 152
R122 A.n26 A.n25 152
R123 A.n24 A.n23 152
R124 A.n20 A.n19 152
R125 A.n18 A.n17 152
R126 A.n16 A.n15 152
R127 A.n14 A.n13 152
R128 A.n7 A.n6 61.346
R129 A.n27 A.n26 49.6611
R130 A.n17 A.n16 49.6611
R131 A.n9 A.n8 43.0884
R132 A.n20 A.n3 37.246
R133 A.n23 A.n2 28.4823
R134 A.n13 A.n10 28.4823
R135 A.n13 A.n12 27.0217
R136 A.n23 A.n22 21.1793
R137 A.n10 A.n5 17.5278
R138 A.n2 A.n1 16.0672
R139 A.n21 A.n20 15.3369
R140 A.n11 A.n9 15.3369
R141 A.n22 A.n21 13.146
R142 A.n27 A.n0 10.955
R143 A.n4 A.n3 10.2247
R144 A.n25 A.n24 10.1214
R145 A.n15 A.n14 10.1214
R146 A.n19 A 9.37724
R147 A.n18 A 9.07957
R148 A A.n28 7.5912
R149 A.n12 A.n11 7.30353
R150 A.n28 A 6.69817
R151 A A.n18 5.2098
R152 A.n26 A.n1 5.11262
R153 A.n19 A 4.91213
R154 A.n8 A.n7 4.38232
R155 A.n16 A.n5 3.65202
R156 A.n25 A 3.42376
R157 A.n17 A.n4 2.19141
R158 A.n15 A 1.04236
R159 A.n24 A 0.744686
R160 Z.n2 Z.n0 340.937
R161 Z.n6 Z.n5 300.733
R162 Z.n2 Z.n1 298.019
R163 Z.n4 Z.n3 298.019
R164 Z.n9 Z.n8 254.819
R165 Z.n9 Z.n7 202.319
R166 Z.n11 Z.n10 185
R167 Z.n13 Z.n12 185
R168 Z.n11 Z.n9 62.7517
R169 Z.n6 Z.n4 59.1064
R170 Z.n4 Z.n2 42.9181
R171 Z.n3 Z.t2 35.1791
R172 Z.n8 Z.t13 34.0546
R173 Z.n8 Z.t15 34.0546
R174 Z.n13 Z.n11 29.8628
R175 Z Z.n14 27.8266
R176 Z.n14 Z.n13 26.4301
R177 Z.n5 Z.t1 26.3844
R178 Z.n5 Z.t0 26.3844
R179 Z.n0 Z.t7 26.3844
R180 Z.n0 Z.t6 26.3844
R181 Z.n1 Z.t5 26.3844
R182 Z.n1 Z.t4 26.3844
R183 Z.n3 Z.t3 26.3844
R184 Z.n12 Z.t11 22.7032
R185 Z.n12 Z.t9 22.7032
R186 Z.n10 Z.t12 22.7032
R187 Z.n10 Z.t10 22.7032
R188 Z.n7 Z.t8 22.7032
R189 Z.n7 Z.t14 22.7032
R190 Z.n14 Z.n6 18.2524
R191 a_239_368.n12 a_239_368.n1 305.901
R192 a_239_368.n13 a_239_368.n0 305.901
R193 a_239_368.n11 a_239_368.n10 302.74
R194 a_239_368.n4 a_239_368.t1 302.459
R195 a_239_368.t11 a_239_368.n13 301.389
R196 a_239_368.n4 a_239_368.n3 223.369
R197 a_239_368.n6 a_239_368.n5 223.369
R198 a_239_368.n7 a_239_368.n2 202.3
R199 a_239_368.n9 a_239_368.n8 189.115
R200 a_239_368.n13 a_239_368.n12 67.7652
R201 a_239_368.n9 a_239_368.n7 64.8587
R202 a_239_368.n11 a_239_368.n9 62.9747
R203 a_239_368.n12 a_239_368.n11 59.1064
R204 a_239_368.n7 a_239_368.n6 57.3481
R205 a_239_368.n6 a_239_368.n4 52.7064
R206 a_239_368.n8 a_239_368.t4 26.3844
R207 a_239_368.n8 a_239_368.t3 26.3844
R208 a_239_368.n2 a_239_368.t0 26.3844
R209 a_239_368.n2 a_239_368.t12 26.3844
R210 a_239_368.n3 a_239_368.t13 26.3844
R211 a_239_368.n3 a_239_368.t14 26.3844
R212 a_239_368.n5 a_239_368.t15 26.3844
R213 a_239_368.n5 a_239_368.t2 26.3844
R214 a_239_368.n10 a_239_368.t6 26.3844
R215 a_239_368.n10 a_239_368.t5 26.3844
R216 a_239_368.n1 a_239_368.t8 26.3844
R217 a_239_368.n1 a_239_368.t7 26.3844
R218 a_239_368.n0 a_239_368.t10 26.3844
R219 a_239_368.n0 a_239_368.t9 26.3844
R220 VPB.t4 VPB.t1 515.861
R221 VPB VPB.t4 283.469
R222 VPB.t0 VPB.t3 280.914
R223 VPB.t7 VPB.t8 255.376
R224 VPB.t16 VPB.t13 255.376
R225 VPB.t14 VPB.t2 255.376
R226 VPB.t1 VPB.t15 255.376
R227 VPB.t11 VPB.t12 229.839
R228 VPB.t10 VPB.t11 229.839
R229 VPB.t9 VPB.t10 229.839
R230 VPB.t8 VPB.t9 229.839
R231 VPB.t6 VPB.t7 229.839
R232 VPB.t5 VPB.t6 229.839
R233 VPB.t3 VPB.t5 229.839
R234 VPB.t13 VPB.t0 229.839
R235 VPB.t2 VPB.t16 229.839
R236 VPB.t15 VPB.t14 229.839
R237 TE_B.n0 TE_B.t6 376.567
R238 TE_B.n7 TE_B.n6 289.538
R239 TE_B.n7 TE_B.t7 221.452
R240 TE_B.n0 TE_B.t0 204.048
R241 TE_B.n1 TE_B.t2 204.048
R242 TE_B.n2 TE_B.t4 204.048
R243 TE_B.n3 TE_B.t5 204.048
R244 TE_B.n4 TE_B.t8 204.048
R245 TE_B.n5 TE_B.t9 204.048
R246 TE_B.n6 TE_B.t1 204.048
R247 TE_B.n8 TE_B.t3 194.674
R248 TE_B TE_B.n8 161.892
R249 TE_B.n2 TE_B.n1 148.49
R250 TE_B.n4 TE_B.n3 148.49
R251 TE_B.n6 TE_B.n5 148.49
R252 TE_B.n1 TE_B.n0 132.423
R253 TE_B.n3 TE_B.n2 132.423
R254 TE_B.n5 TE_B.n4 132.423
R255 TE_B.n8 TE_B.n7 16.5135
R256 VPWR.n8 VPWR.n7 321.365
R257 VPWR.n18 VPWR.t8 258.875
R258 VPWR.n2 VPWR.n1 222.837
R259 VPWR.n11 VPWR.n4 222.837
R260 VPWR.n6 VPWR.n5 222.837
R261 VPWR.n17 VPWR.n16 36.1417
R262 VPWR.n1 VPWR.t0 35.1791
R263 VPWR.n4 VPWR.t3 35.1791
R264 VPWR.n5 VPWR.t5 35.1791
R265 VPWR.n7 VPWR.t2 35.1791
R266 VPWR.n7 VPWR.t7 35.1791
R267 VPWR.n16 VPWR.n2 32.0005
R268 VPWR.n12 VPWR.n11 31.2476
R269 VPWR.n10 VPWR.n6 30.4946
R270 VPWR.n1 VPWR.t6 26.3844
R271 VPWR.n4 VPWR.t1 26.3844
R272 VPWR.n5 VPWR.t4 26.3844
R273 VPWR.n18 VPWR.n17 20.7064
R274 VPWR.n11 VPWR.n10 16.1887
R275 VPWR.n12 VPWR.n2 15.4358
R276 VPWR.n10 VPWR.n9 9.3005
R277 VPWR.n11 VPWR.n3 9.3005
R278 VPWR.n13 VPWR.n12 9.3005
R279 VPWR.n14 VPWR.n2 9.3005
R280 VPWR.n16 VPWR.n15 9.3005
R281 VPWR.n17 VPWR.n0 9.3005
R282 VPWR.n19 VPWR.n18 9.3005
R283 VPWR.n8 VPWR.n6 6.37487
R284 VPWR.n9 VPWR.n8 0.499395
R285 VPWR.n9 VPWR.n3 0.122949
R286 VPWR.n13 VPWR.n3 0.122949
R287 VPWR.n14 VPWR.n13 0.122949
R288 VPWR.n15 VPWR.n14 0.122949
R289 VPWR.n15 VPWR.n0 0.122949
R290 VPWR.n19 VPWR.n0 0.122949
R291 VPWR VPWR.n19 0.0617245
C0 VGND A 0.04842f
C1 TE_B A 0.023013f
C2 VPWR VGND 0.14739f
C3 VPWR TE_B 0.222167f
C4 VPWR A 0.048958f
C5 Z VPB 0.007461f
C6 Z VGND 0.039112f
C7 VGND VPB 0.00886f
C8 Z TE_B 0.011621f
C9 VPB TE_B 0.380308f
C10 Z A 0.704367f
C11 VGND TE_B 0.061303f
C12 VPB A 0.285966f
C13 VPWR Z 0.041745f
C14 VPWR VPB 0.22203f
C15 VGND VNB 1.06114f
C16 Z VNB 0.037725f
C17 VPWR VNB 0.85336f
C18 A VNB 0.86308f
C19 TE_B VNB 0.512007f
C20 VPB VNB 2.1204f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvn_4 VNB VPB VPWR VGND TE_B A Z
X0 a_241_368.t5 A.t0 Z.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Z.t4 A.t1 a_241_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_281_74.t5 A.t2 Z.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_241_368.t7 TE_B.t0 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 a_114_74.t1 TE_B.t1 VPWR.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 VGND.t4 a_114_74.t2 a_281_74.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_114_74.t0 TE_B.t2 VGND.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 Z.t0 A.t3 a_281_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1073 ps=1.03 w=0.74 l=0.15
X8 VPWR.t3 TE_B.t3 a_241_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_241_368.t1 TE_B.t4 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Z.t7 A.t4 a_281_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VGND.t3 a_114_74.t3 a_281_74.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_281_74.t2 A.t5 Z.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t1 TE_B.t5 a_241_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X14 a_281_74.t0 a_114_74.t4 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_281_74.t1 a_114_74.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_241_368.t3 A.t6 Z.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X17 Z.t2 A.t7 a_241_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n3 A.t6 214.758
R1 A.n6 A.t7 214.758
R2 A.n8 A.t0 214.758
R3 A.n7 A.t1 214.645
R4 A A.n10 161.514
R5 A.n2 A.n1 161.067
R6 A.n7 A.t4 154.24
R7 A.n9 A.t5 154.24
R8 A.n5 A.t3 154.24
R9 A.n2 A.t2 154.24
R10 A.n4 A.n0 152
R11 A.n8 A.n7 37.2243
R12 A.n10 A.n9 27.2025
R13 A.n4 A.n3 22.4302
R14 A.n5 A.n4 17.6579
R15 A.n10 A.n6 11.9312
R16 A.n1 A.n0 11.7627
R17 A.n9 A.n8 3.81832
R18 A.n6 A.n5 2.86387
R19 A.n1 A 2.59509
R20 A A.n0 2.24915
R21 A.n3 A.n2 0.954955
R22 Z.n2 Z.n0 251.494
R23 Z.n5 Z.n3 225.673
R24 Z.n2 Z.n1 208.577
R25 Z.n5 Z.n4 185
R26 Z Z.n5 37.2601
R27 Z.n1 Z.t5 26.3844
R28 Z.n1 Z.t4 26.3844
R29 Z.n0 Z.t3 26.3844
R30 Z.n0 Z.t2 26.3844
R31 Z.n4 Z.t6 22.7032
R32 Z.n4 Z.t7 22.7032
R33 Z.n3 Z.t1 22.7032
R34 Z.n3 Z.t0 22.7032
R35 Z Z.n2 8.72777
R36 a_241_368.n5 a_241_368.n4 309.978
R37 a_241_368.n1 a_241_368.t0 303.25
R38 a_241_368.n4 a_241_368.t3 303.128
R39 a_241_368.n1 a_241_368.n0 227.923
R40 a_241_368.n3 a_241_368.n2 185.916
R41 a_241_368.n3 a_241_368.n1 94.7148
R42 a_241_368.n4 a_241_368.n3 90.8293
R43 a_241_368.n2 a_241_368.t4 26.3844
R44 a_241_368.n2 a_241_368.t7 26.3844
R45 a_241_368.n0 a_241_368.t6 26.3844
R46 a_241_368.n0 a_241_368.t1 26.3844
R47 a_241_368.n5 a_241_368.t2 26.3844
R48 a_241_368.t5 a_241_368.n5 26.3844
R49 VPB.t8 VPB.t0 515.861
R50 VPB VPB.t8 288.575
R51 VPB.t6 VPB.t7 255.376
R52 VPB.t2 VPB.t3 229.839
R53 VPB.t5 VPB.t2 229.839
R54 VPB.t4 VPB.t5 229.839
R55 VPB.t7 VPB.t4 229.839
R56 VPB.t1 VPB.t6 229.839
R57 VPB.t0 VPB.t1 229.839
R58 a_281_74.t5 a_281_74.n5 267.104
R59 a_281_74.n1 a_281_74.t7 225.786
R60 a_281_74.n5 a_281_74.n4 185
R61 a_281_74.n1 a_281_74.n0 113.438
R62 a_281_74.n3 a_281_74.n2 88.4224
R63 a_281_74.n3 a_281_74.n1 80.5269
R64 a_281_74.n5 a_281_74.n3 39.5417
R65 a_281_74.n4 a_281_74.t4 23.514
R66 a_281_74.n4 a_281_74.t2 23.514
R67 a_281_74.n2 a_281_74.t3 22.7032
R68 a_281_74.n2 a_281_74.t0 22.7032
R69 a_281_74.n0 a_281_74.t6 22.7032
R70 a_281_74.n0 a_281_74.t1 22.7032
R71 VNB.t6 VNB.t8 2933.33
R72 VNB VNB.t6 1143.31
R73 VNB.t2 VNB.t4 1016.27
R74 VNB.t4 VNB.t5 993.177
R75 VNB.t3 VNB.t2 993.177
R76 VNB.t0 VNB.t3 993.177
R77 VNB.t7 VNB.t0 993.177
R78 VNB.t1 VNB.t7 993.177
R79 VNB.t8 VNB.t1 993.177
R80 TE_B.n0 TE_B.t0 360.5
R81 TE_B.n3 TE_B.n2 289.538
R82 TE_B.n3 TE_B.t1 221.579
R83 TE_B.n0 TE_B.t3 204.048
R84 TE_B.n1 TE_B.t4 204.048
R85 TE_B.n2 TE_B.t5 204.048
R86 TE_B.n4 TE_B.t2 194.952
R87 TE_B TE_B.n4 155.601
R88 TE_B.n1 TE_B.n0 132.423
R89 TE_B.n2 TE_B.n1 132.423
R90 TE_B.n4 TE_B.n3 16.825
R91 VPWR.n8 VPWR.t0 257.433
R92 VPWR.n2 VPWR.n1 232.787
R93 VPWR.n4 VPWR.n3 229.286
R94 VPWR.n7 VPWR.n6 36.1417
R95 VPWR.n3 VPWR.t4 35.1791
R96 VPWR.n6 VPWR.n2 32.7534
R97 VPWR.n1 VPWR.t2 26.3844
R98 VPWR.n1 VPWR.t1 26.3844
R99 VPWR.n3 VPWR.t3 26.3844
R100 VPWR.n8 VPWR.n7 22.2123
R101 VPWR.n6 VPWR.n5 9.3005
R102 VPWR.n7 VPWR.n0 9.3005
R103 VPWR.n9 VPWR.n8 9.3005
R104 VPWR.n4 VPWR.n2 6.59907
R105 VPWR.n5 VPWR.n4 0.518303
R106 VPWR.n5 VPWR.n0 0.122949
R107 VPWR.n9 VPWR.n0 0.122949
R108 VPWR VPWR.n9 0.0617245
R109 a_114_74.n0 a_114_74.t4 281.168
R110 a_114_74.t1 a_114_74.n3 271.154
R111 a_114_74.n3 a_114_74.n2 241.428
R112 a_114_74.n2 a_114_74.t2 142.994
R113 a_114_74.n1 a_114_74.t5 142.994
R114 a_114_74.n0 a_114_74.t3 142.994
R115 a_114_74.n3 a_114_74.t0 141.698
R116 a_114_74.n1 a_114_74.n0 138.173
R117 a_114_74.n2 a_114_74.n1 138.173
R118 VGND.n10 VGND.t0 171.77
R119 VGND.n5 VGND.n4 121.352
R120 VGND.n3 VGND.n2 115.885
R121 VGND.n8 VGND.n1 36.1417
R122 VGND.n9 VGND.n8 36.1417
R123 VGND.n10 VGND.n9 26.7299
R124 VGND.n4 VGND.t2 22.7032
R125 VGND.n4 VGND.t3 22.7032
R126 VGND.n2 VGND.t1 22.7032
R127 VGND.n2 VGND.t4 22.7032
R128 VGND.n3 VGND.n1 10.1652
R129 VGND.n11 VGND.n10 9.3005
R130 VGND.n6 VGND.n1 9.3005
R131 VGND.n8 VGND.n7 9.3005
R132 VGND.n9 VGND.n0 9.3005
R133 VGND.n5 VGND.n3 7.77179
R134 VGND.n6 VGND.n5 1.11297
R135 VGND.n7 VGND.n6 0.122949
R136 VGND.n7 VGND.n0 0.122949
R137 VGND.n11 VGND.n0 0.122949
R138 VGND VGND.n11 0.0617245
C0 VPWR VGND 0.085547f
C1 Z VGND 0.017055f
C2 VPWR VPB 0.14556f
C3 VPWR TE_B 0.142451f
C4 Z VPB 0.005173f
C5 VPWR A 0.025659f
C6 VGND VPB 0.008258f
C7 VGND TE_B 0.0495f
C8 Z A 0.284037f
C9 VGND A 0.026672f
C10 VPB TE_B 0.228346f
C11 VPB A 0.140061f
C12 TE_B A 0.023586f
C13 VPWR Z 0.020156f
C14 VGND VNB 0.662707f
C15 Z VNB 0.019837f
C16 VPWR VNB 0.53574f
C17 A VNB 0.458717f
C18 TE_B VNB 0.357631f
C19 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvn_2 VNB VPB VPWR VGND TE_B A Z
X0 Z.t3 A.t0 a_227_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_227_368.t0 TE_B.t0 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t1 TE_B.t1 a_227_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_231_74.t1 a_115_464.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_115_464.t1 TE_B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1856 pd=1.86 as=0.1856 ps=1.86 w=0.64 l=0.15
X5 a_115_464.t0 TE_B.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X6 VGND.t1 a_115_464.t3 a_231_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 Z.t0 A.t1 a_231_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_231_74.t2 A.t2 Z.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1995 pd=2.08 as=0.10545 ps=1.025 w=0.74 l=0.15
X9 a_227_368.t2 A.t3 Z.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A.n0 A.t0 328.358
R1 A.n2 A.t3 261.62
R2 A A.n2 193.113
R3 A.n0 A.t1 172.779
R4 A.n1 A.t2 154.24
R5 A.n1 A.n0 88.075
R6 A.n2 A.n1 6.57323
R7 a_227_368.n0 a_227_368.t2 316.44
R8 a_227_368.n0 a_227_368.t1 303.375
R9 a_227_368.n1 a_227_368.n0 186.857
R10 a_227_368.n1 a_227_368.t3 26.3844
R11 a_227_368.t0 a_227_368.n1 26.3844
R12 Z Z.n0 202.953
R13 Z.n2 Z.n1 185
R14 Z.n0 Z.t2 26.3844
R15 Z.n0 Z.t3 26.3844
R16 Z.n1 Z.t1 23.514
R17 Z.n1 Z.t0 22.7032
R18 Z Z.n2 12.0649
R19 Z.n2 Z 2.71565
R20 VPB.t0 VPB.t2 513.307
R21 VPB VPB.t0 255.376
R22 VPB.t4 VPB.t3 229.839
R23 VPB.t1 VPB.t4 229.839
R24 VPB.t2 VPB.t1 229.839
R25 TE_B.t2 TE_B.n0 449.868
R26 TE_B.n0 TE_B.t0 348.647
R27 TE_B.n0 TE_B.t1 204.048
R28 TE_B.n1 TE_B.t2 200.673
R29 TE_B.n2 TE_B.t3 195.31
R30 TE_B.n3 TE_B.n2 152
R31 TE_B TE_B.n1 70.0219
R32 TE_B.n2 TE_B.n1 63.9023
R33 TE_B TE_B.n3 8.88521
R34 TE_B.n3 TE_B 2.25932
R35 VPWR.n1 VPWR.t0 389.99
R36 VPWR.n1 VPWR.n0 333.384
R37 VPWR.n0 VPWR.t2 26.3844
R38 VPWR.n0 VPWR.t1 26.3844
R39 VPWR VPWR.n1 0.148859
R40 a_115_464.t1 a_115_464.n1 415.443
R41 a_115_464.n0 a_115_464.t2 324.548
R42 a_115_464.n1 a_115_464.n0 290.173
R43 a_115_464.n1 a_115_464.t0 277.122
R44 a_115_464.n0 a_115_464.t3 186.374
R45 VGND.n1 VGND.t0 261.882
R46 VGND.n1 VGND.n0 214.708
R47 VGND.n0 VGND.t2 22.7032
R48 VGND.n0 VGND.t1 22.7032
R49 VGND VGND.n1 0.151277
R50 a_231_74.n0 a_231_74.t2 268.558
R51 a_231_74.n0 a_231_74.t0 222.797
R52 a_231_74.n1 a_231_74.n0 86.1054
R53 a_231_74.n1 a_231_74.t3 22.7032
R54 a_231_74.t1 a_231_74.n1 22.7032
R55 VNB.t0 VNB.t1 2321.26
R56 VNB VNB.t0 1177.95
R57 VNB.t4 VNB.t3 1004.72
R58 VNB.t2 VNB.t4 993.177
R59 VNB.t1 VNB.t2 993.177
C0 VPB Z 0.006193f
C1 TE_B VPWR 0.119189f
C2 VPB VGND 0.008754f
C3 A VPWR 0.013202f
C4 TE_B Z 0.001289f
C5 TE_B VGND 0.039471f
C6 A Z 0.125476f
C7 A VGND 0.020492f
C8 VPWR Z 0.009856f
C9 VPWR VGND 0.053091f
C10 Z VGND 0.007284f
C11 VPB TE_B 0.243789f
C12 VPB A 0.072118f
C13 TE_B A 0.014859f
C14 VPB VPWR 0.089574f
C15 VGND VNB 0.462814f
C16 Z VNB 0.020825f
C17 VPWR VNB 0.371458f
C18 A VNB 0.296906f
C19 TE_B VNB 0.342922f
C20 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvn_1 VNB VPB VPWR VGND A Z TE_B
X0 VGND.t1 TE_B.t0 a_22_46.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1282 pd=1.18 as=0.1218 ps=1.42 w=0.42 l=0.15
X1 Z.t1 A.t0 a_278_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X2 a_278_368.t1 TE_B.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.194 ps=1.505 w=1.12 l=0.15
X3 VPWR.t0 TE_B.t2 a_22_46.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.505 as=0.1888 ps=1.87 w=0.64 l=0.15
X4 Z.t0 A.t1 a_281_100.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5 a_281_100.t0 a_22_46.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1282 ps=1.18 w=0.74 l=0.15
R0 TE_B.n0 TE_B.t1 338.075
R1 TE_B TE_B.n1 171.201
R2 TE_B.n0 TE_B.t2 157.905
R3 TE_B.n1 TE_B.t0 120.903
R4 TE_B.n1 TE_B.n0 9.85959
R5 a_22_46.n0 a_22_46.t2 443.882
R6 a_22_46.t0 a_22_46.n0 423.901
R7 a_22_46.n0 a_22_46.t1 225
R8 VGND.n3 VGND.n0 202.456
R9 VGND.n3 VGND.n2 185
R10 VGND.n1 VGND.t1 57.6101
R11 VGND.t0 VGND.n0 49.4123
R12 VGND.n2 VGND.t0 42.0005
R13 VGND VGND.n3 31.0211
R14 VGND.n1 VGND.n0 1.76521
R15 VGND.n2 VGND.n1 1.5005
R16 VNB VNB.t2 1893.96
R17 VNB.t2 VNB.t1 1177.95
R18 VNB.t1 VNB.t0 900.788
R19 A.n0 A.t0 250.909
R20 A.n0 A.t1 178.34
R21 A A.n0 158.4
R22 a_278_368.t0 a_278_368.t1 47.4916
R23 Z Z.n0 587.909
R24 Z.n2 Z.n0 585
R25 Z.n1 Z.n0 585
R26 Z.n1 Z.t0 196.612
R27 Z.n0 Z.t1 26.3844
R28 Z Z.n1 6.63323
R29 Z Z.n2 6.16777
R30 Z.n2 Z 2.44414
R31 VPB VPB.t1 398.387
R32 VPB.t1 VPB.t2 273.253
R33 VPB.t2 VPB.t0 214.517
R34 VPWR VPWR.n0 245.413
R35 VPWR.n0 VPWR.t0 72.3364
R36 VPWR.n0 VPWR.t1 29.2942
R37 a_281_100.t0 a_281_100.t1 38.9194
C0 VPB Z 0.022629f
C1 TE_B VPWR 0.071651f
C2 VPB VGND 0.008409f
C3 TE_B Z 0.006729f
C4 A VPWR 0.014235f
C5 TE_B VGND 0.046501f
C6 A Z 0.098211f
C7 A VGND 0.014827f
C8 VPWR Z 0.102031f
C9 VPWR VGND 0.040831f
C10 Z VGND 0.076618f
C11 VPB TE_B 0.100545f
C12 VPB A 0.036841f
C13 VPB VPWR 0.084405f
C14 TE_B A 0.053272f
C15 VGND VNB 0.334572f
C16 Z VNB 0.114651f
C17 VPWR VNB 0.279049f
C18 A VNB 0.12778f
C19 TE_B VNB 0.173506f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__edfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__edfxtp_1 VNB VPB VPWR VGND DE D CLK Q
X0 a_1895_74.t0 a_763_74.t2 a_1794_392.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.3925 ps=1.785 w=1 l=0.15
X1 VPWR.t7 DE.t0 a_159_446.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.14045 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X2 a_1797_74# a_1409_64.t1 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_27_508.t3 a_533_61.t1 a_554_436.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.39 as=0.0504 ps=0.66 w=0.42 l=0.15
X4 a_1382_508.t0 a_763_74.t3 a_1156_90.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.07455 pd=0.775 as=0.063 ps=0.72 w=0.42 l=0.15
X5 a_1156_90.t2 a_958_74.t2 a_27_508.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X6 a_1349_90.t0 a_958_74.t3 a_1156_90.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.17115 ps=1.235 w=0.42 l=0.15
X7 a_554_436.t1 DE.t1 VPWR.t8 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.14045 ps=1.17 w=0.42 l=0.15
X8 a_763_74.t1 CLK.t0 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 VPWR.t4 a_159_446.t2 a_114_508.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.0504 ps=0.66 w=0.42 l=0.15
X10 VGND.t5 DE.t2 a_131_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1176 pd=1.4 as=0.0504 ps=0.66 w=0.42 l=0.15
X11 a_131_74.t0 D.t0 a_27_508.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X12 a_491_87.t1 a_159_446.t3 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 a_958_74.t1 a_763_74.t4 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X14 a_958_74.t0 a_763_74.t5 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2072 ps=2.04 w=0.74 l=0.15
X15 a_533_61.t0 a_1895_74.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.83 as=0.14675 ps=1.2 w=0.64 l=0.15
X16 a_27_508.t2 a_533_61.t2 a_491_87.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_1409_64.t0 a_1156_90.t4 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1469 ps=1.33 w=0.84 l=0.15
X18 a_1997_74# a_763_74.t6 a_1895_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1212 ps=1.1 w=0.42 l=0.15
X19 VGND.t0 a_1895_74.t4 Q.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X20 VPWR.t0 a_533_61.t3 a_2088_502.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.14675 pd=1.2 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND.t4 DE.t3 a_159_446.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X22 a_763_74.t0 CLK.t1 VPWR.t9 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.3136 ps=2.8 w=1.12 l=0.15
X23 a_2088_502.t1 a_958_74.t4 a_1895_74.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1664 ps=1.385 w=0.42 l=0.15
X24 a_1794_392.t1 a_1409_64.t2 VPWR.t5 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3925 pd=1.785 as=0.295 ps=2.59 w=1 l=0.15
X25 a_114_508.t0 D.t1 a_27_508.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X26 VPWR.t1 a_1895_74.t5 Q.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.308 ps=2.79 w=1.12 l=0.15
X27 a_1156_90.t0 a_763_74.t7 a_27_508.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.17115 pd=1.235 as=0.1197 ps=1.41 w=0.42 l=0.15
R0 a_763_74.t0 a_763_74.n5 857.218
R1 a_763_74.n1 a_763_74.n0 582.788
R2 a_763_74.n2 a_763_74.n1 448.17
R3 a_763_74.n0 a_763_74.t6 310.087
R4 a_763_74.n2 a_763_74.t7 295.627
R5 a_763_74.n4 a_763_74.t5 259.93
R6 a_763_74.n0 a_763_74.t2 231.629
R7 a_763_74.n3 a_763_74.t4 204.048
R8 a_763_74.n5 a_763_74.t1 183.421
R9 a_763_74.n4 a_763_74.n3 160.052
R10 a_763_74.n1 a_763_74.t3 150.133
R11 a_763_74.n5 a_763_74.n4 94.0143
R12 a_763_74.n3 a_763_74.n2 89.3225
R13 a_1794_392.t0 a_1794_392.t1 154.645
R14 a_1895_74.n2 a_1895_74.t3 371.389
R15 a_1895_74.n1 a_1895_74.t5 341.685
R16 a_1895_74.n0 a_1895_74.n5 290.077
R17 a_1895_74.n2 a_1895_74.n1 260.281
R18 a_1895_74.n5 a_1895_74.t1 253.12
R19 a_1895_74.n5 a_1895_74.n4 170.619
R20 a_1895_74.n4 a_1895_74.n3 155.964
R21 a_1895_74.n1 a_1895_74.t4 142.994
R22 a_1895_74.n0 a_1895_74.t2 111.816
R23 a_1895_74.n0 a_1895_74.t0 26.9229
R24 a_1895_74.n6 a_1895_74.n0 10.7687
R25 a_1895_74.n4 a_1895_74.n2 10.581
R26 VPB.t15 VPB.t5 689.516
R27 VPB.t10 VPB.t12 577.152
R28 VPB.t6 VPB.t11 536.29
R29 VPB.t11 VPB.t14 515.861
R30 VPB.t5 VPB.t8 497.985
R31 VPB.t0 VPB.t15 497.985
R32 VPB.t4 VPB.t3 495.43
R33 VPB.t14 VPB.t7 477.555
R34 VPB.t1 VPB.t4 362.635
R35 VPB.t12 VPB.t13 347.312
R36 VPB.t7 VPB.t9 273.253
R37 VPB VPB.t2 252.823
R38 VPB.t8 VPB.t6 229.839
R39 VPB.t9 VPB.t1 214.517
R40 VPB.t13 VPB.t0 199.195
R41 VPB.t2 VPB.t10 199.195
R42 a_1409_64.t0 a_1409_64.n4 832.12
R43 a_1409_64.n3 a_1409_64.n1 361.116
R44 a_1409_64.n0 a_1409_64.t2 259.745
R45 a_1409_64.n4 a_1409_64.n3 227.702
R46 a_1409_64.n3 a_1409_64.n2 192.685
R47 a_1409_64.n0 a_1409_64.t1 174.105
R48 a_1409_64.n4 a_1409_64.n0 111.436
R49 VPWR.n34 VPWR.t3 908.659
R50 VPWR.n3 VPWR.t9 900.062
R51 VPWR.n21 VPWR.t5 854.625
R52 VPWR.n27 VPWR.t6 696.476
R53 VPWR.n49 VPWR.t4 685.053
R54 VPWR.n42 VPWR.n41 629.801
R55 VPWR.n14 VPWR.n13 600.17
R56 VPWR.n12 VPWR.t1 266.74
R57 VPWR.n41 VPWR.t7 157.279
R58 VPWR.n13 VPWR.t0 131.333
R59 VPWR.n13 VPWR.t2 109.567
R60 VPWR.n41 VPWR.t8 70.3576
R61 VPWR.n47 VPWR.n1 36.1417
R62 VPWR.n48 VPWR.n47 36.1417
R63 VPWR.n40 VPWR.n39 36.1417
R64 VPWR.n43 VPWR.n40 36.1417
R65 VPWR.n36 VPWR.n35 36.1417
R66 VPWR.n29 VPWR.n28 36.1417
R67 VPWR.n29 VPWR.n6 36.1417
R68 VPWR.n33 VPWR.n6 36.1417
R69 VPWR.n26 VPWR.n9 36.1417
R70 VPWR.n15 VPWR.n11 36.1417
R71 VPWR.n19 VPWR.n11 36.1417
R72 VPWR.n20 VPWR.n19 36.1417
R73 VPWR.n22 VPWR.n20 36.1417
R74 VPWR.n35 VPWR.n34 34.6358
R75 VPWR.n28 VPWR.n27 33.8829
R76 VPWR.n50 VPWR.n49 24.645
R77 VPWR.n34 VPWR.n33 18.824
R78 VPWR.n42 VPWR.n1 16.9417
R79 VPWR.n27 VPWR.n26 13.5534
R80 VPWR.n16 VPWR.n15 9.3005
R81 VPWR.n17 VPWR.n11 9.3005
R82 VPWR.n19 VPWR.n18 9.3005
R83 VPWR.n20 VPWR.n10 9.3005
R84 VPWR.n23 VPWR.n22 9.3005
R85 VPWR.n24 VPWR.n9 9.3005
R86 VPWR.n26 VPWR.n25 9.3005
R87 VPWR.n27 VPWR.n8 9.3005
R88 VPWR.n28 VPWR.n7 9.3005
R89 VPWR.n30 VPWR.n29 9.3005
R90 VPWR.n31 VPWR.n6 9.3005
R91 VPWR.n33 VPWR.n32 9.3005
R92 VPWR.n34 VPWR.n5 9.3005
R93 VPWR.n35 VPWR.n4 9.3005
R94 VPWR.n37 VPWR.n36 9.3005
R95 VPWR.n39 VPWR.n38 9.3005
R96 VPWR.n40 VPWR.n2 9.3005
R97 VPWR.n44 VPWR.n43 9.3005
R98 VPWR.n45 VPWR.n1 9.3005
R99 VPWR.n47 VPWR.n46 9.3005
R100 VPWR.n48 VPWR.n0 9.3005
R101 VPWR.n21 VPWR.n9 7.90638
R102 VPWR.n14 VPWR.n12 7.29491
R103 VPWR.n36 VPWR.n3 6.02403
R104 VPWR.n39 VPWR.n3 5.27109
R105 VPWR.n15 VPWR.n14 3.38874
R106 VPWR.n22 VPWR.n21 3.38874
R107 VPWR.n49 VPWR.n48 0.376971
R108 VPWR.n43 VPWR.n42 0.376971
R109 VPWR.n16 VPWR.n12 0.221392
R110 VPWR VPWR.n50 0.163644
R111 VPWR.n50 VPWR.n0 0.144205
R112 VPWR.n17 VPWR.n16 0.122949
R113 VPWR.n18 VPWR.n17 0.122949
R114 VPWR.n18 VPWR.n10 0.122949
R115 VPWR.n23 VPWR.n10 0.122949
R116 VPWR.n24 VPWR.n23 0.122949
R117 VPWR.n25 VPWR.n24 0.122949
R118 VPWR.n25 VPWR.n8 0.122949
R119 VPWR.n8 VPWR.n7 0.122949
R120 VPWR.n30 VPWR.n7 0.122949
R121 VPWR.n31 VPWR.n30 0.122949
R122 VPWR.n32 VPWR.n31 0.122949
R123 VPWR.n32 VPWR.n5 0.122949
R124 VPWR.n5 VPWR.n4 0.122949
R125 VPWR.n37 VPWR.n4 0.122949
R126 VPWR.n38 VPWR.n37 0.122949
R127 VPWR.n38 VPWR.n2 0.122949
R128 VPWR.n44 VPWR.n2 0.122949
R129 VPWR.n45 VPWR.n44 0.122949
R130 VPWR.n46 VPWR.n45 0.122949
R131 VPWR.n46 VPWR.n0 0.122949
R132 DE.n0 DE.t1 310.087
R133 DE.n1 DE.t2 294.021
R134 DE.n2 DE.n0 277.954
R135 DE DE.n2 155.298
R136 DE.n1 DE.t3 131.748
R137 DE.n0 DE.t0 126.927
R138 DE.n2 DE.n1 36.5157
R139 a_159_446.t1 a_159_446.n1 685.008
R140 a_159_446.n1 a_159_446.t3 434.969
R141 a_159_446.n0 a_159_446.t2 340.074
R142 a_159_446.n0 a_159_446.t0 284.969
R143 a_159_446.n1 a_159_446.n0 39.6891
R144 VGND.n9 VGND.t3 291.312
R145 VGND.n34 VGND.t5 244.976
R146 VGND.n32 VGND.n2 210.018
R147 VGND.n4 VGND.t1 172.618
R148 VGND.n10 VGND.t0 162.621
R149 VGND.n27 VGND.t6 152.814
R150 VGND.n2 VGND.t2 40.0005
R151 VGND.n2 VGND.t4 40.0005
R152 VGND.n13 VGND.n8 36.1417
R153 VGND.n14 VGND.n13 36.1417
R154 VGND.n15 VGND.n6 36.1417
R155 VGND.n19 VGND.n6 36.1417
R156 VGND.n20 VGND.n19 36.1417
R157 VGND.n21 VGND.n20 36.1417
R158 VGND.n26 VGND.n25 36.1417
R159 VGND.n28 VGND.n1 36.1417
R160 VGND.n21 VGND.n4 34.2593
R161 VGND.n28 VGND.n27 30.4946
R162 VGND.n34 VGND.n33 24.8476
R163 VGND.n33 VGND.n32 24.0946
R164 VGND.n32 VGND.n1 23.3417
R165 VGND.n25 VGND.n4 19.2005
R166 VGND.n15 VGND.n14 17.3181
R167 VGND.n9 VGND.n8 15.8123
R168 VGND.n33 VGND.n0 9.3005
R169 VGND.n32 VGND.n31 9.3005
R170 VGND.n30 VGND.n1 9.3005
R171 VGND.n29 VGND.n28 9.3005
R172 VGND.n26 VGND.n3 9.3005
R173 VGND.n25 VGND.n24 9.3005
R174 VGND.n11 VGND.n8 9.3005
R175 VGND.n13 VGND.n12 9.3005
R176 VGND.n14 VGND.n7 9.3005
R177 VGND.n16 VGND.n15 9.3005
R178 VGND.n17 VGND.n6 9.3005
R179 VGND.n19 VGND.n18 9.3005
R180 VGND.n20 VGND.n5 9.3005
R181 VGND.n22 VGND.n21 9.3005
R182 VGND.n23 VGND.n4 9.3005
R183 VGND.n10 VGND.n9 9.15597
R184 VGND.n35 VGND.n34 7.09071
R185 VGND.n27 VGND.n26 5.64756
R186 VGND VGND.n35 0.273695
R187 VGND.n35 VGND.n0 0.157083
R188 VGND.n11 VGND.n10 0.14978
R189 VGND.n12 VGND.n11 0.122949
R190 VGND.n12 VGND.n7 0.122949
R191 VGND.n16 VGND.n7 0.122949
R192 VGND.n17 VGND.n16 0.122949
R193 VGND.n18 VGND.n17 0.122949
R194 VGND.n18 VGND.n5 0.122949
R195 VGND.n22 VGND.n5 0.122949
R196 VGND.n23 VGND.n22 0.122949
R197 VGND.n24 VGND.n23 0.122949
R198 VGND.n24 VGND.n3 0.122949
R199 VGND.n29 VGND.n3 0.122949
R200 VGND.n30 VGND.n29 0.122949
R201 VGND.n31 VGND.n30 0.122949
R202 VGND.n31 VGND.n0 0.122949
R203 VNB.n0 VNB 10601.6
R204 VNB VNB.n1 8498.63
R205 VNB.t4 VNB.t2 5739.63
R206 VNB.t6 VNB.t8 5173.75
R207 VNB.t8 VNB.t4 2309.71
R208 VNB.t5 VNB.t3 2286.61
R209 VNB.t9 VNB.t10 2263.52
R210 VNB.t3 VNB.t6 2228.87
R211 VNB.t11 VNB.n0 2049.32
R212 VNB.n1 VNB.t0 1813.12
R213 VNB.t1 VNB 1339.63
R214 VNB.t7 VNB.t9 993.177
R215 VNB.t10 VNB.t1 900.788
R216 VNB.t0 VNB.t7 831.496
R217 VNB.n1 VNB.t11 518.356
R218 VNB.n0 VNB.t5 288.714
R219 a_533_61.n1 a_533_61.n0 628.207
R220 a_533_61.t0 a_533_61.n3 367.466
R221 a_533_61.n2 a_533_61.t1 225.655
R222 a_533_61.n3 a_533_61.n1 193.244
R223 a_533_61.n2 a_533_61.t2 159.246
R224 a_533_61.n1 a_533_61.t3 138.441
R225 a_533_61.n3 a_533_61.n2 129.281
R226 a_554_436.t0 a_554_436.t1 112.572
R227 a_27_508.n1 a_27_508.t5 721.691
R228 a_27_508.n2 a_27_508.t1 673.095
R229 a_27_508.n0 a_27_508.t3 655.357
R230 a_27_508.t0 a_27_508.n2 338.022
R231 a_27_508.n1 a_27_508.t4 316.529
R232 a_27_508.n0 a_27_508.t2 312.341
R233 a_27_508.n2 a_27_508.n0 307.954
R234 a_27_508.n0 a_27_508.n1 138.436
R235 a_1156_90.n3 a_1156_90.n0 647.39
R236 a_1156_90.n4 a_1156_90.n3 279.495
R237 a_1156_90.n2 a_1156_90.n1 269.921
R238 a_1156_90.n3 a_1156_90.n2 252.177
R239 a_1156_90.n2 a_1156_90.t4 205.922
R240 a_1156_90.t0 a_1156_90.n4 174.286
R241 a_1156_90.n0 a_1156_90.t1 70.3576
R242 a_1156_90.n0 a_1156_90.t2 70.3576
R243 a_1156_90.n4 a_1156_90.t3 58.5719
R244 a_958_74.t1 a_958_74.n4 864.818
R245 a_958_74.n1 a_958_74.t4 565.924
R246 a_958_74.n4 a_958_74.t2 361.568
R247 a_958_74.n1 a_958_74.n0 330.341
R248 a_958_74.n2 a_958_74.t3 285.925
R249 a_958_74.n2 a_958_74.n1 261.635
R250 a_958_74.n3 a_958_74.t0 212.255
R251 a_958_74.n4 a_958_74.n3 117.082
R252 a_958_74.n3 a_958_74.n2 111.059
R253 CLK.n0 CLK.t1 321.973
R254 CLK.n0 CLK.t0 176.03
R255 CLK CLK.n0 158.788
R256 a_114_508.t0 a_114_508.t1 112.572
R257 a_131_74.t0 a_131_74.t1 68.5719
R258 D.n0 D.t1 242.875
R259 D D.n0 160.254
R260 D.n1 D 154.19
R261 D.n1 D.t0 152.633
R262 D.n3 D.n2 152
R263 D.n2 D.n0 49.6611
R264 D.n2 D.n1 49.6611
R265 D.n3 D 9.26366
R266 D D.n3 3.2005
R267 a_491_87.t0 a_491_87.t1 60.0005
R268 Q.n1 Q 589.85
R269 Q.n1 Q.n0 585
R270 Q.n2 Q.n1 585
R271 Q Q.t0 171.577
R272 Q.n1 Q.t1 26.3844
R273 Q Q.n2 12.9944
R274 Q Q.n0 11.249
R275 Q Q.n0 3.10353
R276 Q.n2 Q 1.35808
R277 a_2088_502.t0 a_2088_502.t1 126.644
C0 VGND Q 0.103599f
C1 VPB D 0.090405f
C2 VPB VPWR 0.429191f
C3 a_1797_74# VGND 0.010821f
C4 VPB DE 0.15749f
C5 D VPWR 0.014401f
C6 a_1997_74# VGND 0.006222f
C7 D DE 0.036346f
C8 VPB CLK 0.060061f
C9 VPWR DE 0.020031f
C10 VPB VGND 0.014745f
C11 VPWR CLK 0.011408f
C12 D VGND 0.02154f
C13 VPB Q 0.013186f
C14 DE CLK 9.88e-19
C15 VPWR VGND 0.06855f
C16 VPWR Q 0.128422f
C17 DE VGND 0.035562f
C18 CLK VGND 0.0351f
C19 Q VNB 0.035441f
C20 VGND VNB 1.55592f
C21 CLK VNB 0.144759f
C22 DE VNB 0.294416f
C23 VPWR VNB 1.1995f
C24 D VNB 0.196427f
C25 VPB VNB 2.98771f
.ends

* NGSPICE file created from sky130_fd_sc_hs__edfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__edfxbp_1 VNB VPB VPWR VGND CLK Q D DE Q_N
X0 Q_N.t0 a_575_48.t2 VPWR.t9 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_1198_97.t0 a_818_74.t2 a_27_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
X2 a_527_74.t1 a_161_446.t2 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3 a_818_74.t0 CLK.t0 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 VPWR.t10 a_575_48.t3 a_2206_443.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2459 pd=1.805 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 VPWR.t3 a_1879_74.t3 Q.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 a_2206_443.t0 a_1008_74.t2 a_1879_74.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.17375 ps=1.42 w=0.42 l=0.15
X7 Q_N.t1 a_575_48.t4 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2257 ps=1.35 w=0.74 l=0.15
X8 a_116_508.t1 D.t0 a_27_74.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.1239 ps=1.43 w=0.42 l=0.15
X9 VGND.t6 a_575_48.t5 a_2227_118.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1451 pd=1.145 as=0.0504 ps=0.66 w=0.42 l=0.15
X10 a_575_48.t1 a_1879_74.t4 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2459 ps=1.805 w=1 l=0.15
X11 a_818_74.t1 CLK.t1 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X12 VGND.t2 a_1419_71.t2 a_1334_97.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1388 pd=1.17 as=0.08925 ps=0.845 w=0.42 l=0.15
X13 VPWR.t2 a_1419_71.t3 a_1423_508# VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.188425 pd=1.545 as=0.0756 ps=0.78 w=0.42 l=0.15
X14 VGND.t5 DE.t0 a_161_446.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.1281 ps=1.45 w=0.42 l=0.15
X15 a_1008_74.t1 a_818_74.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X16 a_1879_74.t2 a_818_74.t4 a_2008_392.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.17375 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR.t11 DE.t1 a_161_446.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.14045 pd=1.17 as=0.1888 ps=1.87 w=0.64 l=0.15
X18 a_2227_118.t0 a_818_74.t5 a_1879_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.3739 ps=2.33 w=0.42 l=0.15
X19 a_27_74.t5 a_575_48.t6 a_556_504.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.0504 ps=0.66 w=0.42 l=0.15
X20 a_145_74.t1 D.t1 a_27_74.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1848 ps=1.72 w=0.42 l=0.15
X21 a_1419_71.t1 a_1198_97.t3 VGND.t9 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1388 ps=1.17 w=0.64 l=0.15
X22 a_27_74.t4 a_575_48.t7 a_527_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 a_575_48.t0 a_1879_74.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1451 ps=1.145 w=0.64 l=0.15
X24 a_556_504.t0 DE.t2 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.14045 ps=1.17 w=0.42 l=0.15
X25 a_1334_97.t0 a_1008_74.t3 a_1198_97.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.08925 pd=0.845 as=0.1113 ps=0.95 w=0.42 l=0.15
X26 a_1198_97.t2 a_1008_74.t4 a_27_74.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.206 ps=1.92 w=0.42 l=0.15
X27 VGND.t1 a_1879_74.t6 Q.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=1.35 as=0.2109 ps=2.05 w=0.74 l=0.15
X28 a_1008_74.t0 a_818_74.t6 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X29 a_2008_392.t1 a_1419_71.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X30 VPWR.t7 a_161_446.t3 a_116_508.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.0504 ps=0.66 w=0.42 l=0.15
X31 a_1419_71.t0 a_1198_97.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.188425 ps=1.545 w=0.84 l=0.15
X32 VGND.t10 DE.t3 a_145_74.t0 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_575_48.n1 a_575_48.n0 317.897
R1 a_575_48.n4 a_575_48.t5 297.233
R2 a_575_48.n2 a_575_48.t6 274.089
R3 a_575_48.n0 a_575_48.t2 258.942
R4 a_575_48.t1 a_575_48.n5 252.619
R5 a_575_48.n5 a_575_48.n4 205.374
R6 a_575_48.n0 a_575_48.t4 204.048
R7 a_575_48.n2 a_575_48.t7 192.43
R8 a_575_48.n1 a_575_48.t0 126.035
R9 a_575_48.n4 a_575_48.t3 116.691
R10 a_575_48.n3 a_575_48.n2 65.9123
R11 a_575_48.n5 a_575_48.n3 45.5278
R12 a_575_48.n3 a_575_48.n1 37.6456
R13 VPWR.n42 VPWR.t5 882.111
R14 VPWR.n6 VPWR.t8 860.485
R15 VPWR.n0 VPWR.t7 682.237
R16 VPWR.n30 VPWR.n29 646.139
R17 VPWR.n48 VPWR.n3 612.393
R18 VPWR.n16 VPWR.n15 261.075
R19 VPWR.n22 VPWR.t1 251.806
R20 VPWR.n14 VPWR.n13 239.198
R21 VPWR.n15 VPWR.t10 160.605
R22 VPWR.n3 VPWR.t11 157.279
R23 VPWR.n15 VPWR.t4 149.475
R24 VPWR.n29 VPWR.t2 110.227
R25 VPWR.n29 VPWR.t0 78.566
R26 VPWR.n3 VPWR.t6 70.3576
R27 VPWR.n50 VPWR.n49 36.1417
R28 VPWR.n47 VPWR.n4 36.1417
R29 VPWR.n41 VPWR.n40 36.1417
R30 VPWR.n43 VPWR.n41 36.1417
R31 VPWR.n31 VPWR.n8 36.1417
R32 VPWR.n35 VPWR.n8 36.1417
R33 VPWR.n36 VPWR.n35 36.1417
R34 VPWR.n37 VPWR.n36 36.1417
R35 VPWR.n23 VPWR.n10 36.1417
R36 VPWR.n27 VPWR.n10 36.1417
R37 VPWR.n17 VPWR.n12 36.1417
R38 VPWR.n21 VPWR.n12 36.1417
R39 VPWR.n50 VPWR.n0 35.7652
R40 VPWR.n48 VPWR.n47 35.7652
R41 VPWR.n22 VPWR.n21 31.2476
R42 VPWR.n28 VPWR.n27 30.7716
R43 VPWR.n13 VPWR.t9 26.3844
R44 VPWR.n13 VPWR.t3 26.3844
R45 VPWR.n31 VPWR.n30 23.1854
R46 VPWR.n49 VPWR.n48 17.6946
R47 VPWR.n23 VPWR.n22 16.1887
R48 VPWR.n17 VPWR.n16 16.1887
R49 VPWR.n18 VPWR.n17 9.3005
R50 VPWR.n19 VPWR.n12 9.3005
R51 VPWR.n21 VPWR.n20 9.3005
R52 VPWR.n22 VPWR.n11 9.3005
R53 VPWR.n24 VPWR.n23 9.3005
R54 VPWR.n25 VPWR.n10 9.3005
R55 VPWR.n27 VPWR.n26 9.3005
R56 VPWR.n28 VPWR.n9 9.3005
R57 VPWR.n32 VPWR.n31 9.3005
R58 VPWR.n33 VPWR.n8 9.3005
R59 VPWR.n35 VPWR.n34 9.3005
R60 VPWR.n36 VPWR.n7 9.3005
R61 VPWR.n38 VPWR.n37 9.3005
R62 VPWR.n40 VPWR.n39 9.3005
R63 VPWR.n41 VPWR.n5 9.3005
R64 VPWR.n44 VPWR.n43 9.3005
R65 VPWR.n45 VPWR.n4 9.3005
R66 VPWR.n47 VPWR.n46 9.3005
R67 VPWR.n48 VPWR.n2 9.3005
R68 VPWR.n49 VPWR.n1 9.3005
R69 VPWR.n51 VPWR.n50 9.3005
R70 VPWR.n42 VPWR.n4 8.65932
R71 VPWR.n52 VPWR.n0 6.78023
R72 VPWR.n37 VPWR.n6 6.4005
R73 VPWR.n40 VPWR.n6 4.89462
R74 VPWR.n16 VPWR.n14 4.10254
R75 VPWR.n43 VPWR.n42 2.63579
R76 VPWR.n30 VPWR.n28 1.44956
R77 VPWR VPWR.n52 0.268898
R78 VPWR.n18 VPWR.n14 0.235192
R79 VPWR.n52 VPWR.n51 0.161808
R80 VPWR.n19 VPWR.n18 0.122949
R81 VPWR.n20 VPWR.n19 0.122949
R82 VPWR.n20 VPWR.n11 0.122949
R83 VPWR.n24 VPWR.n11 0.122949
R84 VPWR.n25 VPWR.n24 0.122949
R85 VPWR.n26 VPWR.n25 0.122949
R86 VPWR.n26 VPWR.n9 0.122949
R87 VPWR.n32 VPWR.n9 0.122949
R88 VPWR.n33 VPWR.n32 0.122949
R89 VPWR.n34 VPWR.n33 0.122949
R90 VPWR.n34 VPWR.n7 0.122949
R91 VPWR.n38 VPWR.n7 0.122949
R92 VPWR.n39 VPWR.n38 0.122949
R93 VPWR.n39 VPWR.n5 0.122949
R94 VPWR.n44 VPWR.n5 0.122949
R95 VPWR.n45 VPWR.n44 0.122949
R96 VPWR.n46 VPWR.n45 0.122949
R97 VPWR.n46 VPWR.n2 0.122949
R98 VPWR.n2 VPWR.n1 0.122949
R99 VPWR.n51 VPWR.n1 0.122949
R100 Q_N.n0 Q_N.t0 293.048
R101 Q_N.t1 Q_N.n0 279.738
R102 Q_N.n1 Q_N.t1 279.738
R103 Q_N.n1 Q_N 10.8449
R104 Q_N.n0 Q_N 5.15606
R105 Q_N Q_N.n1 2.31161
R106 VPB.t0 VPB.t2 916.802
R107 VPB.t7 VPB.t12 709.947
R108 VPB.t9 VPB.t16 577.152
R109 VPB.t12 VPB.t10 559.274
R110 VPB.t5 VPB.t4 515.861
R111 VPB.t13 VPB.t7 515.861
R112 VPB.t10 VPB.t3 490.324
R113 VPB.t14 VPB.t5 487.769
R114 VPB.t16 VPB.t8 347.312
R115 VPB.t3 VPB.t0 316.668
R116 VPB.t11 VPB.t1 291.13
R117 VPB VPB.t6 257.93
R118 VPB.t1 VPB.t14 245.161
R119 VPB.t4 VPB.t15 229.839
R120 VPB.t2 VPB.t11 214.517
R121 VPB.t8 VPB.t13 199.195
R122 VPB.t6 VPB.t9 199.195
R123 a_818_74.t1 a_818_74.n6 850.788
R124 a_818_74.n2 a_818_74.n1 636.574
R125 a_818_74.n3 a_818_74.n2 388.813
R126 a_818_74.n1 a_818_74.t5 351.861
R127 a_818_74.n3 a_818_74.t2 292.413
R128 a_818_74.n5 a_818_74.t3 286.88
R129 a_818_74.n1 a_818_74.t4 234.306
R130 a_818_74.n6 a_818_74.t0 218.083
R131 a_818_74.n4 a_818_74.t6 204.048
R132 a_818_74.n6 a_818_74.n5 193.315
R133 a_818_74.n5 a_818_74.n4 146.208
R134 a_818_74.n2 a_818_74.n0 138.441
R135 a_818_74.n4 a_818_74.n3 134.96
R136 a_27_74.n2 a_27_74.t3 810.076
R137 a_27_74.n1 a_27_74.t1 668.691
R138 a_27_74.n0 a_27_74.t5 666.352
R139 a_27_74.n1 a_27_74.t2 354.255
R140 a_27_74.n0 a_27_74.t4 347.435
R141 a_27_74.t0 a_27_74.n2 337.942
R142 a_27_74.n0 a_27_74.n1 271.06
R143 a_27_74.n2 a_27_74.n0 132.798
R144 a_1198_97.n1 a_1198_97.t2 718.845
R145 a_1198_97.n0 a_1198_97.t3 326.154
R146 a_1198_97.n2 a_1198_97.n1 265.188
R147 a_1198_97.n1 a_1198_97.n0 256.32
R148 a_1198_97.n0 a_1198_97.t4 207.261
R149 a_1198_97.t0 a_1198_97.n2 111.43
R150 a_1198_97.n2 a_1198_97.t1 40.0005
R151 VNB.n0 VNB 27633.9
R152 VNB.n1 VNB 13962.2
R153 VNB VNB.n2 11481.8
R154 VNB.t14 VNB.t3 7414.17
R155 VNB.t6 VNB.t11 2459.84
R156 VNB.t0 VNB.t1 2421.16
R157 VNB.t7 VNB.t15 2332.81
R158 VNB.t4 VNB.t5 2205.8
R159 VNB.n2 VNB.t6 2148.03
R160 VNB.t1 VNB.t13 1769.31
R161 VNB.t2 VNB.t14 1570.6
R162 VNB.t8 VNB 1501.31
R163 VNB.t9 VNB.t2 1328.08
R164 VNB.n1 VNB.t9 1270.34
R165 VNB.t10 VNB.t7 1177.95
R166 VNB.t12 VNB.n0 970.08
R167 VNB.t3 VNB.t12 900.788
R168 VNB.t11 VNB.t10 900.788
R169 VNB.t15 VNB.t8 900.788
R170 VNB.n0 VNB.t0 547.091
R171 VNB.t5 VNB.n1 301.848
R172 VNB.n2 VNB.t4 23.1584
R173 a_161_446.t1 a_161_446.n1 660.16
R174 a_161_446.n0 a_161_446.t3 307.954
R175 a_161_446.n1 a_161_446.t2 305.055
R176 a_161_446.n0 a_161_446.t0 295.231
R177 a_161_446.n1 a_161_446.n0 43.5801
R178 VGND.n39 VGND.t3 292.372
R179 VGND.n51 VGND.t10 247.498
R180 VGND.n9 VGND.n8 217.256
R181 VGND.n2 VGND.n1 207.498
R182 VGND.n4 VGND.t4 152.814
R183 VGND.n17 VGND.n16 141.637
R184 VGND.n15 VGND.n14 117.859
R185 VGND.n8 VGND.t9 96.6123
R186 VGND.n14 VGND.t6 88.4533
R187 VGND.n16 VGND.t1 76.2167
R188 VGND.n1 VGND.t5 60.0005
R189 VGND.n1 VGND.t8 42.8576
R190 VGND.n8 VGND.t2 40.0005
R191 VGND.n14 VGND.t0 37.976
R192 VGND.n20 VGND.n13 36.1417
R193 VGND.n21 VGND.n20 36.1417
R194 VGND.n22 VGND.n21 36.1417
R195 VGND.n22 VGND.n11 36.1417
R196 VGND.n28 VGND.n27 36.1417
R197 VGND.n33 VGND.n32 36.1417
R198 VGND.n34 VGND.n33 36.1417
R199 VGND.n34 VGND.n6 36.1417
R200 VGND.n38 VGND.n6 36.1417
R201 VGND.n41 VGND.n40 36.1417
R202 VGND.n45 VGND.n44 36.1417
R203 VGND.n46 VGND.n45 36.1417
R204 VGND.n50 VGND.n49 36.1417
R205 VGND.n26 VGND.n11 33.8829
R206 VGND.n28 VGND.n9 33.8829
R207 VGND.n15 VGND.n13 28.2358
R208 VGND.n16 VGND.t7 22.7032
R209 VGND.n41 VGND.n4 21.0829
R210 VGND.n27 VGND.n26 19.577
R211 VGND.n32 VGND.n9 19.577
R212 VGND.n51 VGND.n50 19.577
R213 VGND.n44 VGND.n4 15.0593
R214 VGND.n46 VGND.n2 10.5417
R215 VGND.n39 VGND.n38 9.41227
R216 VGND.n50 VGND.n0 9.3005
R217 VGND.n49 VGND.n48 9.3005
R218 VGND.n47 VGND.n46 9.3005
R219 VGND.n45 VGND.n3 9.3005
R220 VGND.n44 VGND.n43 9.3005
R221 VGND.n42 VGND.n41 9.3005
R222 VGND.n40 VGND.n5 9.3005
R223 VGND.n38 VGND.n37 9.3005
R224 VGND.n36 VGND.n6 9.3005
R225 VGND.n35 VGND.n34 9.3005
R226 VGND.n33 VGND.n7 9.3005
R227 VGND.n32 VGND.n31 9.3005
R228 VGND.n30 VGND.n9 9.3005
R229 VGND.n29 VGND.n28 9.3005
R230 VGND.n27 VGND.n10 9.3005
R231 VGND.n26 VGND.n25 9.3005
R232 VGND.n24 VGND.n11 9.3005
R233 VGND.n23 VGND.n22 9.3005
R234 VGND.n21 VGND.n12 9.3005
R235 VGND.n20 VGND.n19 9.3005
R236 VGND.n18 VGND.n13 9.3005
R237 VGND.n52 VGND.n51 7.34955
R238 VGND.n17 VGND.n15 6.86979
R239 VGND.n40 VGND.n39 1.88285
R240 VGND.n49 VGND.n2 0.753441
R241 VGND VGND.n52 0.277695
R242 VGND.n18 VGND.n17 0.171944
R243 VGND.n52 VGND.n0 0.153144
R244 VGND.n19 VGND.n18 0.122949
R245 VGND.n19 VGND.n12 0.122949
R246 VGND.n23 VGND.n12 0.122949
R247 VGND.n24 VGND.n23 0.122949
R248 VGND.n25 VGND.n24 0.122949
R249 VGND.n25 VGND.n10 0.122949
R250 VGND.n29 VGND.n10 0.122949
R251 VGND.n30 VGND.n29 0.122949
R252 VGND.n31 VGND.n30 0.122949
R253 VGND.n31 VGND.n7 0.122949
R254 VGND.n35 VGND.n7 0.122949
R255 VGND.n36 VGND.n35 0.122949
R256 VGND.n37 VGND.n36 0.122949
R257 VGND.n37 VGND.n5 0.122949
R258 VGND.n42 VGND.n5 0.122949
R259 VGND.n43 VGND.n42 0.122949
R260 VGND.n43 VGND.n3 0.122949
R261 VGND.n47 VGND.n3 0.122949
R262 VGND.n48 VGND.n47 0.122949
R263 VGND.n48 VGND.n0 0.122949
R264 a_527_74.t0 a_527_74.t1 68.5719
R265 CLK.n0 CLK.t1 267.973
R266 CLK.n0 CLK.t0 160.561
R267 CLK CLK.n0 84.9017
R268 a_2206_443.t0 a_2206_443.t1 154.786
R269 a_1879_74.n7 a_1879_74.n5 645.102
R270 a_1879_74.n8 a_1879_74.n0 611.739
R271 a_1879_74.n6 a_1879_74.n0 585
R272 a_1879_74.n1 a_1879_74.t3 310.639
R273 a_1879_74.n2 a_1879_74.t4 251.177
R274 a_1879_74.n4 a_1879_74.n3 200.802
R275 a_1879_74.n4 a_1879_74.t1 178.575
R276 a_1879_74.n3 a_1879_74.t5 152.163
R277 a_1879_74.n1 a_1879_74.t6 142.994
R278 a_1879_74.n2 a_1879_74.n1 131.113
R279 a_1879_74.n6 a_1879_74.t0 126.644
R280 a_1879_74.n8 a_1879_74.n7 106.847
R281 a_1879_74.n5 a_1879_74.n4 83.828
R282 a_1879_74.n3 a_1879_74.n2 55.2304
R283 a_1879_74.n7 a_1879_74.t2 34.0462
R284 a_1879_74.n5 a_1879_74.n0 13.3823
R285 a_1879_74.n7 a_1879_74.n6 2.34574
R286 Q.n1 Q 588.856
R287 Q.n1 Q.n0 585
R288 Q.n2 Q.n1 585
R289 Q Q.t1 280.824
R290 Q.n1 Q.t0 26.3844
R291 Q Q.n2 10.333
R292 Q Q.n0 8.94508
R293 Q Q.n0 2.46797
R294 Q.n2 Q 1.08002
R295 a_1008_74.t0 a_1008_74.n4 871.251
R296 a_1008_74.n1 a_1008_74.n0 458.873
R297 a_1008_74.n1 a_1008_74.t2 441.981
R298 a_1008_74.n4 a_1008_74.t4 365.815
R299 a_1008_74.n2 a_1008_74.n1 294.651
R300 a_1008_74.n2 a_1008_74.t3 283.272
R301 a_1008_74.n3 a_1008_74.t1 210.272
R302 a_1008_74.n4 a_1008_74.n3 116.707
R303 a_1008_74.n3 a_1008_74.n2 81.1525
R304 D.n0 D.t0 242.167
R305 D D.n0 159.649
R306 D.n1 D 154.03
R307 D.n3 D.n2 152
R308 D.n1 D.t1 151.924
R309 D.n2 D.n0 48.2005
R310 D.n2 D.n1 48.2005
R311 D.n3 D 8.58587
R312 D D.n3 2.96635
R313 a_116_508.t0 a_116_508.t1 112.572
R314 a_2227_118.t0 a_2227_118.t1 68.5719
R315 a_1419_71.t0 a_1419_71.n6 771.303
R316 a_1419_71.n0 a_1419_71.t4 483.608
R317 a_1419_71.n1 a_1419_71.t3 380.197
R318 a_1419_71.n1 a_1419_71.t2 299.087
R319 a_1419_71.n4 a_1419_71.n3 292.055
R320 a_1419_71.n2 a_1419_71.t1 248.522
R321 a_1419_71.n2 a_1419_71.n1 199.876
R322 a_1419_71.n5 a_1419_71.n4 152
R323 a_1419_71.n6 a_1419_71.n0 125.004
R324 a_1419_71.n5 a_1419_71.n2 61.388
R325 a_1419_71.n6 a_1419_71.n5 15.9265
R326 a_1419_71.n4 a_1419_71.n0 10.0721
R327 a_1334_97.t0 a_1334_97.t1 121.43
R328 DE.n0 DE.t2 350.789
R329 DE.n1 DE.t3 287.594
R330 DE.n1 DE.t0 220.113
R331 DE.n0 DE.t1 183.161
R332 DE DE.n2 157.625
R333 DE.n2 DE.n1 154.508
R334 DE.n2 DE.n0 31.2412
R335 a_2008_392.t0 a_2008_392.t1 53.1905
R336 a_556_504.t0 a_556_504.t1 112.572
R337 a_145_74.t0 a_145_74.t1 68.5719
C0 VGND Q 0.009997f
C1 VPB VPWR 0.440885f
C2 VGND Q_N 0.101834f
C3 a_1807_74# VGND 0.007513f
C4 VPB D 0.091875f
C5 Q Q_N 0.003643f
C6 a_1423_508# VPWR 0.004047f
C7 VPB DE 0.188915f
C8 VPWR D 0.013261f
C9 VPWR DE 0.022721f
C10 VPB CLK 0.053526f
C11 D DE 0.033908f
C12 VPWR CLK 0.015875f
C13 VPB VGND 0.015281f
C14 VPB Q 0.0189f
C15 VPWR VGND 0.07784f
C16 D VGND 0.019681f
C17 VPB Q_N 0.016752f
C18 VPWR Q 0.141706f
C19 VPWR Q_N 0.128318f
C20 DE VGND 0.04361f
C21 CLK VGND 0.035833f
C22 Q_N VNB 0.113084f
C23 Q VNB 0.007802f
C24 VGND VNB 1.69426f
C25 CLK VNB 0.161773f
C26 DE VNB 0.314318f
C27 D VNB 0.201141f
C28 VPWR VNB 1.2663f
C29 VPB VNB 3.30214f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ebufn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ebufn_8 VNB VPB VPWR VGND TE_B A Z
X0 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 ad=0.28785 pd=1.76 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Z.t15 a_84_48.t3 a_28_368# VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_28_368# TE_B.t0 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X3 Z.t4 a_84_48.t4 a_27_74.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12395 pd=1.075 as=0.13505 ps=1.105 w=0.74 l=0.15
X4 VGND.t6 a_833_48.t1 a_27_74.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_84_48.t1 A.t0 VPWR.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6 Z.t3 a_84_48.t5 a_27_74.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 a_28_368# TE_B.t1 VPWR.t6 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X8 Z.t14 a_84_48.t6 a_28_368# VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X9 VPWR.t5 TE_B.t2 a_28_368# VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_28_368# a_84_48.t7 Z.t13 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
X11 Z.t2 a_84_48.t8 a_27_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11285 ps=1.045 w=0.74 l=0.15
X12 Z.t1 a_84_48.t9 a_27_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 a_27_74.t12 a_833_48.t2 VGND.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_28_368# a_84_48.t10 Z.t12 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Z.t11 a_84_48.t11 a_28_368# VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VPWR.t2 TE_B.t3 a_833_48.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.5712 ps=3.26 w=1.12 l=0.15
X17 a_27_74.t3 a_84_48.t12 Z.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12395 ps=1.075 w=0.74 l=0.15
X18 a_27_74.t8 a_833_48.t3 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_27_74.t2 a_84_48.t13 Z.t7 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_28_368# a_84_48.t14 Z.t10 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X21 a_27_74.t13 a_833_48.t4 VGND.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_27_74.t10 a_833_48.t5 VGND.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_28_368# TE_B.t4 VPWR.t4 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X25 VPWR.t3 TE_B.t5 a_28_368# VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.1764 ps=1.435 w=1.12 l=0.15
X26 a_27_74.t1 a_84_48.t15 Z.t6 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 Z.t9 a_84_48.t16 a_28_368# VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X28 a_28_368# a_84_48.t17 Z.t8 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 VPWR.t1 A.t1 a_84_48.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.28785 ps=1.76 w=1.12 l=0.15
X31 VGND.t1 a_833_48.t6 a_27_74.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 a_27_74.t0 a_84_48.t18 Z.t5 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.13505 pd=1.105 as=0.1295 ps=1.09 w=0.74 l=0.15
X33 a_84_48.t0 A.t2 VGND.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 TE_B.n9 TE_B.t5 380.781
R1 TE_B.n15 TE_B.n6 204.048
R2 TE_B.n14 TE_B.n7 204.048
R3 TE_B.n13 TE_B.t0 204.048
R4 TE_B.n12 TE_B.n8 204.048
R5 TE_B.n11 TE_B.t4 204.048
R6 TE_B.n10 TE_B.t2 204.048
R7 TE_B.n9 TE_B.t1 204.048
R8 TE_B.n4 TE_B.t3 204.048
R9 TE_B.n15 TE_B.n14 199.227
R10 TE_B.n13 TE_B.n12 176.733
R11 TE_B.n11 TE_B.n10 176.733
R12 TE_B.n3 TE_B.n1 170.595
R13 TE_B.n3 TE_B.n2 152
R14 TE_B.n5 TE_B.n0 152
R15 TE_B.n17 TE_B.n16 152
R16 TE_B.n14 TE_B.n13 144.601
R17 TE_B.n12 TE_B.n11 144.601
R18 TE_B.n10 TE_B.n9 144.601
R19 TE_B.n16 TE_B.n15 138.306
R20 TE_B.n16 TE_B.n5 30.0702
R21 TE_B.n5 TE_B.n4 29.628
R22 TE_B.n17 TE_B.n0 11.7627
R23 TE_B.n2 TE_B 10.8978
R24 TE_B.n2 TE_B 5.70861
R25 TE_B TE_B.n17 3.97888
R26 TE_B TE_B.n0 0.865365
R27 TE_B.n4 TE_B.n3 0.442702
R28 VPWR.n4 VPWR.t7 809.364
R29 VPWR.n9 VPWR.n8 608.662
R30 VPWR.n23 VPWR.n1 604.976
R31 VPWR.n21 VPWR.n3 604.976
R32 VPWR.n7 VPWR.t1 254.802
R33 VPWR.n10 VPWR.n6 36.1417
R34 VPWR.n14 VPWR.n6 36.1417
R35 VPWR.n1 VPWR.t6 35.1791
R36 VPWR.n1 VPWR.t3 35.1791
R37 VPWR.n3 VPWR.t4 35.1791
R38 VPWR.n3 VPWR.t5 35.1791
R39 VPWR.n8 VPWR.t0 35.1791
R40 VPWR.n16 VPWR.n15 33.5064
R41 VPWR.n20 VPWR.n4 27.8593
R42 VPWR.n8 VPWR.t2 26.3844
R43 VPWR.n23 VPWR.n22 25.6005
R44 VPWR.n22 VPWR.n21 24.8476
R45 VPWR.n21 VPWR.n20 22.5887
R46 VPWR.n10 VPWR.n9 21.4593
R47 VPWR.n16 VPWR.n4 19.577
R48 VPWR.n15 VPWR.n14 13.9299
R49 VPWR.n11 VPWR.n10 9.3005
R50 VPWR.n12 VPWR.n6 9.3005
R51 VPWR.n14 VPWR.n13 9.3005
R52 VPWR.n15 VPWR.n5 9.3005
R53 VPWR.n17 VPWR.n16 9.3005
R54 VPWR.n18 VPWR.n4 9.3005
R55 VPWR.n20 VPWR.n19 9.3005
R56 VPWR.n21 VPWR.n2 9.3005
R57 VPWR.n22 VPWR.n0 9.3005
R58 VPWR.n24 VPWR.n23 7.04398
R59 VPWR.n9 VPWR.n7 6.75308
R60 VPWR VPWR.n24 1.13296
R61 VPWR.n11 VPWR.n7 0.636608
R62 VPWR.n24 VPWR.n0 0.159033
R63 VPWR.n12 VPWR.n11 0.122949
R64 VPWR.n13 VPWR.n12 0.122949
R65 VPWR.n13 VPWR.n5 0.122949
R66 VPWR.n17 VPWR.n5 0.122949
R67 VPWR.n18 VPWR.n17 0.122949
R68 VPWR.n19 VPWR.n18 0.122949
R69 VPWR.n19 VPWR.n2 0.122949
R70 VPWR.n2 VPWR.n0 0.122949
R71 VPB.t15 VPB.t12 1172.18
R72 VPB.t11 VPB.t15 510.753
R73 VPB.t13 VPB.t11 280.914
R74 VPB.t10 VPB.t14 280.914
R75 VPB VPB.t1 260.485
R76 VPB.t12 VPB.t8 255.376
R77 VPB.t3 VPB.t0 255.376
R78 VPB.t6 VPB.t5 255.376
R79 VPB.t0 VPB.t2 247.715
R80 VPB.t2 VPB.t10 237.5
R81 VPB.t8 VPB.t9 229.839
R82 VPB.t14 VPB.t13 229.839
R83 VPB.t4 VPB.t3 229.839
R84 VPB.t5 VPB.t4 229.839
R85 VPB.t7 VPB.t6 229.839
R86 VPB.t1 VPB.t7 229.839
R87 a_84_48.n28 a_84_48.n27 492.767
R88 a_84_48.n28 a_84_48.t0 257.301
R89 a_84_48.n1 a_84_48.t7 234.841
R90 a_84_48.n24 a_84_48.t3 234.841
R91 a_84_48.n2 a_84_48.t10 234.841
R92 a_84_48.n18 a_84_48.t11 234.841
R93 a_84_48.n15 a_84_48.t14 234.841
R94 a_84_48.n10 a_84_48.t16 234.841
R95 a_84_48.n7 a_84_48.t17 234.841
R96 a_84_48.n5 a_84_48.t6 234.841
R97 a_84_48.n29 a_84_48.n28 195.736
R98 a_84_48.n5 a_84_48.t9 188.565
R99 a_84_48.n1 a_84_48.t12 188.565
R100 a_84_48.n2 a_84_48.t18 186.374
R101 a_84_48.n6 a_84_48.t15 186.374
R102 a_84_48.n9 a_84_48.t8 186.374
R103 a_84_48.n4 a_84_48.t13 186.374
R104 a_84_48.n17 a_84_48.t5 186.374
R105 a_84_48.n25 a_84_48.t4 186.374
R106 a_84_48.n12 a_84_48.n8 165.189
R107 a_84_48.n12 a_84_48.n11 152
R108 a_84_48.n14 a_84_48.n13 152
R109 a_84_48.n16 a_84_48.n3 152
R110 a_84_48.n20 a_84_48.n19 152
R111 a_84_48.n22 a_84_48.n21 152
R112 a_84_48.n23 a_84_48.n0 152
R113 a_84_48.n27 a_84_48.n26 152
R114 a_84_48.n6 a_84_48.n5 60.6157
R115 a_84_48.n23 a_84_48.n22 49.6611
R116 a_84_48.n11 a_84_48.n4 48.2005
R117 a_84_48.n19 a_84_48.n2 45.2793
R118 a_84_48.n26 a_84_48.n1 40.1672
R119 a_84_48.n16 a_84_48.n15 36.5157
R120 a_84_48.n9 a_84_48.n8 35.055
R121 a_84_48.n26 a_84_48.n25 28.4823
R122 a_84_48.n29 a_84_48.t2 26.3844
R123 a_84_48.t1 a_84_48.n29 26.3844
R124 a_84_48.n8 a_84_48.n7 26.2914
R125 a_84_48.n17 a_84_48.n16 21.9096
R126 a_84_48.n19 a_84_48.n18 20.449
R127 a_84_48.n24 a_84_48.n23 18.9884
R128 a_84_48.n27 a_84_48.n0 13.1884
R129 a_84_48.n21 a_84_48.n0 13.1884
R130 a_84_48.n21 a_84_48.n20 13.1884
R131 a_84_48.n20 a_84_48.n3 13.1884
R132 a_84_48.n13 a_84_48.n3 13.1884
R133 a_84_48.n13 a_84_48.n12 13.1884
R134 a_84_48.n15 a_84_48.n14 13.146
R135 a_84_48.n11 a_84_48.n10 10.2247
R136 a_84_48.n18 a_84_48.n17 7.30353
R137 a_84_48.n7 a_84_48.n6 5.11262
R138 a_84_48.n22 a_84_48.n2 4.38232
R139 a_84_48.n10 a_84_48.n9 4.38232
R140 a_84_48.n25 a_84_48.n24 2.19141
R141 a_84_48.n14 a_84_48.n4 1.46111
R142 Z.n2 Z.n0 251.381
R143 Z.n9 Z.n7 251.083
R144 Z.n2 Z.n1 204.698
R145 Z.n4 Z.n3 204.698
R146 Z.n6 Z.n5 204.025
R147 Z Z.n12 188.103
R148 Z.n9 Z.n8 185
R149 Z.n11 Z.n10 185
R150 Z.n11 Z.n9 58.0584
R151 Z.n6 Z.n4 46.6829
R152 Z.n13 Z.n11 45.5941
R153 Z.n4 Z.n2 42.9181
R154 Z.n3 Z.t9 35.1791
R155 Z.n8 Z.t3 34.0546
R156 Z.n0 Z.t13 32.5407
R157 Z.n7 Z.t4 31.6221
R158 Z.n5 Z.t8 26.3844
R159 Z.n5 Z.t14 26.3844
R160 Z.n0 Z.t15 26.3844
R161 Z.n1 Z.t12 26.3844
R162 Z.n1 Z.t11 26.3844
R163 Z.n3 Z.t10 26.3844
R164 Z.n12 Z.t6 22.7032
R165 Z.n12 Z.t1 22.7032
R166 Z.n10 Z.t7 22.7032
R167 Z.n10 Z.t2 22.7032
R168 Z.n8 Z.t5 22.7032
R169 Z.n7 Z.t0 22.7032
R170 Z Z.n6 13.6584
R171 Z.n13 Z 8.72777
R172 Z Z.n13 5.94575
R173 a_27_74.n1 a_27_74.t8 212.835
R174 a_27_74.n7 a_27_74.t4 212.715
R175 a_27_74.n7 a_27_74.n6 200.435
R176 a_27_74.n9 a_27_74.n8 185
R177 a_27_74.n11 a_27_74.n10 185
R178 a_27_74.n1 a_27_74.t13 167.754
R179 a_27_74.n2 a_27_74.t10 167.754
R180 a_27_74.n3 a_27_74.n0 106.883
R181 a_27_74.n5 a_27_74.n3 88.9784
R182 a_27_74.n5 a_27_74.n4 84.741
R183 a_27_74.n10 a_27_74.n5 83.7028
R184 a_27_74.n9 a_27_74.n7 63.2883
R185 a_27_74.n10 a_27_74.n9 58.0584
R186 a_27_74.n2 a_27_74.n1 45.9299
R187 a_27_74.n3 a_27_74.n2 44.7549
R188 a_27_74.n8 a_27_74.t2 34.0546
R189 a_27_74.n11 a_27_74.t0 34.0546
R190 a_27_74.n6 a_27_74.t5 26.7573
R191 a_27_74.t7 a_27_74.n11 25.1356
R192 a_27_74.n8 a_27_74.t6 22.7032
R193 a_27_74.n6 a_27_74.t1 22.7032
R194 a_27_74.n4 a_27_74.t9 22.7032
R195 a_27_74.n4 a_27_74.t3 22.7032
R196 a_27_74.n0 a_27_74.t11 22.7032
R197 a_27_74.n0 a_27_74.t12 22.7032
R198 VNB.t8 VNB.t12 5497.11
R199 VNB.t14 VNB.t8 1986.35
R200 VNB.t10 VNB.t14 1986.35
R201 VNB.t0 VNB.t7 1189.5
R202 VNB.t6 VNB.t0 1154.86
R203 VNB.t2 VNB.t6 1154.86
R204 VNB VNB.t4 1143.31
R205 VNB.t7 VNB.t3 1120.21
R206 VNB.t1 VNB.t5 1050.92
R207 VNB.t11 VNB.t10 993.177
R208 VNB.t13 VNB.t11 993.177
R209 VNB.t9 VNB.t13 993.177
R210 VNB.t3 VNB.t9 993.177
R211 VNB.t5 VNB.t2 993.177
R212 VNB.t4 VNB.t1 993.177
R213 a_833_48.t0 a_833_48.n8 1279.23
R214 a_833_48.n2 a_833_48.t1 281.168
R215 a_833_48.n2 a_833_48.t2 142.994
R216 a_833_48.n3 a_833_48.t6 142.994
R217 a_833_48.n4 a_833_48.t5 142.994
R218 a_833_48.n5 a_833_48.n1 142.994
R219 a_833_48.n6 a_833_48.t4 142.994
R220 a_833_48.n7 a_833_48.n0 142.994
R221 a_833_48.n8 a_833_48.t3 142.994
R222 a_833_48.n8 a_833_48.n7 138.173
R223 a_833_48.n7 a_833_48.n6 138.173
R224 a_833_48.n6 a_833_48.n5 138.173
R225 a_833_48.n5 a_833_48.n4 138.173
R226 a_833_48.n4 a_833_48.n3 138.173
R227 a_833_48.n3 a_833_48.n2 138.173
R228 VGND.n4 VGND.t4 172.618
R229 VGND.n5 VGND.t3 172.618
R230 VGND.n3 VGND.t0 162.434
R231 VGND.n11 VGND.n1 132.637
R232 VGND.n14 VGND.n13 114.885
R233 VGND.n10 VGND.n2 36.1417
R234 VGND.n14 VGND.n12 31.624
R235 VGND.n6 VGND.n4 29.3652
R236 VGND.n1 VGND.t2 22.7032
R237 VGND.n1 VGND.t1 22.7032
R238 VGND.n13 VGND.t5 22.7032
R239 VGND.n13 VGND.t6 22.7032
R240 VGND.n12 VGND.n11 20.7064
R241 VGND.n6 VGND.n5 16.5652
R242 VGND.n11 VGND.n10 15.4358
R243 VGND.n12 VGND.n0 9.3005
R244 VGND.n10 VGND.n9 9.3005
R245 VGND.n8 VGND.n2 9.3005
R246 VGND.n7 VGND.n6 9.3005
R247 VGND.n4 VGND.n3 7.16629
R248 VGND.n15 VGND.n14 6.63088
R249 VGND VGND.n15 1.12634
R250 VGND.n5 VGND.n2 0.753441
R251 VGND.n15 VGND.n0 0.165546
R252 VGND.n7 VGND.n3 0.158533
R253 VGND.n8 VGND.n7 0.122949
R254 VGND.n9 VGND.n8 0.122949
R255 VGND.n9 VGND.n0 0.122949
R256 A.n2 A.t0 265.271
R257 A.n1 A.t1 261.62
R258 A A.n3 158.788
R259 A.n1 A.n0 154.97
R260 A.n2 A.t2 154.24
R261 A.n3 A.n1 35.7853
R262 A.n3 A.n2 26.2914
C0 VPB VGND 0.012602f
C1 VPB Z 0.013432f
C2 TE_B VPWR 0.120197f
C3 TE_B VGND 0.050412f
C4 VPB A 0.06077f
C5 TE_B Z 0.001453f
C6 VPWR VGND 0.171195f
C7 VPWR Z 0.044335f
C8 TE_B A 0.091099f
C9 Z VGND 0.042696f
C10 VPWR A 0.037654f
C11 A VGND 0.031405f
C12 a_28_368# VPB 0.049268f
C13 a_28_368# TE_B 0.108109f
C14 a_28_368# VPWR 0.986458f
C15 a_28_368# VGND 0.014428f
C16 a_28_368# Z 0.624513f
C17 a_28_368# A 6.68e-20
C18 VPB TE_B 0.390378f
C19 VPB VPWR 0.255402f
C20 VGND VNB 1.20618f
C21 A VNB 0.220618f
C22 Z VNB 0.042575f
C23 VPWR VNB 0.971206f
C24 TE_B VNB 0.489092f
C25 VPB VNB 2.44181f
C26 a_28_368# VNB 0.057131f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ebufn_4 VNB VPB VPWR VGND Z TE_B A
X0 VPWR.t2 A.t0 a_27_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.182 pd=1.445 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t4 a_208_74.t2 a_378_74.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2072 ps=2.04 w=0.74 l=0.15
X2 Z.t3 a_27_368.t2 a_348_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_348_368.t3 a_27_368.t3 Z.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_348_368.t4 a_27_368.t4 Z.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X5 Z.t0 a_27_368.t5 a_348_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_348_368.t5 TE_B.t0 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Z.t7 a_27_368.t6 a_378_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t5 TE_B.t1 a_348_368.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_348_368.t0 TE_B.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_208_74.t1 TE_B.t3 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_208_74.t0 TE_B.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.182 ps=1.445 w=1.12 l=0.15
X12 VGND.t0 A.t1 a_27_368.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 a_378_74.t2 a_27_368.t7 Z.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t4 TE_B.t5 a_348_368.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X15 a_378_74.t6 a_208_74.t3 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_378_74.t0 a_27_368.t8 Z.t5 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.111 ps=1.04 w=0.74 l=0.15
X17 a_378_74.t5 a_208_74.t4 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 Z.t4 a_27_368.t9 a_378_74.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 VGND.t1 a_208_74.t5 a_378_74.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t0 264.298
R1 A.n0 A.t1 204.048
R2 A A.n0 155.201
R3 a_27_368.n11 a_27_368.n10 315.048
R4 a_27_368.n8 a_27_368.t5 242.875
R5 a_27_368.n1 a_27_368.t4 234.841
R6 a_27_368.n3 a_27_368.t2 234.841
R7 a_27_368.n6 a_27_368.t3 234.841
R8 a_27_368.n11 a_27_368.t1 230.691
R9 a_27_368.t0 a_27_368.n11 219.476
R10 a_27_368.n1 a_27_368.t8 188.565
R11 a_27_368.n8 a_27_368.t9 186.374
R12 a_27_368.n5 a_27_368.t7 186.374
R13 a_27_368.n2 a_27_368.t6 186.374
R14 a_27_368.n4 a_27_368.n0 165.189
R15 a_27_368.n10 a_27_368.n9 152
R16 a_27_368.n7 a_27_368.n0 152
R17 a_27_368.n2 a_27_368.n1 63.5369
R18 a_27_368.n9 a_27_368.n7 49.6611
R19 a_27_368.n5 a_27_368.n4 39.4369
R20 a_27_368.n4 a_27_368.n3 21.1793
R21 a_27_368.n10 a_27_368.n0 13.1884
R22 a_27_368.n6 a_27_368.n5 5.11262
R23 a_27_368.n7 a_27_368.n6 5.11262
R24 a_27_368.n9 a_27_368.n8 2.92171
R25 a_27_368.n3 a_27_368.n2 2.19141
R26 VPWR.n4 VPWR.n3 604.588
R27 VPWR.n11 VPWR.n1 603.569
R28 VPWR.n6 VPWR.n5 329.755
R29 VPWR.n9 VPWR.n2 36.1417
R30 VPWR.n10 VPWR.n9 36.1417
R31 VPWR.n1 VPWR.t0 29.0228
R32 VPWR.n1 VPWR.t2 28.1434
R33 VPWR.n3 VPWR.t1 26.3844
R34 VPWR.n3 VPWR.t4 26.3844
R35 VPWR.n5 VPWR.t3 26.3844
R36 VPWR.n5 VPWR.t5 26.3844
R37 VPWR.n11 VPWR.n10 21.0829
R38 VPWR.n6 VPWR.n4 16.708
R39 VPWR.n7 VPWR.n2 9.3005
R40 VPWR.n9 VPWR.n8 9.3005
R41 VPWR.n10 VPWR.n0 9.3005
R42 VPWR.n12 VPWR.n11 7.27223
R43 VPWR.n7 VPWR.n6 1.48647
R44 VPWR.n4 VPWR.n2 0.753441
R45 VPWR VPWR.n12 0.157962
R46 VPWR.n12 VPWR.n0 0.149814
R47 VPWR.n8 VPWR.n7 0.122949
R48 VPWR.n8 VPWR.n0 0.122949
R49 VPB.t0 VPB.t8 577.152
R50 VPB VPB.t6 257.93
R51 VPB.t6 VPB.t0 242.608
R52 VPB.t5 VPB.t3 229.839
R53 VPB.t4 VPB.t5 229.839
R54 VPB.t2 VPB.t4 229.839
R55 VPB.t7 VPB.t2 229.839
R56 VPB.t9 VPB.t7 229.839
R57 VPB.t1 VPB.t9 229.839
R58 VPB.t8 VPB.t1 229.839
R59 a_208_74.t0 a_208_74.n3 893.708
R60 a_208_74.n0 a_208_74.t3 281.168
R61 a_208_74.n3 a_208_74.n2 235.763
R62 a_208_74.n2 a_208_74.t2 142.994
R63 a_208_74.n1 a_208_74.t4 142.994
R64 a_208_74.n0 a_208_74.t5 142.994
R65 a_208_74.n1 a_208_74.n0 138.173
R66 a_208_74.n2 a_208_74.n1 138.173
R67 a_208_74.n3 a_208_74.t1 119.811
R68 a_378_74.n2 a_378_74.t7 232.281
R69 a_378_74.t0 a_378_74.n5 215.946
R70 a_378_74.n5 a_378_74.n0 196.672
R71 a_378_74.n2 a_378_74.n1 107.79
R72 a_378_74.n4 a_378_74.n3 87.0786
R73 a_378_74.n5 a_378_74.n4 78.1586
R74 a_378_74.n4 a_378_74.n2 61.8951
R75 a_378_74.n3 a_378_74.t3 22.7032
R76 a_378_74.n3 a_378_74.t6 22.7032
R77 a_378_74.n1 a_378_74.t4 22.7032
R78 a_378_74.n1 a_378_74.t5 22.7032
R79 a_378_74.n0 a_378_74.t1 22.7032
R80 a_378_74.n0 a_378_74.t2 22.7032
R81 VGND.n5 VGND.n4 224.109
R82 VGND.n3 VGND.n2 115.659
R83 VGND.n11 VGND.n10 115.424
R84 VGND.n8 VGND.n1 36.1417
R85 VGND.n9 VGND.n8 36.1417
R86 VGND.n4 VGND.t3 22.7032
R87 VGND.n4 VGND.t1 22.7032
R88 VGND.n2 VGND.t2 22.7032
R89 VGND.n2 VGND.t4 22.7032
R90 VGND.n10 VGND.t5 22.7032
R91 VGND.n10 VGND.t0 22.7032
R92 VGND.n11 VGND.n9 21.4593
R93 VGND.n3 VGND.n1 10.1652
R94 VGND.n6 VGND.n1 9.3005
R95 VGND.n8 VGND.n7 9.3005
R96 VGND.n9 VGND.n0 9.3005
R97 VGND.n5 VGND.n3 7.67732
R98 VGND.n12 VGND.n11 7.34058
R99 VGND.n6 VGND.n5 1.22444
R100 VGND VGND.n12 0.158861
R101 VGND.n12 VGND.n0 0.148926
R102 VGND.n7 VGND.n6 0.122949
R103 VGND.n7 VGND.n0 0.122949
R104 VNB.t9 VNB.t8 2956.43
R105 VNB VNB.t4 1235.7
R106 VNB.t3 VNB.t1 1039.37
R107 VNB.t2 VNB.t3 993.177
R108 VNB.t0 VNB.t2 993.177
R109 VNB.t7 VNB.t0 993.177
R110 VNB.t5 VNB.t7 993.177
R111 VNB.t6 VNB.t5 993.177
R112 VNB.t8 VNB.t6 993.177
R113 VNB.t4 VNB.t9 993.177
R114 a_348_368.n4 a_348_368.t6 772.996
R115 a_348_368.n2 a_348_368.n1 308.902
R116 a_348_368.n2 a_348_368.t4 294.469
R117 a_348_368.n5 a_348_368.n4 190.346
R118 a_348_368.n3 a_348_368.n0 185.916
R119 a_348_368.n4 a_348_368.n3 99.7247
R120 a_348_368.n3 a_348_368.n2 82.1705
R121 a_348_368.n0 a_348_368.t1 26.3844
R122 a_348_368.n0 a_348_368.t5 26.3844
R123 a_348_368.n1 a_348_368.t2 26.3844
R124 a_348_368.n1 a_348_368.t3 26.3844
R125 a_348_368.n5 a_348_368.t7 26.3844
R126 a_348_368.t0 a_348_368.n5 26.3844
R127 Z.n5 Z.n1 247.617
R128 Z.n4 Z.n2 234.41
R129 Z.n6 Z.n0 193.445
R130 Z.n4 Z.n3 192.952
R131 Z.n5 Z.n4 56.9923
R132 Z.n0 Z.t1 26.3844
R133 Z.n0 Z.t3 26.3844
R134 Z.n1 Z.t2 26.3844
R135 Z.n1 Z.t0 26.3844
R136 Z.n3 Z.t5 25.9464
R137 Z.n3 Z.t7 22.7032
R138 Z.n2 Z.t6 22.7032
R139 Z.n2 Z.t4 22.7032
R140 Z.n6 Z 9.3932
R141 Z Z.n6 4.55261
R142 Z Z.n5 1.7199
R143 TE_B.n0 TE_B.t0 344.433
R144 TE_B.n3 TE_B.n2 273.473
R145 TE_B.n3 TE_B.t4 225.087
R146 TE_B.n0 TE_B.t1 204.048
R147 TE_B.n1 TE_B.t2 204.048
R148 TE_B.n2 TE_B.t5 204.048
R149 TE_B.n4 TE_B.t3 176.964
R150 TE_B TE_B.n4 159.226
R151 TE_B.n1 TE_B.n0 132.423
R152 TE_B.n2 TE_B.n1 132.423
R153 TE_B.n4 TE_B.n3 36.4948
C0 VPB A 0.035421f
C1 VPB TE_B 0.206984f
C2 VPB VPWR 0.147232f
C3 A TE_B 0.089722f
C4 A VPWR 0.017824f
C5 VPB Z 0.008261f
C6 TE_B VPWR 0.073494f
C7 VPB VGND 0.009385f
C8 TE_B Z 5.23e-19
C9 A VGND 0.037699f
C10 TE_B VGND 0.02999f
C11 VPWR Z 0.019756f
C12 VPWR VGND 0.091096f
C13 Z VGND 0.019264f
C14 VGND VNB 0.679955f
C15 Z VNB 0.033442f
C16 VPWR VNB 0.544786f
C17 TE_B VNB 0.283162f
C18 A VNB 0.135414f
C19 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ebufn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ebufn_2 VNB VPB VPWR VGND Z TE_B A
X0 VPWR.t0 TE_B.t0 a_283_48.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.295 ps=2.59 w=1 l=0.15
X1 Z.t2 a_84_48.t2 a_33_368.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t2 TE_B.t1 a_33_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.29075 pd=1.78 as=0.196 ps=1.47 w=1.12 l=0.15
X3 a_27_74.t1 a_283_48.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10545 ps=1.025 w=0.74 l=0.15
X4 VGND.t1 TE_B.t2 a_283_48.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.1824 ps=1.85 w=0.64 l=0.15
X5 a_33_368.t0 TE_B.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.29075 ps=1.78 w=1.12 l=0.15
X6 Z.t0 a_84_48.t3 a_27_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 a_33_368.t2 a_84_48.t4 Z.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X8 VGND.t2 a_283_48.t3 a_27_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.15355 ps=1.155 w=0.74 l=0.15
X9 a_84_48.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1344 ps=1.06 w=0.64 l=0.15
X10 a_27_74.t2 a_84_48.t5 Z.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.15355 pd=1.155 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_84_48.t1 A.t1 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.25 ps=1.5 w=1 l=0.15
R0 TE_B.n0 TE_B.t1 399.06
R1 TE_B.n1 TE_B.n0 254.192
R2 TE_B.n2 TE_B.t2 226.541
R3 TE_B.n1 TE_B.t0 206.433
R4 TE_B.n0 TE_B.t3 204.048
R5 TE_B TE_B.n2 162.667
R6 TE_B.n2 TE_B.n1 24.1005
R7 a_283_48.t1 a_283_48.n1 868.217
R8 a_283_48.n0 a_283_48.t3 282.774
R9 a_283_48.n1 a_283_48.n0 233.698
R10 a_283_48.n0 a_283_48.t2 142.994
R11 a_283_48.n1 a_283_48.t0 133.944
R12 VPWR.n2 VPWR.n0 623.375
R13 VPWR.n2 VPWR.n1 607.322
R14 VPWR.n1 VPWR.t3 54.1755
R15 VPWR.n1 VPWR.t0 44.3255
R16 VPWR.n0 VPWR.t1 41.3353
R17 VPWR.n0 VPWR.t2 41.3353
R18 VPWR VPWR.n2 0.494511
R19 VPB.t2 VPB.t4 515.861
R20 VPB.t4 VPB.t5 331.99
R21 VPB.t3 VPB.t2 316.668
R22 VPB VPB.t0 273.253
R23 VPB.t1 VPB.t3 255.376
R24 VPB.t0 VPB.t1 255.376
R25 a_84_48.n3 a_84_48.n2 378.995
R26 a_84_48.n2 a_84_48.t4 240.197
R27 a_84_48.n0 a_84_48.t2 240.197
R28 a_84_48.t1 a_84_48.n3 224.367
R29 a_84_48.n3 a_84_48.t0 218.056
R30 a_84_48.n0 a_84_48.t3 186.839
R31 a_84_48.n1 a_84_48.t5 179.947
R32 a_84_48.n1 a_84_48.n0 56.9641
R33 a_84_48.n2 a_84_48.n1 16.0672
R34 a_33_368.n0 a_33_368.t0 903.064
R35 a_33_368.n0 a_33_368.t3 390.717
R36 a_33_368.n1 a_33_368.n0 293.027
R37 a_33_368.n1 a_33_368.t2 35.1791
R38 a_33_368.t1 a_33_368.n1 26.3844
R39 Z Z.n2 285.894
R40 Z Z.n0 220.852
R41 Z.n0 Z.t2 35.1791
R42 Z.n1 Z 28.2358
R43 Z.n1 Z 26.6672
R44 Z.n0 Z.t1 26.3844
R45 Z.n2 Z.t3 22.7032
R46 Z.n2 Z.t0 22.7032
R47 Z Z.n1 7.90638
R48 Z.n1 Z 7.46717
R49 VGND.n2 VGND.n1 222.982
R50 VGND.n2 VGND.n0 121.928
R51 VGND.n0 VGND.t0 39.3755
R52 VGND.n0 VGND.t1 39.3755
R53 VGND.n1 VGND.t2 23.514
R54 VGND.n1 VGND.t3 22.7032
R55 VGND VGND.n2 0.441051
R56 a_27_74.n1 a_27_74.t3 220.685
R57 a_27_74.t1 a_27_74.n1 206.113
R58 a_27_74.n1 a_27_74.n0 88.3339
R59 a_27_74.n0 a_27_74.t2 34.0546
R60 a_27_74.n0 a_27_74.t0 33.2437
R61 VNB.t3 VNB.t1 2991.08
R62 VNB.t1 VNB.t0 1316.54
R63 VNB.t4 VNB.t2 1304.99
R64 VNB VNB.t5 1143.31
R65 VNB.t2 VNB.t3 1004.72
R66 VNB.t5 VNB.t4 993.177
R67 A.n0 A.t0 233.576
R68 A.n0 A.t1 229.023
R69 A A.n0 157.507
C0 VPB VPWR 0.120733f
C1 VPB TE_B 0.152138f
C2 A VPB 0.04124f
C3 VPWR TE_B 0.029904f
C4 VPB Z 0.009428f
C5 VGND VPB 0.00948f
C6 A VPWR 0.016207f
C7 VPWR Z 0.021829f
C8 VGND VPWR 0.070578f
C9 A TE_B 0.076442f
C10 TE_B Z 0.014997f
C11 VGND TE_B 0.022531f
C12 A VGND 0.032793f
C13 VGND Z 0.010727f
C14 VGND VNB 0.534103f
C15 A VNB 0.150666f
C16 Z VNB 0.038984f
C17 TE_B VNB 0.227371f
C18 VPWR VNB 0.429305f
C19 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__ebufn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__ebufn_1 VNB VPB VPWR VGND A Z TE_B
X0 Z.t0 a_229_74.t2 a_569_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 VGND.t2 TE_B.t0 a_27_404.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0825 pd=0.85 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 VPWR.t1 TE_B.t1 a_27_404.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.22785 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X3 Z.t1 a_229_74.t3 a_566_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X4 a_566_368.t0 TE_B.t2 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 a_569_74.t0 a_27_404.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_229_74.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.0825 ps=0.85 w=0.55 l=0.15
X7 a_229_74.t1 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2562 pd=2.29 as=0.22785 ps=1.52 w=0.84 l=0.15
R0 a_229_74.t1 a_229_74.n1 848.952
R1 a_229_74.n1 a_229_74.t0 329.64
R2 a_229_74.n0 a_229_74.t3 258.942
R3 a_229_74.n0 a_229_74.t2 210.474
R4 a_229_74.n1 a_229_74.n0 170.72
R5 a_569_74.t0 a_569_74.t1 38.9194
R6 Z.n0 Z.t1 286.86
R7 Z.t0 Z.n0 279.738
R8 Z.n1 Z.t0 279.738
R9 Z.n1 Z 7.63353
R10 Z.n0 Z 2.93628
R11 Z Z.n1 1.05738
R12 VNB.t0 VNB.t1 3926.51
R13 VNB VNB.t3 1432.02
R14 VNB.t3 VNB.t0 1039.37
R15 VNB.t1 VNB.t2 900.788
R16 TE_B.n1 TE_B.t2 839.509
R17 TE_B.n0 TE_B.t0 298.132
R18 TE_B.n0 TE_B.t1 213.246
R19 TE_B.n1 TE_B.n0 152
R20 TE_B TE_B.n1 2.65416
R21 a_27_404.n0 a_27_404.t2 555.986
R22 a_27_404.t1 a_27_404.n0 448.663
R23 a_27_404.n0 a_27_404.t0 232.517
R24 VGND.n1 VGND.t1 298.214
R25 VGND.n1 VGND.n0 219.719
R26 VGND.n0 VGND.t0 32.7278
R27 VGND.n0 VGND.t2 32.7278
R28 VGND VGND.n1 0.220189
R29 VPWR.n1 VPWR.n0 650.564
R30 VPWR.n1 VPWR.t2 254.614
R31 VPWR.n0 VPWR.t0 55.1136
R32 VPWR.n0 VPWR.t1 55.1136
R33 VPWR VPWR.n1 0.218411
R34 VPB.t0 VPB.t1 832.528
R35 VPB.t2 VPB.t0 316.668
R36 VPB VPB.t2 257.93
R37 VPB.t1 VPB.t3 214.517
R38 a_566_368.t0 a_566_368.t1 47.4916
R39 A.n0 A.t0 282.774
R40 A.n0 A.t1 189.855
R41 A.n1 A.n0 90.1298
R42 A.n1 A 10.5475
R43 A A.n1 7.5986
C0 A VGND 0.018531f
C1 Z VGND 0.072515f
C2 VPB VPWR 0.122732f
C3 VPB TE_B 0.293059f
C4 VPB A 0.077243f
C5 VPWR TE_B 0.234879f
C6 VPWR A 0.012191f
C7 VPB Z 0.022895f
C8 VPB VGND 0.009751f
C9 TE_B A 0.140622f
C10 VPWR Z 0.09388f
C11 TE_B Z 0.007947f
C12 VPWR VGND 0.060357f
C13 TE_B VGND 0.019427f
C14 A Z 1.26e-19
C15 VGND VNB 0.513428f
C16 Z VNB 0.122275f
C17 A VNB 0.160851f
C18 TE_B VNB 0.223592f
C19 VPWR VNB 0.39415f
C20 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvp_1 VNB VPB VPWR VGND TE Z A
X0 a_310_392.t0 a_44_549.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.1664 ps=1.385 w=1 l=0.15
X1 VGND.t1 TE.t0 a_44_549.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1138 pd=1.08 as=0.2604 ps=2.08 w=0.42 l=0.15
X2 VPWR.t1 TE.t1 a_44_549.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.2646 ps=2.1 w=0.42 l=0.15
X3 a_318_74.t0 TE.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1138 ps=1.08 w=0.74 l=0.15
X4 Z.t1 A.t0 a_318_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5 Z.t0 A.t1 a_310_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
R0 a_44_549.n0 a_44_549.t2 487.257
R1 a_44_549.n0 a_44_549.t1 397.945
R2 a_44_549.t0 a_44_549.n0 233.912
R3 VPWR VPWR.n0 228.542
R4 VPWR.n0 VPWR.t1 110.227
R5 VPWR.n0 VPWR.t0 29.5505
R6 a_310_392.t0 a_310_392.t1 53.1905
R7 VPB VPB.t2 480.108
R8 VPB.t2 VPB.t0 273.253
R9 VPB.t0 VPB.t1 214.517
R10 TE.n0 TE.t2 366.613
R11 TE.n0 TE.t0 276.348
R12 TE.n1 TE 201.142
R13 TE.n3 TE.n2 152
R14 TE.n1 TE.t1 122.374
R15 TE.n3 TE 11.8593
R16 TE.n2 TE.n0 10.955
R17 TE TE.n3 6.21226
R18 TE.n2 TE.n1 1.46111
R19 VGND VGND.n0 126.648
R20 VGND.n0 VGND.t1 57.8155
R21 VGND.n0 VGND.t0 22.6447
R22 VNB VNB.t1 2367.45
R23 VNB.t1 VNB.t0 1131.76
R24 VNB.t0 VNB.t2 900.788
R25 a_318_74.t0 a_318_74.t1 38.9194
R26 A.n0 A.t1 281.373
R27 A.n0 A.t0 197.82
R28 A A.n0 156.462
R29 Z Z.n0 589.85
R30 Z.n2 Z.n0 585
R31 Z.n1 Z.n0 585
R32 Z.n1 Z.t1 239.53
R33 Z.n0 Z.t0 29.5505
R34 Z Z.n2 8.72777
R35 Z Z.n1 7.95202
R36 Z.n2 Z 5.62474
C0 VGND TE 0.062021f
C1 VPB A 0.052271f
C2 VGND Z 0.084389f
C3 VPB VPWR 0.063567f
C4 VPB TE 0.090212f
C5 A VPWR 0.014046f
C6 A TE 0.046395f
C7 VPB Z 0.018794f
C8 VPWR TE 0.035922f
C9 A Z 0.148412f
C10 VPWR Z 0.094094f
C11 TE Z 0.036956f
C12 VGND VPB 0.007804f
C13 VGND A 0.013556f
C14 VGND VPWR 0.042441f
C15 VGND VNB 0.335537f
C16 Z VNB 0.093702f
C17 TE VNB 0.280054f
C18 VPWR VNB 0.265132f
C19 A VNB 0.16757f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvp_2 VNB VPB VPWR VGND Z A TE
X0 Z.t1 A.t0 a_27_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VGND.t1 TE.t0 a_36_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t0 TE.t1 a_263_323.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1888 pd=1.87 as=0.1856 ps=1.86 w=0.64 l=0.15
X3 VGND.t2 TE.t2 a_263_323.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.1197 ps=1.41 w=0.42 l=0.15
X4 a_36_74.t1 A.t1 Z.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 Z.t2 A.t2 a_36_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_27_368.t2 a_263_323.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VPWR.t1 a_263_323.t3 a_27_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_27_368.t0 A.t3 Z.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_36_74.t2 TE.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t3 261.62
R1 A.n2 A.t0 261.62
R2 A A.n2 193.113
R3 A.n0 A.t1 156.431
R4 A.n1 A.t2 154.24
R5 A.n1 A.n0 60.6157
R6 A.n2 A.n1 5.11262
R7 a_27_368.n0 a_27_368.t2 364.536
R8 a_27_368.n0 a_27_368.t1 339.568
R9 a_27_368.n1 a_27_368.n0 181.875
R10 a_27_368.n1 a_27_368.t3 26.3844
R11 a_27_368.t0 a_27_368.n1 26.3844
R12 Z.n0 Z 595.159
R13 Z.n1 Z.n0 585
R14 Z Z.n2 204.651
R15 Z.n0 Z.t0 26.3844
R16 Z.n0 Z.t1 26.3844
R17 Z.n2 Z.t3 22.7032
R18 Z.n2 Z.t2 22.7032
R19 Z.n1 Z 13.6132
R20 Z Z.n1 1.42272
R21 VPB.t3 VPB.t0 510.753
R22 VPB VPB.t2 257.93
R23 VPB.t4 VPB.t3 229.839
R24 VPB.t1 VPB.t4 229.839
R25 VPB.t2 VPB.t1 229.839
R26 TE.t2 TE.t1 592.861
R27 TE.n1 TE.n0 424.161
R28 TE.n0 TE.t0 281.168
R29 TE TE.n1 154.81
R30 TE.n0 TE.t3 142.994
R31 TE.n1 TE.t2 132.769
R32 a_36_74.n0 a_36_74.t2 244.294
R33 a_36_74.n0 a_36_74.t0 221.048
R34 a_36_74.n1 a_36_74.n0 84.741
R35 a_36_74.n1 a_36_74.t3 22.7032
R36 a_36_74.t1 a_36_74.n1 22.7032
R37 VGND.n1 VGND.t2 274.776
R38 VGND.n1 VGND.n0 121.347
R39 VGND.n0 VGND.t0 22.7032
R40 VGND.n0 VGND.t1 22.7032
R41 VGND VGND.n1 0.476529
R42 VNB.t2 VNB.t3 2355.91
R43 VNB VNB.t0 1247.24
R44 VNB.t4 VNB.t2 993.177
R45 VNB.t1 VNB.t4 993.177
R46 VNB.t0 VNB.t1 993.177
R47 a_263_323.t0 a_263_323.n1 384.2
R48 a_263_323.n1 a_263_323.n0 356.048
R49 a_263_323.n0 a_263_323.t3 348.647
R50 a_263_323.n1 a_263_323.t1 254.868
R51 a_263_323.n0 a_263_323.t2 204.048
R52 VPWR.n1 VPWR.t0 381.534
R53 VPWR.n1 VPWR.n0 238.639
R54 VPWR.n0 VPWR.t2 26.3844
R55 VPWR.n0 VPWR.t1 26.3844
R56 VPWR VPWR.n1 0.476004
C0 TE VPWR 0.033173f
C1 A VGND 0.014918f
C2 Z VPWR 0.010116f
C3 TE VGND 0.149925f
C4 Z VGND 0.008902f
C5 VPWR VGND 0.062087f
C6 VPB A 0.072886f
C7 VPB TE 0.090364f
C8 VPB Z 0.003686f
C9 A TE 0.02211f
C10 A Z 0.094364f
C11 VPB VPWR 0.102762f
C12 VPB VGND 0.010757f
C13 A VPWR 0.012545f
C14 TE Z 0.00115f
C15 VGND VNB 0.46294f
C16 VPWR VNB 0.372671f
C17 Z VNB 0.020262f
C18 TE VNB 0.480836f
C19 A VNB 0.277685f
C20 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvp_4 VNB VPB VPWR VGND TE Z A
X0 VGND.t4 TE.t0 a_27_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 a_27_368.t6 A.t0 Z.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t0 TE.t1 a_473_323.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 Z.t2 A.t1 a_27_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 Z.t1 A.t2 a_27_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.336 ps=2.84 w=1.12 l=0.15
X5 a_27_74.t4 A.t3 Z.t7 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.12025 ps=1.065 w=0.74 l=0.15
X6 a_27_74.t2 TE.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X7 Z.t6 A.t4 a_27_74.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 Z.t5 A.t5 a_27_74.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.13875 ps=1.115 w=0.74 l=0.15
X9 a_27_368.t3 A.t6 Z.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1932 ps=1.465 w=1.12 l=0.15
X10 VPWR.t4 a_473_323.t2 a_27_368.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_27_368.t0 a_473_323.t3 VPWR.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X12 VGND.t2 TE.t3 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_27_368.t1 a_473_323.t4 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1736 ps=1.43 w=1.12 l=0.15
X14 VPWR.t1 a_473_323.t5 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X15 a_27_74.t7 A.t7 Z.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.13875 pd=1.115 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 a_27_74.t0 TE.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X17 VGND.t0 TE.t5 a_473_323.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
R0 TE.n2 TE.t0 339.007
R1 TE.n5 TE.n4 302.947
R2 TE.n1 TE.t1 240.197
R3 TE.n4 TE.n3 183.161
R4 TE.n1 TE.n0 179.374
R5 TE TE.n6 163.249
R6 TE.n2 TE.t4 155.847
R7 TE.n3 TE.t3 155.847
R8 TE.n4 TE.t2 155.847
R9 TE.n5 TE.t5 155.847
R10 TE.n3 TE.n2 138.173
R11 TE.n6 TE.n1 13.0919
R12 TE.n0 TE 11.152
R13 TE.n6 TE.n5 10.7116
R14 TE TE.n0 1.93989
R15 a_27_74.n4 a_27_74.t2 210.839
R16 a_27_74.n1 a_27_74.t5 205.212
R17 a_27_74.n1 a_27_74.n0 185
R18 a_27_74.n5 a_27_74.n4 112.96
R19 a_27_74.n3 a_27_74.n2 88.3339
R20 a_27_74.n4 a_27_74.n3 75.0731
R21 a_27_74.n3 a_27_74.n1 69.4453
R22 a_27_74.n2 a_27_74.t4 34.0546
R23 a_27_74.n0 a_27_74.t7 34.0546
R24 a_27_74.n0 a_27_74.t6 26.7573
R25 a_27_74.n2 a_27_74.t3 22.7032
R26 a_27_74.n5 a_27_74.t1 22.7032
R27 a_27_74.t0 a_27_74.n5 22.7032
R28 VGND.n3 VGND.t0 156.894
R29 VGND.n8 VGND.n7 116.644
R30 VGND.n2 VGND.n1 116.644
R31 VGND.n6 VGND.n5 36.1417
R32 VGND.n1 VGND.t3 34.0546
R33 VGND.n1 VGND.t2 34.0546
R34 VGND.n7 VGND.t1 34.0546
R35 VGND.n7 VGND.t4 34.0546
R36 VGND.n3 VGND.n2 17.7124
R37 VGND.n8 VGND.n6 13.177
R38 VGND.n5 VGND.n4 9.3005
R39 VGND.n6 VGND.n0 9.3005
R40 VGND.n9 VGND.n8 7.58996
R41 VGND.n5 VGND.n2 1.12991
R42 VGND VGND.n9 0.649578
R43 VGND.n4 VGND.n3 0.25103
R44 VGND.n9 VGND.n0 0.15042
R45 VGND.n4 VGND.n0 0.122949
R46 VNB.t3 VNB.t0 2286.61
R47 VNB.t2 VNB.t3 1316.54
R48 VNB.t4 VNB.t1 1316.54
R49 VNB.t8 VNB.t7 1212.6
R50 VNB.t5 VNB.t4 1154.86
R51 VNB.t6 VNB.t8 1154.86
R52 VNB VNB.t6 1143.31
R53 VNB.t7 VNB.t5 1097.11
R54 VNB.t1 VNB.t2 993.177
R55 A.n0 A.t0 292.642
R56 A.n2 A.t1 226.809
R57 A.n4 A.t6 226.809
R58 A.n6 A.t2 226.809
R59 A.n0 A.t3 213.648
R60 A.n6 A.t4 198.204
R61 A.n5 A.t7 196.013
R62 A.n1 A.t5 196.013
R63 A A.n3 156.465
R64 A.n10 A.n9 152
R65 A.n8 A.n7 152
R66 A.n1 A.n0 97.715
R67 A.n9 A.n8 49.6611
R68 A.n4 A.n3 37.9763
R69 A.n3 A.n2 35.055
R70 A.n7 A 12.8005
R71 A.n8 A.n6 10.955
R72 A.n9 A.n5 10.2247
R73 A.n10 A 8.63306
R74 A A.n10 5.65631
R75 A.n2 A.n1 2.19141
R76 A.n7 A 1.48887
R77 A.n5 A.n4 1.46111
R78 Z.n4 Z.n0 344.702
R79 Z.n6 Z.n5 292.596
R80 Z.n3 Z.n1 245.921
R81 Z.n3 Z.n2 195.474
R82 Z.n4 Z.n3 41.7944
R83 Z.n0 Z.t1 34.2996
R84 Z.n1 Z.t6 34.0546
R85 Z.n2 Z.t5 30.0005
R86 Z.n0 Z.t0 26.3844
R87 Z.n5 Z.t3 26.3844
R88 Z.n5 Z.t2 26.3844
R89 Z.n2 Z.t7 22.7032
R90 Z.n1 Z.t4 22.7032
R91 Z Z.n6 5.53007
R92 Z.n6 Z.n4 5.424
R93 a_27_368.n1 a_27_368.n0 305.998
R94 a_27_368.n3 a_27_368.t1 295.81
R95 a_27_368.n1 a_27_368.t4 287.644
R96 a_27_368.n3 a_27_368.n2 219.732
R97 a_27_368.n5 a_27_368.n4 188.054
R98 a_27_368.n4 a_27_368.n1 75.1613
R99 a_27_368.n4 a_27_368.n3 72.4344
R100 a_27_368.n0 a_27_368.t3 35.1791
R101 a_27_368.t6 a_27_368.n5 35.1791
R102 a_27_368.n0 a_27_368.t5 26.3844
R103 a_27_368.n2 a_27_368.t7 26.3844
R104 a_27_368.n2 a_27_368.t0 26.3844
R105 a_27_368.n5 a_27_368.t2 26.3844
R106 VPB.t1 VPB.t8 709.947
R107 VPB VPB.t4 260.485
R108 VPB.t2 VPB.t0 255.376
R109 VPB.t6 VPB.t2 255.376
R110 VPB.t3 VPB.t5 255.376
R111 VPB.t4 VPB.t3 252.823
R112 VPB.t7 VPB.t1 234.946
R113 VPB.t0 VPB.t7 229.839
R114 VPB.t5 VPB.t6 229.839
R115 a_473_323.n0 a_473_323.t5 364.714
R116 a_473_323.n3 a_473_323.n2 253.173
R117 a_473_323.t0 a_473_323.n3 224.252
R118 a_473_323.n2 a_473_323.t4 204.048
R119 a_473_323.n1 a_473_323.t2 204.048
R120 a_473_323.n0 a_473_323.t3 204.048
R121 a_473_323.n3 a_473_323.t1 196.391
R122 a_473_323.n2 a_473_323.n1 147.814
R123 a_473_323.n1 a_473_323.n0 144.601
R124 VPWR.n2 VPWR.t0 266.884
R125 VPWR.n6 VPWR.n1 230.268
R126 VPWR.n4 VPWR.n3 228.922
R127 VPWR.n1 VPWR.t1 35.1791
R128 VPWR.n3 VPWR.t2 27.2639
R129 VPWR.n3 VPWR.t4 27.2639
R130 VPWR.n1 VPWR.t3 26.3844
R131 VPWR.n5 VPWR.n4 25.977
R132 VPWR.n6 VPWR.n5 22.9652
R133 VPWR.n5 VPWR.n0 9.3005
R134 VPWR.n7 VPWR.n6 7.45461
R135 VPWR.n4 VPWR.n2 7.28361
R136 VPWR VPWR.n7 0.647411
R137 VPWR.n2 VPWR.n0 0.167447
R138 VPWR.n7 VPWR.n0 0.152553
C0 VPWR TE 0.05079f
C1 Z VGND 0.020093f
C2 VPWR VGND 0.092373f
C3 TE VGND 0.126072f
C4 VPB A 0.14354f
C5 VPB Z 0.003876f
C6 VPB VPWR 0.153243f
C7 A Z 0.308418f
C8 VPB TE 0.061444f
C9 A VPWR 0.025485f
C10 VPB VGND 0.007633f
C11 A TE 0.019371f
C12 Z VPWR 0.021388f
C13 A VGND 0.026745f
C14 VGND VNB 0.712766f
C15 TE VNB 0.565854f
C16 VPWR VNB 0.583254f
C17 Z VNB 0.023768f
C18 A VNB 0.472671f
C19 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fa_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fa_1 VNB VPB VPWR CIN VGND A B COUT SUM
X0 a_465_249.t2 B.t0 a_936_75.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0768 ps=0.88 w=0.64 l=0.15
X1 a_501_75.t1 A.t0 VGND.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.169075 ps=1.275 w=0.64 l=0.15
X2 a_318_389.t1 B.t1 a_217_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.195875 pd=1.565 as=0.186675 ps=1.46 w=1 l=0.15
X3 VPWR.t6 CIN.t0 a_509_347.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.31 as=0.1775 ps=1.355 w=1 l=0.15
X4 a_69_260.t0 CIN.t1 a_315_75.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
X5 a_501_75.t3 a_465_249.t3 a_69_260.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1152 pd=1 as=0.1248 ps=1.03 w=0.64 l=0.15
X6 VGND.t4 A.t1 a_1100_75.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.212275 pd=1.41 as=0.3596 ps=1.73 w=0.64 l=0.15
X7 VGND.t7 a_69_260.t4 SUM.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.191575 pd=1.395 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VGND.t6 CIN.t2 a_501_75.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1584 pd=1.135 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 a_237_75.t1 A.t2 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.191575 ps=1.395 w=0.64 l=0.15
X10 a_509_347.t1 A.t3 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1775 pd=1.355 as=0.243625 ps=1.64 w=1 l=0.15
X11 COUT.t0 a_465_249.t4 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.3304 ps=2.83 w=1.12 l=0.15
X12 a_465_249.t1 B.t2 a_916_347.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1775 ps=1.355 w=1 l=0.15
X13 VPWR.t5 A.t4 a_1107_347.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.34905 pd=1.76 as=0.2225 ps=1.445 w=1 l=0.15
X14 a_1100_75.t0 B.t3 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.212275 ps=1.41 w=0.64 l=0.15
X15 a_509_347.t3 a_465_249.t5 a_69_260.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1675 pd=1.335 as=0.15 ps=1.3 w=1 l=0.15
X16 a_217_368.t1 A.t5 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.186675 pd=1.46 as=0.199 ps=1.485 w=1 l=0.15
X17 a_916_347.t1 A.t6 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1775 pd=1.355 as=0.155 ps=1.31 w=1 l=0.15
X18 a_936_75.t0 A.t7 VGND.t5 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1584 ps=1.135 w=0.64 l=0.15
X19 a_69_260.t1 CIN.t3 a_318_389.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.195875 ps=1.565 w=1 l=0.15
X20 a_1100_75.t2 CIN.t4 a_465_249.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3596 pd=1.73 as=0.0896 ps=0.92 w=0.64 l=0.15
X21 VPWR.t7 a_69_260.t5 SUM.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.199 pd=1.485 as=0.3192 ps=2.81 w=1.12 l=0.15
X22 VPWR.t0 B.t4 a_509_347.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.243625 pd=1.64 as=0.1675 ps=1.335 w=1 l=0.15
X23 a_1107_347.t0 B.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.335 pd=2.67 as=0.34905 ps=1.76 w=1 l=0.15
X24 a_315_75.t0 B.t6 a_237_75.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.0768 ps=0.88 w=0.64 l=0.15
X25 VGND.t0 B.t7 a_501_75.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.169075 pd=1.275 as=0.1152 ps=1 w=0.64 l=0.15
R0 B.t5 B.n1 801.995
R1 B.n0 B.t1 624.458
R2 B.n1 B.n0 602.5
R3 B.t1 B.t6 554.033
R4 B.t4 B.t7 464.327
R5 B.t2 B.t0 464.327
R6 B.n0 B.t4 275.812
R7 B.n1 B.t2 275.812
R8 B.n2 B.t5 233.463
R9 B.n2 B.t3 218.113
R10 B B.n2 75.9
R11 a_936_75.t0 a_936_75.t1 45.0005
R12 a_465_249.t1 a_465_249.n5 385.529
R13 a_465_249.n5 a_465_249.n0 355.63
R14 a_465_249.n4 a_465_249.n3 289.659
R15 a_465_249.n2 a_465_249.t4 276.767
R16 a_465_249.n4 a_465_249.n2 258.154
R17 a_465_249.n0 a_465_249.t5 231.629
R18 a_465_249.n0 a_465_249.t3 200.833
R19 a_465_249.n2 a_465_249.n1 169.389
R20 a_465_249.n5 a_465_249.n4 129.431
R21 a_465_249.n3 a_465_249.t0 26.2505
R22 a_465_249.n3 a_465_249.t2 26.2505
R23 VNB.t2 VNB.t11 2591.11
R24 VNB.t11 VNB.t5 1772.22
R25 VNB.t8 VNB.t0 1576.67
R26 VNB.t9 VNB.t1 1503.33
R27 VNB.t3 VNB.t10 1442.22
R28 VNB.t7 VNB.t12 1320
R29 VNB.t12 VNB.t3 1246.67
R30 VNB VNB.t9 1210
R31 VNB.t6 VNB.t2 1051.11
R32 VNB.t10 VNB.t8 1051.11
R33 VNB.t0 VNB.t6 953.333
R34 VNB.t4 VNB.t7 953.333
R35 VNB.t1 VNB.t4 953.333
R36 A.n5 A.n3 335.524
R37 A.n2 A.n0 268.889
R38 A.n3 A.t5 266.44
R39 A.n1 A.t6 263.762
R40 A.n4 A.t3 263.762
R41 A.n0 A.t1 254.584
R42 A.n0 A.t4 231.629
R43 A.n3 A.t2 192.8
R44 A.n1 A.t7 162.274
R45 A.n4 A.t0 162.274
R46 A.n5 A.n4 152
R47 A.n2 A.n1 152
R48 A A.n5 62.6917
R49 A A.n2 1.67527
R50 VGND.n6 VGND.n5 236.218
R51 VGND.n11 VGND.n10 205.69
R52 VGND.n1 VGND.n0 203.681
R53 VGND.n8 VGND.n7 199.686
R54 VGND.n5 VGND.t4 66.563
R55 VGND.n7 VGND.t6 52.5005
R56 VGND.n0 VGND.t3 50.6255
R57 VGND.n10 VGND.t2 41.2505
R58 VGND.n10 VGND.t0 41.2505
R59 VGND.n5 VGND.t1 41.2505
R60 VGND.n7 VGND.t5 40.313
R61 VGND.n9 VGND.n8 36.1417
R62 VGND.n16 VGND.n3 36.1417
R63 VGND.n17 VGND.n16 36.1417
R64 VGND.n18 VGND.n17 36.1417
R65 VGND.n12 VGND.n3 33.6699
R66 VGND.n0 VGND.t7 25.524
R67 VGND.n18 VGND.n1 21.2197
R68 VGND.n11 VGND.n9 19.326
R69 VGND.n20 VGND.n1 9.62295
R70 VGND.n19 VGND.n18 9.3005
R71 VGND.n17 VGND.n2 9.3005
R72 VGND.n16 VGND.n15 9.3005
R73 VGND.n14 VGND.n3 9.3005
R74 VGND.n13 VGND.n12 9.3005
R75 VGND.n9 VGND.n4 9.3005
R76 VGND.n8 VGND.n6 4.27169
R77 VGND.n12 VGND.n11 2.97424
R78 VGND.n6 VGND.n4 0.203518
R79 VGND VGND.n20 0.161675
R80 VGND.n20 VGND.n19 0.146149
R81 VGND.n13 VGND.n4 0.122949
R82 VGND.n14 VGND.n13 0.122949
R83 VGND.n15 VGND.n14 0.122949
R84 VGND.n15 VGND.n2 0.122949
R85 VGND.n19 VGND.n2 0.122949
R86 a_501_75.n1 a_501_75.n0 436.305
R87 a_501_75.t0 a_501_75.n1 33.7505
R88 a_501_75.n1 a_501_75.t3 33.7505
R89 a_501_75.n0 a_501_75.t2 26.2505
R90 a_501_75.n0 a_501_75.t1 26.2505
R91 a_217_368.t0 a_217_368.t1 72.8687
R92 a_318_389.n1 a_318_389.n0 78.0571
R93 a_318_389.n0 a_318_389.t1 50.6238
R94 a_318_389.n0 a_318_389.t0 29.1182
R95 VPB.n0 VPB 3820.43
R96 VPB VPB.n1 725.192
R97 VPB.t3 VPB.t7 505.216
R98 VPB.t7 VPB.t1 403.69
R99 VPB.n0 VPB.t12 339.651
R100 VPB.t1 VPB.n0 285.243
R101 VPB.t2 VPB.t8 282.825
R102 VPB.t6 VPB.t10 263.038
R103 VPB.t10 VPB 252.823
R104 VPB.n1 VPB.t6 250.269
R105 VPB.t5 VPB.t3 244.149
R106 VPB.t8 VPB.t9 244.149
R107 VPB.t4 VPB.t0 244.149
R108 VPB.t11 VPB.t2 234.478
R109 VPB.t9 VPB.t5 222.393
R110 VPB.t0 VPB.t11 217.558
R111 VPB.n1 VPB.t4 3.72599
R112 CIN.n2 CIN.t0 231.629
R113 CIN.n4 CIN.t3 231.629
R114 CIN.n1 CIN.n0 231.629
R115 CIN.n2 CIN.t2 200.833
R116 CIN.n4 CIN.t1 200.833
R117 CIN.n1 CIN.t4 200.833
R118 CIN.n3 CIN.n1 185.625
R119 CIN CIN.n4 179.275
R120 CIN.n3 CIN.n2 170.494
R121 CIN CIN.n3 0.0466957
R122 a_509_347.n1 a_509_347.n0 943.649
R123 a_509_347.n0 a_509_347.t2 40.3855
R124 a_509_347.t0 a_509_347.n1 36.4455
R125 a_509_347.n0 a_509_347.t1 29.5505
R126 a_509_347.n1 a_509_347.t3 29.5505
R127 VPWR.n22 VPWR.n4 652.105
R128 VPWR.n16 VPWR.n15 618.359
R129 VPWR.n9 VPWR.n8 290.43
R130 VPWR.n10 VPWR.t8 256.14
R131 VPWR.n29 VPWR.n1 222.153
R132 VPWR.n8 VPWR.t5 63.7716
R133 VPWR.n8 VPWR.t1 55.9756
R134 VPWR.n4 VPWR.t2 43.3405
R135 VPWR.n1 VPWR.t3 42.3555
R136 VPWR.n4 VPWR.t0 42.3555
R137 VPWR.n23 VPWR.n2 36.1417
R138 VPWR.n27 VPWR.n2 36.1417
R139 VPWR.n28 VPWR.n27 36.1417
R140 VPWR.n21 VPWR.n5 36.1417
R141 VPWR.n13 VPWR.n7 36.1417
R142 VPWR.n14 VPWR.n13 36.1417
R143 VPWR.n17 VPWR.n14 36.1417
R144 VPWR.n23 VPWR.n22 33.1299
R145 VPWR.n15 VPWR.t4 31.5205
R146 VPWR.n15 VPWR.t6 29.5505
R147 VPWR.n1 VPWR.t7 27.4811
R148 VPWR.n29 VPWR.n28 23.7181
R149 VPWR.n22 VPWR.n21 14.3064
R150 VPWR.n17 VPWR.n16 9.41227
R151 VPWR.n11 VPWR.n7 9.3005
R152 VPWR.n13 VPWR.n12 9.3005
R153 VPWR.n14 VPWR.n6 9.3005
R154 VPWR.n18 VPWR.n17 9.3005
R155 VPWR.n19 VPWR.n5 9.3005
R156 VPWR.n21 VPWR.n20 9.3005
R157 VPWR.n22 VPWR.n3 9.3005
R158 VPWR.n24 VPWR.n23 9.3005
R159 VPWR.n25 VPWR.n2 9.3005
R160 VPWR.n27 VPWR.n26 9.3005
R161 VPWR.n28 VPWR.n0 9.3005
R162 VPWR.n9 VPWR.n7 9.03579
R163 VPWR.n30 VPWR.n29 7.23624
R164 VPWR.n10 VPWR.n9 5.97509
R165 VPWR.n16 VPWR.n5 1.88285
R166 VPWR.n11 VPWR.n10 0.275151
R167 VPWR VPWR.n30 0.157488
R168 VPWR.n30 VPWR.n0 0.150282
R169 VPWR.n12 VPWR.n11 0.122949
R170 VPWR.n12 VPWR.n6 0.122949
R171 VPWR.n18 VPWR.n6 0.122949
R172 VPWR.n19 VPWR.n18 0.122949
R173 VPWR.n20 VPWR.n19 0.122949
R174 VPWR.n20 VPWR.n3 0.122949
R175 VPWR.n24 VPWR.n3 0.122949
R176 VPWR.n25 VPWR.n24 0.122949
R177 VPWR.n26 VPWR.n25 0.122949
R178 VPWR.n26 VPWR.n0 0.122949
R179 a_315_75.t0 a_315_75.t1 45.0005
R180 a_69_260.n2 a_69_260.n0 338.69
R181 a_69_260.n3 a_69_260.n2 329.421
R182 a_69_260.n1 a_69_260.t5 264.298
R183 a_69_260.n1 a_69_260.t4 204.048
R184 a_69_260.n2 a_69_260.n1 152
R185 a_69_260.n0 a_69_260.t3 46.8755
R186 a_69_260.n3 a_69_260.t2 29.5505
R187 a_69_260.t1 a_69_260.n3 29.5505
R188 a_69_260.n0 a_69_260.t0 26.2505
R189 a_1100_75.t0 a_1100_75.n0 400.389
R190 a_1100_75.n0 a_1100_75.t2 67.2514
R191 a_1100_75.n0 a_1100_75.t1 62.1182
R192 SUM.n0 SUM.t0 299.301
R193 SUM.t1 SUM.n0 279.738
R194 SUM.n1 SUM.t1 279.738
R195 SUM.n1 SUM 14.8576
R196 SUM.n0 SUM 5.71479
R197 SUM SUM.n1 2.05764
R198 a_237_75.t0 a_237_75.t1 45.0005
R199 COUT.n1 COUT 591.274
R200 COUT.n1 COUT.n0 585
R201 COUT.n2 COUT.n1 585
R202 COUT.n1 COUT.t0 26.3844
R203 COUT.n2 COUT 16.8162
R204 COUT.n3 COUT 15.1211
R205 COUT.n0 COUT 14.5574
R206 COUT COUT.n3 13.978
R207 COUT.n0 COUT 4.01619
R208 COUT COUT.n2 1.75736
R209 COUT.n3 COUT 0.105043
R210 a_916_347.t0 a_916_347.t1 69.9355
R211 a_1107_347.t0 a_1107_347.t1 871.835
C0 VPWR COUT 0.121788f
C1 A CIN 0.467379f
C2 A COUT 1.67e-19
C3 CIN COUT 9.18e-20
C4 VPB B 0.627254f
C5 VPB SUM 0.012825f
C6 VPB VGND 0.013021f
C7 B SUM 1.72e-19
C8 VPB VPWR 0.245734f
C9 B VGND 0.040329f
C10 B VPWR 0.219558f
C11 VPB A 0.143253f
C12 SUM VGND 0.037599f
C13 SUM VPWR 0.105041f
C14 B A 0.26846f
C15 VPB CIN 0.123233f
C16 VPWR VGND 0.084645f
C17 VPB COUT 0.014191f
C18 B CIN 0.195912f
C19 SUM A 7.32e-19
C20 A VGND 0.131515f
C21 VPWR A 0.049123f
C22 SUM CIN 4.08e-19
C23 B COUT 0.006875f
C24 CIN VGND 0.137887f
C25 VPWR CIN 0.134937f
C26 COUT VGND 0.074187f
C27 VGND VNB 0.998021f
C28 COUT VNB 0.11284f
C29 CIN VNB 0.315731f
C30 A VNB 0.498853f
C31 VPWR VNB 0.790121f
C32 SUM VNB 0.116945f
C33 B VNB 0.612386f
C34 VPB VNB 2.08861f
.ends

* NGSPICE file created from sky130_fd_sc_hs__einvp_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__einvp_8 VNB VPB VPWR VGND Z TE A
X0 a_27_74.t7 TE.t0 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 VPWR.t6 a_802_323.t2 a_27_368# VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_27_368# A.t0 Z.t7 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_27_74.t13 A.t1 Z.t15 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 Z.t6 A.t2 a_27_368# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_27_74.t14 A.t3 Z.t14 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X6 a_27_74.t6 TE.t1 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 a_27_368# A.t4 Z.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Z.t13 A.t5 a_27_74.t15 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 Z.t4 A.t6 a_27_368# VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_27_74.t5 TE.t2 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VGND.t4 TE.t3 a_27_74.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_27_368# A.t7 Z.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VPWR.t0 TE.t4 a_802_323.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.3192 ps=2.81 w=1.12 l=0.15
X14 Z.t2 A.t8 a_27_368# VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_27_368# A.t9 Z.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 Z.t12 A.t10 a_27_74.t8 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 Z.t11 A.t11 a_27_74.t9 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 VGND.t3 TE.t5 a_27_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 VGND.t2 TE.t6 a_27_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_27_368# a_802_323.t3 VPWR.t5 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_27_74.t10 A.t12 Z.t10 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X22 a_27_74.t11 A.t13 Z.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 VGND.t1 TE.t7 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_27_368# a_802_323.t4 VPWR.t4 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 VPWR.t3 a_802_323.t5 a_27_368# VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 Z.t0 A.t14 a_27_368# VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
X27 a_27_368# a_802_323.t6 VPWR.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 a_27_368# a_802_323.t7 VPWR.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 a_27_74.t0 TE.t8 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 Z.t8 A.t15 a_27_74.t12 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X31 VGND.t8 TE.t9 a_802_323.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2146 ps=2.06 w=0.74 l=0.15
R0 TE.n0 TE.t3 314.908
R1 TE.n7 TE.n6 298.841
R2 TE.n8 TE.t4 285.719
R3 TE.n7 TE.t9 165.196
R4 TE TE.n8 162.44
R5 TE.n6 TE.n5 160.667
R6 TE.n0 TE.t0 154.24
R7 TE.n1 TE.t7 154.24
R8 TE.n2 TE.t8 154.24
R9 TE.n3 TE.t6 154.24
R10 TE.n4 TE.t2 154.24
R11 TE.n5 TE.t5 154.24
R12 TE.n6 TE.t1 154.24
R13 TE.n5 TE.n4 138.173
R14 TE.n4 TE.n3 138.173
R15 TE.n3 TE.n2 138.173
R16 TE.n2 TE.n1 138.173
R17 TE.n1 TE.n0 138.173
R18 TE.n8 TE.n7 13.146
R19 VGND.n4 VGND.t8 151.28
R20 VGND.n16 VGND.n15 116.334
R21 VGND.n6 VGND.n5 116.332
R22 VGND.n9 VGND.n8 116.332
R23 VGND.n13 VGND.n2 116.332
R24 VGND.n5 VGND.t3 34.0546
R25 VGND.n15 VGND.t7 34.0546
R26 VGND.n9 VGND.n7 32.7534
R27 VGND.n13 VGND.n1 25.224
R28 VGND.n16 VGND.n14 22.9652
R29 VGND.n5 VGND.t6 22.7032
R30 VGND.n8 VGND.t5 22.7032
R31 VGND.n8 VGND.t2 22.7032
R32 VGND.n2 VGND.t0 22.7032
R33 VGND.n2 VGND.t1 22.7032
R34 VGND.n15 VGND.t4 22.7032
R35 VGND.n14 VGND.n13 22.2123
R36 VGND.n9 VGND.n1 14.6829
R37 VGND.n7 VGND.n6 12.424
R38 VGND.n7 VGND.n3 9.3005
R39 VGND.n10 VGND.n9 9.3005
R40 VGND.n11 VGND.n1 9.3005
R41 VGND.n13 VGND.n12 9.3005
R42 VGND.n14 VGND.n0 9.3005
R43 VGND.n6 VGND.n4 7.54482
R44 VGND.n17 VGND.n16 7.18706
R45 VGND VGND.n17 1.13525
R46 VGND.n4 VGND.n3 0.219331
R47 VGND.n17 VGND.n0 0.156777
R48 VGND.n10 VGND.n3 0.122949
R49 VGND.n11 VGND.n10 0.122949
R50 VGND.n12 VGND.n11 0.122949
R51 VGND.n12 VGND.n0 0.122949
R52 a_27_74.n10 a_27_74.t6 213.499
R53 a_27_74.n1 a_27_74.t15 193.952
R54 a_27_74.n1 a_27_74.n0 185
R55 a_27_74.n3 a_27_74.n2 185
R56 a_27_74.n5 a_27_74.n4 185
R57 a_27_74.n11 a_27_74.n8 118.709
R58 a_27_74.n10 a_27_74.n9 114.82
R59 a_27_74.n13 a_27_74.n12 114.82
R60 a_27_74.n12 a_27_74.n7 91.568
R61 a_27_74.n7 a_27_74.n5 84.9866
R62 a_27_74.n7 a_27_74.n6 84.741
R63 a_27_74.n3 a_27_74.n1 60.6259
R64 a_27_74.n5 a_27_74.n3 60.6259
R65 a_27_74.n11 a_27_74.n10 58.3534
R66 a_27_74.n12 a_27_74.n11 58.3534
R67 a_27_74.n4 a_27_74.t10 34.0546
R68 a_27_74.n2 a_27_74.t14 34.0546
R69 a_27_74.n0 a_27_74.t11 34.0546
R70 a_27_74.n9 a_27_74.t3 22.7032
R71 a_27_74.n9 a_27_74.t5 22.7032
R72 a_27_74.n8 a_27_74.t2 22.7032
R73 a_27_74.n8 a_27_74.t0 22.7032
R74 a_27_74.n6 a_27_74.t4 22.7032
R75 a_27_74.n6 a_27_74.t13 22.7032
R76 a_27_74.n4 a_27_74.t8 22.7032
R77 a_27_74.n2 a_27_74.t12 22.7032
R78 a_27_74.n0 a_27_74.t9 22.7032
R79 a_27_74.n13 a_27_74.t1 22.7032
R80 a_27_74.t7 a_27_74.n13 22.7032
R81 VNB.t7 VNB.t0 2425.2
R82 VNB.t4 VNB.t7 1154.86
R83 VNB.t5 VNB.t8 1154.86
R84 VNB.t9 VNB.t14 1154.86
R85 VNB.t11 VNB.t9 1154.86
R86 VNB.t13 VNB.t11 1154.86
R87 VNB.t15 VNB.t13 1154.86
R88 VNB.t10 VNB.t15 1154.86
R89 VNB.t12 VNB.t10 1154.86
R90 VNB VNB.t16 1143.31
R91 VNB.t6 VNB.t4 993.177
R92 VNB.t3 VNB.t6 993.177
R93 VNB.t1 VNB.t3 993.177
R94 VNB.t2 VNB.t1 993.177
R95 VNB.t8 VNB.t2 993.177
R96 VNB.t14 VNB.t5 993.177
R97 VNB.t16 VNB.t12 993.177
R98 a_802_323.n2 a_802_323.t2 348.647
R99 a_802_323.n9 a_802_323.n8 247.726
R100 a_802_323.t0 a_802_323.n9 224.657
R101 a_802_323.n8 a_802_323.t3 204.048
R102 a_802_323.n7 a_802_323.n0 204.048
R103 a_802_323.n6 a_802_323.t4 204.048
R104 a_802_323.n5 a_802_323.n1 204.048
R105 a_802_323.n4 a_802_323.t7 204.048
R106 a_802_323.n3 a_802_323.t5 204.048
R107 a_802_323.n2 a_802_323.t6 204.048
R108 a_802_323.n9 a_802_323.t1 192.237
R109 a_802_323.n8 a_802_323.n7 144.601
R110 a_802_323.n7 a_802_323.n6 144.601
R111 a_802_323.n6 a_802_323.n5 144.601
R112 a_802_323.n5 a_802_323.n4 144.601
R113 a_802_323.n4 a_802_323.n3 144.601
R114 a_802_323.n3 a_802_323.n2 144.601
R115 VPWR.n1 VPWR.n0 315.349
R116 VPWR.n5 VPWR.t0 266.916
R117 VPWR.n4 VPWR.t4 258.238
R118 VPWR.n6 VPWR.t5 258.238
R119 VPWR.n12 VPWR.n3 242.582
R120 VPWR.n14 VPWR.n13 36.1417
R121 VPWR.n11 VPWR.n4 33.1299
R122 VPWR.n7 VPWR.n6 28.6123
R123 VPWR.n0 VPWR.t2 26.3844
R124 VPWR.n0 VPWR.t6 26.3844
R125 VPWR.n3 VPWR.t1 26.3844
R126 VPWR.n3 VPWR.t3 26.3844
R127 VPWR.n12 VPWR.n11 22.2123
R128 VPWR.n7 VPWR.n4 20.3299
R129 VPWR.n13 VPWR.n12 13.9299
R130 VPWR.n16 VPWR.n1 13.674
R131 VPWR.n8 VPWR.n7 9.3005
R132 VPWR.n9 VPWR.n4 9.3005
R133 VPWR.n11 VPWR.n10 9.3005
R134 VPWR.n13 VPWR.n2 9.3005
R135 VPWR.n15 VPWR.n14 9.3005
R136 VPWR.n6 VPWR.n5 7.1933
R137 VPWR.n14 VPWR.n1 5.27109
R138 VPWR VPWR.n16 1.01964
R139 VPWR.n8 VPWR.n5 0.169199
R140 VPWR.n16 VPWR.n15 0.149471
R141 VPWR.n9 VPWR.n8 0.122949
R142 VPWR.n10 VPWR.n9 0.122949
R143 VPWR.n10 VPWR.n2 0.122949
R144 VPWR.n15 VPWR.n2 0.122949
R145 VPB.t13 VPB.t0 702.285
R146 VPB.t12 VPB.t13 459.678
R147 VPB.t9 VPB.t12 459.678
R148 VPB VPB.t3 255.376
R149 VPB.t11 VPB.t9 229.839
R150 VPB.t10 VPB.t11 229.839
R151 VPB.t14 VPB.t10 229.839
R152 VPB.t4 VPB.t14 229.839
R153 VPB.t5 VPB.t4 229.839
R154 VPB.t6 VPB.t5 229.839
R155 VPB.t7 VPB.t6 229.839
R156 VPB.t8 VPB.t7 229.839
R157 VPB.t1 VPB.t8 229.839
R158 VPB.t2 VPB.t1 229.839
R159 VPB.t3 VPB.t2 229.839
R160 A.n4 A.t0 261.62
R161 A.n7 A.t2 261.62
R162 A.n10 A.t4 261.62
R163 A.n2 A.t6 261.62
R164 A.n18 A.t7 261.62
R165 A.n24 A.t8 261.62
R166 A.n22 A.t9 261.62
R167 A.n19 A.t14 261.62
R168 A.n4 A.t1 226.833
R169 A.n6 A 160.995
R170 A.n19 A.t5 154.97
R171 A.n21 A.t13 154.24
R172 A.n25 A.t11 154.24
R173 A.n17 A.t3 154.24
R174 A.n11 A.t15 154.24
R175 A.n9 A.t12 154.24
R176 A.n5 A.t10 154.24
R177 A.n8 A.n3 152
R178 A.n13 A.n12 152
R179 A.n15 A.n14 152
R180 A.n16 A.n0 152
R181 A A.n26 152
R182 A.n23 A.n1 152
R183 A.n20 A 75.0379
R184 A.n16 A.n15 49.6611
R185 A.n23 A.n22 44.549
R186 A.n26 A.n18 37.246
R187 A.n8 A.n7 35.7853
R188 A.n20 A.n19 33.2107
R189 A.n5 A.n4 32.8641
R190 A.n12 A.n11 27.752
R191 A.n10 A.n9 25.5611
R192 A.n26 A.n25 24.8308
R193 A.n21 A.n20 22.1183
R194 A.n24 A.n23 21.1793
R195 A.n12 A.n10 19.7187
R196 A.n6 A.n5 18.9884
R197 A.n11 A.n2 18.2581
R198 A.n7 A.n6 13.8763
R199 A.n13 A.n3 11.7627
R200 A A.n0 11.7627
R201 A A.n1 11.7627
R202 A.n18 A.n17 10.955
R203 A.n14 A 9.68699
R204 A.n14 A 6.91942
R205 A A.n0 4.84374
R206 A A.n1 4.84374
R207 A.n9 A.n8 4.38232
R208 A.n15 A.n2 3.65202
R209 A.n25 A.n24 3.65202
R210 A.n22 A.n21 3.65202
R211 A A.n3 2.76807
R212 A A.n13 2.07618
R213 A.n17 A.n16 1.46111
R214 Z.n9 Z.n7 251.495
R215 Z.n2 Z.n0 246.142
R216 Z.n9 Z.n8 208.577
R217 Z.n11 Z.n10 208.577
R218 Z.n13 Z.n12 208.577
R219 Z.n6 Z.n5 191.4
R220 Z.n2 Z.n1 185
R221 Z.n4 Z.n3 185
R222 Z.n4 Z.n2 61.1412
R223 Z.n6 Z.n4 55.7944
R224 Z.n14 Z.n6 43.9563
R225 Z.n11 Z.n9 42.9181
R226 Z.n13 Z.n11 42.9181
R227 Z.n5 Z.t12 34.0546
R228 Z.n3 Z.t8 34.0546
R229 Z.n1 Z.t11 34.0546
R230 Z.n7 Z.t1 26.3844
R231 Z.n7 Z.t0 26.3844
R232 Z.n8 Z.t3 26.3844
R233 Z.n8 Z.t2 26.3844
R234 Z.n10 Z.t5 26.3844
R235 Z.n10 Z.t4 26.3844
R236 Z.n12 Z.t7 26.3844
R237 Z.n12 Z.t6 26.3844
R238 Z.n5 Z.t15 22.7032
R239 Z.n3 Z.t10 22.7032
R240 Z.n1 Z.t14 22.7032
R241 Z.n0 Z.t9 22.7032
R242 Z.n0 Z.t13 22.7032
R243 Z.n14 Z.n13 11.8593
R244 Z Z.n14 7.71815
C0 VPB A 0.267586f
C1 VPB Z 0.015855f
C2 VPB a_27_368# 0.051938f
C3 VPB VPWR 0.225288f
C4 A Z 0.784718f
C5 A a_27_368# 0.14531f
C6 VPB TE 0.047284f
C7 A VPWR 0.04813f
C8 Z a_27_368# 0.73735f
C9 A TE 0.023116f
C10 VPB VGND 0.009263f
C11 Z VPWR 0.044023f
C12 VPWR a_27_368# 1.29105f
C13 Z TE 2.14e-20
C14 A VGND 0.054399f
C15 TE a_27_368# 0.00524f
C16 Z VGND 0.043475f
C17 VPWR TE 0.039131f
C18 VGND a_27_368# 0.019522f
C19 VPWR VGND 0.144305f
C20 TE VGND 0.195169f
C21 VGND VNB 1.0572f
C22 TE VNB 0.781246f
C23 VPWR VNB 0.876472f
C24 Z VNB 0.030757f
C25 A VNB 0.899406f
C26 VPB VNB 2.1204f
C27 a_27_368# VNB 0.081301f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fa_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fa_2 VNB VPB VPWR A VGND CIN B COUT SUM
X0 a_1202_368.t1 B.t0 a_1094_347.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.20235 ps=1.495 w=1 l=0.15
X1 VGND.t7 A.t0 a_27_79.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.18315 pd=1.235 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 a_487_79.t1 B.t1 a_336_347.t2 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 VGND A a_1205_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.25365 pd=1.52 as=0.0888 ps=0.98 w=0.74 l=0.15
X4 a_992_347.t1 a_336_347.t4 a_683_347.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X5 COUT.t1 a_336_347.t5 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2212 pd=1.515 as=0.2277 ps=1.54 w=1.12 l=0.15
X6 a_336_347.t0 CIN.t0 a_27_378.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=1.59 as=0.15 ps=1.3 w=1 l=0.15
X7 VPWR.t7 A.t1 a_484_347.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2125 pd=1.425 as=0.135 ps=1.27 w=1 l=0.15
X8 a_683_347.t2 A.t2 VPWR.t6 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.23355 ps=1.595 w=1 l=0.15
X9 a_701_79.t1 CIN.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=1.27 w=0.74 l=0.15
X10 VGND.t1 a_336_347.t6 COUT.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.251275 pd=1.515 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_27_378.t2 B.t2 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.26355 ps=1.655 w=1 l=0.15
X12 a_484_347.t1 B.t3 a_336_347.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=1.59 w=1 l=0.15
X13 VGND.t3 a_992_347.t3 SUM.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_1094_347.t1 CIN.t2 a_992_347.t2 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.20235 pd=1.495 as=0.18 ps=1.36 w=1 l=0.15
X15 a_992_347.t0 a_336_347.t7 a_701_79.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 VGND.t8 B.t4 a_701_79.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.193975 pd=1.395 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_336_347.t1 CIN.t3 a_27_79.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=1.31 w=0.74 l=0.15
X18 VPWR.t1 a_336_347.t8 COUT.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3024 pd=1.66 as=0.2212 ps=1.515 w=1.12 l=0.15
X19 a_683_347.t1 CIN.t4 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.19105 pd=1.51 as=0.2125 ps=1.425 w=1 l=0.15
X20 COUT.t2 a_336_347.t9 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.25365 ps=1.52 w=0.74 l=0.15
X21 a_701_79.t2 A.t3 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.193975 ps=1.395 w=0.74 l=0.15
X22 SUM.t1 a_992_347.t4 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.251275 ps=1.515 w=0.74 l=0.15
X23 VGND.t5 A.t4 a_487_79.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=1.27 as=0.0888 ps=0.98 w=0.74 l=0.15
X24 a_1205_79# B.t5 a_1119_79# VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 VPWR.t8 B.t6 a_683_347.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.23355 pd=1.595 as=0.19105 ps=1.51 w=1 l=0.15
X26 VPWR.t5 A.t5 a_27_378.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.26355 pd=1.655 as=0.295 ps=2.59 w=1 l=0.15
X27 VPWR.t3 a_992_347.t5 SUM.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X28 VPWR.t4 A.t6 a_1202_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.54 as=0.135 ps=1.27 w=1 l=0.15
X29 a_27_79.t2 B.t7 VGND.t9 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=1.31 as=0.18315 ps=1.235 w=0.74 l=0.15
R0 B.n0 B.t0 861.442
R1 B.t2 B.n1 600.359
R2 B.t6 B.t4 489.767
R3 B.t0 B.t5 476.377
R4 B.t3 B.t1 448.26
R5 B.n1 B.n0 424.161
R6 B.n1 B.t3 275.812
R7 B.n0 B.t6 234.306
R8 B.n2 B.t2 230.526
R9 B B.n2 194.073
R10 B.n2 B.t7 175.169
R11 a_1094_347.t0 a_1094_347.t1 80.5726
R12 a_1202_368.t0 a_1202_368.t1 53.1905
R13 VPB.n0 VPB 3021.1
R14 VPB.t8 VPB.t9 582.259
R15 VPB.n1 VPB 570
R16 VPB.t2 VPB.t11 357.762
R17 VPB VPB.n1 306.998
R18 VPB.t5 VPB.t7 291.13
R19 VPB.t10 VPB.t4 285.243
R20 VPB.t7 VPB.t8 278.361
R21 VPB.t3 VPB.t1 277.99
R22 VPB.t14 VPB.n0 251.399
R23 VPB.n1 VPB.t12 251.399
R24 VPB.t6 VPB.t14 246.565
R25 VPB.t1 VPB.t10 244.149
R26 VPB.n1 VPB.t0 230.304
R27 VPB.t4 VPB.t6 217.558
R28 VPB.t12 VPB.t2 217.558
R29 VPB.t13 VPB.t5 214.517
R30 VPB.t11 VPB.t3 203.054
R31 VPB.n0 VPB.t13 4.96782
R32 A.n6 A.t5 252.192
R33 A.n4 A.t1 231.629
R34 A.n2 A.t2 231.629
R35 A.n1 A.t6 231.629
R36 A.n1 A.n0 212.081
R37 A.n6 A.t0 189.018
R38 A.n4 A.t4 178.34
R39 A.n2 A.t3 178.34
R40 A.n3 A.n2 177.686
R41 A.n5 A.n4 174.436
R42 A.n3 A.n1 169.161
R43 A.n7 A.n6 169.059
R44 A.n7 A.n5 2.04204
R45 A.n5 A.n3 1.18489
R46 A A.n7 0.0466957
R47 a_27_79.n0 a_27_79.t1 404.24
R48 a_27_79.t0 a_27_79.n0 46.2167
R49 a_27_79.n0 a_27_79.t2 46.2167
R50 VGND.n13 VGND.t2 285.272
R51 VGND.n21 VGND.n20 213.966
R52 VGND.n36 VGND.n35 213.417
R53 VGND.n8 VGND.n7 206.952
R54 VGND.n28 VGND.n27 198.554
R55 VGND.n9 VGND.t3 180.136
R56 VGND.n27 VGND.t0 48.6491
R57 VGND.n35 VGND.t9 46.2167
R58 VGND.n7 VGND.t4 45.4059
R59 VGND.n7 VGND.t1 45.4059
R60 VGND.n27 VGND.t5 37.2978
R61 VGND.n12 VGND.n11 36.1417
R62 VGND.n18 VGND.n5 36.1417
R63 VGND.n19 VGND.n18 36.1417
R64 VGND.n22 VGND.n19 36.1417
R65 VGND.n29 VGND.n1 36.1417
R66 VGND.n33 VGND.n1 36.1417
R67 VGND.n34 VGND.n33 36.1417
R68 VGND.n20 VGND.t6 35.6762
R69 VGND.n20 VGND.t8 35.6762
R70 VGND.n14 VGND.n5 35.65
R71 VGND.n35 VGND.t7 34.0546
R72 VGND.n26 VGND.n3 31.6925
R73 VGND.n36 VGND.n34 25.224
R74 VGND.n22 VGND.n21 22.3378
R75 VGND.n28 VGND.n26 21.8358
R76 VGND.n11 VGND.n8 19.0545
R77 VGND.n29 VGND.n28 12.0476
R78 VGND.n34 VGND.n0 9.3005
R79 VGND.n33 VGND.n32 9.3005
R80 VGND.n31 VGND.n1 9.3005
R81 VGND.n30 VGND.n29 9.3005
R82 VGND.n28 VGND.n2 9.3005
R83 VGND.n26 VGND.n25 9.3005
R84 VGND.n24 VGND.n3 9.3005
R85 VGND.n23 VGND.n22 9.3005
R86 VGND.n19 VGND.n4 9.3005
R87 VGND.n18 VGND.n17 9.3005
R88 VGND.n16 VGND.n5 9.3005
R89 VGND.n15 VGND.n14 9.3005
R90 VGND.n12 VGND.n6 9.3005
R91 VGND.n11 VGND.n10 9.3005
R92 VGND.n9 VGND.n8 9.08752
R93 VGND.n13 VGND.n12 8.64396
R94 VGND.n37 VGND.n36 7.43488
R95 VGND.n14 VGND.n13 5.61683
R96 VGND.n21 VGND.n3 1.93989
R97 VGND.n10 VGND.n9 0.539608
R98 VGND VGND.n37 0.160103
R99 VGND.n37 VGND.n0 0.1477
R100 VGND.n10 VGND.n6 0.122949
R101 VGND.n15 VGND.n6 0.122949
R102 VGND.n16 VGND.n15 0.122949
R103 VGND.n17 VGND.n16 0.122949
R104 VGND.n17 VGND.n4 0.122949
R105 VGND.n23 VGND.n4 0.122949
R106 VGND.n24 VGND.n23 0.122949
R107 VGND.n25 VGND.n24 0.122949
R108 VGND.n25 VGND.n2 0.122949
R109 VGND.n30 VGND.n2 0.122949
R110 VGND.n31 VGND.n30 0.122949
R111 VGND.n32 VGND.n31 0.122949
R112 VGND.n32 VGND.n0 0.122949
R113 VNB VNB.n0 13661.9
R114 VNB.t11 VNB.t3 2552.23
R115 VNB.n0 VNB.t2 2187.78
R116 VNB.t6 VNB.t10 1760
R117 VNB.t0 VNB.t7 1662.22
R118 VNB.t1 VNB.t5 1639.9
R119 VNB.t10 VNB.t9 1576.67
R120 VNB.t8 VNB.t12 1442.22
R121 VNB.t2 VNB.t8 1393.33
R122 VNB.t13 VNB.t6 1222.22
R123 VNB.t9 VNB 1210
R124 VNB.t12 VNB.t0 1051.11
R125 VNB.t5 VNB.t4 993.177
R126 VNB.t3 VNB.t1 993.177
R127 VNB.t7 VNB.t13 953.333
R128 VNB.n0 VNB.t11 41.566
R129 a_336_347.n7 a_336_347.n6 735.063
R130 a_336_347.n0 a_336_347.t8 320.531
R131 a_336_347.n4 a_336_347.n2 301.846
R132 a_336_347.n2 a_336_347.t5 276.348
R133 a_336_347.n3 a_336_347.t4 231.629
R134 a_336_347.n6 a_336_347.n4 184.847
R135 a_336_347.n3 a_336_347.t7 178.34
R136 a_336_347.n0 a_336_347.t6 177.537
R137 a_336_347.n1 a_336_347.t9 168.409
R138 a_336_347.n4 a_336_347.n3 167.709
R139 a_336_347.n6 a_336_347.n5 99.193
R140 a_336_347.n1 a_336_347.n0 69.0872
R141 a_336_347.t0 a_336_347.n7 63.0405
R142 a_336_347.n7 a_336_347.t3 53.1905
R143 a_336_347.n5 a_336_347.t1 34.0546
R144 a_336_347.n5 a_336_347.t2 22.7032
R145 a_336_347.n2 a_336_347.n1 13.146
R146 a_487_79.t0 a_487_79.t1 38.9194
R147 a_683_347.n1 a_683_347.n0 1236.48
R148 a_683_347.n0 a_683_347.t3 43.1876
R149 a_683_347.n0 a_683_347.t1 32.9336
R150 a_683_347.t0 a_683_347.n1 29.5505
R151 a_683_347.n1 a_683_347.t2 29.5505
R152 a_992_347.n5 a_992_347.n4 550.751
R153 a_992_347.n4 a_992_347.t0 461.788
R154 a_992_347.n1 a_992_347.t5 303.125
R155 a_992_347.n3 a_992_347.n0 256.63
R156 a_992_347.n1 a_992_347.t3 198.423
R157 a_992_347.n2 a_992_347.t4 188.244
R158 a_992_347.n4 a_992_347.n3 152
R159 a_992_347.n2 a_992_347.n1 80.3338
R160 a_992_347.t1 a_992_347.n5 41.3705
R161 a_992_347.n5 a_992_347.t2 29.5505
R162 a_992_347.n3 a_992_347.n2 11.8854
R163 VPWR.n11 VPWR.t1 736.399
R164 VPWR.n28 VPWR.n4 618.939
R165 VPWR.n6 VPWR.n5 610.078
R166 VPWR.n35 VPWR.n1 608.763
R167 VPWR.n16 VPWR.n10 606.333
R168 VPWR.n12 VPWR.t3 266.233
R169 VPWR.n1 VPWR.t9 65.3355
R170 VPWR.n5 VPWR.t6 58.3414
R171 VPWR.n4 VPWR.t2 54.1755
R172 VPWR.n10 VPWR.t4 53.1905
R173 VPWR.n1 VPWR.t5 37.0978
R174 VPWR.n29 VPWR.n2 36.1417
R175 VPWR.n33 VPWR.n2 36.1417
R176 VPWR.n34 VPWR.n33 36.1417
R177 VPWR.n17 VPWR.n8 36.1417
R178 VPWR.n21 VPWR.n8 36.1417
R179 VPWR.n22 VPWR.n21 36.1417
R180 VPWR.n23 VPWR.n22 36.1417
R181 VPWR.n15 VPWR.n14 36.1417
R182 VPWR.n5 VPWR.t8 33.7157
R183 VPWR.n28 VPWR.n27 33.5064
R184 VPWR.n4 VPWR.t7 29.5505
R185 VPWR.n10 VPWR.t0 26.8503
R186 VPWR.n27 VPWR.n6 22.9652
R187 VPWR.n23 VPWR.n6 20.3299
R188 VPWR.n35 VPWR.n34 14.3064
R189 VPWR.n29 VPWR.n28 13.9299
R190 VPWR.n14 VPWR.n11 11.6354
R191 VPWR.n12 VPWR.n11 9.41126
R192 VPWR.n14 VPWR.n13 9.3005
R193 VPWR.n15 VPWR.n9 9.3005
R194 VPWR.n18 VPWR.n17 9.3005
R195 VPWR.n19 VPWR.n8 9.3005
R196 VPWR.n21 VPWR.n20 9.3005
R197 VPWR.n22 VPWR.n7 9.3005
R198 VPWR.n24 VPWR.n23 9.3005
R199 VPWR.n25 VPWR.n6 9.3005
R200 VPWR.n27 VPWR.n26 9.3005
R201 VPWR.n28 VPWR.n3 9.3005
R202 VPWR.n30 VPWR.n29 9.3005
R203 VPWR.n31 VPWR.n2 9.3005
R204 VPWR.n33 VPWR.n32 9.3005
R205 VPWR.n34 VPWR.n0 9.3005
R206 VPWR.n36 VPWR.n35 7.43488
R207 VPWR.n16 VPWR.n15 7.15344
R208 VPWR.n17 VPWR.n16 4.14168
R209 VPWR.n13 VPWR.n12 0.54513
R210 VPWR VPWR.n36 0.160103
R211 VPWR.n36 VPWR.n0 0.1477
R212 VPWR.n13 VPWR.n9 0.122949
R213 VPWR.n18 VPWR.n9 0.122949
R214 VPWR.n19 VPWR.n18 0.122949
R215 VPWR.n20 VPWR.n19 0.122949
R216 VPWR.n20 VPWR.n7 0.122949
R217 VPWR.n24 VPWR.n7 0.122949
R218 VPWR.n25 VPWR.n24 0.122949
R219 VPWR.n26 VPWR.n25 0.122949
R220 VPWR.n26 VPWR.n3 0.122949
R221 VPWR.n30 VPWR.n3 0.122949
R222 VPWR.n31 VPWR.n30 0.122949
R223 VPWR.n32 VPWR.n31 0.122949
R224 VPWR.n32 VPWR.n0 0.122949
R225 COUT COUT.n1 591.207
R226 COUT COUT.n0 259.861
R227 COUT.n1 COUT.t0 35.1791
R228 COUT.n1 COUT.t1 34.2996
R229 COUT.n0 COUT.t3 22.7032
R230 COUT.n0 COUT.t2 22.7032
R231 CIN.n4 CIN.n3 288.849
R232 CIN CIN.n1 265.281
R233 CIN.n1 CIN.t2 231.629
R234 CIN.n2 CIN.t4 231.629
R235 CIN.n3 CIN.t0 222.534
R236 CIN.n4 CIN.n2 185.506
R237 CIN.n1 CIN.n0 178.34
R238 CIN.n2 CIN.t1 178.34
R239 CIN.n3 CIN.t3 169.246
R240 CIN CIN.n4 3.27492
R241 a_27_378.n0 a_27_378.t1 581.686
R242 a_27_378.t0 a_27_378.n0 29.5505
R243 a_27_378.n0 a_27_378.t2 29.5505
R244 a_484_347.t0 a_484_347.t1 53.1905
R245 a_701_79.n1 a_701_79.n0 436.7
R246 a_701_79.t0 a_701_79.n1 34.0546
R247 a_701_79.n1 a_701_79.t2 34.0546
R248 a_701_79.n0 a_701_79.t3 22.7032
R249 a_701_79.n0 a_701_79.t1 22.7032
R250 SUM.n2 SUM 589.508
R251 SUM.n2 SUM.n0 585
R252 SUM.n3 SUM.n2 585
R253 SUM SUM.n1 158.159
R254 SUM.n2 SUM.t0 26.3844
R255 SUM.n1 SUM.t2 22.7032
R256 SUM.n1 SUM.t1 22.7032
R257 SUM SUM.n3 12.0794
R258 SUM SUM.n0 10.4568
R259 SUM SUM.n0 2.88501
R260 SUM.n3 SUM 1.26247
C0 VPWR CIN 0.105655f
C1 B SUM 1.69e-19
C2 VPB VGND 0.00755f
C3 A COUT 0.007517f
C4 B VGND 0.032701f
C5 A SUM 4.98e-19
C6 VPWR COUT 0.023897f
C7 A VGND 0.241047f
C8 VPWR SUM 0.162442f
C9 CIN COUT 0.00406f
C10 a_1119_79# A 0.001523f
C11 VPWR VGND 0.05691f
C12 CIN SUM 1.34e-19
C13 a_1205_79# A 0.001305f
C14 CIN VGND 0.029937f
C15 COUT SUM 0.001997f
C16 VPB B 0.548733f
C17 a_1119_79# CIN 5.46e-20
C18 COUT VGND 0.010872f
C19 a_1119_79# COUT 1.33e-20
C20 VPB A 0.191678f
C21 SUM VGND 0.105137f
C22 a_1205_79# COUT 1.76e-20
C23 B A 0.346741f
C24 VPB VPWR 0.244133f
C25 a_1119_79# SUM 1.71e-19
C26 a_1205_79# SUM 1.99e-19
C27 a_1119_79# VGND 0.003178f
C28 B VPWR 0.199214f
C29 VPB CIN 0.127913f
C30 A VPWR 0.249947f
C31 VPB COUT 0.004893f
C32 a_1205_79# VGND 0.002504f
C33 B CIN 0.276382f
C34 A CIN 0.393197f
C35 VPB SUM 0.006048f
C36 B COUT 7.04e-19
C37 VGND VNB 1.0947f
C38 SUM VNB 0.030565f
C39 COUT VNB 0.010236f
C40 CIN VNB 0.297887f
C41 VPWR VNB 0.870643f
C42 A VNB 0.483229f
C43 B VNB 0.534382f
C44 VPB VNB 2.18693f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fa_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fa_4 VNB VPB VPWR CIN VGND B COUT SUM A
X0 VPWR.t9 a_1024_74.t4 SUM.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1 SUM.t7 a_1024_74.t5 VGND.t9 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19615 ps=1.41 w=0.74 l=0.15
X2 SUM.t2 a_1024_74.t6 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3 VPWR.t11 A.t0 a_27_392.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.253375 pd=1.725 as=0.295 ps=2.59 w=1 l=0.15
X4 a_737_347.t2 CIN.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X5 VGND.t1 a_418_74.t4 COUT.t7 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 COUT.t3 a_418_74.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7 a_418_74.t1 CIN.t1 a_27_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_27_392.t2 B.t0 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.49065 pd=2.05 as=0.253375 ps=1.725 w=1 l=0.15
X9 VPWR A a_1235_347# VPB sky130_fd_pr__pfet_01v8 ad=0.2152 pd=1.515 as=0.20235 ps=1.495 w=1 l=0.15
X10 a_734_74.t1 A.t1 VGND.t13 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19035 ps=1.37 w=0.74 l=0.15
X11 SUM.t6 a_1024_74.t7 VGND.t8 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19385 ps=1.41 w=0.74 l=0.15
X12 a_737_347.t3 A.t2 VPWR.t13 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.21 ps=1.42 w=1 l=0.15
X13 VGND.t7 a_1024_74.t8 SUM.t5 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.19615 pd=1.41 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VGND.t2 a_418_74.t6 COUT.t6 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VGND.t10 A.t3 a_27_74.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.39435 pd=1.87 as=0.2109 ps=2.05 w=0.74 l=0.15
X16 a_1238_74.t1 B.t1 a_1160_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X17 a_535_347.t1 B.t2 a_418_74.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.15 ps=1.3 w=1 l=0.15
X18 VPWR.t7 a_1024_74.t9 SUM.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_1160_74.t0 CIN.t2 a_1024_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1961 ps=1.27 w=0.74 l=0.15
X20 COUT.t5 a_418_74.t7 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19615 ps=1.41 w=0.74 l=0.15
X21 a_418_74.t2 CIN.t3 a_27_392.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.49065 ps=2.05 w=1 l=0.15
X22 VPWR.t10 A.t4 a_535_347.t0 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X23 SUM.t0 a_1024_74.t10 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2152 ps=1.515 w=1.12 l=0.15
X24 a_532_74.t1 B.t3 a_418_74.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1554 ps=1.16 w=0.74 l=0.15
X25 VGND.t11 A.t5 a_532_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1443 ps=1.13 w=0.74 l=0.15
X26 VPWR.t2 a_418_74.t8 COUT.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X27 VGND.t12 A.t6 a_1238_74.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.19385 pd=1.41 as=0.1332 ps=1.1 w=0.74 l=0.15
X28 COUT.t4 a_418_74.t9 VGND.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 VGND.t14 B.t4 a_734_74.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.19035 pd=1.37 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 a_1141_347.t0 CIN.t4 a_1024_74.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X31 COUT.t1 a_418_74.t10 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X32 VPWR.t0 B.t5 a_737_347.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.15 ps=1.3 w=1 l=0.15
X33 a_734_74.t0 CIN.t5 VGND.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1184 ps=1.06 w=0.74 l=0.15
X34 VPWR.t4 a_418_74.t11 COUT.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X35 VGND.t6 a_1024_74.t11 SUM.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.19615 pd=1.41 as=0.1036 ps=1.02 w=0.74 l=0.15
X36 a_27_74.t0 B.t6 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.39435 ps=1.87 w=0.74 l=0.15
X37 a_1024_74.t0 a_418_74.t12 a_734_74.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=1.27 as=0.1036 ps=1.02 w=0.74 l=0.15
X38 a_1024_74.t1 a_418_74.t13 a_737_347.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
R0 a_1024_74.n12 a_1024_74.n11 419.726
R1 a_1024_74.n11 a_1024_74.n1 303.829
R2 a_1024_74.n8 a_1024_74.t10 233.868
R3 a_1024_74.n3 a_1024_74.t4 229.487
R4 a_1024_74.n5 a_1024_74.t6 229.487
R5 a_1024_74.n0 a_1024_74.t9 229.487
R6 a_1024_74.n3 a_1024_74.t8 194.304
R7 a_1024_74.n8 a_1024_74.t7 179.947
R8 a_1024_74.n0 a_1024_74.t11 179.947
R9 a_1024_74.n4 a_1024_74.t5 179.947
R10 a_1024_74.n6 a_1024_74.n2 165.189
R11 a_1024_74.n10 a_1024_74.n9 152
R12 a_1024_74.n7 a_1024_74.n2 152
R13 a_1024_74.n1 a_1024_74.t0 63.2437
R14 a_1024_74.n4 a_1024_74.n3 51.1217
R15 a_1024_74.n9 a_1024_74.n7 49.6611
R16 a_1024_74.n0 a_1024_74.n6 43.0884
R17 a_1024_74.t1 a_1024_74.n12 39.4005
R18 a_1024_74.n12 a_1024_74.t3 29.5505
R19 a_1024_74.n6 a_1024_74.n5 28.4823
R20 a_1024_74.n1 a_1024_74.t2 22.7032
R21 a_1024_74.n5 a_1024_74.n4 14.6066
R22 a_1024_74.n10 a_1024_74.n2 13.1884
R23 a_1024_74.n11 a_1024_74.n10 10.4732
R24 a_1024_74.n9 a_1024_74.n8 6.57323
R25 a_1024_74.n7 a_1024_74.n0 6.57323
R26 SUM.n7 SUM.n6 585
R27 SUM.n6 SUM.n0 291.017
R28 SUM.n5 SUM.n1 253.302
R29 SUM.n4 SUM.n3 234.921
R30 SUM.n4 SUM.n2 187.304
R31 SUM.n5 SUM.n4 39.0308
R32 SUM.n6 SUM.t3 26.3844
R33 SUM.n6 SUM.t2 26.3844
R34 SUM.n1 SUM.t1 26.3844
R35 SUM.n1 SUM.t0 26.3844
R36 SUM.n3 SUM.t4 22.7032
R37 SUM.n3 SUM.t6 22.7032
R38 SUM.n2 SUM.t5 22.7032
R39 SUM.n2 SUM.t7 22.7032
R40 SUM SUM.n7 12.2187
R41 SUM SUM.n0 8.85027
R42 SUM.n0 SUM 5.40377
R43 SUM.n7 SUM 2.13383
R44 SUM SUM.n5 0.970197
R45 VPWR.n45 VPWR.n1 634.318
R46 VPWR.n32 VPWR.n7 608.681
R47 VPWR.n25 VPWR.t6 350.255
R48 VPWR.n37 VPWR.n4 325.221
R49 VPWR.n15 VPWR.n14 325.01
R50 VPWR.n11 VPWR.n10 324.764
R51 VPWR.n16 VPWR.t4 266.036
R52 VPWR.n19 VPWR.n13 232.787
R53 VPWR.n1 VPWR.t12 84.0359
R54 VPWR.n7 VPWR.t0 46.2955
R55 VPWR.n4 VPWR.t5 39.4005
R56 VPWR.n7 VPWR.t13 36.4455
R57 VPWR.n39 VPWR.n38 36.1417
R58 VPWR.n39 VPWR.n2 36.1417
R59 VPWR.n43 VPWR.n2 36.1417
R60 VPWR.n44 VPWR.n43 36.1417
R61 VPWR.n36 VPWR.n5 36.1417
R62 VPWR.n26 VPWR.n8 36.1417
R63 VPWR.n30 VPWR.n8 36.1417
R64 VPWR.n31 VPWR.n30 36.1417
R65 VPWR.n45 VPWR.n44 35.3887
R66 VPWR.n32 VPWR.n31 35.3887
R67 VPWR.n10 VPWR.t8 35.1791
R68 VPWR.n13 VPWR.t3 35.1791
R69 VPWR.n14 VPWR.t1 35.1791
R70 VPWR.n1 VPWR.t11 33.5313
R71 VPWR.n25 VPWR.n24 29.7417
R72 VPWR.n4 VPWR.t10 29.5505
R73 VPWR.n19 VPWR.n18 28.9887
R74 VPWR.n20 VPWR.n11 28.2358
R75 VPWR.n10 VPWR.t7 26.3844
R76 VPWR.n13 VPWR.t9 26.3844
R77 VPWR.n14 VPWR.t2 26.3844
R78 VPWR.n24 VPWR.n11 25.224
R79 VPWR.n20 VPWR.n19 24.4711
R80 VPWR.n26 VPWR.n25 23.7181
R81 VPWR.n18 VPWR.n15 23.7181
R82 VPWR.n18 VPWR.n17 9.3005
R83 VPWR.n19 VPWR.n12 9.3005
R84 VPWR.n21 VPWR.n20 9.3005
R85 VPWR.n22 VPWR.n11 9.3005
R86 VPWR.n24 VPWR.n23 9.3005
R87 VPWR.n25 VPWR.n9 9.3005
R88 VPWR.n27 VPWR.n26 9.3005
R89 VPWR.n28 VPWR.n8 9.3005
R90 VPWR.n30 VPWR.n29 9.3005
R91 VPWR.n31 VPWR.n6 9.3005
R92 VPWR.n33 VPWR.n32 9.3005
R93 VPWR.n34 VPWR.n5 9.3005
R94 VPWR.n36 VPWR.n35 9.3005
R95 VPWR.n38 VPWR.n3 9.3005
R96 VPWR.n40 VPWR.n39 9.3005
R97 VPWR.n41 VPWR.n2 9.3005
R98 VPWR.n43 VPWR.n42 9.3005
R99 VPWR.n44 VPWR.n0 9.3005
R100 VPWR.n46 VPWR.n45 8.45673
R101 VPWR.n37 VPWR.n36 7.52991
R102 VPWR.n16 VPWR.n15 6.99053
R103 VPWR.n32 VPWR.n5 6.77697
R104 VPWR.n38 VPWR.n37 3.76521
R105 VPWR.n17 VPWR.n16 0.569506
R106 VPWR VPWR.n46 0.163644
R107 VPWR.n46 VPWR.n0 0.144205
R108 VPWR.n17 VPWR.n12 0.122949
R109 VPWR.n21 VPWR.n12 0.122949
R110 VPWR.n22 VPWR.n21 0.122949
R111 VPWR.n23 VPWR.n22 0.122949
R112 VPWR.n23 VPWR.n9 0.122949
R113 VPWR.n27 VPWR.n9 0.122949
R114 VPWR.n28 VPWR.n27 0.122949
R115 VPWR.n29 VPWR.n28 0.122949
R116 VPWR.n29 VPWR.n6 0.122949
R117 VPWR.n33 VPWR.n6 0.122949
R118 VPWR.n34 VPWR.n33 0.122949
R119 VPWR.n35 VPWR.n34 0.122949
R120 VPWR.n35 VPWR.n3 0.122949
R121 VPWR.n40 VPWR.n3 0.122949
R122 VPWR.n41 VPWR.n40 0.122949
R123 VPWR.n42 VPWR.n41 0.122949
R124 VPWR.n42 VPWR.n0 0.122949
R125 VPB.n0 VPB 3381.18
R126 VPB.t16 VPB.t7 481.043
R127 VPB.t8 VPB.n0 478.627
R128 VPB VPB.n1 306.998
R129 VPB.n0 VPB.t10 288.575
R130 VPB.t0 VPB.t17 275.574
R131 VPB.t15 VPB 257.93
R132 VPB.t2 VPB.t1 255.376
R133 VPB.t13 VPB.t3 255.376
R134 VPB.t11 VPB.t12 255.376
R135 VPB.n1 VPB.t16 251.399
R136 VPB.t9 VPB.t14 246.565
R137 VPB.t5 VPB.t8 241.731
R138 VPB.t17 VPB.t5 241.731
R139 VPB.t14 VPB.t6 241.731
R140 VPB.t1 VPB.t4 229.839
R141 VPB.t3 VPB.t2 229.839
R142 VPB.t12 VPB.t13 229.839
R143 VPB.t10 VPB.t11 229.839
R144 VPB.t6 VPB.t0 217.558
R145 VPB.t7 VPB.t9 217.558
R146 VPB.n1 VPB.t15 66.3984
R147 VGND.n21 VGND.n20 220.173
R148 VGND.n18 VGND.n17 220.173
R149 VGND.n13 VGND.n12 218.024
R150 VGND.n29 VGND.n28 216.772
R151 VGND.n42 VGND.n41 206.333
R152 VGND.n6 VGND.n5 203.621
R153 VGND.n1 VGND.n0 196.02
R154 VGND.n14 VGND.t2 172.269
R155 VGND.n0 VGND.t0 100.541
R156 VGND.n0 VGND.t10 51.8924
R157 VGND.n28 VGND.t8 42.0185
R158 VGND.n30 VGND.n8 36.1417
R159 VGND.n34 VGND.n8 36.1417
R160 VGND.n35 VGND.n34 36.1417
R161 VGND.n36 VGND.n35 36.1417
R162 VGND.n40 VGND.n39 36.1417
R163 VGND.n43 VGND.n3 36.1417
R164 VGND.n47 VGND.n3 36.1417
R165 VGND.n48 VGND.n47 36.1417
R166 VGND.n49 VGND.n48 36.1417
R167 VGND.n5 VGND.t13 35.6762
R168 VGND.n5 VGND.t14 35.6762
R169 VGND.n20 VGND.t9 35.6762
R170 VGND.n20 VGND.t6 35.6762
R171 VGND.n17 VGND.t3 35.6762
R172 VGND.n17 VGND.t7 35.6762
R173 VGND.n22 VGND.n19 31.9397
R174 VGND.n27 VGND.n26 29.9622
R175 VGND.n41 VGND.t5 29.1897
R176 VGND.n26 VGND.n10 28.9735
R177 VGND.n16 VGND.n13 28.2358
R178 VGND.n22 VGND.n21 26.4789
R179 VGND.n30 VGND.n29 24.973
R180 VGND.n28 VGND.t12 24.0248
R181 VGND.n12 VGND.t4 22.7032
R182 VGND.n12 VGND.t1 22.7032
R183 VGND.n41 VGND.t11 22.7032
R184 VGND.n18 VGND.n16 21.9613
R185 VGND.n51 VGND.n1 11.9502
R186 VGND.n49 VGND.n1 10.2413
R187 VGND.n36 VGND.n6 9.91422
R188 VGND.n39 VGND.n6 9.91422
R189 VGND.n50 VGND.n49 9.3005
R190 VGND.n48 VGND.n2 9.3005
R191 VGND.n47 VGND.n46 9.3005
R192 VGND.n45 VGND.n3 9.3005
R193 VGND.n44 VGND.n43 9.3005
R194 VGND.n40 VGND.n4 9.3005
R195 VGND.n39 VGND.n38 9.3005
R196 VGND.n37 VGND.n36 9.3005
R197 VGND.n35 VGND.n7 9.3005
R198 VGND.n34 VGND.n33 9.3005
R199 VGND.n32 VGND.n8 9.3005
R200 VGND.n31 VGND.n30 9.3005
R201 VGND.n27 VGND.n9 9.3005
R202 VGND.n26 VGND.n25 9.3005
R203 VGND.n24 VGND.n10 9.3005
R204 VGND.n23 VGND.n22 9.3005
R205 VGND.n19 VGND.n11 9.3005
R206 VGND.n16 VGND.n15 9.3005
R207 VGND.n42 VGND.n40 7.15344
R208 VGND.n14 VGND.n13 6.70714
R209 VGND.n43 VGND.n42 4.14168
R210 VGND.n19 VGND.n18 2.06919
R211 VGND.n29 VGND.n27 1.03484
R212 VGND.n15 VGND.n14 0.645862
R213 VGND.n21 VGND.n10 0.517672
R214 VGND VGND.n51 0.161675
R215 VGND.n51 VGND.n50 0.146149
R216 VGND.n15 VGND.n11 0.122949
R217 VGND.n23 VGND.n11 0.122949
R218 VGND.n24 VGND.n23 0.122949
R219 VGND.n25 VGND.n24 0.122949
R220 VGND.n25 VGND.n9 0.122949
R221 VGND.n31 VGND.n9 0.122949
R222 VGND.n32 VGND.n31 0.122949
R223 VGND.n33 VGND.n32 0.122949
R224 VGND.n33 VGND.n7 0.122949
R225 VGND.n37 VGND.n7 0.122949
R226 VGND.n38 VGND.n37 0.122949
R227 VGND.n38 VGND.n4 0.122949
R228 VGND.n44 VGND.n4 0.122949
R229 VGND.n45 VGND.n44 0.122949
R230 VGND.n46 VGND.n45 0.122949
R231 VGND.n46 VGND.n2 0.122949
R232 VGND.n50 VGND.n2 0.122949
R233 VNB.t0 VNB.t7 2664.44
R234 VNB.t5 VNB.t2 1662.22
R235 VNB.t10 VNB.t12 1442.22
R236 VNB.t11 VNB.t4 1393.33
R237 VNB.t8 VNB.t11 1320
R238 VNB.n0 VNB.t6 1234.44
R239 VNB.t7 VNB 1210
R240 VNB.t3 VNB.t8 1148.89
R241 VNB.t2 VNB.t10 1051.11
R242 VNB.t12 VNB.t3 1051.11
R243 VNB.t4 VNB.t0 1051.11
R244 VNB.t6 VNB.t5 953.333
R245 VNB VNB.n0 625.163
R246 VNB.t9 VNB.t1 38.1784
R247 VNB.n0 VNB.t9 10.6225
R248 A.t0 A.n3 994.794
R249 A.n2 A.n1 835.735
R250 A.n1 A.t6 506.101
R251 A.t2 A.t1 454.954
R252 A.t4 A.t5 454.954
R253 A.n3 A.n2 430.587
R254 A.n2 A.t2 275.812
R255 A.n3 A.t4 275.812
R256 A.n4 A.t0 267.779
R257 A.n6 A.n5 181.942
R258 A.n4 A.n0 170.258
R259 A.n5 A.t3 162.274
R260 A.n6 A.n0 8.13508
R261 A A.n6 3.23041
R262 A.n5 A.n4 1.46111
R263 A.n0 A 0.120126
R264 a_27_392.n0 a_27_392.t1 708.056
R265 a_27_392.t0 a_27_392.n0 83.7255
R266 a_27_392.n0 a_27_392.t2 82.7405
R267 CIN.n3 CIN.t3 238.322
R268 CIN.n0 CIN.t4 238.322
R269 CIN.n1 CIN.t0 231.629
R270 CIN.n1 CIN.t5 186.374
R271 CIN.n2 CIN.n1 179.79
R272 CIN.n3 CIN.t1 178.34
R273 CIN.n0 CIN.t2 178.34
R274 CIN.n2 CIN.n0 167.321
R275 CIN.n4 CIN.n3 165.567
R276 CIN.n4 CIN.n2 0.756323
R277 CIN CIN.n4 0.0466957
R278 a_737_347.n1 a_737_347.n0 648.753
R279 a_737_347.n0 a_737_347.t3 39.4005
R280 a_737_347.n0 a_737_347.t1 29.5505
R281 a_737_347.t0 a_737_347.n1 29.5505
R282 a_737_347.n1 a_737_347.t2 29.5505
R283 a_418_74.n15 a_418_74.n14 826.011
R284 a_418_74.n12 a_418_74.n11 391.615
R285 a_418_74.n10 a_418_74.t10 245.797
R286 a_418_74.n0 a_418_74.t13 238.322
R287 a_418_74.n2 a_418_74.t11 234.841
R288 a_418_74.n4 a_418_74.t5 234.841
R289 a_418_74.n7 a_418_74.t8 234.841
R290 a_418_74.n2 a_418_74.t6 183.369
R291 a_418_74.n14 a_418_74.n12 181.505
R292 a_418_74.n0 a_418_74.t12 178.34
R293 a_418_74.n9 a_418_74.t7 173.52
R294 a_418_74.n6 a_418_74.t4 173.52
R295 a_418_74.n3 a_418_74.t9 173.52
R296 a_418_74.n12 a_418_74.n0 166.869
R297 a_418_74.n5 a_418_74.n1 165.189
R298 a_418_74.n11 a_418_74.n10 152
R299 a_418_74.n8 a_418_74.n1 152
R300 a_418_74.n14 a_418_74.n13 96.3134
R301 a_418_74.n3 a_418_74.n2 54.0429
R302 a_418_74.n9 a_418_74.n8 35.7853
R303 a_418_74.n13 a_418_74.t3 34.0546
R304 a_418_74.n13 a_418_74.t1 34.0546
R305 a_418_74.t0 a_418_74.n15 29.5505
R306 a_418_74.n15 a_418_74.t2 29.5505
R307 a_418_74.n5 a_418_74.n4 28.4823
R308 a_418_74.n6 a_418_74.n5 22.6399
R309 a_418_74.n7 a_418_74.n6 21.9096
R310 a_418_74.n10 a_418_74.n9 13.8763
R311 a_418_74.n11 a_418_74.n1 13.1884
R312 a_418_74.n4 a_418_74.n3 11.6853
R313 a_418_74.n8 a_418_74.n7 5.11262
R314 COUT.n7 COUT.n6 585
R315 COUT.n6 COUT.n0 290.969
R316 COUT.n5 COUT.n1 253.506
R317 COUT.n4 COUT.n2 147.721
R318 COUT.n4 COUT.n3 100.68
R319 COUT.n6 COUT.t0 26.3844
R320 COUT.n6 COUT.t3 26.3844
R321 COUT.n1 COUT.t2 26.3844
R322 COUT.n1 COUT.t1 26.3844
R323 COUT COUT.n4 25.2996
R324 COUT.n3 COUT.t6 22.7032
R325 COUT.n3 COUT.t4 22.7032
R326 COUT.n2 COUT.t7 22.7032
R327 COUT.n2 COUT.t5 22.7032
R328 COUT.n5 COUT 14.5783
R329 COUT COUT.n7 12.6123
R330 COUT COUT.n0 8.39965
R331 COUT.n0 COUT 5.43122
R332 COUT COUT.n5 1.69462
R333 COUT.n7 COUT 1.31815
R334 a_27_74.n0 a_27_74.t2 406.637
R335 a_27_74.n0 a_27_74.t1 22.7032
R336 a_27_74.t0 a_27_74.n0 22.7032
R337 B.n0 B.t0 259.38
R338 B.n2 B.n0 257.286
R339 B.n6 B.n5 231.629
R340 B.n1 B.t2 231.629
R341 B.n3 B.t5 231.629
R342 B.n6 B.t1 186.374
R343 B.n1 B.t3 186.374
R344 B.n3 B.t4 186.374
R345 B.n0 B.t6 173.228
R346 B.n2 B.n1 168.292
R347 B.n4 B.n3 168.292
R348 B.n7 B.n6 152
R349 B B.n4 138.406
R350 B.n4 B.n2 85.8358
R351 B.n7 B 8.32871
R352 B B.n7 6.73353
R353 a_734_74.n1 a_734_74.n0 432.514
R354 a_734_74.n0 a_734_74.t3 22.7032
R355 a_734_74.n0 a_734_74.t1 22.7032
R356 a_734_74.n1 a_734_74.t2 22.7032
R357 a_734_74.t0 a_734_74.n1 22.7032
R358 a_1160_74.t0 a_1160_74.t1 38.9194
R359 a_1238_74.t0 a_1238_74.t1 58.3789
R360 a_535_347.t0 a_535_347.t1 70.9205
R361 a_532_74.t0 a_532_74.t1 63.2437
C0 a_1235_347# VGND 0.001918f
C1 VPWR CIN 0.113535f
C2 a_1235_347# VPWR 0.012151f
C3 B CIN 0.590746f
C4 a_1235_347# B 0.003844f
C5 SUM COUT 0.003502f
C6 VPB SUM 0.01249f
C7 SUM VGND 0.025756f
C8 VPB COUT 0.012766f
C9 A SUM 0.001593f
C10 COUT VGND 0.233401f
C11 VPWR SUM 0.387019f
C12 A COUT 1.73e-19
C13 VPB VGND 0.014225f
C14 VPB A 0.665324f
C15 VPWR COUT 0.433771f
C16 B SUM 3.23e-19
C17 A VGND 0.043996f
C18 VPB VPWR 0.289443f
C19 B COUT 4.71e-20
C20 VPWR VGND 0.13659f
C21 CIN SUM 1.69e-19
C22 VPB B 0.171778f
C23 A VPWR 0.242469f
C24 a_1235_347# SUM 6.64e-19
C25 B VGND 0.031811f
C26 CIN COUT 4.59e-20
C27 VPB CIN 0.104143f
C28 A B 0.260282f
C29 CIN VGND 0.16227f
C30 VPWR B 0.096631f
C31 A CIN 0.114814f
C32 VGND VNB 1.28118f
C33 COUT VNB 0.034317f
C34 SUM VNB 0.0106f
C35 CIN VNB 0.301431f
C36 B VNB 0.411469f
C37 VPWR VNB 1.03388f
C38 A VNB 0.681688f
C39 VPB VNB 2.62435f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fah_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fah_1 VNB VPB VPWR VGND A CI SUM COUT B
X0 VPWR.t3 a_83_21.t4 SUM.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.28225 pd=1.65 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_1849_374.t2 B.t0 a_811_379.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.660675 pd=2.395 as=0.147 ps=1.19 w=0.84 l=0.15
X2 a_83_21.t2 a_811_379.t4 a_231_132.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.11875 pd=1.08 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 a_644_104.t2 a_1023_379.t3 a_83_21.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.11875 ps=1.08 w=0.64 l=0.15
X4 a_410_58.t3 a_811_379.t5 a_879_55# VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.131975 pd=1.205 as=0.28315 ps=3.17 w=0.64 l=0.15
X5 a_83_21.t3 a_811_379.t6 a_644_104.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3822 pd=1.75 as=0.27935 ps=1.635 w=0.84 l=0.15
X6 a_811_379.t2 a_879_55# a_1660_374.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X7 a_1660_374.t3 B.t1 a_811_379.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.3264 ps=1.66 w=0.64 l=0.15
X8 VGND.t7 A.t0 a_1849_374.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1216 pd=1.02 as=0.208 ps=1.93 w=0.64 l=0.15
X9 VPWR B a_879_55# VPB sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.2018 ps=1.505 w=1.12 l=0.15
X10 VPWR.t1 a_2342_48.t2 a_1660_374.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.31 as=0.1862 ps=1.475 w=1.12 l=0.15
X11 a_2342_48.t1 A.t1 VPWR.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X12 a_2342_48.t0 A.t2 VGND.t6 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1216 ps=1.02 w=0.64 l=0.15
X13 VGND.t4 B.t2 a_879_55# VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.3136 pd=2.51 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 a_644_104.t1 a_231_132.t6 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.23505 pd=2.02 as=0.29265 ps=1.61 w=0.64 l=0.15
X15 a_879_55# a_1023_379.t4 a_410_58.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2018 pd=1.505 as=0.2541 ps=1.445 w=0.84 l=0.15
X16 a_231_132.t2 CI.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.28225 ps=1.65 w=1 l=0.15
X17 VGND.t5 a_410_58.t4 COUT.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.29265 pd=1.61 as=0.2072 ps=2.04 w=0.74 l=0.15
X18 a_1849_374.t1 B.t3 a_1023_379.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1524 pd=1.16 as=0.24825 ps=1.49 w=0.64 l=0.15
X19 a_1660_374.t2 B.t4 a_1023_379.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.126 ps=1.14 w=0.84 l=0.15
X20 VPWR.t5 a_410_58.t5 COUT.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.30565 pd=1.85 as=0.46765 ps=3.29 w=1.12 l=0.15
X21 VGND.t0 a_2342_48.t3 a_1660_374.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2875 pd=2.33 as=0.12945 ps=1.1 w=0.74 l=0.15
X22 VGND.t2 a_83_21.t5 SUM.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1924 pd=1.41 as=0.2072 ps=2.04 w=0.74 l=0.15
X23 VPWR.t4 A.t3 a_1849_374.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X24 a_231_132.t0 a_1023_379.t5 a_410_58.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.131975 ps=1.205 w=0.64 l=0.15
X25 a_644_104.t0 a_231_132.t7 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.27935 pd=1.635 as=0.30565 ps=1.85 w=1 l=0.15
X26 a_231_132.t1 a_1023_379.t6 a_83_21.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.4066 pd=2.01 as=0.3822 ps=1.75 w=0.84 l=0.15
X27 a_231_132.t5 CI.t1 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2016 pd=1.91 as=0.1924 ps=1.41 w=0.64 l=0.15
X28 a_1023_379.t2 a_879_55# a_1660_374.t4 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.24825 pd=1.49 as=0.2568 ps=2.17 w=0.64 l=0.15
X29 a_811_379.t3 a_879_55# a_1849_374.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.3264 pd=1.66 as=0.1524 ps=1.16 w=0.64 l=0.15
X30 a_410_58.t2 a_811_379.t7 a_231_132.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2541 pd=1.445 as=0.4066 ps=2.01 w=0.84 l=0.15
R0 a_83_21.n1 a_83_21.t5 1117.31
R1 a_83_21.n1 a_83_21.n0 566.254
R2 a_83_21.n2 a_83_21.n1 454.404
R3 a_83_21.t5 a_83_21.t4 451.474
R4 a_83_21.t0 a_83_21.n2 178.238
R5 a_83_21.n0 a_83_21.t2 40.416
R6 a_83_21.n2 a_83_21.t3 35.1791
R7 a_83_21.n0 a_83_21.t1 25.1433
R8 SUM.n1 SUM 589.777
R9 SUM.n1 SUM.n0 585
R10 SUM.n2 SUM.n1 585
R11 SUM SUM.t1 146.988
R12 SUM.n1 SUM.t0 26.3844
R13 SUM SUM.n2 12.8005
R14 SUM SUM.n0 11.0811
R15 SUM SUM.n0 3.05722
R16 SUM.n2 SUM 1.33781
R17 VPWR.n45 VPWR.n44 677.768
R18 VPWR.n52 VPWR.n1 331.58
R19 VPWR.n14 VPWR.t1 258.358
R20 VPWR.n15 VPWR.n13 236.706
R21 VPWR.n1 VPWR.t0 74.7789
R22 VPWR.n44 VPWR.t2 58.1155
R23 VPWR.n13 VPWR.t6 39.4005
R24 VPWR.n46 VPWR.n2 36.1417
R25 VPWR.n50 VPWR.n2 36.1417
R26 VPWR.n51 VPWR.n50 36.1417
R27 VPWR.n31 VPWR.n30 36.1417
R28 VPWR.n32 VPWR.n31 36.1417
R29 VPWR.n32 VPWR.n6 36.1417
R30 VPWR.n36 VPWR.n6 36.1417
R31 VPWR.n37 VPWR.n36 36.1417
R32 VPWR.n38 VPWR.n37 36.1417
R33 VPWR.n38 VPWR.n4 36.1417
R34 VPWR.n42 VPWR.n4 36.1417
R35 VPWR.n18 VPWR.n12 36.1417
R36 VPWR.n19 VPWR.n18 36.1417
R37 VPWR.n20 VPWR.n19 36.1417
R38 VPWR.n20 VPWR.n10 36.1417
R39 VPWR.n24 VPWR.n10 36.1417
R40 VPWR.n25 VPWR.n24 36.1417
R41 VPWR.n26 VPWR.n25 36.1417
R42 VPWR.n52 VPWR.n51 35.3887
R43 VPWR.n44 VPWR.t5 32.577
R44 VPWR.n26 VPWR.n8 30.1181
R45 VPWR.n13 VPWR.t4 29.5505
R46 VPWR.n43 VPWR.n42 28.1772
R47 VPWR.n46 VPWR.n45 27.19
R48 VPWR.n1 VPWR.t3 25.5754
R49 VPWR.n30 VPWR.n8 17.3181
R50 VPWR.n14 VPWR.n12 14.3064
R51 VPWR.n16 VPWR.n12 9.3005
R52 VPWR.n18 VPWR.n17 9.3005
R53 VPWR.n19 VPWR.n11 9.3005
R54 VPWR.n21 VPWR.n20 9.3005
R55 VPWR.n22 VPWR.n10 9.3005
R56 VPWR.n24 VPWR.n23 9.3005
R57 VPWR.n25 VPWR.n9 9.3005
R58 VPWR.n27 VPWR.n26 9.3005
R59 VPWR.n28 VPWR.n8 9.3005
R60 VPWR.n30 VPWR.n29 9.3005
R61 VPWR.n31 VPWR.n7 9.3005
R62 VPWR.n33 VPWR.n32 9.3005
R63 VPWR.n34 VPWR.n6 9.3005
R64 VPWR.n36 VPWR.n35 9.3005
R65 VPWR.n37 VPWR.n5 9.3005
R66 VPWR.n39 VPWR.n38 9.3005
R67 VPWR.n40 VPWR.n4 9.3005
R68 VPWR.n42 VPWR.n41 9.3005
R69 VPWR.n43 VPWR.n3 9.3005
R70 VPWR.n47 VPWR.n46 9.3005
R71 VPWR.n48 VPWR.n2 9.3005
R72 VPWR.n50 VPWR.n49 9.3005
R73 VPWR.n51 VPWR.n0 9.3005
R74 VPWR.n53 VPWR.n52 8.45673
R75 VPWR.n15 VPWR.n14 7.19259
R76 VPWR.n16 VPWR.n15 0.467758
R77 VPWR.n45 VPWR.n43 0.284944
R78 VPWR VPWR.n53 0.163644
R79 VPWR.n53 VPWR.n0 0.144205
R80 VPWR.n17 VPWR.n16 0.122949
R81 VPWR.n17 VPWR.n11 0.122949
R82 VPWR.n21 VPWR.n11 0.122949
R83 VPWR.n22 VPWR.n21 0.122949
R84 VPWR.n23 VPWR.n22 0.122949
R85 VPWR.n23 VPWR.n9 0.122949
R86 VPWR.n27 VPWR.n9 0.122949
R87 VPWR.n28 VPWR.n27 0.122949
R88 VPWR.n29 VPWR.n28 0.122949
R89 VPWR.n29 VPWR.n7 0.122949
R90 VPWR.n33 VPWR.n7 0.122949
R91 VPWR.n34 VPWR.n33 0.122949
R92 VPWR.n35 VPWR.n34 0.122949
R93 VPWR.n35 VPWR.n5 0.122949
R94 VPWR.n39 VPWR.n5 0.122949
R95 VPWR.n40 VPWR.n39 0.122949
R96 VPWR.n41 VPWR.n40 0.122949
R97 VPWR.n41 VPWR.n3 0.122949
R98 VPWR.n47 VPWR.n3 0.122949
R99 VPWR.n48 VPWR.n47 0.122949
R100 VPWR.n49 VPWR.n48 0.122949
R101 VPWR.n49 VPWR.n0 0.122949
R102 VPB.n0 VPB 6358.87
R103 VPB.n1 VPB 4528.02
R104 VPB.n2 VPB 2740.86
R105 VPB VPB.t5 2492.25
R106 VPB.n1 VPB.t8 864.071
R107 VPB.t12 VPB.t2 819.759
R108 VPB.t0 VPB.t11 816.058
R109 VPB.t5 VPB.t1 630.841
R110 VPB.t6 VPB.t0 374.543
R111 VPB.n2 VPB.t6 369.582
R112 VPB.t5 VPB.t4 362.635
R113 VPB.t2 VPB.t9 347.312
R114 VPB.t4 VPB.t12 329.435
R115 VPB.t3 VPB.n0 310.303
R116 VPB.t9 VPB 257.93
R117 VPB.t10 VPB.t13 255.376
R118 VPB.t11 VPB.t7 248.042
R119 VPB.t8 VPB.t3 241.081
R120 VPB.n0 VPB.t10 234.946
R121 VPB.t1 VPB.n2 192.405
R122 VPB.t7 VPB.n1 156.267
R123 B.n2 B.n1 909.374
R124 B.n2 B.t4 890.093
R125 B.t4 B.t1 449.05
R126 B.n1 B.t2 263.493
R127 B.t0 B.n2 256.8
R128 B.n3 B.t0 245.114
R129 B.n1 B.n0 221.72
R130 B.n3 B.t3 168.117
R131 B B.n3 158.788
R132 a_811_379.t4 a_811_379.t5 811.367
R133 a_811_379.t5 a_811_379.t6 568.76
R134 a_811_379.n2 a_811_379.n0 442.517
R135 a_811_379.n3 a_811_379.n2 287.779
R136 a_811_379.n1 a_811_379.t7 287.447
R137 a_811_379.n2 a_811_379.n1 213.18
R138 a_811_379.n1 a_811_379.t4 162.274
R139 a_811_379.n0 a_811_379.t0 103.126
R140 a_811_379.n0 a_811_379.t3 88.1255
R141 a_811_379.n3 a_811_379.t2 46.9053
R142 a_811_379.t1 a_811_379.n3 35.1791
R143 a_1849_374.n2 a_1849_374.t0 254.96
R144 a_1849_374.t3 a_1849_374.n2 234.393
R145 a_1849_374.n1 a_1849_374.n0 216.428
R146 a_1849_374.n1 a_1849_374.t2 192.227
R147 a_1849_374.n0 a_1849_374.t4 41.2505
R148 a_1849_374.n0 a_1849_374.t1 41.2505
R149 a_1849_374.n2 a_1849_374.n1 18.7367
R150 a_231_132.t2 a_231_132.n6 775.322
R151 a_231_132.t2 a_231_132.n5 698.525
R152 a_231_132.n3 a_231_132.n1 473.649
R153 a_231_132.n6 a_231_132.t5 332.243
R154 a_231_132.n3 a_231_132.n2 313.933
R155 a_231_132.n4 a_231_132.n0 245.547
R156 a_231_132.n5 a_231_132.n4 236.976
R157 a_231_132.n0 a_231_132.t7 218.239
R158 a_231_132.n0 a_231_132.t6 202.548
R159 a_231_132.n2 a_231_132.t4 157.768
R160 a_231_132.n4 a_231_132.n3 33.4153
R161 a_231_132.n2 a_231_132.t1 30.6533
R162 a_231_132.n1 a_231_132.t3 26.2505
R163 a_231_132.n1 a_231_132.t0 26.2505
R164 a_231_132.n6 a_231_132.n5 16.6405
R165 VNB.n0 VNB 23512.1
R166 VNB VNB.n1 13140.5
R167 VNB.t6 VNB.t3 3891.86
R168 VNB.t4 VNB.t10 3210.81
R169 VNB.t12 VNB.t11 2900.28
R170 VNB.t1 VNB.t2 2751.55
R171 VNB.t10 VNB.t13 2735.14
R172 VNB.t14 VNB.t8 2413.65
R173 VNB.t3 VNB.t14 2355.91
R174 VNB.t13 VNB.n0 1712.43
R175 VNB.t9 VNB.t12 1462.54
R176 VNB.t8 VNB.t5 1362.73
R177 VNB.t2 VNB.t15 1313.8
R178 VNB.t11 VNB.t1 1264.23
R179 VNB.t7 VNB.t4 1189.19
R180 VNB.t0 VNB.t6 1166.4
R181 VNB.t5 VNB 1131.76
R182 VNB.n1 VNB.t7 570.812
R183 VNB.n1 VNB.t0 438.846
R184 VNB.n0 VNB.t9 36.4143
R185 a_1023_379.t4 a_1023_379.t6 974.98
R186 a_1023_379.t6 a_1023_379.t5 488.836
R187 a_1023_379.n2 a_1023_379.n0 447.06
R188 a_1023_379.t0 a_1023_379.n2 418.736
R189 a_1023_379.n1 a_1023_379.t3 334.188
R190 a_1023_379.n1 a_1023_379.t4 300.447
R191 a_1023_379.n2 a_1023_379.n1 138.237
R192 a_1023_379.n0 a_1023_379.t1 56.2505
R193 a_1023_379.n0 a_1023_379.t2 56.2505
R194 a_644_104.n1 a_644_104.n0 646.797
R195 a_644_104.n0 a_644_104.t2 290.933
R196 a_644_104.n0 a_644_104.t1 264.865
R197 a_644_104.n1 a_644_104.t3 79.5435
R198 a_644_104.t0 a_644_104.n1 39.174
R199 a_410_58.n3 a_410_58.n2 752.073
R200 a_410_58.n2 a_410_58.n0 378.712
R201 a_410_58.n0 a_410_58.t4 299.132
R202 a_410_58.n0 a_410_58.t5 254.571
R203 a_410_58.n2 a_410_58.n1 185
R204 a_410_58.t1 a_410_58.n3 106.709
R205 a_410_58.n1 a_410_58.t0 48.5543
R206 a_410_58.n3 a_410_58.t2 35.1791
R207 a_410_58.n1 a_410_58.t3 26.2505
R208 a_1660_374.n1 a_1660_374.t5 375.505
R209 a_1660_374.n1 a_1660_374.t4 342.481
R210 a_1660_374.n3 a_1660_374.n2 287.495
R211 a_1660_374.n2 a_1660_374.n1 254.59
R212 a_1660_374.n2 a_1660_374.n0 144.109
R213 a_1660_374.n0 a_1660_374.t3 41.0701
R214 a_1660_374.n3 a_1660_374.t2 41.0422
R215 a_1660_374.t1 a_1660_374.n3 38.0348
R216 a_1660_374.n0 a_1660_374.t0 21.1849
R217 A.n1 A.t0 252.832
R218 A.n0 A.t2 252.832
R219 A.n0 A.t1 207.529
R220 A.n1 A.t3 207.529
R221 A A.n2 68.5569
R222 A.n2 A.n0 34.0952
R223 A.n2 A.n1 32.2145
R224 VGND.n7 VGND.t4 322.87
R225 VGND.n52 VGND.n51 271.474
R226 VGND.n12 VGND.t0 238.325
R227 VGND.n44 VGND.n43 221.142
R228 VGND.n43 VGND.t1 136.875
R229 VGND.n14 VGND.n13 121.409
R230 VGND.n51 VGND.t3 48.7505
R231 VGND.n13 VGND.t6 39.3755
R232 VGND.n17 VGND.n11 36.1417
R233 VGND.n18 VGND.n17 36.1417
R234 VGND.n19 VGND.n18 36.1417
R235 VGND.n19 VGND.n9 36.1417
R236 VGND.n23 VGND.n9 36.1417
R237 VGND.n24 VGND.n23 36.1417
R238 VGND.n25 VGND.n24 36.1417
R239 VGND.n30 VGND.n29 36.1417
R240 VGND.n31 VGND.n30 36.1417
R241 VGND.n31 VGND.n5 36.1417
R242 VGND.n35 VGND.n5 36.1417
R243 VGND.n36 VGND.n35 36.1417
R244 VGND.n37 VGND.n36 36.1417
R245 VGND.n37 VGND.n3 36.1417
R246 VGND.n41 VGND.n3 36.1417
R247 VGND.n42 VGND.n41 36.1417
R248 VGND.n45 VGND.n42 36.1417
R249 VGND.n49 VGND.n1 36.1417
R250 VGND.n50 VGND.n49 36.1417
R251 VGND.n13 VGND.t7 31.8755
R252 VGND.n25 VGND.n7 24.4711
R253 VGND.n51 VGND.t2 24.4533
R254 VGND.n29 VGND.n7 22.9652
R255 VGND.n45 VGND.n44 22.5887
R256 VGND.n43 VGND.t5 21.3263
R257 VGND.n52 VGND.n50 18.824
R258 VGND.n44 VGND.n1 13.5534
R259 VGND.n12 VGND.n11 11.6711
R260 VGND.n50 VGND.n0 9.3005
R261 VGND.n49 VGND.n48 9.3005
R262 VGND.n47 VGND.n1 9.3005
R263 VGND.n46 VGND.n45 9.3005
R264 VGND.n42 VGND.n2 9.3005
R265 VGND.n41 VGND.n40 9.3005
R266 VGND.n39 VGND.n3 9.3005
R267 VGND.n38 VGND.n37 9.3005
R268 VGND.n36 VGND.n4 9.3005
R269 VGND.n35 VGND.n34 9.3005
R270 VGND.n33 VGND.n5 9.3005
R271 VGND.n32 VGND.n31 9.3005
R272 VGND.n30 VGND.n6 9.3005
R273 VGND.n29 VGND.n28 9.3005
R274 VGND.n27 VGND.n7 9.3005
R275 VGND.n26 VGND.n25 9.3005
R276 VGND.n24 VGND.n8 9.3005
R277 VGND.n23 VGND.n22 9.3005
R278 VGND.n21 VGND.n9 9.3005
R279 VGND.n20 VGND.n19 9.3005
R280 VGND.n18 VGND.n10 9.3005
R281 VGND.n17 VGND.n16 9.3005
R282 VGND.n15 VGND.n11 9.3005
R283 VGND.n53 VGND.n52 7.44972
R284 VGND.n14 VGND.n12 7.26981
R285 VGND.n15 VGND.n14 0.49428
R286 VGND VGND.n53 0.160299
R287 VGND.n53 VGND.n0 0.147507
R288 VGND.n16 VGND.n15 0.122949
R289 VGND.n16 VGND.n10 0.122949
R290 VGND.n20 VGND.n10 0.122949
R291 VGND.n21 VGND.n20 0.122949
R292 VGND.n22 VGND.n21 0.122949
R293 VGND.n22 VGND.n8 0.122949
R294 VGND.n26 VGND.n8 0.122949
R295 VGND.n27 VGND.n26 0.122949
R296 VGND.n28 VGND.n27 0.122949
R297 VGND.n28 VGND.n6 0.122949
R298 VGND.n32 VGND.n6 0.122949
R299 VGND.n33 VGND.n32 0.122949
R300 VGND.n34 VGND.n33 0.122949
R301 VGND.n34 VGND.n4 0.122949
R302 VGND.n38 VGND.n4 0.122949
R303 VGND.n39 VGND.n38 0.122949
R304 VGND.n40 VGND.n39 0.122949
R305 VGND.n40 VGND.n2 0.122949
R306 VGND.n46 VGND.n2 0.122949
R307 VGND.n47 VGND.n46 0.122949
R308 VGND.n48 VGND.n47 0.122949
R309 VGND.n48 VGND.n0 0.122949
R310 a_2342_48.n1 a_2342_48.n0 315.81
R311 a_2342_48.t1 a_2342_48.n1 290.519
R312 a_2342_48.n0 a_2342_48.t2 261.62
R313 a_2342_48.n0 a_2342_48.t3 156.431
R314 a_2342_48.n1 a_2342_48.t0 145.043
R315 CI.n0 CI.t0 231.629
R316 CI.n0 CI.t1 162.274
R317 CI CI.n0 153.904
R318 COUT COUT.t1 1205.32
R319 COUT COUT.t0 293.647
C0 VPWR a_879_55# 0.144353f
C1 A VPB 0.095587f
C2 CI VGND 0.004883f
C3 B VGND 0.022609f
C4 a_879_55# VPB 0.124621f
C5 B A 4.45e-19
C6 VGND A 0.037797f
C7 B a_879_55# 0.295285f
C8 VPWR COUT 0.296356f
C9 VPWR VPB 0.288227f
C10 VGND a_879_55# 0.473096f
C11 VPWR SUM 0.093807f
C12 COUT VPB 0.024669f
C13 A a_879_55# 3.93e-20
C14 VPWR CI 0.005662f
C15 COUT SUM 0.108446f
C16 SUM VPB 0.012746f
C17 COUT CI 0.088625f
C18 VPWR B 0.13705f
C19 CI VPB 0.045353f
C20 SUM CI 0.001369f
C21 COUT B 1e-20
C22 VPWR VGND 0.076148f
C23 B VPB 0.577107f
C24 VPWR A 0.07081f
C25 SUM B 1.59e-20
C26 COUT VGND 0.152105f
C27 VGND VPB 0.010769f
C28 SUM VGND 0.031501f
C29 A VNB 0.255571f
C30 VGND VNB 1.55565f
C31 B VNB 0.477834f
C32 CI VNB 0.091932f
C33 SUM VNB 0.100548f
C34 COUT VNB 0.019941f
C35 VPWR VNB 1.21655f
C36 VPB VNB 3.21845f
C37 a_879_55# VNB 0.330235f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fah_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fah_2 VNB VPB VPWR VGND A CI SUM COUT B
X0 VGND.t6 A.t0 a_81_260.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2272 ps=1.99 w=0.64 l=0.15
X1 SUM.t1 a_1895_424# VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_2052_424.t2 a_514_424.t4 a_1895_424# VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.23645 ps=1.45 w=0.64 l=0.15
X3 VPWR.t6 a_1451_424# COUT.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_849_424.t1 a_481_379.t2 a_114_368.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.5649 pd=2.185 as=0.1932 ps=1.3 w=0.84 l=0.15
X5 a_1689_424.t3 a_514_424.t5 a_1451_424# VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2176 pd=1.32 as=0.28 ps=1.515 w=0.64 l=0.15
X6 a_413_392.t0 B.t0 a_849_424.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.2394 pd=2.25 as=0.5649 ps=2.185 w=0.84 l=0.15
X7 a_1689_424.t2 CI.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0.2957 ps=1.73 w=1 l=0.15
X8 COUT.t0 a_1451_424# VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.303 ps=2.81 w=1.12 l=0.15
X9 SUM.t3 a_1895_424# VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 VPWR.t9 A.t1 a_81_260.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.285 ps=2.57 w=1 l=0.15
X11 a_481_379.t1 B.t1 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.31405 ps=2.87 w=0.74 l=0.15
X12 a_413_392.t4 A.t2 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1703 pd=1.355 as=0.18 ps=1.36 w=1 l=0.15
X13 COUT.t2 a_1451_424# VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2739 ps=2.27 w=0.74 l=0.15
X14 a_413_392.t5 A.t3 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 a_114_368.t2 a_481_379.t3 a_514_424.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.272 pd=1.49 as=0.1952 ps=1.25 w=0.64 l=0.15
X16 a_114_368.t5 B.t2 a_514_424.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.3 as=0.3843 ps=1.755 w=0.84 l=0.15
X17 a_114_368.t4 a_81_260.t2 VGND.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.222 ps=2.08 w=0.74 l=0.15
X18 VPWR.t1 a_1895_424# SUM.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.1736 ps=1.43 w=1.12 l=0.15
X19 VGND a_1451_424# COUT VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_514_424.t0 B.t3 a_413_392.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1952 pd=1.25 as=0.0896 ps=0.92 w=0.64 l=0.15
X21 VPWR.t0 a_1689_424.t4 a_2052_424.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2957 pd=1.73 as=0.2459 ps=1.535 w=1 l=0.15
X22 a_481_379.t0 B.t4 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1974 pd=1.495 as=0.3192 ps=2.81 w=1.12 l=0.15
X23 a_114_368.t3 a_81_260.t3 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.3192 ps=2.81 w=1.12 l=0.15
X24 a_514_424.t2 a_481_379.t4 a_413_392.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3843 pd=1.755 as=0.1703 ps=1.355 w=0.84 l=0.15
X25 a_849_424.t0 B.t5 a_114_368.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2224 pd=1.335 as=0.272 ps=1.49 w=0.64 l=0.15
X26 a_1895_424# a_849_424.t4 a_1689_424.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.23645 pd=1.45 as=0.2176 ps=1.32 w=0.64 l=0.15
X27 a_413_392.t2 a_481_379.t5 a_849_424.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2455 pd=2.38 as=0.2224 ps=1.335 w=0.64 l=0.15
X28 a_1689_424.t1 a_849_424.t5 a_1451_424# VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3696 pd=1.72 as=0.4368 ps=1.88 w=0.84 l=0.15
X29 VGND.t1 a_1895_424# SUM.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1073 ps=1.03 w=0.74 l=0.15
X30 VGND.t0 a_1689_424.t5 a_2052_424.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1826 pd=1.32 as=0.1344 ps=1.06 w=0.64 l=0.15
X31 a_2052_424.t3 a_849_424.t6 a_1895_424# VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.2459 pd=1.535 as=0.2667 ps=1.475 w=0.84 l=0.15
R0 A.n1 A.t1 306.12
R1 A.n0 A.t2 255.728
R2 A.n0 A.t3 181.7
R3 A A.n2 160.359
R4 A.n1 A.t0 142.994
R5 A.n2 A.n1 13.146
R6 A.n2 A.n0 10.955
R7 a_81_260.t1 a_81_260.n1 262.358
R8 a_81_260.n0 a_81_260.t3 253.343
R9 a_81_260.n1 a_81_260.n0 210.424
R10 a_81_260.n0 a_81_260.t2 179.947
R11 a_81_260.n1 a_81_260.t0 154.114
R12 VGND.n35 VGND.t7 401.108
R13 VGND.n11 VGND.t0 305.168
R14 VGND.n14 VGND.t1 300.62
R15 VGND.n17 VGND.t3 239.101
R16 VGND.n56 VGND.t4 230.849
R17 VGND.n49 VGND.n48 219.56
R18 VGND.n13 VGND.t2 155.272
R19 VGND.n23 VGND.n22 36.1417
R20 VGND.n24 VGND.n23 36.1417
R21 VGND.n24 VGND.n9 36.1417
R22 VGND.n28 VGND.n9 36.1417
R23 VGND.n29 VGND.n28 36.1417
R24 VGND.n30 VGND.n29 36.1417
R25 VGND.n30 VGND.n7 36.1417
R26 VGND.n34 VGND.n7 36.1417
R27 VGND.n36 VGND.n5 36.1417
R28 VGND.n40 VGND.n5 36.1417
R29 VGND.n41 VGND.n40 36.1417
R30 VGND.n42 VGND.n41 36.1417
R31 VGND.n42 VGND.n3 36.1417
R32 VGND.n46 VGND.n3 36.1417
R33 VGND.n47 VGND.n46 36.1417
R34 VGND.n50 VGND.n47 36.1417
R35 VGND.n54 VGND.n1 36.1417
R36 VGND.n55 VGND.n54 36.1417
R37 VGND.n18 VGND.n11 30.4946
R38 VGND.n48 VGND.t5 26.2505
R39 VGND.n48 VGND.t6 26.2505
R40 VGND.n36 VGND.n35 25.224
R41 VGND.n17 VGND.n16 23.7181
R42 VGND.n18 VGND.n17 23.7181
R43 VGND.n22 VGND.n11 22.9652
R44 VGND.n16 VGND.n13 22.2123
R45 VGND.n35 VGND.n34 22.2123
R46 VGND.n49 VGND.n1 14.6829
R47 VGND.n56 VGND.n55 13.9299
R48 VGND.n57 VGND.n56 9.3005
R49 VGND.n55 VGND.n0 9.3005
R50 VGND.n54 VGND.n53 9.3005
R51 VGND.n52 VGND.n1 9.3005
R52 VGND.n51 VGND.n50 9.3005
R53 VGND.n47 VGND.n2 9.3005
R54 VGND.n46 VGND.n45 9.3005
R55 VGND.n44 VGND.n3 9.3005
R56 VGND.n43 VGND.n42 9.3005
R57 VGND.n41 VGND.n4 9.3005
R58 VGND.n40 VGND.n39 9.3005
R59 VGND.n38 VGND.n5 9.3005
R60 VGND.n37 VGND.n36 9.3005
R61 VGND.n35 VGND.n6 9.3005
R62 VGND.n34 VGND.n33 9.3005
R63 VGND.n32 VGND.n7 9.3005
R64 VGND.n31 VGND.n30 9.3005
R65 VGND.n29 VGND.n8 9.3005
R66 VGND.n28 VGND.n27 9.3005
R67 VGND.n26 VGND.n9 9.3005
R68 VGND.n25 VGND.n24 9.3005
R69 VGND.n23 VGND.n10 9.3005
R70 VGND.n22 VGND.n21 9.3005
R71 VGND.n20 VGND.n11 9.3005
R72 VGND.n19 VGND.n18 9.3005
R73 VGND.n17 VGND.n12 9.3005
R74 VGND.n16 VGND.n15 9.3005
R75 VGND.n14 VGND.n13 6.70714
R76 VGND.n50 VGND.n49 2.63579
R77 VGND.n15 VGND.n14 0.645862
R78 VGND.n15 VGND.n12 0.122949
R79 VGND.n19 VGND.n12 0.122949
R80 VGND.n20 VGND.n19 0.122949
R81 VGND.n21 VGND.n20 0.122949
R82 VGND.n21 VGND.n10 0.122949
R83 VGND.n25 VGND.n10 0.122949
R84 VGND.n26 VGND.n25 0.122949
R85 VGND.n27 VGND.n26 0.122949
R86 VGND.n27 VGND.n8 0.122949
R87 VGND.n31 VGND.n8 0.122949
R88 VGND.n32 VGND.n31 0.122949
R89 VGND.n33 VGND.n32 0.122949
R90 VGND.n33 VGND.n6 0.122949
R91 VGND.n37 VGND.n6 0.122949
R92 VGND.n38 VGND.n37 0.122949
R93 VGND.n39 VGND.n38 0.122949
R94 VGND.n39 VGND.n4 0.122949
R95 VGND.n43 VGND.n4 0.122949
R96 VGND.n44 VGND.n43 0.122949
R97 VGND.n45 VGND.n44 0.122949
R98 VGND.n45 VGND.n2 0.122949
R99 VGND.n51 VGND.n2 0.122949
R100 VGND.n52 VGND.n51 0.122949
R101 VGND.n53 VGND.n52 0.122949
R102 VGND.n53 VGND.n0 0.122949
R103 VGND.n57 VGND.n0 0.122949
R104 VGND VGND.n57 0.0617245
R105 VNB.t8 VNB.t13 4238.32
R106 VNB.t1 VNB.t9 3880.31
R107 VNB.t13 VNB.t5 3464.57
R108 VNB.t10 VNB.t12 2864.04
R109 VNB.t7 VNB.t0 2309.71
R110 VNB.t9 VNB.t3 2148.03
R111 VNB.t0 VNB.t8 1951.71
R112 VNB.t14 VNB.t4 1917.06
R113 VNB.t5 VNB.t14 1917.06
R114 VNB.t6 VNB.t7 1755.38
R115 VNB VNB.t10 1351.18
R116 VNB.t4 VNB.t1 1316.54
R117 VNB.t3 VNB.t2 1016.27
R118 VNB.t11 VNB.t6 993.177
R119 VNB.t12 VNB.t11 993.177
R120 VPWR.n39 VPWR.t4 846.165
R121 VPWR.n21 VPWR.t5 802.049
R122 VPWR.n13 VPWR.n12 622.663
R123 VPWR.n17 VPWR.n16 605.365
R124 VPWR.n58 VPWR.t7 350.757
R125 VPWR.n18 VPWR.t1 268.866
R126 VPWR.n2 VPWR.n1 222.361
R127 VPWR.n12 VPWR.t3 51.2205
R128 VPWR.n12 VPWR.t0 51.2205
R129 VPWR.n1 VPWR.t8 41.3705
R130 VPWR.n57 VPWR.n56 36.1417
R131 VPWR.n40 VPWR.n6 36.1417
R132 VPWR.n44 VPWR.n6 36.1417
R133 VPWR.n45 VPWR.n44 36.1417
R134 VPWR.n46 VPWR.n45 36.1417
R135 VPWR.n46 VPWR.n4 36.1417
R136 VPWR.n50 VPWR.n4 36.1417
R137 VPWR.n51 VPWR.n50 36.1417
R138 VPWR.n52 VPWR.n51 36.1417
R139 VPWR.n27 VPWR.n26 36.1417
R140 VPWR.n28 VPWR.n27 36.1417
R141 VPWR.n28 VPWR.n10 36.1417
R142 VPWR.n32 VPWR.n10 36.1417
R143 VPWR.n33 VPWR.n32 36.1417
R144 VPWR.n34 VPWR.n33 36.1417
R145 VPWR.n34 VPWR.n8 36.1417
R146 VPWR.n38 VPWR.n8 36.1417
R147 VPWR.n23 VPWR.n22 30.5818
R148 VPWR.n1 VPWR.t9 29.5505
R149 VPWR.n22 VPWR.n21 28.6123
R150 VPWR.n39 VPWR.n38 27.4829
R151 VPWR.n58 VPWR.n57 27.1064
R152 VPWR.n16 VPWR.t2 26.3844
R153 VPWR.n16 VPWR.t6 26.3844
R154 VPWR.n56 VPWR.n2 25.6005
R155 VPWR.n20 VPWR.n17 24.0946
R156 VPWR.n52 VPWR.n2 21.8358
R157 VPWR.n26 VPWR.n13 21.3087
R158 VPWR.n40 VPWR.n39 19.9534
R159 VPWR.n21 VPWR.n20 18.824
R160 VPWR.n20 VPWR.n19 9.3005
R161 VPWR.n21 VPWR.n15 9.3005
R162 VPWR.n22 VPWR.n14 9.3005
R163 VPWR.n24 VPWR.n23 9.3005
R164 VPWR.n26 VPWR.n25 9.3005
R165 VPWR.n27 VPWR.n11 9.3005
R166 VPWR.n29 VPWR.n28 9.3005
R167 VPWR.n30 VPWR.n10 9.3005
R168 VPWR.n32 VPWR.n31 9.3005
R169 VPWR.n33 VPWR.n9 9.3005
R170 VPWR.n35 VPWR.n34 9.3005
R171 VPWR.n36 VPWR.n8 9.3005
R172 VPWR.n38 VPWR.n37 9.3005
R173 VPWR.n39 VPWR.n7 9.3005
R174 VPWR.n41 VPWR.n40 9.3005
R175 VPWR.n42 VPWR.n6 9.3005
R176 VPWR.n44 VPWR.n43 9.3005
R177 VPWR.n45 VPWR.n5 9.3005
R178 VPWR.n47 VPWR.n46 9.3005
R179 VPWR.n48 VPWR.n4 9.3005
R180 VPWR.n50 VPWR.n49 9.3005
R181 VPWR.n51 VPWR.n3 9.3005
R182 VPWR.n53 VPWR.n52 9.3005
R183 VPWR.n54 VPWR.n2 9.3005
R184 VPWR.n56 VPWR.n55 9.3005
R185 VPWR.n57 VPWR.n0 9.3005
R186 VPWR.n59 VPWR.n58 9.3005
R187 VPWR.n18 VPWR.n17 6.68184
R188 VPWR.n23 VPWR.n13 2.02155
R189 VPWR.n19 VPWR.n18 0.590726
R190 VPWR.n19 VPWR.n15 0.122949
R191 VPWR.n15 VPWR.n14 0.122949
R192 VPWR.n24 VPWR.n14 0.122949
R193 VPWR.n25 VPWR.n24 0.122949
R194 VPWR.n25 VPWR.n11 0.122949
R195 VPWR.n29 VPWR.n11 0.122949
R196 VPWR.n30 VPWR.n29 0.122949
R197 VPWR.n31 VPWR.n30 0.122949
R198 VPWR.n31 VPWR.n9 0.122949
R199 VPWR.n35 VPWR.n9 0.122949
R200 VPWR.n36 VPWR.n35 0.122949
R201 VPWR.n37 VPWR.n36 0.122949
R202 VPWR.n37 VPWR.n7 0.122949
R203 VPWR.n41 VPWR.n7 0.122949
R204 VPWR.n42 VPWR.n41 0.122949
R205 VPWR.n43 VPWR.n42 0.122949
R206 VPWR.n43 VPWR.n5 0.122949
R207 VPWR.n47 VPWR.n5 0.122949
R208 VPWR.n48 VPWR.n47 0.122949
R209 VPWR.n49 VPWR.n48 0.122949
R210 VPWR.n49 VPWR.n3 0.122949
R211 VPWR.n53 VPWR.n3 0.122949
R212 VPWR.n54 VPWR.n53 0.122949
R213 VPWR.n55 VPWR.n54 0.122949
R214 VPWR.n55 VPWR.n0 0.122949
R215 VPWR.n59 VPWR.n0 0.122949
R216 VPWR VPWR.n59 0.0617245
R217 SUM SUM.n0 241.684
R218 SUM.n2 SUM.n1 107.85
R219 SUM.n0 SUM.t0 27.2639
R220 SUM.n0 SUM.t1 27.2639
R221 SUM.n1 SUM.t2 23.514
R222 SUM.n1 SUM.t3 23.514
R223 SUM.n2 SUM 3.29747
R224 SUM SUM.n2 1.79699
R225 VPB.t14 VPB.t15 927.016
R226 VPB.t4 VPB.t14 875.942
R227 VPB.t11 VPB.t12 763.576
R228 VPB.t5 VPB.t13 543.952
R229 VPB.t3 VPB.t6 505.646
R230 VPB.t12 VPB.t4 505.646
R231 VPB.t8 VPB.t10 503.091
R232 VPB.t15 VPB.t0 349.866
R233 VPB.t0 VPB.t3 342.204
R234 VPB.t13 VPB.t11 311.56
R235 VPB.t10 VPB.t9 260.485
R236 VPB.t9 VPB.t5 257.93
R237 VPB VPB.t8 252.823
R238 VPB.t2 VPB.t1 234.946
R239 VPB.t7 VPB.t2 229.839
R240 VPB.t6 VPB.t7 229.839
R241 a_514_424.n9 a_514_424.n8 601.679
R242 a_514_424.n7 a_514_424.n0 585
R243 a_514_424.n3 a_514_424.t4 568.905
R244 a_514_424.n4 a_514_424.t5 420.295
R245 a_514_424.n6 a_514_424.n5 381.351
R246 a_514_424.n3 a_514_424.n2 357.921
R247 a_514_424.n7 a_514_424.n6 311.584
R248 a_514_424.n8 a_514_424.n1 282.13
R249 a_514_424.n4 a_514_424.n3 134.4
R250 a_514_424.n9 a_514_424.n0 132.506
R251 a_514_424.n6 a_514_424.n4 126.118
R252 a_514_424.n1 a_514_424.t0 88.1255
R253 a_514_424.n0 a_514_424.t3 46.9053
R254 a_514_424.t2 a_514_424.n9 35.1791
R255 a_514_424.n1 a_514_424.t1 26.2505
R256 a_514_424.n8 a_514_424.n7 5.23686
R257 a_2052_424.n1 a_2052_424.n0 881.461
R258 a_2052_424.n3 a_2052_424.n2 59.4722
R259 a_2052_424.n1 a_2052_424.t3 55.1136
R260 a_2052_424.n0 a_2052_424.t1 50.6255
R261 a_2052_424.n2 a_2052_424.n1 38.6969
R262 a_2052_424.n2 a_2052_424.t0 28.1368
R263 a_2052_424.n0 a_2052_424.t2 28.1255
R264 COUT COUT.n0 587.293
R265 COUT COUT.t2 177.347
R266 COUT.n0 COUT.t1 26.3844
R267 COUT.n0 COUT.t0 26.3844
R268 a_481_379.t0 a_481_379.n3 767.322
R269 a_481_379.n0 a_481_379.t4 626.601
R270 a_481_379.n1 a_481_379.n0 379.173
R271 a_481_379.n2 a_481_379.n1 300.594
R272 a_481_379.n3 a_481_379.n2 260.048
R273 a_481_379.n3 a_481_379.t1 256.26
R274 a_481_379.n2 a_481_379.t5 206.238
R275 a_481_379.n1 a_481_379.t2 172.45
R276 a_481_379.n0 a_481_379.t3 126.927
R277 a_481_379.n4 a_481_379.t0 73.5472
R278 a_114_368.n2 a_114_368.n0 648.513
R279 a_114_368.t3 a_114_368.n3 267.704
R280 a_114_368.n2 a_114_368.n1 196.933
R281 a_114_368.n3 a_114_368.t4 171.637
R282 a_114_368.n1 a_114_368.t2 103.126
R283 a_114_368.n1 a_114_368.t0 56.2505
R284 a_114_368.n0 a_114_368.t1 53.941
R285 a_114_368.n0 a_114_368.t5 53.941
R286 a_114_368.n3 a_114_368.n2 26.1209
R287 a_849_424.n1 a_849_424.t6 555.908
R288 a_849_424.n2 a_849_424.n1 467.219
R289 a_849_424.n5 a_849_424.n3 393.252
R290 a_849_424.n6 a_849_424.n5 322.245
R291 a_849_424.n3 a_849_424.n0 237.389
R292 a_849_424.n5 a_849_424.n4 197.607
R293 a_849_424.n6 a_849_424.t3 189.536
R294 a_849_424.n1 a_849_424.t4 168.701
R295 a_849_424.n2 a_849_424.t5 159.06
R296 a_849_424.n3 a_849_424.n2 128.489
R297 a_849_424.t1 a_849_424.n6 110.907
R298 a_849_424.n4 a_849_424.t0 76.8755
R299 a_849_424.n4 a_849_424.t2 53.438
R300 a_1689_424.t2 a_1689_424.n3 872.015
R301 a_1689_424.n1 a_1689_424.t1 541.304
R302 a_1689_424.n2 a_1689_424.t5 259.897
R303 a_1689_424.n2 a_1689_424.t4 224.817
R304 a_1689_424.n3 a_1689_424.n1 209.498
R305 a_1689_424.n3 a_1689_424.n2 152
R306 a_1689_424.n1 a_1689_424.n0 89.2272
R307 a_1689_424.n0 a_1689_424.t0 88.1255
R308 a_1689_424.n0 a_1689_424.t3 39.3755
R309 B.n3 B.t2 429.452
R310 B.n2 B.t5 365.474
R311 B.n4 B.t3 339.981
R312 B.n1 B.t0 311.846
R313 B.n0 B.t1 291.036
R314 B.n2 B.n1 290.656
R315 B.n0 B.t4 204.048
R316 B.n4 B.n3 113.882
R317 B.n3 B.n2 56.8476
R318 B.n1 B.n0 56.4634
R319 B B.n4 2.25932
R320 a_413_392.n2 a_413_392.t0 903.068
R321 a_413_392.n1 a_413_392.t2 593.846
R322 a_413_392.n3 a_413_392.n2 287.077
R323 a_413_392.n2 a_413_392.n1 100.555
R324 a_413_392.n1 a_413_392.n0 89.0318
R325 a_413_392.n3 a_413_392.t3 46.9053
R326 a_413_392.t4 a_413_392.n3 33.07
R327 a_413_392.n0 a_413_392.t1 26.2505
R328 a_413_392.n0 a_413_392.t5 26.2505
R329 CI.n1 CI.n0 250.133
R330 CI.n1 CI.t0 236.983
R331 CI CI.n1 154.327
C0 VPB SUM 0.007201f
C1 VPWR COUT 0.016694f
C2 B COUT 5.74e-21
C3 VGND CI 0.009119f
C4 VPWR SUM 0.175941f
C5 B SUM 1.15e-20
C6 VGND COUT 0.121234f
C7 a_1451_424# VPB 0.095689f
C8 VGND SUM 0.164261f
C9 CI COUT 0.007622f
C10 a_1451_424# VPWR 0.138598f
C11 a_1895_424# VPB 0.098514f
C12 a_1451_424# B 0.001115f
C13 CI SUM 1.65e-19
C14 a_1451_424# A 4.97e-20
C15 a_1895_424# VPWR 0.331944f
C16 a_1895_424# B 2.19e-20
C17 a_1451_424# VGND 0.357318f
C18 COUT SUM 0.005173f
C19 a_1451_424# CI 0.045712f
C20 a_1895_424# VGND 0.059662f
C21 a_1451_424# COUT 0.122983f
C22 a_1895_424# CI 0.010847f
C23 VPB VPWR 0.376624f
C24 VPB B 0.209313f
C25 a_1451_424# SUM 0.002956f
C26 a_1895_424# COUT 0.087189f
C27 VPB A 0.103699f
C28 VPWR B 0.034751f
C29 VPB VGND 0.012324f
C30 a_1895_424# SUM 0.186339f
C31 VPWR A 0.077919f
C32 A B 0.041622f
C33 VPWR VGND 0.098499f
C34 VPB CI 0.05308f
C35 B VGND 0.060112f
C36 a_1451_424# a_1895_424# 0.131326f
C37 A VGND 0.034339f
C38 VPB COUT 0.00684f
C39 VPWR CI 0.012179f
C40 SUM VNB 0.055793f
C41 COUT VNB 0.009295f
C42 CI VNB 0.128363f
C43 VGND VNB 1.65023f
C44 B VNB 0.523791f
C45 A VNB 0.221836f
C46 VPWR VNB 1.33635f
C47 VPB VNB 3.2989f
C48 a_1895_424# VNB 0.239357f
C49 a_1451_424# VNB 0.278532f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fah_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fah_4 VNB VPB VPWR VGND SUM COUT B A CI
X0 VPWR.t3 a_1278_102.t4 SUM.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1736 ps=1.43 w=1.12 l=0.15
X1 a_586_257.t0 B.t0 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.05 as=0.27675 ps=2.42 w=0.74 l=0.15
X2 VPWR.t9 A.t0 a_27_74.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X3 a_1278_102.t2 a_528_362.t4 a_1378_125.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.336 pd=1.64 as=0.22505 ps=1.55 w=0.84 l=0.15
X4 a_1278_102.t3 a_528_362.t5 a_1183_102.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.12205 pd=1.105 as=0.208 ps=1.93 w=0.64 l=0.15
X5 a_200_74.t0 a_586_257.t4 a_536_114.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1222 pd=1.08 as=0.0896 ps=0.92 w=0.64 l=0.15
X6 a_536_114.t2 B.t1 a_427_362.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1165 ps=1.065 w=0.64 l=0.15
X7 a_528_362.t2 B.t2 a_200_74.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1222 ps=1.08 w=0.64 l=0.15
X8 a_1378_125.t1 a_536_114.t4 a_1278_102.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.12205 ps=1.105 w=0.64 l=0.15
X9 a_427_362.t4 a_27_74.t2 VGND.t7 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.418 ps=2.8 w=0.74 l=0.15
X10 VGND.t11 A.t1 a_27_74.t0 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X11 a_1265_379.t2 a_528_362.t6 a_586_257.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1869 pd=1.285 as=0.202175 ps=1.505 w=0.84 l=0.15
X12 a_1378_125.t2 a_536_114.t5 a_1265_379.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.22505 pd=1.55 as=0.1869 ps=1.285 w=0.84 l=0.15
X13 a_586_257.t1 B.t3 VPWR.t12 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.202175 pd=1.505 as=0.3304 ps=2.83 w=1.12 l=0.15
X14 VGND.t2 a_1278_102.t5 SUM.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_1265_379.t3 a_528_362.t7 a_1378_125.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.118425 pd=1.09 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 VPWR.t5 a_1378_125.t6 a_1183_102.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.4505 pd=2.05 as=0.19535 ps=1.5 w=1 l=0.15
X17 VPWR.t4 a_1265_379.t4 COUT.t5 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.8914 pd=4.04 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_528_362.t3 B.t4 a_427_362.t3 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.1281 pd=1.145 as=0.1862 ps=1.475 w=0.84 l=0.15
X19 VGND.t4 a_1265_379.t5 COUT.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.36 pd=2.83 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 COUT.t4 a_1265_379.t6 VPWR.t7 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.297275 ps=1.825 w=1.12 l=0.15
X21 COUT.t1 a_1265_379.t7 VGND.t9 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.3311 ps=1.9 w=0.74 l=0.15
X22 SUM.t5 a_1278_102.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.20925 ps=1.5 w=0.74 l=0.15
X23 VPWR.t2 a_1278_102.t7 SUM.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_200_74.t5 A.t2 VPWR.t10 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X25 a_427_362.t5 a_27_74.t3 VPWR.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.5163 ps=3.55 w=1.12 l=0.15
X26 a_200_74.t1 a_586_257.t5 a_528_362.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.23945 pd=1.6 as=0.1281 ps=1.145 w=0.84 l=0.15
X27 SUM.t1 a_1278_102.t8 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2382 ps=1.555 w=1.12 l=0.15
X28 a_1183_102.t2 a_536_114.t6 a_1278_102.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.19535 pd=1.5 as=0.336 ps=1.64 w=0.84 l=0.15
X29 a_200_74.t4 A.t3 VGND.t8 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X30 SUM.t0 a_1278_102.t9 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.2184 ps=1.51 w=1.12 l=0.15
X31 a_427_362.t0 a_586_257.t6 a_536_114.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X32 a_536_114.t3 B.t5 a_200_74.t2 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.23945 ps=1.6 w=0.84 l=0.15
X33 VGND.t5 a_1378_125.t7 a_1183_102.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.3311 pd=1.9 as=0.23505 ps=2.02 w=0.64 l=0.15
X34 VGND.t3 CI.t0 a_1378_125.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.20925 pd=1.5 as=0.1824 ps=1.85 w=0.64 l=0.15
X35 VGND.t0 a_1278_102.t10 SUM.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X36 a_586_257.t2 a_536_114.t7 a_1265_379.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.356425 pd=3.14 as=0.118425 ps=1.09 w=0.64 l=0.15
X37 VGND.t10 a_1265_379.t8 COUT.t0 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.18675 pd=1.45 as=0.1036 ps=1.02 w=0.74 l=0.15
X38 a_427_362.t1 a_586_257.t7 a_528_362.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1024 ps=0.96 w=0.64 l=0.15
X39 COUT.t3 a_1265_379.t9 VPWR.t8 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4505 ps=2.05 w=1.12 l=0.15
X40 VPWR.t11 CI.t1 a_1378_125.t5 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.295 ps=2.59 w=1 l=0.15
R0 a_1278_102.n13 a_1278_102.n12 679.894
R1 a_1278_102.n12 a_1278_102.n11 626.389
R2 a_1278_102.n9 a_1278_102.t8 244.335
R3 a_1278_102.n3 a_1278_102.t4 228.69
R4 a_1278_102.n5 a_1278_102.t9 226.809
R5 a_1278_102.n1 a_1278_102.t7 226.809
R6 a_1278_102.n6 a_1278_102.n0 165.189
R7 a_1278_102.n3 a_1278_102.t5 154.24
R8 a_1278_102.n8 a_1278_102.t6 154.24
R9 a_1278_102.n7 a_1278_102.t10 154.24
R10 a_1278_102.n4 a_1278_102.n2 154.24
R11 a_1278_102.n13 a_1278_102.t2 152.44
R12 a_1278_102.n10 a_1278_102.n9 152
R13 a_1278_102.n1 a_1278_102.n0 152
R14 a_1278_102.n12 a_1278_102.n10 140.252
R15 a_1278_102.n4 a_1278_102.n3 62.8066
R16 a_1278_102.n8 a_1278_102.n1 44.549
R17 a_1278_102.n11 a_1278_102.t0 39.2856
R18 a_1278_102.t1 a_1278_102.n13 35.1791
R19 a_1278_102.n7 a_1278_102.n6 32.8641
R20 a_1278_102.n6 a_1278_102.n5 27.752
R21 a_1278_102.n11 a_1278_102.t3 26.3721
R22 a_1278_102.n1 a_1278_102.n7 18.2581
R23 a_1278_102.n10 a_1278_102.n0 13.1884
R24 a_1278_102.n9 a_1278_102.n8 3.65202
R25 a_1278_102.n5 a_1278_102.n4 2.19141
R26 SUM.n5 SUM.n4 585
R27 SUM.n6 SUM.n5 291.087
R28 SUM.n3 SUM.n0 256.964
R29 SUM.n2 SUM.n1 153.055
R30 SUM.n2 SUM.t6 146.25
R31 SUM.n3 SUM.n2 41.9043
R32 SUM.n5 SUM.t0 28.1434
R33 SUM.n5 SUM.t3 26.3844
R34 SUM.n0 SUM.t2 26.3844
R35 SUM.n0 SUM.t1 26.3844
R36 SUM.n1 SUM.t4 22.7032
R37 SUM.n1 SUM.t5 22.7032
R38 SUM.n4 SUM 11.6542
R39 SUM.n6 SUM 8.81684
R40 SUM SUM.n6 5.22933
R41 SUM.n4 SUM 2.48408
R42 SUM SUM.n3 0.573634
R43 VPWR.n2 VPWR.t6 949.956
R44 VPWR.n31 VPWR.t7 874.068
R45 VPWR.n25 VPWR.t4 772.279
R46 VPWR.n34 VPWR.n33 651.006
R47 VPWR.n6 VPWR.t12 342.973
R48 VPWR.n18 VPWR.n17 316.87
R49 VPWR.n16 VPWR.t3 266.057
R50 VPWR.n64 VPWR.n1 230.78
R51 VPWR.n15 VPWR.n14 223.121
R52 VPWR.n33 VPWR.t5 78.8005
R53 VPWR.n14 VPWR.t11 46.2955
R54 VPWR.n33 VPWR.t8 42.5041
R55 VPWR.n52 VPWR.n51 36.1417
R56 VPWR.n53 VPWR.n52 36.1417
R57 VPWR.n53 VPWR.n4 36.1417
R58 VPWR.n57 VPWR.n4 36.1417
R59 VPWR.n58 VPWR.n57 36.1417
R60 VPWR.n59 VPWR.n58 36.1417
R61 VPWR.n40 VPWR.n39 36.1417
R62 VPWR.n41 VPWR.n40 36.1417
R63 VPWR.n41 VPWR.n8 36.1417
R64 VPWR.n45 VPWR.n8 36.1417
R65 VPWR.n46 VPWR.n45 36.1417
R66 VPWR.n47 VPWR.n46 36.1417
R67 VPWR.n35 VPWR.n32 36.1417
R68 VPWR.n30 VPWR.n12 36.1417
R69 VPWR.n24 VPWR.n23 36.1417
R70 VPWR.n14 VPWR.t1 35.2408
R71 VPWR.n17 VPWR.t2 35.1791
R72 VPWR.n17 VPWR.t0 33.4201
R73 VPWR.n19 VPWR.n15 32.377
R74 VPWR.n63 VPWR.n62 31.256
R75 VPWR.n1 VPWR.t10 29.5505
R76 VPWR.n1 VPWR.t9 29.5505
R77 VPWR.n64 VPWR.n63 28.9887
R78 VPWR.n47 VPWR.n6 25.977
R79 VPWR.n39 VPWR.n10 24.4387
R80 VPWR.n26 VPWR.n12 23.4834
R81 VPWR.n59 VPWR.n2 23.3374
R82 VPWR.n51 VPWR.n6 21.4593
R83 VPWR.n35 VPWR.n34 19.5163
R84 VPWR.n19 VPWR.n18 18.0711
R85 VPWR.n25 VPWR.n24 17.3303
R86 VPWR.n23 VPWR.n15 15.0593
R87 VPWR.n32 VPWR.n31 12.4483
R88 VPWR.n20 VPWR.n19 9.3005
R89 VPWR.n21 VPWR.n15 9.3005
R90 VPWR.n23 VPWR.n22 9.3005
R91 VPWR.n24 VPWR.n13 9.3005
R92 VPWR.n27 VPWR.n26 9.3005
R93 VPWR.n28 VPWR.n12 9.3005
R94 VPWR.n30 VPWR.n29 9.3005
R95 VPWR.n32 VPWR.n11 9.3005
R96 VPWR.n36 VPWR.n35 9.3005
R97 VPWR.n37 VPWR.n10 9.3005
R98 VPWR.n39 VPWR.n38 9.3005
R99 VPWR.n40 VPWR.n9 9.3005
R100 VPWR.n42 VPWR.n41 9.3005
R101 VPWR.n43 VPWR.n8 9.3005
R102 VPWR.n45 VPWR.n44 9.3005
R103 VPWR.n46 VPWR.n7 9.3005
R104 VPWR.n48 VPWR.n47 9.3005
R105 VPWR.n49 VPWR.n6 9.3005
R106 VPWR.n51 VPWR.n50 9.3005
R107 VPWR.n52 VPWR.n5 9.3005
R108 VPWR.n54 VPWR.n53 9.3005
R109 VPWR.n55 VPWR.n4 9.3005
R110 VPWR.n57 VPWR.n56 9.3005
R111 VPWR.n58 VPWR.n3 9.3005
R112 VPWR.n60 VPWR.n59 9.3005
R113 VPWR.n62 VPWR.n61 9.3005
R114 VPWR.n63 VPWR.n0 9.3005
R115 VPWR.n31 VPWR.n30 7.93067
R116 VPWR.n65 VPWR.n64 7.27223
R117 VPWR.n18 VPWR.n16 6.97636
R118 VPWR.n62 VPWR.n2 1.87016
R119 VPWR.n26 VPWR.n25 1.37684
R120 VPWR.n34 VPWR.n10 1.10158
R121 VPWR.n20 VPWR.n16 0.569174
R122 VPWR VPWR.n65 0.157962
R123 VPWR.n65 VPWR.n0 0.149814
R124 VPWR.n21 VPWR.n20 0.122949
R125 VPWR.n22 VPWR.n21 0.122949
R126 VPWR.n22 VPWR.n13 0.122949
R127 VPWR.n27 VPWR.n13 0.122949
R128 VPWR.n28 VPWR.n27 0.122949
R129 VPWR.n29 VPWR.n28 0.122949
R130 VPWR.n29 VPWR.n11 0.122949
R131 VPWR.n36 VPWR.n11 0.122949
R132 VPWR.n37 VPWR.n36 0.122949
R133 VPWR.n38 VPWR.n37 0.122949
R134 VPWR.n38 VPWR.n9 0.122949
R135 VPWR.n42 VPWR.n9 0.122949
R136 VPWR.n43 VPWR.n42 0.122949
R137 VPWR.n44 VPWR.n43 0.122949
R138 VPWR.n44 VPWR.n7 0.122949
R139 VPWR.n48 VPWR.n7 0.122949
R140 VPWR.n49 VPWR.n48 0.122949
R141 VPWR.n50 VPWR.n49 0.122949
R142 VPWR.n50 VPWR.n5 0.122949
R143 VPWR.n54 VPWR.n5 0.122949
R144 VPWR.n55 VPWR.n54 0.122949
R145 VPWR.n56 VPWR.n55 0.122949
R146 VPWR.n56 VPWR.n3 0.122949
R147 VPWR.n60 VPWR.n3 0.122949
R148 VPWR.n61 VPWR.n60 0.122949
R149 VPWR.n61 VPWR.n0 0.122949
R150 VPB.n0 VPB 4290.32
R151 VPB.n1 VPB 3713.16
R152 VPB.t9 VPB.t20 816.799
R153 VPB.t4 VPB.t17 727.823
R154 VPB VPB.n2 711.244
R155 VPB.t14 VPB.t13 546.505
R156 VPB.t10 VPB.n0 481.579
R157 VPB.t5 VPB.t14 439.248
R158 VPB.n2 VPB.t12 324.207
R159 VPB.t8 VPB.t18 311.64
R160 VPB.t11 VPB.t6 299.075
R161 VPB.t17 VPB.t1 298.791
R162 VPB.t2 VPB.t0 275.807
R163 VPB.t7 VPB.t5 273.253
R164 VPB.t20 VPB.t11 268.916
R165 VPB.t15 VPB 257.93
R166 VPB.t12 VPB.t19 253.837
R167 VPB.t0 VPB.t3 234.946
R168 VPB.n2 VPB.t16 234.946
R169 VPB.t1 VPB.t2 229.839
R170 VPB.t13 VPB.t4 229.839
R171 VPB.t16 VPB.t15 229.839
R172 VPB.t19 VPB.t8 228.704
R173 VPB.n1 VPB.t10 226.316
R174 VPB.t18 VPB.t9 226.19
R175 VPB.t6 VPB.n1 105.556
R176 VPB.n0 VPB.t7 9.0728
R177 B.n0 B.t4 545.731
R178 B.t4 B.t1 410.425
R179 B.n3 B.t3 401.668
R180 B.t5 B.t2 384.488
R181 B.n1 B.n0 367.358
R182 B.n0 B.t5 258.139
R183 B.n4 B.t0 171.344
R184 B.n5 B.n4 169.409
R185 B B.n1 153.468
R186 B.n7 B.n6 152
R187 B.n5 B.n2 152
R188 B.n9 B.n8 152
R189 B.n8 B.n1 35.2435
R190 B.n8 B.n7 35.2435
R191 B.n7 B.n2 35.2435
R192 B.n4 B.n3 31.6156
R193 B.n6 B.n5 17.4085
R194 B.n6 B 12.3205
R195 B B.n9 7.6005
R196 B.n3 B.n2 3.62846
R197 B.n9 B 2.26717
R198 VGND.n26 VGND.t10 388.195
R199 VGND.n22 VGND.t4 387.914
R200 VGND.n48 VGND.t6 335.967
R201 VGND.n29 VGND.n28 310.269
R202 VGND.n59 VGND.t7 302.2
R203 VGND.n16 VGND.t0 285.01
R204 VGND.n14 VGND.n13 283
R205 VGND.n15 VGND.t2 166.399
R206 VGND.n28 VGND.t5 126.562
R207 VGND.n62 VGND.n61 122.001
R208 VGND.n13 VGND.t3 48.7505
R209 VGND.n30 VGND.n27 36.1417
R210 VGND.n34 VGND.n9 36.1417
R211 VGND.n35 VGND.n34 36.1417
R212 VGND.n36 VGND.n35 36.1417
R213 VGND.n36 VGND.n7 36.1417
R214 VGND.n40 VGND.n7 36.1417
R215 VGND.n41 VGND.n40 36.1417
R216 VGND.n42 VGND.n41 36.1417
R217 VGND.n42 VGND.n5 36.1417
R218 VGND.n46 VGND.n5 36.1417
R219 VGND.n47 VGND.n46 36.1417
R220 VGND.n49 VGND.n3 36.1417
R221 VGND.n53 VGND.n3 36.1417
R222 VGND.n54 VGND.n53 36.1417
R223 VGND.n55 VGND.n54 36.1417
R224 VGND.n55 VGND.n1 36.1417
R225 VGND.n26 VGND.n11 35.0123
R226 VGND.n22 VGND.n21 32.0005
R227 VGND.n62 VGND.n60 30.4946
R228 VGND.n59 VGND.n1 27.4829
R229 VGND.n21 VGND.n20 27.3284
R230 VGND.n17 VGND.n14 26.6849
R231 VGND.n61 VGND.t8 26.2505
R232 VGND.n61 VGND.t11 26.2505
R233 VGND.n13 VGND.t1 25.2248
R234 VGND.n60 VGND.n59 25.224
R235 VGND.n28 VGND.t9 24.317
R236 VGND.n17 VGND.n16 22.9652
R237 VGND.n29 VGND.n9 16.9417
R238 VGND.n22 VGND.n11 15.4358
R239 VGND.n27 VGND.n26 12.424
R240 VGND.n48 VGND.n47 9.41227
R241 VGND.n60 VGND.n0 9.3005
R242 VGND.n59 VGND.n58 9.3005
R243 VGND.n57 VGND.n1 9.3005
R244 VGND.n56 VGND.n55 9.3005
R245 VGND.n54 VGND.n2 9.3005
R246 VGND.n53 VGND.n52 9.3005
R247 VGND.n51 VGND.n3 9.3005
R248 VGND.n50 VGND.n49 9.3005
R249 VGND.n47 VGND.n4 9.3005
R250 VGND.n46 VGND.n45 9.3005
R251 VGND.n44 VGND.n5 9.3005
R252 VGND.n43 VGND.n42 9.3005
R253 VGND.n41 VGND.n6 9.3005
R254 VGND.n40 VGND.n39 9.3005
R255 VGND.n38 VGND.n7 9.3005
R256 VGND.n37 VGND.n36 9.3005
R257 VGND.n35 VGND.n8 9.3005
R258 VGND.n34 VGND.n33 9.3005
R259 VGND.n32 VGND.n9 9.3005
R260 VGND.n31 VGND.n30 9.3005
R261 VGND.n27 VGND.n10 9.3005
R262 VGND.n26 VGND.n25 9.3005
R263 VGND.n24 VGND.n11 9.3005
R264 VGND.n23 VGND.n22 9.3005
R265 VGND.n21 VGND.n12 9.3005
R266 VGND.n20 VGND.n19 9.3005
R267 VGND.n18 VGND.n17 9.3005
R268 VGND.n63 VGND.n62 7.19894
R269 VGND.n16 VGND.n15 6.6595
R270 VGND.n49 VGND.n48 1.88285
R271 VGND.n18 VGND.n15 0.655456
R272 VGND.n30 VGND.n29 0.376971
R273 VGND VGND.n63 0.156997
R274 VGND.n63 VGND.n0 0.150766
R275 VGND.n19 VGND.n18 0.122949
R276 VGND.n19 VGND.n12 0.122949
R277 VGND.n23 VGND.n12 0.122949
R278 VGND.n24 VGND.n23 0.122949
R279 VGND.n25 VGND.n24 0.122949
R280 VGND.n25 VGND.n10 0.122949
R281 VGND.n31 VGND.n10 0.122949
R282 VGND.n32 VGND.n31 0.122949
R283 VGND.n33 VGND.n32 0.122949
R284 VGND.n33 VGND.n8 0.122949
R285 VGND.n37 VGND.n8 0.122949
R286 VGND.n38 VGND.n37 0.122949
R287 VGND.n39 VGND.n38 0.122949
R288 VGND.n39 VGND.n6 0.122949
R289 VGND.n43 VGND.n6 0.122949
R290 VGND.n44 VGND.n43 0.122949
R291 VGND.n45 VGND.n44 0.122949
R292 VGND.n45 VGND.n4 0.122949
R293 VGND.n50 VGND.n4 0.122949
R294 VGND.n51 VGND.n50 0.122949
R295 VGND.n52 VGND.n51 0.122949
R296 VGND.n52 VGND.n2 0.122949
R297 VGND.n56 VGND.n2 0.122949
R298 VGND.n57 VGND.n56 0.122949
R299 VGND.n58 VGND.n57 0.122949
R300 VGND.n58 VGND.n0 0.122949
R301 VGND.n20 VGND.n14 0.109902
R302 a_586_257.n1 a_586_257.n6 336.543
R303 a_586_257.n4 a_586_257.t2 617.585
R304 a_586_257.n2 a_586_257.t4 505.233
R305 a_586_257.t4 a_586_257.t5 406.488
R306 a_586_257.t7 a_586_257.t6 375.024
R307 a_586_257.n1 a_586_257.n0 15.8645
R308 a_586_257.n3 a_586_257.n2 221.556
R309 a_586_257.n5 a_586_257.n4 188.244
R310 a_586_257.n6 a_586_257.n5 188.244
R311 a_586_257.n2 a_586_257.t7 156.046
R312 a_586_257.n0 a_586_257.t3 55.1136
R313 a_586_257.n0 a_586_257.t1 28.9519
R314 a_586_257.n5 a_586_257.t0 21.0816
R315 a_586_257.n7 a_586_257.n1 54.6316
R316 a_586_257.n4 a_586_257.n3 12.1811
R317 a_586_257.n6 a_586_257.n3 1.85856
R318 VNB VNB.n0 16295
R319 VNB.t13 VNB.t8 3903.41
R320 VNB.t14 VNB.t11 3027.2
R321 VNB.t15 VNB.t16 2827.73
R322 VNB.t7 VNB.t6 2471.39
R323 VNB.t11 VNB.t4 2370.13
R324 VNB.t8 VNB.t17 2309.71
R325 VNB.t18 VNB.t7 2263.52
R326 VNB.t0 VNB.t2 1986.35
R327 VNB.t6 VNB.t1 1385.83
R328 VNB.t9 VNB.t5 1196.8
R329 VNB.t12 VNB.t14 1173.33
R330 VNB.t19 VNB 1161.6
R331 VNB.t3 VNB.t13 1131.76
R332 VNB.t10 VNB.t15 1114.67
R333 VNB.t4 VNB.t9 1102.93
R334 VNB.t5 VNB.t10 1009.07
R335 VNB.t16 VNB.t19 1009.07
R336 VNB.t1 VNB.t0 993.177
R337 VNB.t17 VNB.t18 993.177
R338 VNB.n0 VNB.t12 563.201
R339 VNB.n0 VNB.t3 438.846
R340 A.n2 A.t1 252.101
R341 A.n1 A.t3 250.641
R342 A.n0 A.t2 211.179
R343 A.n2 A.t0 184.768
R344 A A.n0 165.022
R345 A A.n3 153.987
R346 A.n3 A.n1 48.9308
R347 A.n3 A.n2 12.4157
R348 A.n1 A.n0 0.730803
R349 a_27_74.n1 a_27_74.n0 384.983
R350 a_27_74.t1 a_27_74.n1 291.841
R351 a_27_74.n0 a_27_74.t3 275.009
R352 a_27_74.n0 a_27_74.t2 176.733
R353 a_27_74.n1 a_27_74.t0 151.053
R354 a_528_362.t6 a_528_362.t4 780.304
R355 a_528_362.n3 a_528_362.n2 618.518
R356 a_528_362.t4 a_528_362.t7 490.168
R357 a_528_362.n2 a_528_362.n0 353.846
R358 a_528_362.n0 a_528_362.t6 278.221
R359 a_528_362.n2 a_528_362.n1 155.115
R360 a_528_362.n0 a_528_362.t5 147.814
R361 a_528_362.t1 a_528_362.n3 36.3517
R362 a_528_362.n3 a_528_362.t3 35.1791
R363 a_528_362.n1 a_528_362.t2 33.7505
R364 a_528_362.n1 a_528_362.t0 26.2505
R365 a_1378_125.n3 a_1378_125.n2 589.477
R366 a_1378_125.n3 a_1378_125.n1 413.844
R367 a_1378_125.n5 a_1378_125.n4 355.113
R368 a_1378_125.n5 a_1378_125.t0 352.577
R369 a_1378_125.n0 a_1378_125.t7 258.966
R370 a_1378_125.n4 a_1378_125.n0 247.37
R371 a_1378_125.t5 a_1378_125.n5 220.232
R372 a_1378_125.n0 a_1378_125.t6 215.561
R373 a_1378_125.n2 a_1378_125.t2 83.1649
R374 a_1378_125.n2 a_1378_125.t3 46.9053
R375 a_1378_125.n1 a_1378_125.t4 26.2505
R376 a_1378_125.n1 a_1378_125.t1 26.2505
R377 a_1378_125.n4 a_1378_125.n3 21.3948
R378 a_1183_102.n2 a_1183_102.n1 619.053
R379 a_1183_102.n1 a_1183_102.t0 260.132
R380 a_1183_102.n1 a_1183_102.t3 211.643
R381 a_1183_102.n2 a_1183_102.n0 76.7971
R382 a_1183_102.n0 a_1183_102.t2 59.0942
R383 a_1183_102.n0 a_1183_102.t1 32.062
R384 a_1183_102.n3 a_1183_102.n2 16.6954
R385 a_536_114.t4 a_536_114.t7 774.413
R386 a_536_114.t7 a_536_114.t6 604.107
R387 a_536_114.n3 a_536_114.n2 603.336
R388 a_536_114.n1 a_536_114.t5 205.922
R389 a_536_114.n2 a_536_114.n0 191.07
R390 a_536_114.n2 a_536_114.n1 187.671
R391 a_536_114.n1 a_536_114.t4 171.913
R392 a_536_114.t1 a_536_114.n3 35.1791
R393 a_536_114.n3 a_536_114.t3 35.1791
R394 a_536_114.n0 a_536_114.t0 26.2505
R395 a_536_114.n0 a_536_114.t2 26.2505
R396 a_200_74.n3 a_200_74.n2 783.641
R397 a_200_74.n1 a_200_74.n0 328.745
R398 a_200_74.t5 a_200_74.n3 273.807
R399 a_200_74.n1 a_200_74.t4 170.482
R400 a_200_74.n3 a_200_74.n1 122.73
R401 a_200_74.n2 a_200_74.t2 55.1136
R402 a_200_74.n2 a_200_74.t1 55.1136
R403 a_200_74.n0 a_200_74.t3 42.0902
R404 a_200_74.n0 a_200_74.t0 23.133
R405 a_427_362.n0 a_427_362.t1 329.933
R406 a_427_362.n0 a_427_362.t0 326.019
R407 a_427_362.n3 a_427_362.n2 288.673
R408 a_427_362.n2 a_427_362.n1 266.445
R409 a_427_362.n2 a_427_362.n0 144.679
R410 a_427_362.n5 a_427_362.n4 104.076
R411 a_427_362.n3 a_427_362.t3 35.1791
R412 a_427_362.n1 a_427_362.t4 31.0986
R413 a_427_362.n4 a_427_362.t5 26.5935
R414 a_427_362.n1 a_427_362.t2 26.2505
R415 a_427_362.n4 a_427_362.n3 17.5898
R416 a_1265_379.n15 a_1265_379.n14 725.09
R417 a_1265_379.n11 a_1265_379.t9 237.762
R418 a_1265_379.n5 a_1265_379.t6 226.809
R419 a_1265_379.n9 a_1265_379.n1 226.809
R420 a_1265_379.n4 a_1265_379.t4 225.47
R421 a_1265_379.n3 a_1265_379.t5 216.109
R422 a_1265_379.n14 a_1265_379.n12 213.34
R423 a_1265_379.n14 a_1265_379.n13 185
R424 a_1265_379.n7 a_1265_379.n0 165.189
R425 a_1265_379.n3 a_1265_379.n2 154.24
R426 a_1265_379.n8 a_1265_379.t7 154.24
R427 a_1265_379.n6 a_1265_379.t8 154.24
R428 a_1265_379.n12 a_1265_379.n11 152
R429 a_1265_379.n10 a_1265_379.n0 152
R430 a_1265_379.n15 a_1265_379.t2 69.185
R431 a_1265_379.n5 a_1265_379.n4 65.5316
R432 a_1265_379.n11 a_1265_379.n10 49.6611
R433 a_1265_379.n7 a_1265_379.n6 39.4369
R434 a_1265_379.n13 a_1265_379.t3 39.0791
R435 a_1265_379.t1 a_1265_379.n15 35.1791
R436 a_1265_379.n13 a_1265_379.t0 24.2636
R437 a_1265_379.n8 a_1265_379.n7 23.3702
R438 a_1265_379.n9 a_1265_379.n8 21.1793
R439 a_1265_379.n12 a_1265_379.n0 13.1884
R440 a_1265_379.n4 a_1265_379.n3 7.91393
R441 a_1265_379.n6 a_1265_379.n5 6.57323
R442 a_1265_379.n10 a_1265_379.n9 5.11262
R443 COUT.n1 COUT.t3 884.154
R444 COUT.n1 COUT.n0 586.178
R445 COUT.n3 COUT.t2 292.95
R446 COUT.n3 COUT.n2 210.272
R447 COUT.n0 COUT.t5 26.3844
R448 COUT.n0 COUT.t4 26.3844
R449 COUT.n2 COUT.t0 22.7032
R450 COUT.n2 COUT.t1 22.7032
R451 COUT COUT.n3 13.0948
R452 COUT COUT.n1 11.6235
R453 CI.n0 CI.t1 231.629
R454 CI.n0 CI.t0 162.274
R455 CI CI.n0 157.358
C0 VPWR SUM 0.429116f
C1 VGND COUT 0.025909f
C2 VGND CI 0.007425f
C3 VGND SUM 0.220466f
C4 VPB VPWR 0.379799f
C5 COUT SUM 3.97e-19
C6 VPB A 0.0931f
C7 CI SUM 0.003483f
C8 VPWR A 0.071123f
C9 VPB B 0.53524f
C10 VPWR B 0.181603f
C11 VPB VGND 0.017669f
C12 VPWR VGND 0.163649f
C13 A B 0.001626f
C14 VPB COUT 0.009015f
C15 A VGND 0.034924f
C16 VPWR COUT 0.035786f
C17 VPB CI 0.046608f
C18 VPWR CI 0.02744f
C19 B VGND 0.022633f
C20 VPB SUM 0.012378f
C21 SUM VNB 0.031847f
C22 CI VNB 0.111806f
C23 COUT VNB 0.007579f
C24 VGND VNB 1.75894f
C25 B VNB 0.415395f
C26 A VNB 0.253311f
C27 VPWR VNB 1.3796f
C28 VPB VNB 3.52459f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fahcin_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fahcin_1 VNB VPB VPWR VGND COUT B A CIN SUM
X0 a_1854_368.t2 a_430_418.t4 a_2004_136.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.43155 pd=3.07 as=0.126 ps=1.14 w=0.84 l=0.15
X1 a_2004_136.t0 a_608_74.t4 a_1967_384.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 a_1197_368.t1 a_492_48.t2 VGND.t6 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1981 ps=1.32 w=0.64 l=0.15
X3 a_1595_400.t0 a_608_74.t5 COUT.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.4528 ps=2.055 w=0.64 l=0.15
X4 a_1197_368.t2 a_492_48.t3 VPWR.t6 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2063 pd=1.435 as=0.227 ps=1.535 w=1 l=0.15
X5 a_1967_384.t3 a_430_418.t5 a_2004_136.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1404 pd=1.145 as=0.2544 ps=1.435 w=0.64 l=0.15
X6 VPWR.t3 B.t0 a_492_48.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.227 pd=1.535 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 a_256_368.t3 a_492_48.t4 a_430_418.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.18 as=0.273 ps=2.33 w=0.84 l=0.15
X8 VGND.t4 A.t0 a_28_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.26095 pd=1.5 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_28_74.t3 a_492_48.t5 a_430_418.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X10 VPWR.t5 A.t1 a_28_74.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2877 pd=1.66 as=0.3304 ps=2.83 w=1.12 l=0.15
X11 VGND.t1 B.t1 a_492_48.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1981 pd=1.32 as=0.222 ps=2.08 w=0.74 l=0.15
X12 a_256_368.t0 a_28_74.t6 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.26095 ps=1.5 w=0.64 l=0.15
X13 a_608_74.t0 B.t2 a_28_74.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.17015 pd=1.395 as=0.0896 ps=0.92 w=0.64 l=0.15
X14 VPWR.t7 CIN.t0 a_1595_400.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2952 pd=1.675 as=0.2128 ps=1.44 w=1 l=0.15
X15 a_1854_368.t0 CIN.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2952 ps=1.675 w=1.12 l=0.15
X16 VPWR.t2 a_1854_368.t4 a_1967_384.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2827 pd=1.65 as=0.295 ps=2.59 w=1 l=0.15
X17 a_256_368.t1 a_28_74.t7 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2877 ps=1.66 w=1 l=0.15
X18 a_608_74.t3 B.t3 a_256_368.t4 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.17875 pd=1.42 as=0.1428 ps=1.18 w=0.84 l=0.15
X19 a_28_74.t2 a_492_48.t6 a_608_74.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2373 pd=1.405 as=0.17875 ps=1.42 w=0.84 l=0.15
X20 SUM.t1 a_2004_136.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2827 ps=1.65 w=1.12 l=0.15
X21 COUT.t0 a_608_74.t6 a_1197_368.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.5271 pd=2.095 as=0.2063 ps=1.435 w=0.84 l=0.15
X22 a_256_368.t2 a_492_48.t7 a_608_74.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1632 pd=1.15 as=0.17015 ps=1.395 w=0.64 l=0.15
X23 a_1854_368.t3 CIN.t2 VGND.t7 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.2372 ps=1.65 w=0.74 l=0.15
X24 VGND.t3 a_1854_368.t5 a_1967_384.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.29825 pd=1.59 as=0.1404 ps=1.145 w=0.64 l=0.15
X25 SUM.t0 a_2004_136.t5 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.29825 ps=1.59 w=0.74 l=0.15
X26 a_430_418.t3 B.t4 a_28_74.t5 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.2604 pd=2.3 as=0.2373 ps=1.405 w=0.84 l=0.15
X27 VGND.t5 CIN.t3 a_1595_400.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2372 pd=1.65 as=0.112 ps=0.99 w=0.64 l=0.15
X28 a_430_418.t0 B.t5 a_256_368.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1952 pd=1.89 as=0.1632 ps=1.15 w=0.64 l=0.15
X29 a_2004_136.t1 a_608_74.t7 a_1854_368.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2544 pd=1.435 as=0.1165 ps=1.065 w=0.64 l=0.15
R0 a_430_418.t2 a_430_418.n7 732.891
R1 a_430_418.n3 a_430_418.n1 389.897
R2 a_430_418.n5 a_430_418.t3 383.443
R3 a_430_418.n3 a_430_418.n2 319.699
R4 a_430_418.n7 a_430_418.t1 273.099
R5 a_430_418.n5 a_430_418.t0 271.774
R6 a_430_418.n0 a_430_418.t4 199.494
R7 a_430_418.n4 a_430_418.n0 181.266
R8 a_430_418.n0 a_430_418.t5 155.847
R9 a_430_418.n4 a_430_418.n3 92.5163
R10 a_430_418.n7 a_430_418.n6 11.342
R11 a_430_418.n6 a_430_418.n5 9.3005
R12 a_430_418.n6 a_430_418.n4 2.47061
R13 a_2004_136.n5 a_2004_136.n4 626.216
R14 a_2004_136.n1 a_2004_136.n0 332.005
R15 a_2004_136.n0 a_2004_136.t4 245.522
R16 a_2004_136.n0 a_2004_136.t5 172.953
R17 a_2004_136.n4 a_2004_136.n3 96.3159
R18 a_2004_136.n2 a_2004_136.n1 92.5005
R19 a_2004_136.n3 a_2004_136.n2 82.5005
R20 a_2004_136.n3 a_2004_136.t1 40.313
R21 a_2004_136.n5 a_2004_136.t2 35.1791
R22 a_2004_136.t0 a_2004_136.n5 35.1791
R23 a_2004_136.n2 a_2004_136.t3 26.2505
R24 a_2004_136.n4 a_2004_136.n1 7.01588
R25 a_1854_368.n2 a_1854_368.t2 879.98
R26 a_1854_368.n2 a_1854_368.n1 313.825
R27 a_1854_368.n1 a_1854_368.t4 224.272
R28 a_1854_368.t0 a_1854_368.n3 217.018
R29 a_1854_368.n3 a_1854_368.n0 163.715
R30 a_1854_368.n1 a_1854_368.t5 154.917
R31 a_1854_368.n3 a_1854_368.n2 102.168
R32 a_1854_368.n0 a_1854_368.t3 29.2236
R33 a_1854_368.n0 a_1854_368.t1 28.1255
R34 VPB.t6 VPB.t13 1018.95
R35 VPB.t8 VPB.t10 686.962
R36 VPB.t7 VPB.t2 572.043
R37 VPB.t12 VPB.t3 538.845
R38 VPB.t0 VPB.t5 515.861
R39 VPB.t4 VPB.t12 365.188
R40 VPB.t13 VPB.t0 360.082
R41 VPB.t9 VPB.t8 352.42
R42 VPB.t2 VPB.t1 347.312
R43 VPB.t14 VPB.t6 298.791
R44 VPB.t3 VPB.t14 288.575
R45 VPB.t11 VPB.t4 273.253
R46 VPB VPB.t9 263.038
R47 VPB.t10 VPB.t11 250.269
R48 VPB.t5 VPB.t7 229.839
R49 a_608_74.n0 a_608_74.t7 547.532
R50 a_608_74.t7 a_608_74.t4 441.031
R51 a_608_74.n0 a_608_74.t5 429.935
R52 a_608_74.n1 a_608_74.t6 407.647
R53 a_608_74.n5 a_608_74.n3 292.344
R54 a_608_74.n3 a_608_74.n1 288.753
R55 a_608_74.n3 a_608_74.n2 170.143
R56 a_608_74.n1 a_608_74.n0 105.043
R57 a_608_74.n2 a_608_74.t0 98.9813
R58 a_608_74.n4 a_608_74.t3 64.1585
R59 a_608_74.n6 a_608_74.n5 49.3499
R60 a_608_74.n4 a_608_74.t2 35.1094
R61 a_608_74.n2 a_608_74.t1 20.1094
R62 a_608_74.n5 a_608_74.n4 16.5209
R63 a_1967_384.t1 a_1967_384.n2 802.034
R64 a_1967_384.t1 a_1967_384.n0 744.169
R65 a_1967_384.n0 a_1967_384.t2 474.099
R66 a_1967_384.n2 a_1967_384.n1 173.715
R67 a_1967_384.n1 a_1967_384.t3 55.7673
R68 a_1967_384.n1 a_1967_384.t0 22.9459
R69 a_1967_384.n2 a_1967_384.n0 13.6732
R70 a_492_48.t1 a_492_48.n5 876.952
R71 a_492_48.n3 a_492_48.n2 345.88
R72 a_492_48.n0 a_492_48.t4 252.782
R73 a_492_48.n4 a_492_48.t3 249.197
R74 a_492_48.n0 a_492_48.t5 224.257
R75 a_492_48.n1 a_492_48.t6 188.517
R76 a_492_48.n4 a_492_48.t2 186.537
R77 a_492_48.n1 a_492_48.n0 171.275
R78 a_492_48.n5 a_492_48.n4 152
R79 a_492_48.n2 a_492_48.t7 149.421
R80 a_492_48.n3 a_492_48.t0 114.453
R81 a_492_48.n5 a_492_48.n3 62.6504
R82 a_492_48.n2 a_492_48.n1 10.2247
R83 VGND.n38 VGND.n37 211.183
R84 VGND.n10 VGND.n9 210.852
R85 VGND.n23 VGND.n6 198.941
R86 VGND.n11 VGND.t7 126.504
R87 VGND.n12 VGND.n11 120.123
R88 VGND.n9 VGND.t3 104.062
R89 VGND.n37 VGND.t0 103.126
R90 VGND.n6 VGND.t6 56.2505
R91 VGND.n6 VGND.t1 48.9111
R92 VGND.n11 VGND.t5 38.2907
R93 VGND.n13 VGND.n8 36.1417
R94 VGND.n17 VGND.n8 36.1417
R95 VGND.n18 VGND.n17 36.1417
R96 VGND.n19 VGND.n18 36.1417
R97 VGND.n19 VGND.n5 36.1417
R98 VGND.n25 VGND.n24 36.1417
R99 VGND.n25 VGND.n3 36.1417
R100 VGND.n29 VGND.n3 36.1417
R101 VGND.n30 VGND.n29 36.1417
R102 VGND.n31 VGND.n30 36.1417
R103 VGND.n31 VGND.n1 36.1417
R104 VGND.n35 VGND.n1 36.1417
R105 VGND.n36 VGND.n35 36.1417
R106 VGND.n9 VGND.t2 33.1513
R107 VGND.n24 VGND.n23 32.0005
R108 VGND.n37 VGND.t4 30.6984
R109 VGND.n13 VGND.n12 22.9652
R110 VGND.n38 VGND.n36 18.824
R111 VGND.n36 VGND.n0 9.3005
R112 VGND.n35 VGND.n34 9.3005
R113 VGND.n33 VGND.n1 9.3005
R114 VGND.n32 VGND.n31 9.3005
R115 VGND.n30 VGND.n2 9.3005
R116 VGND.n29 VGND.n28 9.3005
R117 VGND.n27 VGND.n3 9.3005
R118 VGND.n26 VGND.n25 9.3005
R119 VGND.n24 VGND.n4 9.3005
R120 VGND.n23 VGND.n22 9.3005
R121 VGND.n21 VGND.n5 9.3005
R122 VGND.n20 VGND.n19 9.3005
R123 VGND.n18 VGND.n7 9.3005
R124 VGND.n17 VGND.n16 9.3005
R125 VGND.n15 VGND.n8 9.3005
R126 VGND.n14 VGND.n13 9.3005
R127 VGND.n39 VGND.n38 7.44972
R128 VGND.n12 VGND.n10 7.14797
R129 VGND.n23 VGND.n5 2.25932
R130 VGND VGND.n39 0.160299
R131 VGND.n14 VGND.n10 0.157483
R132 VGND.n39 VGND.n0 0.147507
R133 VGND.n15 VGND.n14 0.122949
R134 VGND.n16 VGND.n15 0.122949
R135 VGND.n16 VGND.n7 0.122949
R136 VGND.n20 VGND.n7 0.122949
R137 VGND.n21 VGND.n20 0.122949
R138 VGND.n22 VGND.n21 0.122949
R139 VGND.n22 VGND.n4 0.122949
R140 VGND.n26 VGND.n4 0.122949
R141 VGND.n27 VGND.n26 0.122949
R142 VGND.n28 VGND.n27 0.122949
R143 VGND.n28 VGND.n2 0.122949
R144 VGND.n32 VGND.n2 0.122949
R145 VGND.n33 VGND.n32 0.122949
R146 VGND.n34 VGND.n33 0.122949
R147 VGND.n34 VGND.n0 0.122949
R148 a_1197_368.n0 a_1197_368.t1 790.404
R149 a_1197_368.n0 a_1197_368.t0 66.8398
R150 a_1197_368.t2 a_1197_368.n0 30.7494
R151 VNB.t13 VNB.t7 4607.87
R152 VNB.t1 VNB.t12 2598.43
R153 VNB.t3 VNB.t2 2436.75
R154 VNB.t5 VNB.t4 2309.71
R155 VNB.t6 VNB.t9 2182.68
R156 VNB.t8 VNB.t1 2101.84
R157 VNB.t10 VNB.t14 2044.09
R158 VNB.t2 VNB.t13 1686.09
R159 VNB.t0 VNB.t11 1570.6
R160 VNB.t11 VNB.t3 1524.41
R161 VNB.t9 VNB.t5 1328.08
R162 VNB.t7 VNB.t10 1154.86
R163 VNB VNB.t8 1154.86
R164 VNB.t14 VNB.t6 1097.11
R165 VNB.t12 VNB.t0 993.177
R166 COUT.n2 COUT.t0 496.632
R167 COUT.n3 COUT.n1 185
R168 COUT.n6 COUT.n1 185
R169 COUT.n1 COUT.n0 185
R170 COUT.n4 COUT.n1 185
R171 COUT.n5 COUT.n3 185
R172 COUT.n6 COUT.n5 185
R173 COUT.n5 COUT.n0 185
R174 COUT.n5 COUT.n4 185
R175 COUT.t1 COUT.n1 14.8415
R176 COUT.n5 COUT.t1 13.9934
R177 COUT COUT.n0 7.5161
R178 COUT.n6 COUT.n2 7.1638
R179 COUT COUT.n6 4.58032
R180 COUT COUT.n0 3.7583
R181 COUT.n3 COUT.n2 1.17481
R182 COUT.n4 COUT 0.822518
R183 a_1595_400.n1 a_1595_400.n0 466.841
R184 a_1595_400.n2 a_1595_400.n1 40.6504
R185 a_1595_400.n0 a_1595_400.t0 39.3755
R186 a_1595_400.n1 a_1595_400.t2 38.1157
R187 a_1595_400.n0 a_1595_400.t1 26.2505
R188 VPWR.n26 VPWR.n7 603.312
R189 VPWR.n14 VPWR.n13 336.709
R190 VPWR.n12 VPWR.n11 239.141
R191 VPWR.n40 VPWR.n1 231.048
R192 VPWR.n13 VPWR.t7 79.7855
R193 VPWR.n1 VPWR.t4 76.8305
R194 VPWR.n11 VPWR.t2 74.8605
R195 VPWR.n7 VPWR.t6 49.2505
R196 VPWR.n14 VPWR.n12 37.0149
R197 VPWR.n28 VPWR.n27 36.1417
R198 VPWR.n28 VPWR.n4 36.1417
R199 VPWR.n32 VPWR.n4 36.1417
R200 VPWR.n33 VPWR.n32 36.1417
R201 VPWR.n34 VPWR.n33 36.1417
R202 VPWR.n34 VPWR.n2 36.1417
R203 VPWR.n38 VPWR.n2 36.1417
R204 VPWR.n39 VPWR.n38 36.1417
R205 VPWR.n15 VPWR.n10 36.1417
R206 VPWR.n19 VPWR.n10 36.1417
R207 VPWR.n20 VPWR.n19 36.1417
R208 VPWR.n21 VPWR.n20 36.1417
R209 VPWR.n21 VPWR.n8 36.1417
R210 VPWR.n25 VPWR.n8 36.1417
R211 VPWR.n7 VPWR.t3 29.1741
R212 VPWR.n40 VPWR.n39 28.2358
R213 VPWR.n27 VPWR.n26 27.4829
R214 VPWR.n1 VPWR.t5 27.0196
R215 VPWR.n13 VPWR.t0 26.8503
R216 VPWR.n11 VPWR.t1 26.8503
R217 VPWR.n26 VPWR.n25 17.6946
R218 VPWR.n16 VPWR.n15 9.3005
R219 VPWR.n17 VPWR.n10 9.3005
R220 VPWR.n19 VPWR.n18 9.3005
R221 VPWR.n20 VPWR.n9 9.3005
R222 VPWR.n22 VPWR.n21 9.3005
R223 VPWR.n23 VPWR.n8 9.3005
R224 VPWR.n25 VPWR.n24 9.3005
R225 VPWR.n26 VPWR.n6 9.3005
R226 VPWR.n27 VPWR.n5 9.3005
R227 VPWR.n29 VPWR.n28 9.3005
R228 VPWR.n30 VPWR.n4 9.3005
R229 VPWR.n32 VPWR.n31 9.3005
R230 VPWR.n33 VPWR.n3 9.3005
R231 VPWR.n35 VPWR.n34 9.3005
R232 VPWR.n36 VPWR.n2 9.3005
R233 VPWR.n38 VPWR.n37 9.3005
R234 VPWR.n39 VPWR.n0 9.3005
R235 VPWR.n41 VPWR.n40 7.30699
R236 VPWR.n15 VPWR.n14 6.77697
R237 VPWR VPWR.n41 0.158419
R238 VPWR.n16 VPWR.n12 0.149714
R239 VPWR.n41 VPWR.n0 0.149362
R240 VPWR.n17 VPWR.n16 0.122949
R241 VPWR.n18 VPWR.n17 0.122949
R242 VPWR.n18 VPWR.n9 0.122949
R243 VPWR.n22 VPWR.n9 0.122949
R244 VPWR.n23 VPWR.n22 0.122949
R245 VPWR.n24 VPWR.n23 0.122949
R246 VPWR.n24 VPWR.n6 0.122949
R247 VPWR.n6 VPWR.n5 0.122949
R248 VPWR.n29 VPWR.n5 0.122949
R249 VPWR.n30 VPWR.n29 0.122949
R250 VPWR.n31 VPWR.n30 0.122949
R251 VPWR.n31 VPWR.n3 0.122949
R252 VPWR.n35 VPWR.n3 0.122949
R253 VPWR.n36 VPWR.n35 0.122949
R254 VPWR.n37 VPWR.n36 0.122949
R255 VPWR.n37 VPWR.n0 0.122949
R256 B.n1 B.n0 708.54
R257 B.n2 B.t2 570.367
R258 B.n3 B.n2 546.534
R259 B.n0 B.t3 541.715
R260 B.n1 B.t0 332.58
R261 B.n0 B.t4 250.105
R262 B.n1 B.t1 225.202
R263 B.n2 B.t5 212.081
R264 B B.n3 160.145
R265 B.n3 B.n1 14.7283
R266 a_256_368.t1 a_256_368.n4 822.068
R267 a_256_368.t1 a_256_368.n3 738.593
R268 a_256_368.n2 a_256_368.n0 398.425
R269 a_256_368.n2 a_256_368.n1 288.375
R270 a_256_368.n4 a_256_368.t0 269.396
R271 a_256_368.n3 a_256_368.n2 72.0832
R272 a_256_368.n0 a_256_368.t5 69.3755
R273 a_256_368.n1 a_256_368.t3 44.56
R274 a_256_368.n1 a_256_368.t4 35.1791
R275 a_256_368.n0 a_256_368.t2 26.2505
R276 a_256_368.n4 a_256_368.n3 15.2821
R277 A.n0 A.t1 244.482
R278 A.n0 A.t0 213.688
R279 A A.n0 154.233
R280 a_28_74.n2 a_28_74.n0 909.861
R281 a_28_74.n4 a_28_74.n3 347.522
R282 a_28_74.t1 a_28_74.n5 276.291
R283 a_28_74.n1 a_28_74.t7 242.411
R284 a_28_74.n1 a_28_74.t6 185.375
R285 a_28_74.n2 a_28_74.n1 152
R286 a_28_74.n5 a_28_74.t0 149.143
R287 a_28_74.n0 a_28_74.t5 85.6017
R288 a_28_74.n0 a_28_74.t2 46.9053
R289 a_28_74.n5 a_28_74.n4 41.7887
R290 a_28_74.n3 a_28_74.t4 26.2505
R291 a_28_74.n3 a_28_74.t3 26.2505
R292 a_28_74.n4 a_28_74.n2 14.0075
R293 CIN.n0 CIN.t1 283.041
R294 CIN.n1 CIN.t0 255.419
R295 CIN.n0 CIN.t2 202.44
R296 CIN CIN.n2 156.268
R297 CIN.n1 CIN.t3 138.173
R298 CIN.n2 CIN.n0 42.8861
R299 CIN.n2 CIN.n1 35.2236
R300 SUM.n2 SUM 591.4
R301 SUM.n2 SUM.n1 585
R302 SUM.n3 SUM.n2 585
R303 SUM.n4 SUM.t0 279.738
R304 SUM.t0 SUM.n0 273.421
R305 SUM.n2 SUM.t1 26.3844
R306 SUM.n3 SUM 17.1525
R307 SUM.n1 SUM 14.8485
R308 SUM SUM.n4 13.0565
R309 SUM.n0 SUM 7.3702
R310 SUM SUM.n0 6.98232
R311 SUM.n4 SUM 5.8885
R312 SUM.n1 SUM 4.0965
R313 SUM SUM.n3 1.7925
C0 B CIN 9.83e-19
C1 VPWR CIN 0.020973f
C2 B COUT 0.001694f
C3 A VGND 0.017779f
C4 B VGND 0.072031f
C5 VPWR COUT 0.017192f
C6 VPWR VGND 0.068676f
C7 B SUM 4.08e-20
C8 CIN COUT 3.78e-19
C9 A VPB 0.04646f
C10 CIN VGND 0.057073f
C11 VPWR SUM 0.11908f
C12 B VPB 0.405813f
C13 COUT VGND 0.119427f
C14 CIN SUM 2.7e-20
C15 VPWR VPB 0.282215f
C16 CIN VPB 0.09758f
C17 VGND SUM 0.064496f
C18 COUT VPB 0.008106f
C19 A B 2.03e-19
C20 VGND VPB 0.0166f
C21 A VPWR 0.04892f
C22 SUM VPB 0.013084f
C23 B VPWR 0.063608f
C24 SUM VNB 0.106358f
C25 VGND VNB 1.44768f
C26 COUT VNB 0.028588f
C27 CIN VNB 0.265737f
C28 VPWR VNB 1.138f
C29 B VNB 0.676278f
C30 A VNB 0.151477f
C31 VPB VNB 2.97749f
.ends

* NGSPICE file created from sky130_fd_sc_hs__fahcon_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fahcon_1 VNB VPB VPWR VGND CI B A SUM COUT_N
X0 a_1261_421.t1 a_369_365.t4 COUT_N.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.4706 pd=2.07 as=0.2121 ps=1.345 w=0.84 l=0.15
X1 SUM.t1 a_1744_94.t3 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.29915 ps=1.69 w=0.74 l=0.15
X2 a_241_368.t2 B.t0 a_374_120.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2436 pd=2.26 as=0.2114 ps=1.43 w=0.84 l=0.15
X3 a_241_368.t1 B.t1 a_369_365.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1456 ps=1.095 w=0.64 l=0.15
X4 a_27_100.t1 B.t2 a_374_120.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.150225 ps=1.145 w=0.64 l=0.15
X5 a_1744_94.t2 a_369_365.t5 a_1719_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.4033 ps=3.02 w=0.84 l=0.15
X6 VPWR.t5 A.t0 a_27_100.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 a_241_368.t4 a_27_100.t6 VGND.t6 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.24615 ps=1.46 w=0.64 l=0.15
X8 a_1719_368.t3 a_374_120.t4 a_1744_94.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1632 pd=1.15 as=0.2112 ps=1.3 w=0.64 l=0.15
X9 VGND.t5 A.t1 a_27_100.t4 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.24615 pd=1.46 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 a_1606_368.t2 CI.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1934 ps=1.475 w=1.12 l=0.15
X11 a_1261_421.t0 a_374_120.t5 COUT_N.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.176 pd=1.19 as=0.1792 ps=1.2 w=0.64 l=0.15
X12 a_369_365.t0 a_336_263.t2 a_241_368.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.26 as=0.229925 ps=1.505 w=0.84 l=0.15
X13 SUM.t0 a_1744_94.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1934 ps=1.475 w=1.12 l=0.15
X14 COUT_N.t3 a_369_365.t6 a_1023_389.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1792 pd=1.2 as=0.2496 ps=1.42 w=0.64 l=0.15
X15 a_1606_368.t1 CI.t1 VGND.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.1277 ps=1.1 w=0.74 l=0.15
X16 a_374_120.t3 a_336_263.t3 a_27_100.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2114 pd=1.43 as=0.126 ps=1.14 w=0.84 l=0.15
X17 a_27_100.t0 B.t3 a_369_365.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1764 ps=1.26 w=0.84 l=0.15
X18 VPWR.t6 CI.t2 a_1261_421.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.4706 ps=2.07 w=1 l=0.15
X19 a_374_120.t0 a_336_263.t4 a_241_368.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.150225 pd=1.145 as=0.0896 ps=0.92 w=0.64 l=0.15
X20 a_1744_94.t1 a_369_365.t7 a_1606_368.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2112 pd=1.3 as=0.12945 ps=1.1 w=0.64 l=0.15
X21 a_1023_389.t0 B.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2496 pd=1.42 as=0.1165 ps=1.065 w=0.64 l=0.15
X22 VPWR.t7 a_1606_368.t3 a_1719_368.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.295 ps=2.59 w=1 l=0.15
X23 VPWR.t0 B.t5 a_336_263.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2482 pd=1.575 as=0.3304 ps=2.83 w=1.12 l=0.15
X24 a_369_365.t3 a_336_263.t5 a_27_100.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1456 pd=1.095 as=0.0928 ps=0.93 w=0.64 l=0.15
X25 VGND.t4 B.t6 a_336_263.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.4662 ps=2.74 w=0.74 l=0.15
X26 VGND.t7 a_1606_368.t4 a_1719_368.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.29915 pd=1.69 as=0.1632 ps=1.15 w=0.64 l=0.15
X27 a_1023_389.t1 B.t7 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1853 pd=1.385 as=0.2482 ps=1.575 w=1 l=0.15
X28 a_241_368.t5 a_27_100.t7 VPWR.t4 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.229925 pd=1.505 as=0.2382 ps=1.555 w=1 l=0.15
X29 COUT_N.t1 a_374_120.t6 a_1023_389.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2121 pd=1.345 as=0.1853 ps=1.385 w=0.84 l=0.15
X30 VGND.t2 CI.t3 a_1261_421.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1277 pd=1.1 as=0.176 ps=1.19 w=0.64 l=0.15
R0 a_369_365.n5 a_369_365.n4 674.771
R1 a_369_365.n2 a_369_365.t6 293.269
R2 a_369_365.n1 a_369_365.t5 278.245
R3 a_369_365.n2 a_369_365.t4 216.149
R4 a_369_365.n1 a_369_365.t7 187.981
R5 a_369_365.n3 a_369_365.n1 179.982
R6 a_369_365.n3 a_369_365.n2 163.715
R7 a_369_365.n4 a_369_365.n0 115.66
R8 a_369_365.t0 a_369_365.n5 63.3219
R9 a_369_365.n0 a_369_365.t1 45.938
R10 a_369_365.n0 a_369_365.t3 39.3755
R11 a_369_365.n5 a_369_365.t2 35.1791
R12 a_369_365.n4 a_369_365.n3 12.1992
R13 COUT_N.n2 COUT_N.n0 396.844
R14 COUT_N.n2 COUT_N.n1 89.2272
R15 COUT_N.n0 COUT_N.t1 71.5303
R16 COUT_N.n1 COUT_N.t0 68.438
R17 COUT_N.n0 COUT_N.t2 46.9053
R18 COUT_N.n1 COUT_N.t3 36.563
R19 COUT_N COUT_N.n2 8.29409
R20 a_1261_421.n1 a_1261_421.n0 257.247
R21 a_1261_421.n1 a_1261_421.t1 105.775
R22 a_1261_421.n0 a_1261_421.t0 76.8755
R23 a_1261_421.n2 a_1261_421.n1 71.5237
R24 a_1261_421.n3 a_1261_421.n2 55.7552
R25 a_1261_421.n0 a_1261_421.t2 26.2505
R26 a_1261_421.n2 a_1261_421.t3 26.2144
R27 VPB VPB.n1 633.333
R28 VPB.t10 VPB.t5 524.4
R29 VPB.t9 VPB.t10 309.067
R30 VPB.t5 VPB.n0 304
R31 VPB.t11 VPB.t8 298.791
R32 VPB.t0 VPB.t4 288.8
R33 VPB.t8 VPB 278.361
R34 VPB.n1 VPB.t0 263.467
R35 VPB.t4 VPB.t9 228
R36 VPB.n0 VPB 70.4499
R37 VPB.n1 VPB.t11 61.2908
R38 VPB.t3 VPB.t2 19.9256
R39 VPB.n0 VPB.t1 9.25144
R40 VPB.t7 VPB.t1 9.25144
R41 VPB.t6 VPB.t3 6.40499
R42 VPB.n0 VPB.t6 2.53383
R43 VPB.t6 VPB.t7 2.13533
R44 a_1744_94.t2 a_1744_94.n2 842.13
R45 a_1744_94.n2 a_1744_94.n0 364.485
R46 a_1744_94.n0 a_1744_94.t4 264.298
R47 a_1744_94.n0 a_1744_94.t3 204.048
R48 a_1744_94.n2 a_1744_94.n1 89.2272
R49 a_1744_94.n1 a_1744_94.t0 82.5005
R50 a_1744_94.n1 a_1744_94.t1 41.2505
R51 VGND.n13 VGND.n12 235.595
R52 VGND.n36 VGND.n1 220.608
R53 VGND.n22 VGND.n7 218.536
R54 VGND.n11 VGND.n10 122.118
R55 VGND.n1 VGND.t6 105.939
R56 VGND.n12 VGND.t7 101.251
R57 VGND.n10 VGND.t2 39.3755
R58 VGND.n37 VGND.n36 38.6652
R59 VGND.n16 VGND.n9 36.1417
R60 VGND.n17 VGND.n16 36.1417
R61 VGND.n18 VGND.n17 36.1417
R62 VGND.n18 VGND.n6 36.1417
R63 VGND.n24 VGND.n23 36.1417
R64 VGND.n24 VGND.n4 36.1417
R65 VGND.n28 VGND.n4 36.1417
R66 VGND.n29 VGND.n28 36.1417
R67 VGND.n30 VGND.n29 36.1417
R68 VGND.n30 VGND.n2 36.1417
R69 VGND.n34 VGND.n2 36.1417
R70 VGND.n35 VGND.n34 36.1417
R71 VGND.n7 VGND.t4 31.0986
R72 VGND.n22 VGND.n6 27.4829
R73 VGND.n12 VGND.t3 26.548
R74 VGND.n7 VGND.t0 26.2505
R75 VGND.n23 VGND.n22 25.977
R76 VGND.n10 VGND.t1 24.5361
R77 VGND.n11 VGND.n9 22.9652
R78 VGND.n1 VGND.t5 22.6604
R79 VGND.n14 VGND.n9 9.3005
R80 VGND.n16 VGND.n15 9.3005
R81 VGND.n17 VGND.n8 9.3005
R82 VGND.n19 VGND.n18 9.3005
R83 VGND.n20 VGND.n6 9.3005
R84 VGND.n22 VGND.n21 9.3005
R85 VGND.n23 VGND.n5 9.3005
R86 VGND.n25 VGND.n24 9.3005
R87 VGND.n26 VGND.n4 9.3005
R88 VGND.n28 VGND.n27 9.3005
R89 VGND.n29 VGND.n3 9.3005
R90 VGND.n31 VGND.n30 9.3005
R91 VGND.n32 VGND.n2 9.3005
R92 VGND.n34 VGND.n33 9.3005
R93 VGND.n35 VGND.n0 9.3005
R94 VGND.n13 VGND.n11 7.45414
R95 VGND.n36 VGND.n35 6.77697
R96 VGND.n14 VGND.n13 0.153023
R97 VGND.n15 VGND.n14 0.122949
R98 VGND.n15 VGND.n8 0.122949
R99 VGND.n19 VGND.n8 0.122949
R100 VGND.n20 VGND.n19 0.122949
R101 VGND.n21 VGND.n20 0.122949
R102 VGND.n21 VGND.n5 0.122949
R103 VGND.n25 VGND.n5 0.122949
R104 VGND.n26 VGND.n25 0.122949
R105 VGND.n27 VGND.n26 0.122949
R106 VGND.n27 VGND.n3 0.122949
R107 VGND.n31 VGND.n3 0.122949
R108 VGND.n32 VGND.n31 0.122949
R109 VGND.n33 VGND.n32 0.122949
R110 VGND.n33 VGND.n0 0.122949
R111 VGND.n37 VGND.n0 0.122949
R112 VGND VGND.n37 0.0617245
R113 SUM.n1 SUM 589.444
R114 SUM.n1 SUM.n0 585
R115 SUM.n2 SUM.n1 585
R116 SUM SUM.t1 208.948
R117 SUM.n1 SUM.t0 26.3844
R118 SUM SUM.n2 11.9116
R119 SUM SUM.n0 10.3116
R120 SUM SUM.n0 2.84494
R121 SUM.n2 SUM 1.24494
R122 VNB VNB.n0 11629.4
R123 VNB.t1 VNB.t5 2148.03
R124 VNB.t12 VNB.t9 2101.84
R125 VNB.t4 VNB.t2 1870.87
R126 VNB.t5 VNB.t3 1639.9
R127 VNB.t3 VNB.t8 1616.8
R128 VNB.t2 VNB.t12 1524.41
R129 VNB.t7 VNB.t4 1177.95
R130 VNB.t8 VNB.t7 1177.95
R131 VNB.n0 VNB 589.475
R132 VNB.n0 VNB.t1 577.428
R133 VNB.t10 VNB.t11 109.475
R134 VNB.t0 VNB.t6 54.7373
R135 VNB.t11 VNB.t0 42.1058
R136 VNB.n0 VNB.t10 33.6847
R137 B.n2 B.n1 751.92
R138 B.n1 B.t3 540.912
R139 B.t0 B.t1 393.757
R140 B.t3 B.t2 383.88
R141 B.n2 B.t5 277.687
R142 B.n0 B.t7 270.457
R143 B.n1 B.t0 258.139
R144 B.n0 B.t4 233.26
R145 B B.n4 166.703
R146 B.n3 B.t6 154.24
R147 B.n3 B.n2 78.435
R148 B.n4 B.n0 20.449
R149 B.n4 B.n3 13.146
R150 a_374_120.n5 a_374_120.n4 793.299
R151 a_374_120.n0 a_374_120.t6 488.851
R152 a_374_120.n0 a_374_120.t5 280.911
R153 a_374_120.n3 a_374_120.n2 227.71
R154 a_374_120.n0 a_374_120.n3 200.861
R155 a_374_120.n3 a_374_120.t4 172.816
R156 a_374_120.n4 a_374_120.n1 92.1043
R157 a_374_120.t2 a_374_120.n5 53.941
R158 a_374_120.n5 a_374_120.t3 53.941
R159 a_374_120.n1 a_374_120.t0 34.2897
R160 a_374_120.n1 a_374_120.t1 33.7396
R161 a_374_120.n4 a_374_120.n0 17.2076
R162 a_241_368.n5 a_241_368.n4 585
R163 a_241_368.n1 a_241_368.t2 380.942
R164 a_241_368.n3 a_241_368.n0 289.24
R165 a_241_368.n4 a_241_368.n1 184.631
R166 a_241_368.n1 a_241_368.t1 172.018
R167 a_241_368.n3 a_241_368.n2 149.755
R168 a_241_368.n0 a_241_368.t3 78.0706
R169 a_241_368.n6 a_241_368.n5 36.7293
R170 a_241_368.n0 a_241_368.t5 29.861
R171 a_241_368.n2 a_241_368.t0 26.2505
R172 a_241_368.n2 a_241_368.t4 26.2505
R173 a_241_368.n5 a_241_368.n0 21.2283
R174 a_241_368.n4 a_241_368.n3 19.7093
R175 a_1606_368.n1 a_1606_368.t3 340.37
R176 a_1606_368.n2 a_1606_368.n1 288.882
R177 a_1606_368.t2 a_1606_368.n2 219.55
R178 a_1606_368.n1 a_1606_368.t4 175.127
R179 a_1606_368.n2 a_1606_368.n0 171.671
R180 a_1606_368.n0 a_1606_368.t0 41.2505
R181 a_1606_368.n0 a_1606_368.t1 21.3263
R182 a_27_100.n3 a_27_100.n1 623.174
R183 a_27_100.t3 a_27_100.n5 295.327
R184 a_27_100.n0 a_27_100.t7 222.677
R185 a_27_100.n4 a_27_100.n3 182.959
R186 a_27_100.n4 a_27_100.n0 179.161
R187 a_27_100.n0 a_27_100.t6 153.322
R188 a_27_100.n5 a_27_100.t4 137.47
R189 a_27_100.n3 a_27_100.n2 89.3175
R190 a_27_100.n5 a_27_100.n4 39.0405
R191 a_27_100.n1 a_27_100.t5 35.1791
R192 a_27_100.n1 a_27_100.t0 35.1791
R193 a_27_100.n2 a_27_100.t1 28.1255
R194 a_27_100.n2 a_27_100.t2 26.2505
R195 a_1719_368.n1 a_1719_368.t0 1028.62
R196 a_1719_368.n1 a_1719_368.n0 326.404
R197 a_1719_368.t2 a_1719_368.n1 216.885
R198 a_1719_368.n0 a_1719_368.t3 69.3755
R199 a_1719_368.n0 a_1719_368.t1 26.2505
R200 A.n0 A.t0 250.909
R201 A.n0 A.t1 178.34
R202 A A.n0 154.828
R203 VPWR.n12 VPWR.n11 332.481
R204 VPWR.n10 VPWR.n9 241.621
R205 VPWR.n22 VPWR.n6 224.279
R206 VPWR.n34 VPWR.n1 222.359
R207 VPWR.n6 VPWR.t1 50.2355
R208 VPWR.n1 VPWR.t4 46.2955
R209 VPWR.n9 VPWR.t6 40.3855
R210 VPWR.n11 VPWR.t3 38.3857
R211 VPWR.n26 VPWR.n4 36.1417
R212 VPWR.n27 VPWR.n26 36.1417
R213 VPWR.n28 VPWR.n27 36.1417
R214 VPWR.n28 VPWR.n2 36.1417
R215 VPWR.n32 VPWR.n2 36.1417
R216 VPWR.n33 VPWR.n32 36.1417
R217 VPWR.n15 VPWR.n14 36.1417
R218 VPWR.n16 VPWR.n15 36.1417
R219 VPWR.n16 VPWR.n7 36.1417
R220 VPWR.n20 VPWR.n7 36.1417
R221 VPWR.n21 VPWR.n20 36.1417
R222 VPWR.n1 VPWR.t5 35.4615
R223 VPWR.n6 VPWR.t0 35.4615
R224 VPWR.n22 VPWR.n4 35.0123
R225 VPWR.n11 VPWR.t7 29.5505
R226 VPWR.n9 VPWR.t2 27.5507
R227 VPWR.n12 VPWR.n10 21.9561
R228 VPWR.n14 VPWR.n10 21.8358
R229 VPWR.n34 VPWR.n33 16.1887
R230 VPWR.n22 VPWR.n21 12.424
R231 VPWR.n14 VPWR.n13 9.3005
R232 VPWR.n15 VPWR.n8 9.3005
R233 VPWR.n17 VPWR.n16 9.3005
R234 VPWR.n18 VPWR.n7 9.3005
R235 VPWR.n20 VPWR.n19 9.3005
R236 VPWR.n21 VPWR.n5 9.3005
R237 VPWR.n23 VPWR.n22 9.3005
R238 VPWR.n24 VPWR.n4 9.3005
R239 VPWR.n26 VPWR.n25 9.3005
R240 VPWR.n27 VPWR.n3 9.3005
R241 VPWR.n29 VPWR.n28 9.3005
R242 VPWR.n30 VPWR.n2 9.3005
R243 VPWR.n32 VPWR.n31 9.3005
R244 VPWR.n33 VPWR.n0 9.3005
R245 VPWR.n35 VPWR.n34 7.54736
R246 VPWR VPWR.n35 0.161584
R247 VPWR.n13 VPWR.n12 0.149745
R248 VPWR.n35 VPWR.n0 0.146238
R249 VPWR.n13 VPWR.n8 0.122949
R250 VPWR.n17 VPWR.n8 0.122949
R251 VPWR.n18 VPWR.n17 0.122949
R252 VPWR.n19 VPWR.n18 0.122949
R253 VPWR.n19 VPWR.n5 0.122949
R254 VPWR.n23 VPWR.n5 0.122949
R255 VPWR.n24 VPWR.n23 0.122949
R256 VPWR.n25 VPWR.n24 0.122949
R257 VPWR.n25 VPWR.n3 0.122949
R258 VPWR.n29 VPWR.n3 0.122949
R259 VPWR.n30 VPWR.n29 0.122949
R260 VPWR.n31 VPWR.n30 0.122949
R261 VPWR.n31 VPWR.n0 0.122949
R262 CI.n1 CI.t2 337.546
R263 CI.n0 CI.t0 264.832
R264 CI.n0 CI.t1 203.756
R265 CI.n1 CI.t3 170.308
R266 CI CI.n2 158.788
R267 CI.n2 CI.n1 31.4035
R268 CI.n2 CI.n0 14.6066
R269 a_336_263.n0 a_336_263.t4 530.157
R270 a_336_263.t4 a_336_263.t2 400.356
R271 a_336_263.t5 a_336_263.t3 381.048
R272 a_336_263.t1 a_336_263.n1 302.466
R273 a_336_263.n1 a_336_263.n0 234.565
R274 a_336_263.n0 a_336_263.t5 159.963
R275 a_336_263.n1 a_336_263.t0 81.3655
R276 a_1023_389.n1 a_1023_389.n0 388.252
R277 a_1023_389.n0 a_1023_389.t2 68.3447
R278 a_1023_389.n0 a_1023_389.t0 60.8835
R279 a_1023_389.n1 a_1023_389.t3 55.1136
R280 a_1023_389.t1 a_1023_389.n1 30.7494
C0 COUT_N VGND 0.041359f
C1 CI SUM 1.8e-20
C2 B VGND 0.052336f
C3 B SUM 5.35e-20
C4 VPB VPWR 0.281584f
C5 VGND SUM 0.038108f
C6 VPB CI 0.088204f
C7 A VPWR 0.038539f
C8 VPB COUT_N 0.012142f
C9 VPB B 0.460373f
C10 VPB VGND 0.00937f
C11 A B 0.001178f
C12 VPB SUM 0.014597f
C13 A VGND 0.015002f
C14 VPWR CI 0.031389f
C15 VPWR COUT_N 0.042787f
C16 B VPWR 0.123175f
C17 VPWR VGND 0.0685f
C18 VPB A 0.040695f
C19 B CI 7.09e-20
C20 CI VGND 0.052394f
C21 VPWR SUM 0.114949f
C22 B COUT_N 0.00104f
C23 SUM VNB 0.113646f
C24 VGND VNB 1.28532f
C25 COUT_N VNB 0.017905f
C26 CI VNB 0.230765f
C27 VPWR VNB 1.03358f
C28 B VNB 0.529991f
C29 A VNB 0.125928f
C30 VPB VNB 2.66289f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkdlyinv3sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkdlyinv3sd2_1 VNB VPB VPWR VGND A Y
X0 a_288_74.t1 a_28_74.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X1 Y.t0 a_288_74.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X2 Y.t1 a_288_74.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.308 ps=2.79 w=1.12 l=0.15
X3 VGND.t0 A.t0 a_28_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VPWR.t0 A.t1 a_28_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3284 pd=1.745 as=0.3136 ps=2.8 w=1.12 l=0.15
X5 a_288_74.t0 a_28_74.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3284 ps=1.745 w=1 l=0.25
R0 a_28_74.t0 a_28_74.n1 448.507
R1 a_28_74.n1 a_28_74.t1 289.522
R2 a_28_74.n0 a_28_74.t3 183.161
R3 a_28_74.n0 a_28_74.t2 163.185
R4 a_28_74.n1 a_28_74.n0 152
R5 VGND.n1 VGND.t2 253.761
R6 VGND.n1 VGND.n0 212.68
R7 VGND.n0 VGND.t1 145.714
R8 VGND.n0 VGND.t0 55.7148
R9 VGND VGND.n1 0.263065
R10 a_288_74.n0 a_288_74.t3 265.637
R11 a_288_74.n1 a_288_74.t1 262.938
R12 a_288_74.n0 a_288_74.t2 253.853
R13 a_288_74.t0 a_288_74.n1 253.458
R14 a_288_74.n1 a_288_74.n0 177.794
R15 VNB.t1 VNB.t2 2228.87
R16 VNB.t0 VNB.t1 2009.45
R17 VNB VNB.t0 1108.66
R18 Y.n1 Y 589.268
R19 Y.n1 Y.n0 585
R20 Y.n2 Y.n1 585
R21 Y.n3 Y.t0 225
R22 Y.n1 Y.t1 27.2639
R23 Y.n2 Y 11.9116
R24 Y Y.n3 9.97283
R25 Y.n0 Y 9.24494
R26 Y.n3 Y 4.26717
R27 Y.n0 Y 3.91161
R28 Y Y.n2 1.24494
R29 VPWR.n1 VPWR.n0 321.021
R30 VPWR.n1 VPWR.t2 256.077
R31 VPWR.n0 VPWR.t1 89.6355
R32 VPWR.n0 VPWR.t0 31.6309
R33 VPWR VPWR.n1 0.260042
R34 VPB.t1 VPB.t2 513.307
R35 VPB.t0 VPB.t1 421.372
R36 VPB VPB.t0 252.823
R37 A.n0 A.t1 293.752
R38 A.n0 A.t0 220.113
R39 A A.n0 159.929
C0 VPB Y 0.019107f
C1 Y VGND 0.073742f
C2 VPB VGND 0.006768f
C3 A VPWR 0.021274f
C4 VPB A 0.04065f
C5 A VGND 0.01746f
C6 VPWR Y 0.14736f
C7 VPB VPWR 0.093331f
C8 VPWR VGND 0.049819f
C9 VGND VNB 0.393996f
C10 Y VNB 0.124951f
C11 VPWR VNB 0.311757f
C12 A VNB 0.205416f
C13 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkdlyinv3sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkdlyinv3sd3_1 VNB VPB VPWR VGND A Y
X0 a_288_74.t0 a_28_74.t2 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X1 Y.t1 a_288_74.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X2 Y.t0 a_288_74.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.308 ps=2.79 w=1.12 l=0.15
X3 VGND.t2 A.t0 a_28_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VPWR.t2 A.t1 a_28_74.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2034 pd=1.495 as=0.3136 ps=2.8 w=1.12 l=0.15
X5 a_288_74.t1 a_28_74.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.2034 ps=1.495 w=1 l=0.5
R0 a_28_74.t1 a_28_74.n1 448.507
R1 a_28_74.n1 a_28_74.t0 289.522
R2 a_28_74.n0 a_28_74.t2 163.185
R3 a_28_74.n1 a_28_74.n0 152
R4 a_28_74.n0 a_28_74.t3 112.306
R5 VGND.n1 VGND.t0 253.761
R6 VGND.n1 VGND.n0 212.68
R7 VGND.n0 VGND.t1 145.714
R8 VGND.n0 VGND.t2 55.7148
R9 VGND VGND.n1 0.263065
R10 a_288_74.n0 a_288_74.t3 265.637
R11 a_288_74.t0 a_288_74.n1 262.938
R12 a_288_74.n0 a_288_74.t2 253.853
R13 a_288_74.n1 a_288_74.t1 253.458
R14 a_288_74.n1 a_288_74.n0 177.794
R15 VNB.t0 VNB.t1 2228.87
R16 VNB.t2 VNB.t0 2009.45
R17 VNB VNB.t2 1108.66
R18 Y.n1 Y 589.268
R19 Y.n1 Y.n0 585
R20 Y.n2 Y.n1 585
R21 Y.n3 Y.t1 225
R22 Y.n1 Y.t0 27.2639
R23 Y.n2 Y 11.9116
R24 Y Y.n3 9.97283
R25 Y.n0 Y 9.24494
R26 Y.n3 Y 4.26717
R27 Y.n0 Y 3.91161
R28 Y Y.n2 1.24494
R29 VPWR.n1 VPWR.n0 321.021
R30 VPWR.n1 VPWR.t1 256.077
R31 VPWR.n0 VPWR.t0 40.3855
R32 VPWR.n0 VPWR.t2 31.6309
R33 VPWR VPWR.n1 0.260042
R34 VPB.t0 VPB.t1 577.152
R35 VPB.t2 VPB.t0 357.527
R36 VPB VPB.t2 252.823
R37 A.n0 A.t1 293.752
R38 A.n0 A.t0 220.113
R39 A A.n0 159.929
C0 VPWR Y 0.14736f
C1 A VGND 0.01746f
C2 VPWR VGND 0.048788f
C3 Y VGND 0.073742f
C4 VPB A 0.038386f
C5 VPB VPWR 0.09135f
C6 VPB Y 0.019107f
C7 A VPWR 0.021264f
C8 VPB VGND 0.006575f
C9 VGND VNB 0.393996f
C10 Y VNB 0.124951f
C11 VPWR VNB 0.312379f
C12 A VNB 0.205416f
C13 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkdlyinv5sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkdlyinv5sd1_1 VNB VPB VPWR VGND A Y
X0 VPWR.t2 a_549_74.t2 a_682_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.254 pd=1.595 as=0.61 ps=3.22 w=1 l=0.15
X1 Y.t0 a_682_74.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.254 ps=1.595 w=1.12 l=0.15
X2 a_549_74.t1 a_288_74.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.2604 ps=2.08 w=0.42 l=0.15
X3 a_288_74.t0 a_28_74.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3784 ps=1.845 w=1 l=0.15
X4 VGND.t2 A.t0 a_28_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.15435 pd=1.155 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VGND.t1 a_549_74.t3 a_682_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0966 pd=0.88 as=0.2583 ps=2.07 w=0.42 l=0.15
X6 a_549_74.t0 a_288_74.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.265 pd=2.53 as=0.62 ps=3.24 w=1 l=0.15
X7 Y.t1 a_682_74.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X8 VPWR.t4 A.t1 a_28_74.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3784 pd=1.845 as=0.3136 ps=2.8 w=1.12 l=0.15
X9 a_288_74.t1 a_28_74.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.15435 ps=1.155 w=0.42 l=0.15
R0 a_549_74.n0 a_549_74.t2 366.32
R1 a_549_74.t0 a_549_74.n1 290.661
R2 a_549_74.n1 a_549_74.t1 273.188
R3 a_549_74.n1 a_549_74.n0 245.94
R4 a_549_74.n0 a_549_74.t3 235.922
R5 a_682_74.n1 a_682_74.t1 440.281
R6 a_682_74.t0 a_682_74.n1 405.103
R7 a_682_74.n0 a_682_74.t2 265.637
R8 a_682_74.n0 a_682_74.t3 253.853
R9 a_682_74.n1 a_682_74.n0 152
R10 VPWR.n2 VPWR.t0 318.418
R11 VPWR.n8 VPWR.n1 315.245
R12 VPWR.n4 VPWR.n3 229.972
R13 VPWR.n1 VPWR.t1 109.335
R14 VPWR.n3 VPWR.t2 64.0255
R15 VPWR.n7 VPWR.n6 36.1417
R16 VPWR.n1 VPWR.t4 31.6309
R17 VPWR.n3 VPWR.t3 27.3314
R18 VPWR.n8 VPWR.n7 22.2123
R19 VPWR.n6 VPWR.n2 17.6946
R20 VPWR.n6 VPWR.n5 9.3005
R21 VPWR.n7 VPWR.n0 9.3005
R22 VPWR.n4 VPWR.n2 7.36044
R23 VPWR.n9 VPWR.n8 7.30699
R24 VPWR VPWR.n9 0.158419
R25 VPWR.n5 VPWR.n4 0.15618
R26 VPWR.n9 VPWR.n0 0.149362
R27 VPWR.n5 VPWR.n0 0.122949
R28 VPB.t0 VPB.t2 727.823
R29 VPB.t1 VPB.t0 663.98
R30 VPB.t4 VPB.t1 446.909
R31 VPB.t2 VPB.t3 319.221
R32 VPB VPB.t4 252.823
R33 Y.n1 Y 589.268
R34 Y.n1 Y.n0 585
R35 Y.n2 Y.n1 585
R36 Y.n3 Y.t1 225
R37 Y.n1 Y.t0 27.2639
R38 Y Y.n3 9.97283
R39 Y.n2 Y 9.06717
R40 Y.n0 Y 8.53383
R41 Y.n0 Y 4.62272
R42 Y.n3 Y 4.26717
R43 Y Y.n2 4.08939
R44 a_288_74.n0 a_288_74.t3 334.026
R45 a_288_74.t0 a_288_74.n1 260.805
R46 a_288_74.n1 a_288_74.t1 254.839
R47 a_288_74.n0 a_288_74.t2 195.853
R48 a_288_74.n1 a_288_74.n0 183.613
R49 VGND.n1 VGND.t0 346.212
R50 VGND.n3 VGND.n2 214.043
R51 VGND.n8 VGND.n7 206.916
R52 VGND.n7 VGND.t3 154.286
R53 VGND.n2 VGND.t1 91.4291
R54 VGND.n7 VGND.t2 55.7148
R55 VGND.n2 VGND.t4 40.0005
R56 VGND.n6 VGND.n5 36.1417
R57 VGND.n8 VGND.n6 21.4593
R58 VGND.n5 VGND.n1 17.6946
R59 VGND.n6 VGND.n0 9.3005
R60 VGND.n5 VGND.n4 9.3005
R61 VGND.n3 VGND.n1 7.36044
R62 VGND.n9 VGND.n8 7.34058
R63 VGND VGND.n9 0.158861
R64 VGND.n4 VGND.n3 0.15618
R65 VGND.n9 VGND.n0 0.148926
R66 VGND.n4 VGND.n0 0.122949
R67 VNB.t0 VNB.t1 3302.89
R68 VNB.t3 VNB.t0 3014.17
R69 VNB.t2 VNB.t3 2044.09
R70 VNB.t1 VNB.t4 1408.92
R71 VNB VNB.t2 1108.66
R72 a_28_74.t1 a_28_74.n1 448.507
R73 a_28_74.n0 a_28_74.t2 337.24
R74 a_28_74.n1 a_28_74.t0 289.522
R75 a_28_74.n0 a_28_74.t3 192.639
R76 a_28_74.n1 a_28_74.n0 152
R77 A.n0 A.t1 293.752
R78 A.n0 A.t0 220.113
R79 A A.n0 159.929
C0 VPB Y 0.019328f
C1 A VPWR 0.021277f
C2 VPB VGND 0.013934f
C3 VPWR Y 0.147313f
C4 A VGND 0.017461f
C5 VPWR VGND 0.092753f
C6 Y VGND 0.068148f
C7 VPB A 0.04205f
C8 VPB VPWR 0.171078f
C9 VGND VNB 0.675472f
C10 Y VNB 0.121065f
C11 VPWR VNB 0.525514f
C12 A VNB 0.208436f
C13 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkdlyinv5sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkdlyinv5sd2_1 VNB VPB VPWR VGND A Y
X0 a_288_74.t1 a_28_74.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X1 Y.t1 a_682_74.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.254 ps=1.595 w=1.12 l=0.15
X2 VGND.t4 a_549_74.t2 a_682_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0966 pd=0.88 as=0.2457 ps=2.01 w=0.42 l=0.18
X3 VPWR.t0 a_549_74.t3 a_682_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.254 pd=1.595 as=0.51 ps=3.02 w=1 l=0.25
X4 VGND.t3 A.t0 a_28_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 a_549_74.t0 a_288_74.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.2478 ps=2.02 w=0.42 l=0.18
X6 Y.t0 a_682_74.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X7 VPWR.t4 A.t1 a_28_74.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3284 pd=1.745 as=0.3136 ps=2.8 w=1.12 l=0.15
X8 a_549_74.t1 a_288_74.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.265 pd=2.53 as=0.52 ps=3.04 w=1 l=0.25
X9 a_288_74.t0 a_28_74.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3284 ps=1.745 w=1 l=0.25
R0 a_28_74.t1 a_28_74.n1 448.507
R1 a_28_74.n1 a_28_74.t0 289.522
R2 a_28_74.n0 a_28_74.t3 208.707
R3 a_28_74.n0 a_28_74.t2 163.185
R4 a_28_74.n1 a_28_74.n0 152
R5 VGND.n1 VGND.t2 337.64
R6 VGND.n3 VGND.n2 214.043
R7 VGND.n8 VGND.n7 206.916
R8 VGND.n7 VGND.t1 145.714
R9 VGND.n2 VGND.t4 91.4291
R10 VGND.n7 VGND.t3 55.7148
R11 VGND.n2 VGND.t0 40.0005
R12 VGND.n6 VGND.n5 36.1417
R13 VGND.n8 VGND.n6 21.4593
R14 VGND.n5 VGND.n1 17.6946
R15 VGND.n6 VGND.n0 9.3005
R16 VGND.n5 VGND.n4 9.3005
R17 VGND.n3 VGND.n1 7.36044
R18 VGND.n9 VGND.n8 7.34058
R19 VGND VGND.n9 0.158861
R20 VGND.n4 VGND.n3 0.15618
R21 VGND.n9 VGND.n0 0.148926
R22 VGND.n4 VGND.n0 0.122949
R23 a_288_74.t0 a_288_74.n1 260.805
R24 a_288_74.n1 a_288_74.t1 254.839
R25 a_288_74.n0 a_288_74.t3 206.779
R26 a_288_74.n1 a_288_74.n0 183.613
R27 a_288_74.n0 a_288_74.t2 165.863
R28 VNB.t2 VNB.t4 3302.89
R29 VNB.t1 VNB.t2 3014.17
R30 VNB.t3 VNB.t1 2009.45
R31 VNB.t4 VNB.t0 1443.57
R32 VNB VNB.t3 1108.66
R33 a_682_74.n1 a_682_74.t1 431.709
R34 a_682_74.t0 a_682_74.n1 385.402
R35 a_682_74.n0 a_682_74.t2 265.637
R36 a_682_74.n0 a_682_74.t3 253.853
R37 a_682_74.n1 a_682_74.n0 152
R38 VPWR.n8 VPWR.n1 315.245
R39 VPWR.n2 VPWR.t2 298.717
R40 VPWR.n4 VPWR.n3 229.972
R41 VPWR.n1 VPWR.t1 89.6355
R42 VPWR.n3 VPWR.t0 64.0255
R43 VPWR.n7 VPWR.n6 36.1417
R44 VPWR.n1 VPWR.t4 31.6309
R45 VPWR.n3 VPWR.t3 27.3314
R46 VPWR.n8 VPWR.n7 22.2123
R47 VPWR.n6 VPWR.n2 17.6946
R48 VPWR.n6 VPWR.n5 9.3005
R49 VPWR.n7 VPWR.n0 9.3005
R50 VPWR.n4 VPWR.n2 7.36044
R51 VPWR.n9 VPWR.n8 7.30699
R52 VPWR VPWR.n9 0.158419
R53 VPWR.n5 VPWR.n4 0.15618
R54 VPWR.n9 VPWR.n0 0.149362
R55 VPWR.n5 VPWR.n0 0.122949
R56 Y.n1 Y 589.268
R57 Y.n1 Y.n0 585
R58 Y.n2 Y.n1 585
R59 Y.n3 Y.t0 225
R60 Y.n1 Y.t1 27.2639
R61 Y Y.n3 9.97283
R62 Y.n2 Y 9.06717
R63 Y.n0 Y 8.53383
R64 Y.n0 Y 4.62272
R65 Y.n3 Y 4.26717
R66 Y Y.n2 4.08939
R67 VPB.t2 VPB.t0 727.823
R68 VPB.t1 VPB.t2 663.98
R69 VPB.t4 VPB.t1 421.372
R70 VPB.t0 VPB.t3 344.759
R71 VPB VPB.t4 252.823
R72 a_549_74.t1 a_549_74.n1 290.661
R73 a_549_74.n1 a_549_74.t0 273.188
R74 a_549_74.n1 a_549_74.n0 245.94
R75 a_549_74.n0 a_549_74.t3 225.302
R76 a_549_74.n0 a_549_74.t2 201.266
R77 A.n0 A.t1 293.752
R78 A.n0 A.t0 220.113
R79 A A.n0 159.929
C0 Y VGND 0.068148f
C1 VPWR VPB 0.168162f
C2 VPB A 0.041283f
C3 Y VPB 0.019111f
C4 VPWR A 0.021274f
C5 VPWR Y 0.147313f
C6 VGND VPB 0.013227f
C7 VPWR VGND 0.091457f
C8 VGND A 0.01746f
C9 VGND VNB 0.67447f
C10 Y VNB 0.12103f
C11 VPWR VNB 0.525306f
C12 A VNB 0.20756f
C13 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkdlyinv5sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkdlyinv5sd3_1 VNB VPB VPWR VGND A Y
X0 a_288_74.t1 a_28_74.t2 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.14805 ps=1.125 w=0.42 l=0.18
X1 a_549_74.t0 a_288_74.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.265 pd=2.53 as=0.27 ps=2.54 w=1 l=0.5
X2 Y.t0 a_682_74.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.254 ps=1.595 w=1.12 l=0.15
X3 VGND.t3 a_549_74.t2 a_682_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0966 pd=0.88 as=0.2457 ps=2.01 w=0.42 l=0.18
X4 VGND.t0 A.t0 a_28_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VPWR.t2 a_549_74.t3 a_682_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.254 pd=1.595 as=0.26 ps=2.52 w=1 l=0.5
X6 a_549_74.t1 a_288_74.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.2478 ps=2.02 w=0.42 l=0.18
X7 Y.t1 a_682_74.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X8 VPWR.t3 A.t1 a_28_74.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2034 pd=1.495 as=0.3136 ps=2.8 w=1.12 l=0.15
X9 a_288_74.t0 a_28_74.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.2034 ps=1.495 w=1 l=0.5
R0 a_28_74.t1 a_28_74.n1 448.507
R1 a_28_74.n1 a_28_74.t0 289.522
R2 a_28_74.n0 a_28_74.t2 163.185
R3 a_28_74.n1 a_28_74.n0 152
R4 a_28_74.n0 a_28_74.t3 112.306
R5 VGND.n1 VGND.t1 337.64
R6 VGND.n3 VGND.n2 214.043
R7 VGND.n8 VGND.n7 206.916
R8 VGND.n7 VGND.t2 145.714
R9 VGND.n2 VGND.t3 91.4291
R10 VGND.n7 VGND.t0 55.7148
R11 VGND.n2 VGND.t4 40.0005
R12 VGND.n6 VGND.n5 36.1417
R13 VGND.n8 VGND.n6 21.4593
R14 VGND.n5 VGND.n1 17.6946
R15 VGND.n6 VGND.n0 9.3005
R16 VGND.n5 VGND.n4 9.3005
R17 VGND.n3 VGND.n1 7.36044
R18 VGND.n9 VGND.n8 7.34058
R19 VGND VGND.n9 0.158861
R20 VGND.n4 VGND.n3 0.15618
R21 VGND.n9 VGND.n0 0.148926
R22 VGND.n4 VGND.n0 0.122949
R23 a_288_74.n1 a_288_74.t0 260.807
R24 a_288_74.t1 a_288_74.n1 254.839
R25 a_288_74.n1 a_288_74.n0 183.613
R26 a_288_74.n0 a_288_74.t3 165.863
R27 a_288_74.n0 a_288_74.t2 111.343
R28 VNB.t2 VNB.t3 3302.89
R29 VNB.t1 VNB.t2 3014.17
R30 VNB.t0 VNB.t1 2009.45
R31 VNB.t3 VNB.t4 1443.57
R32 VNB VNB.t0 1108.66
R33 VPWR.n8 VPWR.n1 315.245
R34 VPWR.n2 VPWR.t1 249.468
R35 VPWR.n4 VPWR.n3 229.972
R36 VPWR.n3 VPWR.t2 64.0255
R37 VPWR.n1 VPWR.t0 40.3855
R38 VPWR.n7 VPWR.n6 36.1417
R39 VPWR.n1 VPWR.t3 31.6309
R40 VPWR.n3 VPWR.t4 27.3314
R41 VPWR.n8 VPWR.n7 22.2123
R42 VPWR.n6 VPWR.n2 17.6946
R43 VPWR.n6 VPWR.n5 9.3005
R44 VPWR.n7 VPWR.n0 9.3005
R45 VPWR.n4 VPWR.n2 7.36044
R46 VPWR.n9 VPWR.n8 7.30699
R47 VPWR VPWR.n9 0.158419
R48 VPWR.n5 VPWR.n4 0.15618
R49 VPWR.n9 VPWR.n0 0.149362
R50 VPWR.n5 VPWR.n0 0.122949
R51 a_549_74.n1 a_549_74.t0 290.661
R52 a_549_74.t1 a_549_74.n1 273.188
R53 a_549_74.n1 a_549_74.n0 223.906
R54 a_549_74.n0 a_549_74.t2 202.23
R55 a_549_74.n0 a_549_74.t3 111.343
R56 VPB.t1 VPB.t2 727.823
R57 VPB.t0 VPB.t1 663.98
R58 VPB.t2 VPB.t4 408.603
R59 VPB.t3 VPB.t0 357.527
R60 VPB VPB.t3 252.823
R61 a_682_74.t1 a_682_74.n1 431.709
R62 a_682_74.n1 a_682_74.t0 336.152
R63 a_682_74.n0 a_682_74.t2 265.637
R64 a_682_74.n0 a_682_74.t3 253.853
R65 a_682_74.n1 a_682_74.n0 152
R66 Y.n1 Y 589.268
R67 Y.n1 Y.n0 585
R68 Y.n2 Y.n1 585
R69 Y.n3 Y.t1 225
R70 Y.n1 Y.t0 27.2639
R71 Y Y.n3 9.97283
R72 Y.n2 Y 9.06717
R73 Y.n0 Y 8.53383
R74 Y.n0 Y 4.62272
R75 Y.n3 Y 4.26717
R76 Y Y.n2 4.08939
R77 A.n0 A.t1 293.752
R78 A.n0 A.t0 220.113
R79 A A.n0 159.929
C0 VPB A 0.038386f
C1 VPB VPWR 0.159762f
C2 VPB Y 0.018631f
C3 A VPWR 0.021264f
C4 VPB VGND 0.011698f
C5 VPWR Y 0.147313f
C6 A VGND 0.01746f
C7 VPWR VGND 0.08908f
C8 Y VGND 0.068148f
C9 VGND VNB 0.673773f
C10 Y VNB 0.12103f
C11 VPWR VNB 0.525147f
C12 A VNB 0.205416f
C13 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkinv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkinv_1 VNB VPB VPWR VGND A Y
X0 Y.t2 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2394 ps=2.25 w=0.84 l=0.15
X1 Y.t0 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.22535 pd=2.17 as=0.1491 ps=1.55 w=0.42 l=0.15
X2 VPWR.t0 A.t2 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2394 pd=2.25 as=0.126 ps=1.14 w=0.84 l=0.15
R0 A.n0 A.t0 189.855
R1 A.n0 A.t2 189.855
R2 A.n2 A 156.294
R3 A A.n1 155.76
R4 A.n4 A.n3 152
R5 A.n2 A.t1 121.877
R6 A.n3 A.n1 26.0132
R7 A.n3 A.n2 26.0132
R8 A.n1 A.n0 12.6243
R9 A.n4 A 4.36875
R10 A A.n4 3.14971
R11 VPWR.n0 VPWR.t0 785.482
R12 VPWR.n0 VPWR.t1 427.678
R13 VPWR VPWR.n0 0.548572
R14 Y Y.n0 312.115
R15 Y.n1 Y.t0 166.948
R16 Y.n0 Y.t1 35.1791
R17 Y.n0 Y.t2 35.1791
R18 Y Y.n1 11.382
R19 Y.n1 Y 0.638642
R20 VPB VPB.t1 252.823
R21 VPB.t1 VPB.t0 229.839
R22 VGND VGND.t0 273.411
R23 VNB VNB.t0 1402.2
C0 VPB Y 0.016222f
C1 VPB A 0.108102f
C2 A Y 0.157415f
C3 VPB VPWR 0.059044f
C4 VPWR Y 0.168788f
C5 VPB VGND 0.005214f
C6 Y VGND 0.101926f
C7 A VPWR 0.053008f
C8 A VGND 0.045583f
C9 VPWR VGND 0.024853f
C10 VGND VNB 0.248987f
C11 Y VNB 0.111995f
C12 VPWR VNB 0.233559f
C13 A VNB 0.335814f
C14 VPB VNB 0.406224f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkinv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkinv_2 VNB VPB VPWR VGND Y A
X0 VPWR.t2 A.t0 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t4 A.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X2 VPWR.t1 A.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t0 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t0 A.t4 Y.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
R0 A.n2 A.t1 239.978
R1 A.n0 A.t4 239.978
R2 A.n0 A.t2 226.809
R3 A.n1 A.t3 226.809
R4 A.n2 A.t0 226.809
R5 A.n6 A.n5 152
R6 A.n4 A.n3 152
R7 A.n1 A.n0 65.7278
R8 A.n5 A.n4 49.6611
R9 A.n3 A 12.8005
R10 A.n4 A.n2 10.955
R11 A.n6 A 8.63306
R12 A A.n6 5.65631
R13 A.n5 A.n1 5.11262
R14 A.n3 A 1.48887
R15 Y.n1 Y.t2 274.788
R16 Y.n1 Y.n0 205.487
R17 Y Y.n2 103.124
R18 Y.n2 Y.t4 101.141
R19 Y.n2 Y.t3 99.6658
R20 Y Y.n1 62.1018
R21 Y.n0 Y.t1 26.3844
R22 Y.n0 Y.t0 26.3844
R23 VPWR.n1 VPWR.t1 356.945
R24 VPWR.n1 VPWR.n0 338.455
R25 VPWR.n0 VPWR.t0 26.3844
R26 VPWR.n0 VPWR.t2 26.3844
R27 VPWR VPWR.n1 0.523201
R28 VPB VPB.t2 260.485
R29 VPB.t0 VPB.t1 229.839
R30 VPB.t2 VPB.t0 229.839
R31 VGND.n0 VGND.t0 255.834
R32 VGND.n0 VGND.t1 255.541
R33 VGND VGND.n0 0.194407
R34 VNB.t1 VNB.t0 2148.03
R35 VNB VNB.t1 1143.31
C0 Y VGND 0.150699f
C1 VPWR VGND 0.032998f
C2 VPB A 0.10582f
C3 VPB Y 0.020369f
C4 VPB VPWR 0.064032f
C5 A Y 0.301411f
C6 VPB VGND 0.005125f
C7 A VPWR 0.047227f
C8 A VGND 0.055255f
C9 Y VPWR 0.302645f
C10 VGND VNB 0.336195f
C11 VPWR VNB 0.254588f
C12 Y VNB 0.136442f
C13 A VNB 0.413442f
C14 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkinv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkinv_4 VNB VPB VPWR VGND Y A
X0 Y.t9 A.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t4 A.t1 Y.t8 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t3 A.t2 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1386 pd=1.5 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 Y.t7 A.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 VPWR.t2 A.t4 Y.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5 Y.t5 A.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t0 A.t6 Y.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t2 A.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.06405 pd=0.725 as=0.0882 ps=0.84 w=0.42 l=0.15
X8 VGND.t1 A.t8 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.14805 ps=1.125 w=0.42 l=0.15
X9 Y.t0 A.t9 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14805 pd=1.125 as=0.3066 ps=2.3 w=0.42 l=0.15
R0 A.n3 A.t0 344.606
R1 A.n0 A.t2 239.978
R2 A.n3 A.t9 237.787
R3 A.n2 A.t8 237.787
R4 A.n15 A.t7 237.787
R5 A.n0 A.t1 226.809
R6 A.n14 A.t3 226.809
R7 A.n1 A.t4 226.809
R8 A.n9 A.t5 226.809
R9 A.n4 A.t6 226.809
R10 A.n17 A.n16 152
R11 A.n13 A.n12 152
R12 A.n11 A.n10 152
R13 A.n8 A.n7 152
R14 A.n6 A.n5 152
R15 A.n16 A.n0 60.6157
R16 A.n8 A.n5 49.6611
R17 A.n14 A.n13 44.549
R18 A.n10 A.n9 44.549
R19 A.n13 A.n1 28.4823
R20 A.n10 A.n2 12.4157
R21 A.n6 A 11.7586
R22 A.n5 A.n4 10.955
R23 A.n12 A.n11 10.1214
R24 A.n17 A 9.37724
R25 A.n2 A.n1 8.76414
R26 A.n7 A 7.5912
R27 A.n7 A 6.69817
R28 A.n9 A.n8 5.11262
R29 A A.n17 4.91213
R30 A.n16 A.n15 3.65202
R31 A.n11 A 3.42376
R32 A A.n6 2.53073
R33 A.n4 A.n3 2.19141
R34 A.n15 A.n14 1.46111
R35 A.n12 A 0.744686
R36 VPWR.n5 VPWR.t4 357.81
R37 VPWR.n11 VPWR.t5 349.788
R38 VPWR.n9 VPWR.n1 331.5
R39 VPWR.n4 VPWR.n3 323.406
R40 VPWR.n8 VPWR.n2 36.1417
R41 VPWR.n3 VPWR.t3 35.1791
R42 VPWR.n10 VPWR.n9 34.6358
R43 VPWR.n11 VPWR.n10 26.7299
R44 VPWR.n1 VPWR.t1 26.3844
R45 VPWR.n1 VPWR.t0 26.3844
R46 VPWR.n3 VPWR.t2 26.3844
R47 VPWR.n4 VPWR.n2 23.7181
R48 VPWR.n6 VPWR.n2 9.3005
R49 VPWR.n8 VPWR.n7 9.3005
R50 VPWR.n10 VPWR.n0 9.3005
R51 VPWR.n12 VPWR.n11 9.3005
R52 VPWR.n5 VPWR.n4 6.96039
R53 VPWR.n9 VPWR.n8 1.50638
R54 VPWR.n6 VPWR.n5 0.594857
R55 VPWR.n7 VPWR.n6 0.122949
R56 VPWR.n7 VPWR.n0 0.122949
R57 VPWR.n12 VPWR.n0 0.122949
R58 VPWR VPWR.n12 0.0617245
R59 Y.n11 Y.n2 203.812
R60 Y.n5 Y.n4 203.333
R61 Y.n1 Y.n0 203.333
R62 Y.n6 Y.n3 203.333
R63 Y.n8 Y.n7 185
R64 Y.n10 Y.n9 185
R65 Y.n7 Y.n6 125.266
R66 Y.n9 Y.n8 121.43
R67 Y Y.n1 65.49
R68 Y.n11 Y.n10 53.3607
R69 Y.n2 Y.t3 47.1434
R70 Y.n5 Y.n1 46.6829
R71 Y.n6 Y.n5 42.9181
R72 Y.n9 Y.t1 40.0005
R73 Y.n8 Y.t0 40.0005
R74 Y.n2 Y.t2 40.0005
R75 Y.n3 Y.t4 26.3844
R76 Y.n3 Y.t9 26.3844
R77 Y.n4 Y.t6 26.3844
R78 Y.n4 Y.t5 26.3844
R79 Y.n0 Y.t8 26.3844
R80 Y.n0 Y.t7 26.3844
R81 Y Y.n11 25.977
R82 Y.n10 Y.n7 7.50395
R83 VPB VPB.t5 257.93
R84 VPB.t2 VPB.t3 255.376
R85 VPB.t3 VPB.t4 229.839
R86 VPB.t1 VPB.t2 229.839
R87 VPB.t0 VPB.t1 229.839
R88 VPB.t5 VPB.t0 229.839
R89 VGND.n4 VGND.t3 268.223
R90 VGND.n3 VGND.n2 208.661
R91 VGND.n9 VGND.t0 171.857
R92 VGND.n2 VGND.t2 60.0005
R93 VGND.n2 VGND.t1 60.0005
R94 VGND.n7 VGND.n1 36.1417
R95 VGND.n8 VGND.n7 30.2223
R96 VGND.n3 VGND.n1 17.6946
R97 VGND.n10 VGND.n9 13.5956
R98 VGND.n8 VGND.n0 9.3005
R99 VGND.n5 VGND.n1 9.3005
R100 VGND.n7 VGND.n6 9.3005
R101 VGND.n4 VGND.n3 6.96039
R102 VGND.n9 VGND.n8 3.35927
R103 VGND.n5 VGND.n4 0.594857
R104 VGND.n6 VGND.n5 0.122949
R105 VGND.n6 VGND.n0 0.122949
R106 VGND.n10 VGND.n0 0.122949
R107 VGND VGND.n10 0.0617245
R108 VNB VNB.t0 2171.13
R109 VNB.t0 VNB.t1 1974.8
R110 VNB.t1 VNB.t2 1316.54
R111 VNB.t2 VNB.t3 1050.92
C0 VPB A 0.216943f
C1 VPWR VPB 0.105959f
C2 Y VPB 0.02307f
C3 VPWR A 0.10147f
C4 VGND VPB 0.006199f
C5 Y A 0.668108f
C6 VPWR Y 0.577601f
C7 VGND A 0.073278f
C8 VPWR VGND 0.061084f
C9 Y VGND 0.34967f
C10 VGND VNB 0.487769f
C11 Y VNB 0.17386f
C12 VPWR VNB 0.398785f
C13 A VNB 0.693837f
C14 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfrbp_2 VNB VPB VPWR RESET_B VGND Q Q_N D CLK
X0 a_70_74.t2 D.t0 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1449 ps=1.53 w=0.42 l=0.15
X1 VGND.t5 a_1586_149# Q_N.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_298_294.t0 a_728_331.t1 a_683_485.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 VGND.t7 RESET_B.t0 a_156_74.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1135 pd=1.09 as=0.0504 ps=0.66 w=0.42 l=0.15
X4 a_683_485.t1 a_331_392# VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.141475 ps=1.12 w=0.42 l=0.15
X5 VPWR.t7 RESET_B.t1 a_298_294.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.141475 pd=1.12 as=0.1176 ps=1.4 w=0.42 l=0.15
X6 a_614_81.t1 a_818_418.t2 a_298_294.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2184 pd=1.88 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND.t10 a_728_331.t2 a_818_418.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.3983 pd=2.005 as=0.1998 ps=2.02 w=0.74 l=0.15
X8 Q_N.t0 a_1586_149# VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_728_331.t0 CLK.t0 VPWR.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.372225 ps=1.805 w=1.12 l=0.15
X10 a_1974_74.t1 RESET_B.t2 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 VGND.t0 a_2363_352.t2 Q.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_614_81.t0 a_331_392# a_536_81.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1281 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 a_331_392# a_818_418.t3 a_1586_149# VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.31255 pd=2.62 as=0.10825 ps=1.065 w=0.74 l=0.15
X14 a_2363_352.t0 a_1586_149# VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1728 pd=1.82 as=0.1165 ps=1.065 w=0.64 l=0.15
X15 a_1800_291.t1 RESET_B.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1426 ps=1.155 w=0.42 l=0.15
X16 a_156_74.t1 D.t1 a_70_74.t3 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1176 ps=1.4 w=0.42 l=0.15
X17 a_2363_352.t1 a_1586_149# VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0.2102 ps=1.505 w=1 l=0.15
X18 VGND.t3 a_1800_291.t2 a_1499_149.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1155 ps=1.39 w=0.42 l=0.15
X19 Q.t0 a_2363_352.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1998 ps=2.02 w=0.74 l=0.15
X20 VPWR.t2 RESET_B.t4 a_70_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.385725 pd=2.7 as=0.063 ps=0.72 w=0.42 l=0.15
X21 a_1586_149# a_728_331.t3 a_1499_149.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.10825 pd=1.065 as=0.1197 ps=1.41 w=0.42 l=0.15
X22 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_1800_291.t0 a_1586_149# a_1974_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 Q_N.t2 a_1586_149# VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.181325 ps=1.505 w=1.12 l=0.15
X25 a_331_392# a_298_294.t5 VGND.t9 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1135 ps=1.09 w=0.74 l=0.15
X26 VPWR.t8 a_728_331.t4 a_818_418.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.372225 pd=1.805 as=0.3304 ps=2.83 w=1.12 l=0.15
X27 a_536_81.t1 RESET_B.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1281 ps=1.45 w=0.42 l=0.15
X28 Q.t2 a_2363_352.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X29 a_298_294.t1 a_728_331.t5 a_70_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1456 ps=1.63 w=0.42 l=0.15
X30 a_331_392# a_298_294.t6 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.385725 ps=2.7 w=1 l=0.15
X31 a_70_74.t4 a_818_418.t4 a_298_294.t4 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.2793 pd=2.17 as=0.063 ps=0.72 w=0.42 l=0.15
R0 D.n0 D.t0 192.161
R1 D D.n0 158.4
R2 D.n2 D.n1 152
R3 D.n1 D.t1 121.898
R4 D.n1 D.n0 33.4454
R5 D.n2 D 7.38512
R6 D D.n2 4.75947
R7 VPWR.n56 VPWR.n55 838.287
R8 VPWR.n23 VPWR.t1 788.779
R9 VPWR.n1 VPWR.t10 704.572
R10 VPWR.n7 VPWR.n6 612.649
R11 VPWR.n4 VPWR.n3 585
R12 VPWR.n55 VPWR.n54 585
R13 VPWR.n35 VPWR.n34 585
R14 VPWR.n15 VPWR.t4 348.618
R15 VPWR.n17 VPWR.t3 273.654
R16 VPWR.n3 VPWR.n2 265.587
R17 VPWR.n16 VPWR.t0 264.767
R18 VPWR.n55 VPWR.n3 253.286
R19 VPWR.n2 VPWR.t2 219.339
R20 VPWR.n6 VPWR.t7 178.238
R21 VPWR.n2 VPWR.t5 164.718
R22 VPWR.n6 VPWR.t6 110.227
R23 VPWR.n34 VPWR.t9 57.1657
R24 VPWR.n34 VPWR.t8 57.1657
R25 VPWR.n48 VPWR.n47 36.1417
R26 VPWR.n49 VPWR.n48 36.1417
R27 VPWR.n37 VPWR.n9 36.1417
R28 VPWR.n41 VPWR.n9 36.1417
R29 VPWR.n42 VPWR.n41 36.1417
R30 VPWR.n43 VPWR.n42 36.1417
R31 VPWR.n27 VPWR.n13 36.1417
R32 VPWR.n28 VPWR.n27 36.1417
R33 VPWR.n29 VPWR.n28 36.1417
R34 VPWR.n29 VPWR.n11 36.1417
R35 VPWR.n22 VPWR.n21 36.1417
R36 VPWR.n37 VPWR.n36 35.5857
R37 VPWR.n33 VPWR.n11 35.0296
R38 VPWR.n18 VPWR.n17 35.0123
R39 VPWR.n43 VPWR.n7 30.4946
R40 VPWR.n23 VPWR.n13 28.9887
R41 VPWR.n49 VPWR.n4 23.1409
R42 VPWR.n47 VPWR.n7 22.9652
R43 VPWR.n23 VPWR.n22 16.1887
R44 VPWR.n54 VPWR.n52 12.0894
R45 VPWR.n53 VPWR.n1 11.6627
R46 VPWR.n57 VPWR.n56 10.4383
R47 VPWR.n19 VPWR.n18 9.3005
R48 VPWR.n21 VPWR.n20 9.3005
R49 VPWR.n22 VPWR.n14 9.3005
R50 VPWR.n24 VPWR.n23 9.3005
R51 VPWR.n25 VPWR.n13 9.3005
R52 VPWR.n27 VPWR.n26 9.3005
R53 VPWR.n28 VPWR.n12 9.3005
R54 VPWR.n30 VPWR.n29 9.3005
R55 VPWR.n31 VPWR.n11 9.3005
R56 VPWR.n33 VPWR.n32 9.3005
R57 VPWR.n36 VPWR.n10 9.3005
R58 VPWR.n38 VPWR.n37 9.3005
R59 VPWR.n39 VPWR.n9 9.3005
R60 VPWR.n41 VPWR.n40 9.3005
R61 VPWR.n42 VPWR.n8 9.3005
R62 VPWR.n44 VPWR.n43 9.3005
R63 VPWR.n45 VPWR.n7 9.3005
R64 VPWR.n47 VPWR.n46 9.3005
R65 VPWR.n48 VPWR.n5 9.3005
R66 VPWR.n50 VPWR.n49 9.3005
R67 VPWR.n52 VPWR.n51 9.3005
R68 VPWR.n53 VPWR.n0 9.3005
R69 VPWR.n18 VPWR.n15 7.90638
R70 VPWR.n17 VPWR.n16 6.20914
R71 VPWR.n36 VPWR.n35 4.82512
R72 VPWR.n35 VPWR.n33 4.62819
R73 VPWR.n21 VPWR.n15 3.38874
R74 VPWR.n52 VPWR.n4 1.99161
R75 VPWR.n54 VPWR.n53 1.56494
R76 VPWR.n56 VPWR.n1 0.853833
R77 VPWR.n19 VPWR.n16 0.28297
R78 VPWR.n20 VPWR.n19 0.122949
R79 VPWR.n20 VPWR.n14 0.122949
R80 VPWR.n24 VPWR.n14 0.122949
R81 VPWR.n25 VPWR.n24 0.122949
R82 VPWR.n26 VPWR.n25 0.122949
R83 VPWR.n26 VPWR.n12 0.122949
R84 VPWR.n30 VPWR.n12 0.122949
R85 VPWR.n31 VPWR.n30 0.122949
R86 VPWR.n32 VPWR.n31 0.122949
R87 VPWR.n32 VPWR.n10 0.122949
R88 VPWR.n38 VPWR.n10 0.122949
R89 VPWR.n39 VPWR.n38 0.122949
R90 VPWR.n40 VPWR.n39 0.122949
R91 VPWR.n40 VPWR.n8 0.122949
R92 VPWR.n44 VPWR.n8 0.122949
R93 VPWR.n45 VPWR.n44 0.122949
R94 VPWR.n46 VPWR.n45 0.122949
R95 VPWR.n46 VPWR.n5 0.122949
R96 VPWR.n50 VPWR.n5 0.122949
R97 VPWR.n51 VPWR.n50 0.122949
R98 VPWR.n51 VPWR.n0 0.122949
R99 VPWR.n57 VPWR.n0 0.122949
R100 VPWR VPWR.n57 0.0617245
R101 a_70_74.n1 a_70_74.n0 585
R102 a_70_74.n2 a_70_74.t4 426.834
R103 a_70_74.n2 a_70_74.n1 357.135
R104 a_70_74.n3 a_70_74.n2 348.959
R105 a_70_74.n1 a_70_74.t3 346.7
R106 a_70_74.n0 a_70_74.t0 70.3576
R107 a_70_74.n0 a_70_74.t2 70.3576
R108 a_70_74.n3 a_70_74.t1 21.2663
R109 VPB.n0 VPB 6325.67
R110 VPB.n1 VPB 5011.98
R111 VPB.n2 VPB 2655.91
R112 VPB VPB.n3 2253.92
R113 VPB.t10 VPB.t1 1596.1
R114 VPB.t12 VPB.n2 760
R115 VPB.t7 VPB.t5 508.2
R116 VPB.t3 VPB.t4 482.346
R117 VPB.t9 VPB.t10 408.603
R118 VPB.t8 VPB.t12 335.295
R119 VPB.n2 VPB.t9 329.435
R120 VPB.t11 VPB 316.668
R121 VPB.t4 VPB.n0 315.851
R122 VPB.t6 VPB.t8 290.589
R123 VPB.n0 VPB.t0 270.7
R124 VPB.t5 VPB.t2 260.485
R125 VPB.n1 VPB.t3 254.639
R126 VPB.t1 VPB.n1 237.5
R127 VPB.n3 VPB.t6 234.707
R128 VPB.n3 VPB.t7 229.839
R129 VPB.t2 VPB.t11 229.839
R130 CLK.n1 CLK.t0 248.883
R131 CLK.n1 CLK.n0 174.707
R132 CLK CLK.n1 163.107
R133 VGND.n5 VGND.t10 316.409
R134 VGND.n1 VGND.t2 254.57
R135 VGND.n55 VGND.n54 210.018
R136 VGND.n25 VGND.n24 206.528
R137 VGND.n18 VGND.n17 204.388
R138 VGND.n14 VGND.t0 180.232
R139 VGND.n11 VGND.t4 176.839
R140 VGND.n13 VGND.t1 174.405
R141 VGND.n54 VGND.t9 44.5565
R142 VGND.n24 VGND.t8 40.0005
R143 VGND.n24 VGND.t3 40.0005
R144 VGND.n54 VGND.t7 40.0005
R145 VGND.n23 VGND.n22 36.1417
R146 VGND.n26 VGND.n23 36.1417
R147 VGND.n30 VGND.n9 36.1417
R148 VGND.n31 VGND.n30 36.1417
R149 VGND.n32 VGND.n31 36.1417
R150 VGND.n32 VGND.n7 36.1417
R151 VGND.n36 VGND.n7 36.1417
R152 VGND.n37 VGND.n36 36.1417
R153 VGND.n38 VGND.n37 36.1417
R154 VGND.n42 VGND.n41 36.1417
R155 VGND.n43 VGND.n42 36.1417
R156 VGND.n43 VGND.n3 36.1417
R157 VGND.n47 VGND.n3 36.1417
R158 VGND.n48 VGND.n47 36.1417
R159 VGND.n49 VGND.n48 36.1417
R160 VGND.n53 VGND.n52 36.1417
R161 VGND.n17 VGND.t6 33.7505
R162 VGND.n16 VGND.n13 29.3652
R163 VGND.n19 VGND.n11 26.3534
R164 VGND.n19 VGND.n18 25.977
R165 VGND.n17 VGND.t5 23.5986
R166 VGND.n18 VGND.n16 20.7064
R167 VGND.n55 VGND.n53 15.4358
R168 VGND.n38 VGND.n5 10.9181
R169 VGND.n22 VGND.n11 9.78874
R170 VGND.n53 VGND.n0 9.3005
R171 VGND.n52 VGND.n51 9.3005
R172 VGND.n50 VGND.n49 9.3005
R173 VGND.n48 VGND.n2 9.3005
R174 VGND.n47 VGND.n46 9.3005
R175 VGND.n45 VGND.n3 9.3005
R176 VGND.n44 VGND.n43 9.3005
R177 VGND.n42 VGND.n4 9.3005
R178 VGND.n41 VGND.n40 9.3005
R179 VGND.n39 VGND.n38 9.3005
R180 VGND.n37 VGND.n6 9.3005
R181 VGND.n36 VGND.n35 9.3005
R182 VGND.n34 VGND.n7 9.3005
R183 VGND.n33 VGND.n32 9.3005
R184 VGND.n31 VGND.n8 9.3005
R185 VGND.n30 VGND.n29 9.3005
R186 VGND.n28 VGND.n9 9.3005
R187 VGND.n27 VGND.n26 9.3005
R188 VGND.n23 VGND.n10 9.3005
R189 VGND.n22 VGND.n21 9.3005
R190 VGND.n20 VGND.n19 9.3005
R191 VGND.n18 VGND.n12 9.3005
R192 VGND.n16 VGND.n15 9.3005
R193 VGND.n49 VGND.n1 7.90638
R194 VGND.n56 VGND.n55 7.51398
R195 VGND.n26 VGND.n25 7.15344
R196 VGND.n14 VGND.n13 6.7255
R197 VGND.n41 VGND.n5 6.4005
R198 VGND.n25 VGND.n9 4.14168
R199 VGND.n52 VGND.n1 3.38874
R200 VGND.n15 VGND.n14 0.585846
R201 VGND VGND.n56 0.280236
R202 VGND.n56 VGND.n0 0.150642
R203 VGND.n15 VGND.n12 0.122949
R204 VGND.n20 VGND.n12 0.122949
R205 VGND.n21 VGND.n20 0.122949
R206 VGND.n21 VGND.n10 0.122949
R207 VGND.n27 VGND.n10 0.122949
R208 VGND.n28 VGND.n27 0.122949
R209 VGND.n29 VGND.n28 0.122949
R210 VGND.n29 VGND.n8 0.122949
R211 VGND.n33 VGND.n8 0.122949
R212 VGND.n34 VGND.n33 0.122949
R213 VGND.n35 VGND.n34 0.122949
R214 VGND.n35 VGND.n6 0.122949
R215 VGND.n39 VGND.n6 0.122949
R216 VGND.n40 VGND.n39 0.122949
R217 VGND.n40 VGND.n4 0.122949
R218 VGND.n44 VGND.n4 0.122949
R219 VGND.n45 VGND.n44 0.122949
R220 VGND.n46 VGND.n45 0.122949
R221 VGND.n46 VGND.n2 0.122949
R222 VGND.n50 VGND.n2 0.122949
R223 VGND.n51 VGND.n50 0.122949
R224 VGND.n51 VGND.n0 0.122949
R225 a_728_331.t2 a_728_331.t5 976.854
R226 a_728_331.t0 a_728_331.n3 822.068
R227 a_728_331.t5 a_728_331.t1 355.877
R228 a_728_331.n3 a_728_331.n1 313.37
R229 a_728_331.n1 a_728_331.t3 245.821
R230 a_728_331.n1 a_728_331.n0 237.787
R231 a_728_331.n2 a_728_331.t4 235.892
R232 a_728_331.n2 a_728_331.t2 201.458
R233 a_728_331.n3 a_728_331.n2 127.882
R234 VNB.n0 VNB 24676.2
R235 VNB.n1 VNB 12010.5
R236 VNB.t6 VNB.t5 5497.11
R237 VNB.t16 VNB.t3 2390.55
R238 VNB.t2 VNB.t14 2332.81
R239 VNB.t8 VNB.t1 2314.52
R240 VNB.n0 VNB.t9 2193.97
R241 VNB.t15 VNB 1628.35
R242 VNB.n1 VNB.t4 1345.29
R243 VNB VNB.t11 1244.14
R244 VNB.t14 VNB.t12 1154.86
R245 VNB.t10 VNB.t8 1145.21
R246 VNB.t5 VNB.t16 1097.11
R247 VNB.t1 VNB.t0 1036.71
R248 VNB.t9 VNB.t10 1036.71
R249 VNB.t3 VNB.t13 993.177
R250 VNB.t11 VNB.t2 900.788
R251 VNB.t12 VNB.t15 900.788
R252 VNB.t13 VNB.t7 831.496
R253 VNB.n1 VNB.t6 635.172
R254 VNB.t7 VNB.n0 184.778
R255 VNB.t11 VNB.n1 50.1906
R256 Q_N Q_N.t2 284.916
R257 Q_N.n1 Q_N.n0 95.3607
R258 Q_N.n0 Q_N.t1 22.7032
R259 Q_N.n0 Q_N.t0 22.7032
R260 Q_N.n2 Q_N 21.3338
R261 Q_N.n2 Q_N 10.2405
R262 Q_N.n2 Q_N.n1 4.84248
R263 Q_N Q_N.n2 2.89861
R264 Q_N.n1 Q_N 1.18364
R265 a_683_485.t0 a_683_485.t1 112.572
R266 a_298_294.n1 a_298_294.t2 683.005
R267 a_298_294.n3 a_298_294.n2 605.946
R268 a_298_294.n0 a_298_294.t5 234.573
R269 a_298_294.n1 a_298_294.n0 227.274
R270 a_298_294.n4 a_298_294.n3 215.249
R271 a_298_294.n0 a_298_294.t6 209.72
R272 a_298_294.n3 a_298_294.n1 102.025
R273 a_298_294.n2 a_298_294.t4 70.3576
R274 a_298_294.n2 a_298_294.t0 70.3576
R275 a_298_294.n4 a_298_294.t3 40.0005
R276 a_298_294.t1 a_298_294.n4 40.0005
R277 RESET_B.n3 RESET_B.t0 303.661
R278 RESET_B.n0 RESET_B.t2 303.661
R279 RESET_B.n1 RESET_B.t5 290.808
R280 RESET_B.n1 RESET_B.t1 269.652
R281 RESET_B.n2 RESET_B.n0 172.864
R282 RESET_B RESET_B.n3 165.736
R283 RESET_B.n2 RESET_B.n1 164.792
R284 RESET_B.n3 RESET_B.t4 143.798
R285 RESET_B.n0 RESET_B.t3 139.78
R286 RESET_B RESET_B.n2 0.0466957
R287 a_156_74.t0 a_156_74.t1 68.5719
R288 a_818_418.n4 a_818_418.n3 461.644
R289 a_818_418.n1 a_818_418.t0 314.286
R290 a_818_418.n1 a_818_418.n0 240.421
R291 a_818_418.n0 a_818_418.t2 231.361
R292 a_818_418.t1 a_818_418.n4 220.516
R293 a_818_418.n3 a_818_418.n2 198.327
R294 a_818_418.n3 a_818_418.t3 173.157
R295 a_818_418.n0 a_818_418.t4 148.35
R296 a_818_418.n4 a_818_418.n1 16.1872
R297 a_614_81.t0 a_614_81.t1 664.804
R298 a_1800_291.n2 a_1800_291.t1 655.357
R299 a_1800_291.t0 a_1800_291.n2 358.241
R300 a_1800_291.n1 a_1800_291.t2 281.998
R301 a_1800_291.n2 a_1800_291.n1 214.548
R302 a_1800_291.n1 a_1800_291.n0 138.441
R303 a_1974_74.t0 a_1974_74.t1 60.0005
R304 a_2363_352.t1 a_2363_352.n4 265.079
R305 a_2363_352.n1 a_2363_352.n0 240.197
R306 a_2363_352.n3 a_2363_352.t4 240.197
R307 a_2363_352.n1 a_2363_352.t2 193.53
R308 a_2363_352.n4 a_2363_352.n3 188.968
R309 a_2363_352.n2 a_2363_352.t3 179.947
R310 a_2363_352.n4 a_2363_352.t0 153.954
R311 a_2363_352.n2 a_2363_352.n1 51.852
R312 a_2363_352.n3 a_2363_352.n2 13.8763
R313 Q.n0 Q.t2 295.44
R314 Q Q.n1 198.382
R315 Q.n1 Q.n0 185
R316 Q.n1 Q.t1 22.7032
R317 Q.n1 Q.t0 22.7032
R318 Q Q.n0 4.26717
R319 a_536_81.t0 a_536_81.t1 68.5719
R320 a_1499_149.t0 a_1499_149.t1 570.667
C0 RESET_B a_331_392# 0.326751f
C1 a_1586_149# a_1755_389# 0.005754f
C2 a_1755_389# VPWR 0.002336f
C3 D VGND 0.018385f
C4 RESET_B CLK 0.023276f
C5 CLK a_331_392# 0.046774f
C6 RESET_B VGND 0.311586f
C7 VGND a_331_392# 0.875174f
C8 D VPB 0.053679f
C9 CLK VGND 0.005514f
C10 RESET_B Q_N 5.85e-19
C11 RESET_B VPB 0.225939f
C12 D VPWR 0.037005f
C13 a_331_392# VPB 0.064039f
C14 RESET_B Q 6.09e-20
C15 CLK Q_N 6.51e-21
C16 RESET_B a_1586_149# 0.203947f
C17 RESET_B VPWR 0.284808f
C18 CLK VPB 0.045764f
C19 a_331_392# a_1586_149# 0.01045f
C20 a_331_392# VPWR 0.027692f
C21 VGND Q_N 0.166762f
C22 CLK Q 4.2e-21
C23 VGND VPB 0.015108f
C24 CLK VPWR 0.011558f
C25 VGND Q 0.171292f
C26 VGND a_1586_149# 0.126924f
C27 VGND VPWR 0.098673f
C28 Q_N VPB 0.006858f
C29 Q_N a_1586_149# 0.120434f
C30 RESET_B a_1755_389# 0.001608f
C31 Q VPB 0.007224f
C32 Q_N VPWR 0.192372f
C33 a_1586_149# VPB 0.210327f
C34 VPB VPWR 0.459204f
C35 Q a_1586_149# 5.73e-19
C36 Q VPWR 0.231274f
C37 a_1586_149# VPWR 0.10175f
C38 D RESET_B 0.086808f
C39 Q VNB 0.03021f
C40 Q_N VNB 0.00928f
C41 VGND VNB 1.63023f
C42 CLK VNB 0.129475f
C43 RESET_B VNB 0.43112f
C44 D VNB 0.235825f
C45 VPWR VNB 1.30116f
C46 VPB VNB 3.05971f
C47 a_1586_149# VNB 0.513304f
C48 a_331_392# VNB 0.342236f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfrbp_1 VNB VPB VPWR RESET_B VGND Q CLK D Q_N
X0 a_796_463.t1 a_319_360.t2 a_706_463.t4 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1 a_841_401.t2 a_706_463.t5 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1611 pd=1.22 as=0.1601 ps=1.27 w=0.64 l=0.15
X2 a_706_463.t2 a_498_360.t2 a_38_78.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3 a_706_463.t3 a_319_360.t3 a_38_78.t4 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4 Q_N a_1224_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_498_360.t0 a_319_360.t4 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X6 a_38_78.t0 D.t0 VPWR.t9 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X7 a_1624_74.t0 RESET_B.t0 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0861 ps=0.83 w=0.42 l=0.15
X8 a_1224_74# a_498_360.t3 a_841_401.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2165 pd=1.54 as=0.1611 ps=1.22 w=0.64 l=0.15
X9 a_706_463.t1 RESET_B.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.139975 ps=1.155 w=0.42 l=0.15
X10 VGND.t1 RESET_B.t2 a_910_118.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1601 pd=1.27 as=0.0504 ps=0.66 w=0.42 l=0.15
X11 VGND.t4 a_1482_48.t2 a_1434_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0861 pd=0.83 as=0.0504 ps=0.66 w=0.42 l=0.15
X12 a_910_118.t1 a_841_401.t3 a_832_118.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 VPWR.t7 a_1224_74# a_1482_48.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1729 pd=1.485 as=0.063 ps=0.72 w=0.42 l=0.15
X14 Q.t1 a_2026_424.t2 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1918 ps=1.485 w=1.12 l=0.15
X15 VPWR.t0 a_1482_48.t3 a_1465_471.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_498_360.t1 a_319_360.t5 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X17 VPWR.t2 CLK.t0 a_319_360.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X18 Q.t0 a_2026_424.t3 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.122375 ps=1.09 w=0.74 l=0.15
X19 a_1465_471.t1 a_498_360.t4 a_1224_74# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.19385 ps=1.6 w=0.42 l=0.15
X20 a_1482_48.t0 a_1224_74# a_1624_74.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X21 a_125_78.t1 D.t1 a_38_78.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X22 Q_N.t0 a_1224_74# VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.6888 pd=3.47 as=0.1729 ps=1.485 w=1.12 l=0.15
X23 VPWR.t4 RESET_B.t3 a_38_78.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X24 VGND.t3 CLK.t1 a_319_360.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X25 a_832_118.t0 a_498_360.t5 a_706_463.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X26 VPWR.t5 a_1224_74# a_2026_424.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1918 pd=1.485 as=0.2478 ps=2.27 w=0.84 l=0.15
X27 a_1434_74.t1 a_319_360.t6 a_1224_74# VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.2165 ps=1.54 w=0.42 l=0.15
X28 VGND.t7 a_1224_74# a_2026_424.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.122375 pd=1.09 as=0.15675 ps=1.67 w=0.55 l=0.15
X29 VPWR.t10 a_841_401.t4 a_796_463.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.139975 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X30 a_841_401.t1 a_706_463.t6 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X31 VGND.t6 RESET_B.t4 a_125_78.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1365 pd=1.49 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_319_360.n1 a_319_360.n0 1064.68
R1 a_319_360.t1 a_319_360.n5 902.143
R2 a_319_360.n2 a_319_360.n1 772.808
R3 a_319_360.n0 a_319_360.t6 651.236
R4 a_319_360.n2 a_319_360.t3 318.385
R5 a_319_360.n3 a_319_360.t5 267.416
R6 a_319_360.n5 a_319_360.n4 204.329
R7 a_319_360.n1 a_319_360.t2 182.625
R8 a_319_360.n5 a_319_360.t0 145.559
R9 a_319_360.n3 a_319_360.t4 142.994
R10 a_319_360.n4 a_319_360.n2 42.9183
R11 a_319_360.n4 a_319_360.n3 9.24434
R12 a_706_463.n1 a_706_463.t1 667.779
R13 a_706_463.n3 a_706_463.n2 610.035
R14 a_706_463.n0 a_706_463.t6 371.433
R15 a_706_463.n4 a_706_463.n3 295.904
R16 a_706_463.n1 a_706_463.n0 232.941
R17 a_706_463.n0 a_706_463.t5 215.293
R18 a_706_463.n2 a_706_463.t4 70.3576
R19 a_706_463.n2 a_706_463.t2 70.3576
R20 a_706_463.n3 a_706_463.n1 64.4891
R21 a_706_463.n4 a_706_463.t3 60.0005
R22 a_706_463.t0 a_706_463.n4 40.0005
R23 a_796_463.t0 a_796_463.t1 112.572
R24 VPB.n0 VPB 3605.91
R25 VPB VPB.n1 707.5
R26 VPB.t10 VPB.t9 692.071
R27 VPB.t2 VPB.t7 580
R28 VPB.t12 VPB.t4 520
R29 VPB.t0 VPB.t11 490.324
R30 VPB.t7 VPB.n0 485
R31 VPB.t3 VPB.t2 317.5
R32 VPB.n1 VPB.t6 275
R33 VPB.t9 VPB.t14 263.038
R34 VPB.t11 VPB.t10 263.038
R35 VPB.t1 VPB 257.93
R36 VPB.n1 VPB.t8 234.946
R37 VPB.t8 VPB.t1 229.839
R38 VPB.t4 VPB.t13 225
R39 VPB.t6 VPB.t12 225
R40 VPB.t5 VPB.t0 214.517
R41 VPB.t13 VPB.t3 195
R42 VPB.n0 VPB.t5 97.0435
R43 VGND.n33 VGND.t6 267.149
R44 VGND.n20 VGND.n19 222.713
R45 VGND.n31 VGND.n2 207.304
R46 VGND.n11 VGND.n8 200.444
R47 VGND.n10 VGND.n9 134.626
R48 VGND.n19 VGND.t1 72.8576
R49 VGND.n8 VGND.t0 58.5719
R50 VGND.n8 VGND.t4 58.5719
R51 VGND.n9 VGND.t7 44.6103
R52 VGND.n13 VGND.n12 36.1417
R53 VGND.n13 VGND.n6 36.1417
R54 VGND.n17 VGND.n6 36.1417
R55 VGND.n18 VGND.n17 36.1417
R56 VGND.n25 VGND.n4 36.1417
R57 VGND.n26 VGND.n25 36.1417
R58 VGND.n27 VGND.n26 36.1417
R59 VGND.n27 VGND.n1 36.1417
R60 VGND.n19 VGND.t5 34.688
R61 VGND.n2 VGND.t8 34.0546
R62 VGND.n2 VGND.t3 34.0546
R63 VGND.n21 VGND.n4 33.9171
R64 VGND.n32 VGND.n31 30.8711
R65 VGND.n33 VGND.n32 30.1181
R66 VGND.n9 VGND.t2 23.1911
R67 VGND.n20 VGND.n18 18.9495
R68 VGND.n31 VGND.n1 16.5652
R69 VGND.n32 VGND.n0 9.3005
R70 VGND.n31 VGND.n30 9.3005
R71 VGND.n29 VGND.n1 9.3005
R72 VGND.n28 VGND.n27 9.3005
R73 VGND.n26 VGND.n3 9.3005
R74 VGND.n25 VGND.n24 9.3005
R75 VGND.n23 VGND.n4 9.3005
R76 VGND.n22 VGND.n21 9.3005
R77 VGND.n18 VGND.n5 9.3005
R78 VGND.n17 VGND.n16 9.3005
R79 VGND.n15 VGND.n6 9.3005
R80 VGND.n14 VGND.n13 9.3005
R81 VGND.n12 VGND.n7 9.3005
R82 VGND.n11 VGND.n10 7.45275
R83 VGND.n12 VGND.n11 7.15344
R84 VGND.n34 VGND.n33 7.13181
R85 VGND.n21 VGND.n20 3.10353
R86 VGND VGND.n34 0.27433
R87 VGND.n34 VGND.n0 0.156458
R88 VGND.n10 VGND.n7 0.153541
R89 VGND.n14 VGND.n7 0.122949
R90 VGND.n15 VGND.n14 0.122949
R91 VGND.n16 VGND.n15 0.122949
R92 VGND.n16 VGND.n5 0.122949
R93 VGND.n22 VGND.n5 0.122949
R94 VGND.n23 VGND.n22 0.122949
R95 VGND.n24 VGND.n23 0.122949
R96 VGND.n24 VGND.n3 0.122949
R97 VGND.n28 VGND.n3 0.122949
R98 VGND.n29 VGND.n28 0.122949
R99 VGND.n30 VGND.n29 0.122949
R100 VGND.n30 VGND.n0 0.122949
R101 a_841_401.t1 a_841_401.n2 314.072
R102 a_841_401.n0 a_841_401.t3 264.659
R103 a_841_401.n2 a_841_401.n1 185
R104 a_841_401.n2 a_841_401.n0 182.793
R105 a_841_401.n0 a_841_401.t4 160.649
R106 a_841_401.n1 a_841_401.t0 41.2505
R107 a_841_401.n1 a_841_401.t2 41.2505
R108 VNB.n0 VNB 16306.6
R109 VNB VNB.n1 13542.2
R110 VNB.t11 VNB.t10 4804.2
R111 VNB.t4 VNB.n0 2481.11
R112 VNB.t14 VNB.t13 2465.42
R113 VNB.t6 VNB.t9 2430.03
R114 VNB.t8 VNB.t3 1391.96
R115 VNB.t13 VNB.t6 1344.77
R116 VNB.t0 VNB 1297.59
R117 VNB.t7 VNB.t2 1293.44
R118 VNB.n1 VNB.t4 1234.44
R119 VNB.t1 VNB.t14 1179.62
R120 VNB.t10 VNB.t5 1154.86
R121 VNB.t3 VNB.t15 920.107
R122 VNB.t15 VNB.t1 920.107
R123 VNB.t9 VNB.t0 920.107
R124 VNB.t2 VNB.t11 900.788
R125 VNB.t12 VNB.t7 900.788
R126 VNB.n1 VNB.t8 200.536
R127 VNB.n0 VNB.t12 41.566
R128 a_498_360.t1 a_498_360.n3 871.173
R129 a_498_360.n0 a_498_360.t3 442.447
R130 a_498_360.n2 a_498_360.t5 378.353
R131 a_498_360.n0 a_498_360.t4 359.974
R132 a_498_360.n1 a_498_360.n0 277.142
R133 a_498_360.n1 a_498_360.t0 254.475
R134 a_498_360.n2 a_498_360.t2 205.387
R135 a_498_360.n3 a_498_360.n2 165.77
R136 a_498_360.n3 a_498_360.n1 63.8392
R137 a_38_78.n0 a_38_78.t2 660.4
R138 a_38_78.n2 a_38_78.n1 601.726
R139 a_38_78.t1 a_38_78.n2 367.041
R140 a_38_78.n0 a_38_78.t4 355.188
R141 a_38_78.n2 a_38_78.n0 163.388
R142 a_38_78.n1 a_38_78.t3 70.3576
R143 a_38_78.n1 a_38_78.t0 70.3576
R144 Q_N.n1 Q_N.n0 585
R145 Q_N.n3 Q_N.n0 585
R146 Q_N.n4 Q_N.n1 585
R147 Q_N.n4 Q_N.n3 585
R148 Q_N.n2 Q_N 280.596
R149 Q_N.n2 Q_N.n1 28.4487
R150 Q_N.n3 Q_N.n2 28.4487
R151 Q_N.n1 Q_N.t0 26.3844
R152 Q_N Q_N.n4 6.21499
R153 Q_N Q_N.n0 5.38021
R154 Q_N Q_N.n0 1.48456
R155 Q_N.n4 Q_N 0.649775
R156 D.n3 D.t0 182.476
R157 D D.n0 153.458
R158 D.n2 D.n1 152
R159 D.n4 D.n3 152
R160 D.n0 D.t1 148.171
R161 D.n3 D.n2 40.4647
R162 D.n2 D.n0 40.4647
R163 D.n1 D 9.55999
R164 D.n4 D 8.58784
R165 D D.n4 3.40303
R166 D.n1 D 2.43088
R167 VPWR.n10 VPWR.t0 710.604
R168 VPWR.n40 VPWR.t9 685.053
R169 VPWR.n38 VPWR.t4 681.726
R170 VPWR.n27 VPWR.n7 671
R171 VPWR.n3 VPWR.n2 607.303
R172 VPWR.n14 VPWR.n13 333.747
R173 VPWR.n8 VPWR.t3 271.959
R174 VPWR.n12 VPWR.n11 240.456
R175 VPWR.n7 VPWR.t1 114.918
R176 VPWR.n7 VPWR.t10 112.572
R177 VPWR.n13 VPWR.t7 103.12
R178 VPWR.n11 VPWR.t5 46.074
R179 VPWR.n31 VPWR.n5 36.1417
R180 VPWR.n32 VPWR.n31 36.1417
R181 VPWR.n33 VPWR.n32 36.1417
R182 VPWR.n26 VPWR.n25 36.1417
R183 VPWR.n20 VPWR.n19 36.1417
R184 VPWR.n21 VPWR.n20 36.1417
R185 VPWR.n11 VPWR.t11 34.8232
R186 VPWR.n21 VPWR.n8 33.8829
R187 VPWR.n15 VPWR.n14 30.8711
R188 VPWR.n19 VPWR.n10 29.7417
R189 VPWR.n13 VPWR.t6 28.9789
R190 VPWR.n39 VPWR.n38 28.2358
R191 VPWR.n27 VPWR.n5 27.1064
R192 VPWR.n40 VPWR.n39 26.7299
R193 VPWR.n2 VPWR.t8 26.3844
R194 VPWR.n2 VPWR.t2 26.3844
R195 VPWR.n37 VPWR.n3 25.977
R196 VPWR.n15 VPWR.n10 25.6005
R197 VPWR.n38 VPWR.n37 25.224
R198 VPWR.n33 VPWR.n3 21.4593
R199 VPWR.n25 VPWR.n8 19.577
R200 VPWR.n27 VPWR.n26 19.2005
R201 VPWR.n16 VPWR.n15 9.3005
R202 VPWR.n17 VPWR.n10 9.3005
R203 VPWR.n19 VPWR.n18 9.3005
R204 VPWR.n20 VPWR.n9 9.3005
R205 VPWR.n22 VPWR.n21 9.3005
R206 VPWR.n23 VPWR.n8 9.3005
R207 VPWR.n25 VPWR.n24 9.3005
R208 VPWR.n26 VPWR.n6 9.3005
R209 VPWR.n28 VPWR.n27 9.3005
R210 VPWR.n29 VPWR.n5 9.3005
R211 VPWR.n31 VPWR.n30 9.3005
R212 VPWR.n32 VPWR.n4 9.3005
R213 VPWR.n34 VPWR.n33 9.3005
R214 VPWR.n35 VPWR.n3 9.3005
R215 VPWR.n37 VPWR.n36 9.3005
R216 VPWR.n38 VPWR.n1 9.3005
R217 VPWR.n39 VPWR.n0 9.3005
R218 VPWR.n41 VPWR.n40 9.3005
R219 VPWR.n14 VPWR.n12 7.21245
R220 VPWR.n16 VPWR.n12 0.168377
R221 VPWR.n17 VPWR.n16 0.122949
R222 VPWR.n18 VPWR.n17 0.122949
R223 VPWR.n18 VPWR.n9 0.122949
R224 VPWR.n22 VPWR.n9 0.122949
R225 VPWR.n23 VPWR.n22 0.122949
R226 VPWR.n24 VPWR.n23 0.122949
R227 VPWR.n24 VPWR.n6 0.122949
R228 VPWR.n28 VPWR.n6 0.122949
R229 VPWR.n29 VPWR.n28 0.122949
R230 VPWR.n30 VPWR.n29 0.122949
R231 VPWR.n30 VPWR.n4 0.122949
R232 VPWR.n34 VPWR.n4 0.122949
R233 VPWR.n35 VPWR.n34 0.122949
R234 VPWR.n36 VPWR.n35 0.122949
R235 VPWR.n36 VPWR.n1 0.122949
R236 VPWR.n1 VPWR.n0 0.122949
R237 VPWR.n41 VPWR.n0 0.122949
R238 VPWR VPWR.n41 0.0617245
R239 RESET_B.n1 RESET_B.t0 427.373
R240 RESET_B.n2 RESET_B.t2 319.509
R241 RESET_B.n3 RESET_B.n2 234.067
R242 RESET_B.n4 RESET_B.t3 222.054
R243 RESET_B.n4 RESET_B.t4 219.34
R244 RESET_B.n3 RESET_B.n1 171.681
R245 RESET_B.n1 RESET_B.n0 146.475
R246 RESET_B.n2 RESET_B.t1 114.341
R247 RESET_B.n5 RESET_B.n4 58.2296
R248 RESET_B.n5 RESET_B.n3 3.75632
R249 RESET_B RESET_B.n5 0.0466957
R250 a_1624_74.t0 a_1624_74.t1 68.5719
R251 a_910_118.t0 a_910_118.t1 68.5719
R252 a_1482_48.n1 a_1482_48.t1 772.643
R253 a_1482_48.n0 a_1482_48.t3 395.471
R254 a_1482_48.t0 a_1482_48.n1 235.69
R255 a_1482_48.n1 a_1482_48.n0 212.988
R256 a_1482_48.n0 a_1482_48.t2 125.55
R257 a_1434_74.t0 a_1434_74.t1 68.5719
R258 a_832_118.t0 a_832_118.t1 68.5719
R259 a_2026_424.t1 a_2026_424.n1 422.212
R260 a_2026_424.n0 a_2026_424.t2 264.298
R261 a_2026_424.n1 a_2026_424.t0 249.338
R262 a_2026_424.n0 a_2026_424.t3 204.048
R263 a_2026_424.n1 a_2026_424.n0 177.213
R264 Q.t0 Q.n0 279.738
R265 Q.n1 Q.t0 279.738
R266 Q Q.t1 230.639
R267 Q.n0 Q 62.2838
R268 Q.n1 Q 11.2437
R269 Q.n0 Q 4.32482
R270 Q Q.n1 1.55726
R271 a_1465_471.t0 a_1465_471.t1 126.644
R272 CLK.n0 CLK.t0 250.909
R273 CLK.n0 CLK.t1 207.261
R274 CLK CLK.n0 156.849
R275 a_125_78.t0 a_125_78.t1 68.5719
C0 a_1224_74# Q 0.003395f
C1 RESET_B VGND 0.222513f
C2 VPB Q 0.014591f
C3 VGND Q_N 0.119544f
C4 RESET_B Q_N 0.001194f
C5 VGND Q 0.106015f
C6 RESET_B Q 1.43e-19
C7 a_1224_74# VPWR 0.154651f
C8 VPB VPWR 0.362201f
C9 VPWR CLK 0.01695f
C10 a_1224_74# VPB 0.26807f
C11 VPB CLK 0.037766f
C12 D VPWR 0.039803f
C13 VPWR VGND 0.078022f
C14 VPB D 0.102354f
C15 a_1224_74# VGND 0.157652f
C16 RESET_B VPWR 0.396054f
C17 VPB VGND 0.020012f
C18 CLK VGND 0.015912f
C19 VPWR Q_N 0.143311f
C20 a_1224_74# RESET_B 0.235844f
C21 VPB RESET_B 0.357821f
C22 a_1224_74# Q_N 0.082234f
C23 D VGND 0.015719f
C24 RESET_B CLK 0.042357f
C25 VPB Q_N 0.019209f
C26 VPWR Q 0.136987f
C27 D RESET_B 0.131765f
C28 Q VNB 0.112976f
C29 Q_N VNB 0.014245f
C30 VGND VNB 1.34005f
C31 CLK VNB 0.110268f
C32 VPWR VNB 1.04737f
C33 RESET_B VNB 0.388084f
C34 D VNB 0.245673f
C35 VPB VNB 2.69503f
C36 a_1224_74# VNB 0.521526f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfbbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfbbp_1 VNB VPB VPWR VGND Q CLK D RESET_B Q_N SET_B
X0 a_422_125.t0 D.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.2604 ps=2.08 w=0.42 l=0.15
X1 a_520_87.t0 a_27_74.t2 a_422_125.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.088025 ps=0.95 w=0.42 l=0.15
X2 VPWR.t6 CLK.t0 a_27_74.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2408 pd=1.55 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_671_93.t2 SET_B.t0 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.23 as=0.14805 ps=1.28 w=0.84 l=0.15
X4 VPWR.t5 a_1062_93.t2 a_1814_392.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.1325 ps=1.265 w=1 l=0.15
X5 a_1318_119.t1 a_671_93.t4 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.05775 pd=0.76 as=0.26105 ps=2.28 w=0.55 l=0.15
X6 VPWR.t8 RESET_B.t0 a_1062_93.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1828 pd=1.485 as=0.176 ps=1.83 w=0.64 l=0.15
X7 Q.t0 a_2320_410.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.10825 ps=1.065 w=0.74 l=0.15
X8 VPWR.t9 a_1062_93.t3 a_1017_379.t0 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.2 as=0.1134 ps=1.11 w=0.84 l=0.15
X9 a_872_119.t0 a_1062_93.t4 a_671_93.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.26245 pd=2.29 as=0.077 ps=0.83 w=0.55 l=0.15
X10 a_1017_379.t1 a_520_87.t4 a_671_93.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.1638 ps=1.23 w=0.84 l=0.15
X11 a_606_87.t0 a_214_74.t2 a_520_87.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.08225 pd=0.905 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 a_872_119.t2 SET_B.t1 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.192025 pd=1.335 as=0.237825 ps=1.52 w=0.55 l=0.15
X13 VPWR.t10 a_671_93.t5 a_713_379.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.14805 pd=1.28 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 VPWR.t3 a_1474_446.t2 a_2320_410.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1918 pd=1.485 as=0.231 ps=2.23 w=0.84 l=0.15
X15 a_1474_446.t1 a_1311_424# a_1708_74# VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 VGND.t5 CLK.t1 a_27_74.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X17 a_1814_392.t1 a_1311_424# a_1474_446.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1325 pd=1.265 as=0.1825 ps=1.365 w=1 l=0.15
X18 Q_N.t1 a_1474_446.t3 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1828 ps=1.485 w=1.12 l=0.15
X19 a_713_379.t0 a_27_74.t3 a_520_87.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.11445 ps=1.21 w=0.42 l=0.15
X20 a_1418_508.t0 a_214_74.t3 a_1311_424# VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.1428 ps=1.225 w=0.42 l=0.15
X21 a_1708_74# SET_B.t2 VGND.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1212 ps=1.1 w=0.74 l=0.15
X22 a_214_74.t1 a_27_74.t4 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.2408 ps=1.55 w=1.12 l=0.15
X23 Q_N.t0 a_1474_446.t4 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1303 ps=1.17 w=0.74 l=0.15
X24 a_214_74.t0 a_27_74.t5 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X25 a_422_125.t1 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.088025 pd=0.95 as=0.1197 ps=1.41 w=0.42 l=0.15
X26 a_1498_74.t0 a_27_74.t6 a_1311_424# VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.11585 ps=1.165 w=0.42 l=0.15
X27 VGND.t7 a_1474_446.t5 a_1498_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X28 VGND.t10 a_671_93.t6 a_606_87.t1 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.237825 pd=1.52 as=0.08225 ps=0.905 w=0.42 l=0.15
X29 a_671_93.t0 a_520_87.t5 a_872_119.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.192025 ps=1.335 w=0.55 l=0.15
X30 a_1311_424# a_214_74.t4 a_1318_119.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.11585 pd=1.165 as=0.05775 ps=0.76 w=0.55 l=0.15
X31 Q.t1 a_2320_410.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1918 ps=1.485 w=1.12 l=0.15
X32 VGND.t8 RESET_B.t1 a_1062_93.t1 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1303 pd=1.17 as=0.1197 ps=1.41 w=0.42 l=0.15
X33 a_520_87.t3 a_214_74.t5 a_422_125.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.11445 pd=1.21 as=0.063 ps=0.72 w=0.42 l=0.15
R0 D.n0 D.t1 331.265
R1 D.n0 D.t0 203.512
R2 D D.n0 153.94
R3 VPWR.n20 VPWR.t5 820.029
R4 VPWR.n33 VPWR.t9 761.087
R5 VPWR.n5 VPWR.n4 645.417
R6 VPWR.n14 VPWR.n13 611.795
R7 VPWR.n2 VPWR.t0 415.945
R8 VPWR.n16 VPWR.n15 243.05
R9 VPWR.n47 VPWR.n1 221.764
R10 VPWR.n4 VPWR.t7 104.364
R11 VPWR.n4 VPWR.t10 70.3576
R12 VPWR.n13 VPWR.t8 69.2583
R13 VPWR.n15 VPWR.t3 51.1307
R14 VPWR.n1 VPWR.t2 40.4559
R15 VPWR.n46 VPWR.n45 36.1417
R16 VPWR.n40 VPWR.n39 36.1417
R17 VPWR.n41 VPWR.n40 36.1417
R18 VPWR.n35 VPWR.n34 36.1417
R19 VPWR.n28 VPWR.n27 36.1417
R20 VPWR.n28 VPWR.n8 36.1417
R21 VPWR.n32 VPWR.n8 36.1417
R22 VPWR.n21 VPWR.n11 36.1417
R23 VPWR.n19 VPWR.n18 36.1417
R24 VPWR.n1 VPWR.t6 35.1791
R25 VPWR.n25 VPWR.n11 34.9704
R26 VPWR.n34 VPWR.n33 34.6358
R27 VPWR.n15 VPWR.t1 28.4473
R28 VPWR.n35 VPWR.n5 27.8593
R29 VPWR.n39 VPWR.n5 25.6005
R30 VPWR.n13 VPWR.t4 24.6255
R31 VPWR.n18 VPWR.n14 20.3299
R32 VPWR.n27 VPWR.n26 18.5533
R33 VPWR.n41 VPWR.n2 17.3181
R34 VPWR.n47 VPWR.n46 12.424
R35 VPWR.n33 VPWR.n32 9.78874
R36 VPWR.n45 VPWR.n2 9.41227
R37 VPWR.n26 VPWR.n10 9.31381
R38 VPWR.n18 VPWR.n17 9.3005
R39 VPWR.n19 VPWR.n12 9.3005
R40 VPWR.n22 VPWR.n21 9.3005
R41 VPWR.n23 VPWR.n11 9.3005
R42 VPWR.n25 VPWR.n24 9.3005
R43 VPWR.n27 VPWR.n9 9.3005
R44 VPWR.n29 VPWR.n28 9.3005
R45 VPWR.n30 VPWR.n8 9.3005
R46 VPWR.n32 VPWR.n31 9.3005
R47 VPWR.n33 VPWR.n7 9.3005
R48 VPWR.n34 VPWR.n6 9.3005
R49 VPWR.n36 VPWR.n35 9.3005
R50 VPWR.n37 VPWR.n5 9.3005
R51 VPWR.n39 VPWR.n38 9.3005
R52 VPWR.n40 VPWR.n3 9.3005
R53 VPWR.n42 VPWR.n41 9.3005
R54 VPWR.n43 VPWR.n2 9.3005
R55 VPWR.n45 VPWR.n44 9.3005
R56 VPWR.n46 VPWR.n0 9.3005
R57 VPWR.n21 VPWR.n20 8.28285
R58 VPWR.n26 VPWR.n25 7.99755
R59 VPWR.n48 VPWR.n47 7.67022
R60 VPWR.n16 VPWR.n14 7.24846
R61 VPWR.n20 VPWR.n19 3.01226
R62 VPWR.n17 VPWR.n16 0.218731
R63 VPWR VPWR.n48 0.163202
R64 VPWR.n48 VPWR.n0 0.144642
R65 VPWR.n17 VPWR.n12 0.122949
R66 VPWR.n22 VPWR.n12 0.122949
R67 VPWR.n23 VPWR.n22 0.122949
R68 VPWR.n24 VPWR.n23 0.122949
R69 VPWR.n24 VPWR.n10 0.122949
R70 VPWR.n10 VPWR.n9 0.122949
R71 VPWR.n29 VPWR.n9 0.122949
R72 VPWR.n30 VPWR.n29 0.122949
R73 VPWR.n31 VPWR.n30 0.122949
R74 VPWR.n31 VPWR.n7 0.122949
R75 VPWR.n7 VPWR.n6 0.122949
R76 VPWR.n36 VPWR.n6 0.122949
R77 VPWR.n37 VPWR.n36 0.122949
R78 VPWR.n38 VPWR.n37 0.122949
R79 VPWR.n38 VPWR.n3 0.122949
R80 VPWR.n42 VPWR.n3 0.122949
R81 VPWR.n43 VPWR.n42 0.122949
R82 VPWR.n44 VPWR.n43 0.122949
R83 VPWR.n44 VPWR.n0 0.122949
R84 a_422_125.n1 a_422_125.n0 917.688
R85 a_422_125.n1 a_422_125.t2 74.8452
R86 a_422_125.n0 a_422_125.t3 70.3576
R87 a_422_125.n0 a_422_125.t0 70.3576
R88 a_422_125.n3 a_422_125.n2 43.0194
R89 a_422_125.n2 a_422_125.t1 7.99026
R90 a_422_125.n2 a_422_125.n1 5.21789
R91 VPB.t9 VPB.t5 1011.29
R92 VPB.t14 VPB.t9 809.543
R93 VPB.t4 VPB.t1 686.962
R94 VPB.t8 VPB.t13 538.845
R95 VPB.t7 VPB.t6 495.43
R96 VPB VPB.t10 303.899
R97 VPB.t15 VPB.t11 301.344
R98 VPB.t10 VPB.t4 296.238
R99 VPB.t11 VPB.t0 275.807
R100 VPB.t12 VPB.t3 265.591
R101 VPB.t6 VPB.t2 263.038
R102 VPB.t13 VPB.t7 263.038
R103 VPB.t1 VPB.t12 229.839
R104 VPB.t0 VPB.t14 214.517
R105 VPB.t5 VPB.t8 211.963
R106 VPB.t3 VPB.t15 199.195
R107 a_27_74.n2 a_27_74.n1 1124.67
R108 a_27_74.n1 a_27_74.n0 1092.8
R109 a_27_74.n0 a_27_74.t6 812.904
R110 a_27_74.n2 a_27_74.t2 782.447
R111 a_27_74.n1 a_27_74.t3 295.091
R112 a_27_74.n4 a_27_74.t4 261.692
R113 a_27_74.t0 a_27_74.n5 232.942
R114 a_27_74.n5 a_27_74.n4 210.73
R115 a_27_74.n5 a_27_74.t1 197.76
R116 a_27_74.n3 a_27_74.t5 189.718
R117 a_27_74.n3 a_27_74.n2 83.5472
R118 a_27_74.n4 a_27_74.n3 11.7248
R119 a_520_87.n2 a_520_87.n1 604.306
R120 a_520_87.n2 a_520_87.n0 293.479
R121 a_520_87.n3 a_520_87.n2 273.057
R122 a_520_87.n0 a_520_87.t4 246.089
R123 a_520_87.n1 a_520_87.t3 177.22
R124 a_520_87.n0 a_520_87.t5 147.814
R125 a_520_87.n1 a_520_87.t1 70.3576
R126 a_520_87.n3 a_520_87.t2 40.0005
R127 a_520_87.t0 a_520_87.n3 40.0005
R128 VNB.t6 VNB.t17 3395.28
R129 VNB.t8 VNB.t1 3383.73
R130 VNB.t14 VNB.t15 2609.97
R131 VNB.t3 VNB.t0 2402.1
R132 VNB.t16 VNB.t9 1974.8
R133 VNB.t9 VNB.t5 1547.51
R134 VNB.t17 VNB.t8 1339.63
R135 VNB.t2 VNB.t7 1247.24
R136 VNB.t12 VNB.t2 1247.24
R137 VNB.t7 VNB.t13 1177.95
R138 VNB.t13 VNB.t6 1154.86
R139 VNB.t11 VNB.t3 1154.86
R140 VNB VNB.t11 1143.31
R141 VNB.t0 VNB.t4 1131.76
R142 VNB.t10 VNB.t16 1097.11
R143 VNB.t5 VNB.t14 993.177
R144 VNB.t4 VNB.t10 993.177
R145 VNB.t15 VNB.t12 831.496
R146 CLK.n0 CLK.t0 285.719
R147 CLK.n0 CLK.t1 178.34
R148 CLK CLK.n0 157.895
R149 SET_B SET_B.n2 699.643
R150 SET_B.n1 SET_B.t2 258.673
R151 SET_B.n1 SET_B.n0 231.629
R152 SET_B.n2 SET_B.t0 215.256
R153 SET_B.n2 SET_B.t1 181.784
R154 SET_B SET_B.n1 154.619
R155 a_671_93.n6 a_671_93.n5 404.423
R156 a_671_93.n2 a_671_93.n0 278.909
R157 a_671_93.n4 a_671_93.n3 246.089
R158 a_671_93.n0 a_671_93.t5 244.75
R159 a_671_93.n4 a_671_93.t4 238.371
R160 a_671_93.n2 a_671_93.n1 185
R161 a_671_93.n5 a_671_93.n4 152
R162 a_671_93.n0 a_671_93.t6 126.197
R163 a_671_93.n5 a_671_93.n2 75.1132
R164 a_671_93.n6 a_671_93.t2 56.2862
R165 a_671_93.t1 a_671_93.n6 35.1791
R166 a_671_93.n1 a_671_93.t3 30.546
R167 a_671_93.n1 a_671_93.t0 30.546
R168 a_1062_93.t0 a_1062_93.n4 739.515
R169 a_1062_93.n3 a_1062_93.t2 342.757
R170 a_1062_93.n1 a_1062_93.t1 264.077
R171 a_1062_93.n0 a_1062_93.t3 246.089
R172 a_1062_93.n4 a_1062_93.n3 243.581
R173 a_1062_93.n1 a_1062_93.n0 179.204
R174 a_1062_93.n3 a_1062_93.n2 174.323
R175 a_1062_93.n0 a_1062_93.t4 147.814
R176 a_1062_93.n4 a_1062_93.n1 3.24557
R177 a_1814_392.t0 a_1814_392.t1 52.2055
R178 a_1474_446.n1 a_1474_446.t5 468.74
R179 a_1474_446.n6 a_1474_446.n5 320.195
R180 a_1474_446.n6 a_1474_446.t1 292.454
R181 a_1474_446.n3 a_1474_446.t2 292.413
R182 a_1474_446.n3 a_1474_446.n2 284.38
R183 a_1474_446.n5 a_1474_446.t3 234.841
R184 a_1474_446.t0 a_1474_446.n7 227.647
R185 a_1474_446.n7 a_1474_446.n1 193.642
R186 a_1474_446.n4 a_1474_446.t4 186.374
R187 a_1474_446.n1 a_1474_446.n0 181.018
R188 a_1474_446.n4 a_1474_446.n3 101.513
R189 a_1474_446.n7 a_1474_446.n6 14.6496
R190 a_1474_446.n5 a_1474_446.n4 5.11262
R191 VGND.n48 VGND.t0 267.752
R192 VGND.n12 VGND.t1 258.368
R193 VGND.n14 VGND.n13 207.498
R194 VGND.n24 VGND.n21 199.739
R195 VGND.n24 VGND.n23 185
R196 VGND.n4 VGND.n3 185
R197 VGND.n32 VGND.t9 158.286
R198 VGND.n51 VGND.n50 116.29
R199 VGND.n3 VGND.t10 69.6043
R200 VGND.n3 VGND.t4 62.9003
R201 VGND.n13 VGND.t8 62.8576
R202 VGND.n22 VGND.t7 61.4291
R203 VGND.t3 VGND.n21 52.5005
R204 VGND.n13 VGND.t6 44.5565
R205 VGND.n23 VGND.t3 40.0005
R206 VGND.n16 VGND.n15 36.1417
R207 VGND.n16 VGND.n10 36.1417
R208 VGND.n20 VGND.n10 36.1417
R209 VGND.n26 VGND.n8 36.1417
R210 VGND.n30 VGND.n8 36.1417
R211 VGND.n31 VGND.n30 36.1417
R212 VGND.n33 VGND.n6 36.1417
R213 VGND.n37 VGND.n6 36.1417
R214 VGND.n38 VGND.n37 36.1417
R215 VGND.n44 VGND.n43 36.1417
R216 VGND.n44 VGND.n1 36.1417
R217 VGND.n25 VGND.n20 35.0123
R218 VGND.n49 VGND.n48 34.2593
R219 VGND.n50 VGND.t5 34.0546
R220 VGND.n43 VGND.n42 33.9237
R221 VGND.n39 VGND.n38 31.983
R222 VGND.n50 VGND.t2 22.7032
R223 VGND.n25 VGND.n24 19.2005
R224 VGND.n48 VGND.n1 19.2005
R225 VGND.n51 VGND.n49 19.2005
R226 VGND.n15 VGND.n14 18.4476
R227 VGND.n26 VGND.n25 12.424
R228 VGND.n15 VGND.n11 9.3005
R229 VGND.n17 VGND.n16 9.3005
R230 VGND.n18 VGND.n10 9.3005
R231 VGND.n20 VGND.n19 9.3005
R232 VGND.n25 VGND.n9 9.3005
R233 VGND.n27 VGND.n26 9.3005
R234 VGND.n28 VGND.n8 9.3005
R235 VGND.n30 VGND.n29 9.3005
R236 VGND.n31 VGND.n7 9.3005
R237 VGND.n34 VGND.n33 9.3005
R238 VGND.n35 VGND.n6 9.3005
R239 VGND.n37 VGND.n36 9.3005
R240 VGND.n38 VGND.n5 9.3005
R241 VGND.n40 VGND.n39 9.3005
R242 VGND.n42 VGND.n41 9.3005
R243 VGND.n43 VGND.n2 9.3005
R244 VGND.n45 VGND.n44 9.3005
R245 VGND.n46 VGND.n1 9.3005
R246 VGND.n48 VGND.n47 9.3005
R247 VGND.n49 VGND.n0 9.3005
R248 VGND.n52 VGND.n51 7.43488
R249 VGND.n14 VGND.n12 7.32935
R250 VGND.n42 VGND.n4 5.06097
R251 VGND.n33 VGND.n32 4.51815
R252 VGND.n39 VGND.n4 4.46562
R253 VGND.n32 VGND.n31 3.76521
R254 VGND.n22 VGND.n21 1.8755
R255 VGND.n23 VGND.n22 1.42907
R256 VGND.n12 VGND.n11 0.217704
R257 VGND VGND.n52 0.160103
R258 VGND.n52 VGND.n0 0.1477
R259 VGND.n17 VGND.n11 0.122949
R260 VGND.n18 VGND.n17 0.122949
R261 VGND.n19 VGND.n18 0.122949
R262 VGND.n19 VGND.n9 0.122949
R263 VGND.n27 VGND.n9 0.122949
R264 VGND.n28 VGND.n27 0.122949
R265 VGND.n29 VGND.n28 0.122949
R266 VGND.n29 VGND.n7 0.122949
R267 VGND.n34 VGND.n7 0.122949
R268 VGND.n35 VGND.n34 0.122949
R269 VGND.n36 VGND.n35 0.122949
R270 VGND.n36 VGND.n5 0.122949
R271 VGND.n40 VGND.n5 0.122949
R272 VGND.n41 VGND.n40 0.122949
R273 VGND.n41 VGND.n2 0.122949
R274 VGND.n45 VGND.n2 0.122949
R275 VGND.n46 VGND.n45 0.122949
R276 VGND.n47 VGND.n46 0.122949
R277 VGND.n47 VGND.n0 0.122949
R278 a_1318_119.t0 a_1318_119.t1 45.8187
R279 RESET_B.n0 RESET_B.t0 203.815
R280 RESET_B.n0 RESET_B.t1 173.57
R281 RESET_B RESET_B.n0 68.3813
R282 a_2320_410.t0 a_2320_410.n0 609.908
R283 a_2320_410.n0 a_2320_410.t2 267.252
R284 a_2320_410.n0 a_2320_410.t1 180.493
R285 Q.n3 Q 589.777
R286 Q.n3 Q.n0 585
R287 Q.n4 Q.n3 585
R288 Q.n2 Q.t0 285
R289 Q.t0 Q.n1 285
R290 Q.n3 Q.t1 26.3844
R291 Q Q.n4 12.8005
R292 Q.n1 Q 12.4184
R293 Q Q.n0 11.0811
R294 Q Q.n2 9.36169
R295 Q.n2 Q 4.77662
R296 Q Q.n0 3.05722
R297 Q.n1 Q 1.7199
R298 Q.n4 Q 1.33781
R299 a_1017_379.t0 a_1017_379.t1 63.3219
R300 a_872_119.t0 a_872_119.n0 607.861
R301 a_872_119.n0 a_872_119.t1 56.7278
R302 a_872_119.n0 a_872_119.t2 56.7278
R303 a_214_74.t2 a_214_74.t4 1582.57
R304 a_214_74.t4 a_214_74.t3 593.586
R305 a_214_74.n0 a_214_74.t5 335.259
R306 a_214_74.n1 a_214_74.n0 290.541
R307 a_214_74.t1 a_214_74.n1 253.284
R308 a_214_74.n0 a_214_74.t2 216.097
R309 a_214_74.n1 a_214_74.t0 160.589
R310 a_606_87.t0 a_606_87.t1 106.044
R311 a_713_379.t0 a_713_379.t1 112.572
R312 Q_N.n1 Q_N 589.707
R313 Q_N.n1 Q_N.n0 585
R314 Q_N.n2 Q_N.n1 585
R315 Q_N Q_N.t0 205.617
R316 Q_N.n1 Q_N.t1 26.3844
R317 Q_N Q_N.n2 12.6123
R318 Q_N Q_N.n0 10.9181
R319 Q_N Q_N.n0 3.01226
R320 Q_N.n2 Q_N 1.31815
R321 a_1498_74.t0 a_1498_74.t1 111.43
C0 a_1708_74# VPWR 6.98e-19
C1 VGND RESET_B 0.023956f
C2 RESET_B Q 7.57e-20
C3 D a_1311_424# 2.42e-21
C4 a_1708_74# D 2.66e-21
C5 VPB CLK 0.035267f
C6 VGND Q_N 0.084379f
C7 SET_B a_1311_424# 0.334354f
C8 VPB VPWR 0.373217f
C9 a_1708_74# SET_B 0.00616f
C10 RESET_B Q_N 0.014657f
C11 VPWR a_1203_379# 0.003601f
C12 VGND a_1311_424# 0.052576f
C13 VPB D 0.097316f
C14 a_1708_74# VGND 0.196023f
C15 CLK VPWR 0.019154f
C16 RESET_B a_1311_424# 1.42e-20
C17 VPB SET_B 0.136988f
C18 a_1708_74# RESET_B 0.001207f
C19 Q_N a_1311_424# 4.72e-20
C20 SET_B a_1203_379# 0.018413f
C21 VPWR D 0.039138f
C22 VPB VGND 0.022412f
C23 VPB Q 0.014259f
C24 VGND a_1203_379# 0.00176f
C25 VPWR SET_B 0.577555f
C26 CLK VGND 0.039479f
C27 VPB RESET_B 0.043744f
C28 a_1708_74# a_1311_424# 0.04868f
C29 VPWR VGND 0.138559f
C30 VPB Q_N 0.015351f
C31 VPWR Q 0.127503f
C32 VPWR RESET_B 0.006114f
C33 D VGND 0.009821f
C34 VPB a_1311_424# 0.051202f
C35 a_1708_74# VPB 8.38e-19
C36 SET_B VGND 0.026611f
C37 VPWR Q_N 0.074696f
C38 a_1311_424# a_1203_379# 0.004582f
C39 SET_B RESET_B 2.28e-20
C40 VGND Q 0.074385f
C41 VPWR a_1311_424# 0.021164f
C42 Q VNB 0.111702f
C43 Q_N VNB 0.01767f
C44 RESET_B VNB 0.152177f
C45 VGND VNB 1.44937f
C46 SET_B VNB 0.19908f
C47 D VNB 0.090599f
C48 VPWR VNB 1.15705f
C49 CLK VNB 0.137231f
C50 VPB VNB 2.97749f
C51 a_1708_74# VNB 0.014797f
C52 a_1311_424# VNB 0.138259f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfbbn_2 VNB VPB VPWR VGND SET_B RESET_B D CLK_N Q_N Q
X0 a_1312_424.t0 a_473_405.t4 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.2352 ps=2.24 w=0.84 l=0.15
X1 a_473_405.t0 a_601_119.t4 a_867_125.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.15675 ps=1.67 w=0.55 l=0.15
X2 a_601_119.t0 a_27_74.t2 a_529_119.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND.t6 SET_B.t0 a_867_125.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.09625 ps=0.9 w=0.55 l=0.15
X4 a_1832_74.t1 a_1335_112.t3 a_1555_410# VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2907 pd=2.39 as=0.1184 ps=1.06 w=0.74 l=0.15
X5 VPWR SET_B a_1555_410# VPB sky130_fd_pr__pfet_01v8 ad=0.269075 pd=1.705 as=0.295 ps=2.59 w=1 l=0.15
X6 a_1555_410# a_975_322.t2 a_1832_74.t2 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t9 a_975_322.t3 a_930_424.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.2 as=0.1134 ps=1.11 w=0.84 l=0.15
X8 VGND.t3 D.t0 a_311_119.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.13355 pd=1.08 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 a_200_74.t0 a_27_74.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t7 CLK_N.t0 a_27_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 a_473_405.t2 SET_B.t1 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=2.24 as=0.1512 ps=1.2 w=0.84 l=0.15
X12 a_529_119.t0 a_473_405.t5 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.13355 ps=1.08 w=0.42 l=0.15
X13 VPWR.t7 RESET_B.t0 a_975_322.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1884 pd=1.495 as=0.1792 ps=1.84 w=0.64 l=0.15
X14 a_1640_138.t0 a_200_74.t2 a_1335_112.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.305 ps=1.925 w=0.42 l=0.15
X15 a_601_119.t2 a_200_74.t3 a_536_503.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_867_125.t2 a_975_322.t4 a_473_405.t3 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.077 ps=0.83 w=0.55 l=0.15
X17 a_311_119.t0 a_27_74.t4 a_601_119.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1653 pd=1.7 as=0.0756 ps=0.78 w=0.42 l=0.15
X18 a_311_119.t3 a_200_74.t4 a_601_119.t3 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.38115 pd=2.52 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VPWR.t3 D.t1 a_311_119.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.09345 pd=0.865 as=0.17805 ps=1.75 w=0.42 l=0.15
X20 a_930_424.t1 a_601_119.t5 a_473_405.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1134 pd=1.11 as=0.2352 ps=2.24 w=0.84 l=0.15
X21 VPWR.t11 a_1555_410# a_2516_368.t0 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.2018 pd=1.49 as=0.28 ps=2.56 w=1 l=0.15
X22 Q.t3 a_2516_368.t2 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1165 ps=1.065 w=0.74 l=0.15
X23 VPWR.t10 a_1555_410# a_1504_508.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.22775 pd=2.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 Q_N.t3 a_1555_410# VGND.t10 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.237375 ps=2.01 w=0.74 l=0.15
X25 VGND.t12 a_1555_410# a_2516_368.t1 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.1824 ps=1.85 w=0.64 l=0.15
X26 VGND.t11 a_1555_410# Q_N.t2 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.222 pd=2.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 VPWR.t4 CLK_N.t1 a_27_74.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X28 a_1504_508.t0 a_27_74.t5 a_1335_112.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.14385 ps=1.23 w=0.42 l=0.15
X29 a_200_74.t1 a_27_74.t6 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 VGND.t0 a_2516_368.t3 Q.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 a_536_503.t0 a_473_405.t6 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.09345 ps=0.865 w=0.42 l=0.15
X32 a_1240_125.t0 a_473_405.t7 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.09505 pd=0.94 as=0.09625 ps=0.9 w=0.55 l=0.15
X33 VGND.t9 RESET_B.t1 a_975_322.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.237375 pd=2.01 as=0.1176 ps=1.4 w=0.42 l=0.15
X34 VPWR.t12 a_1555_410# Q_N.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X35 Q_N.t0 a_1555_410# VPWR.t13 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1884 ps=1.495 w=1.12 l=0.15
X36 a_1335_112.t2 a_200_74.t5 a_1312_424.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.14385 pd=1.23 as=0.1134 ps=1.11 w=0.84 l=0.15
X37 VPWR.t8 a_2516_368.t4 Q.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X38 a_1832_74.t0 SET_B.t2 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1338 ps=1.16 w=0.74 l=0.15
X39 Q.t0 a_2516_368.t5 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2018 ps=1.49 w=1.12 l=0.15
X40 VGND.t13 a_1555_410# a_1640_138.t1 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1338 pd=1.16 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_473_405.n0 a_473_405.t5 416.127
R1 a_473_405.n2 a_473_405.t2 331.601
R2 a_473_405.t1 a_473_405.n5 324.553
R3 a_473_405.n5 a_473_405.n0 322.752
R4 a_473_405.n4 a_473_405.n3 285.243
R5 a_473_405.n1 a_473_405.t7 247.72
R6 a_473_405.n1 a_473_405.t4 221.257
R7 a_473_405.n2 a_473_405.n1 187.332
R8 a_473_405.n0 a_473_405.t6 138.441
R9 a_473_405.n4 a_473_405.n2 60.2358
R10 a_473_405.n3 a_473_405.t3 30.546
R11 a_473_405.n3 a_473_405.t0 30.546
R12 a_473_405.n5 a_473_405.n4 6.33257
R13 VPWR.n39 VPWR.t2 775.191
R14 VPWR.n32 VPWR.t10 759.761
R15 VPWR.n54 VPWR.n53 623.024
R16 VPWR.n24 VPWR.n14 607.417
R17 VPWR.n45 VPWR.n6 606.333
R18 VPWR.n16 VPWR.t8 359.115
R19 VPWR.n15 VPWR.t12 343.255
R20 VPWR.n61 VPWR.n1 331.5
R21 VPWR.n18 VPWR.n17 237.327
R22 VPWR.n53 VPWR.t3 138.369
R23 VPWR.n14 VPWR.t7 70.7974
R24 VPWR.n53 VPWR.t1 70.3576
R25 VPWR.n6 VPWR.t6 49.2505
R26 VPWR.n17 VPWR.t11 43.3405
R27 VPWR.n47 VPWR.n46 36.1417
R28 VPWR.n47 VPWR.n4 36.1417
R29 VPWR.n51 VPWR.n4 36.1417
R30 VPWR.n52 VPWR.n51 36.1417
R31 VPWR.n55 VPWR.n52 36.1417
R32 VPWR.n59 VPWR.n2 36.1417
R33 VPWR.n60 VPWR.n59 36.1417
R34 VPWR.n61 VPWR.n60 36.1417
R35 VPWR.n44 VPWR.n7 36.1417
R36 VPWR.n37 VPWR.n9 36.1417
R37 VPWR.n38 VPWR.n37 36.1417
R38 VPWR.n40 VPWR.n38 36.1417
R39 VPWR.n33 VPWR.n31 36.1417
R40 VPWR.n26 VPWR.n25 36.1417
R41 VPWR.n26 VPWR.n11 36.1417
R42 VPWR.n6 VPWR.t9 35.1791
R43 VPWR.n30 VPWR.n11 32.6519
R44 VPWR.n19 VPWR.n15 28.2358
R45 VPWR.n17 VPWR.t5 27.2944
R46 VPWR.n1 VPWR.t0 26.3844
R47 VPWR.n1 VPWR.t4 26.3844
R48 VPWR.n19 VPWR.n18 25.977
R49 VPWR.n14 VPWR.t13 25.505
R50 VPWR.n31 VPWR.n30 24.2765
R51 VPWR.n25 VPWR.n24 23.7181
R52 VPWR.n24 VPWR.n23 23.7181
R53 VPWR.n55 VPWR.n54 19.577
R54 VPWR.n23 VPWR.n15 19.2005
R55 VPWR.n54 VPWR.n2 16.5652
R56 VPWR.n32 VPWR.n9 11.523
R57 VPWR.n45 VPWR.n44 10.1652
R58 VPWR.n20 VPWR.n19 9.3005
R59 VPWR.n21 VPWR.n15 9.3005
R60 VPWR.n23 VPWR.n22 9.3005
R61 VPWR.n24 VPWR.n13 9.3005
R62 VPWR.n25 VPWR.n12 9.3005
R63 VPWR.n27 VPWR.n26 9.3005
R64 VPWR.n28 VPWR.n11 9.3005
R65 VPWR.n30 VPWR.n29 9.3005
R66 VPWR.n31 VPWR.n10 9.3005
R67 VPWR.n34 VPWR.n33 9.3005
R68 VPWR.n35 VPWR.n9 9.3005
R69 VPWR.n37 VPWR.n36 9.3005
R70 VPWR.n38 VPWR.n8 9.3005
R71 VPWR.n41 VPWR.n40 9.3005
R72 VPWR.n42 VPWR.n7 9.3005
R73 VPWR.n44 VPWR.n43 9.3005
R74 VPWR.n46 VPWR.n5 9.3005
R75 VPWR.n48 VPWR.n47 9.3005
R76 VPWR.n49 VPWR.n4 9.3005
R77 VPWR.n51 VPWR.n50 9.3005
R78 VPWR.n52 VPWR.n3 9.3005
R79 VPWR.n56 VPWR.n55 9.3005
R80 VPWR.n57 VPWR.n2 9.3005
R81 VPWR.n59 VPWR.n58 9.3005
R82 VPWR.n60 VPWR.n0 9.3005
R83 VPWR.n33 VPWR.n32 9.26421
R84 VPWR.n62 VPWR.n61 7.70379
R85 VPWR.n39 VPWR.n7 7.15344
R86 VPWR.n18 VPWR.n16 6.92649
R87 VPWR.n40 VPWR.n39 4.14168
R88 VPWR.n46 VPWR.n45 1.12991
R89 VPWR.n20 VPWR.n16 0.547078
R90 VPWR VPWR.n62 0.163644
R91 VPWR.n62 VPWR.n0 0.144205
R92 VPWR.n21 VPWR.n20 0.122949
R93 VPWR.n22 VPWR.n21 0.122949
R94 VPWR.n22 VPWR.n13 0.122949
R95 VPWR.n13 VPWR.n12 0.122949
R96 VPWR.n27 VPWR.n12 0.122949
R97 VPWR.n28 VPWR.n27 0.122949
R98 VPWR.n29 VPWR.n28 0.122949
R99 VPWR.n29 VPWR.n10 0.122949
R100 VPWR.n34 VPWR.n10 0.122949
R101 VPWR.n35 VPWR.n34 0.122949
R102 VPWR.n36 VPWR.n35 0.122949
R103 VPWR.n36 VPWR.n8 0.122949
R104 VPWR.n41 VPWR.n8 0.122949
R105 VPWR.n42 VPWR.n41 0.122949
R106 VPWR.n43 VPWR.n42 0.122949
R107 VPWR.n43 VPWR.n5 0.122949
R108 VPWR.n48 VPWR.n5 0.122949
R109 VPWR.n49 VPWR.n48 0.122949
R110 VPWR.n50 VPWR.n49 0.122949
R111 VPWR.n50 VPWR.n3 0.122949
R112 VPWR.n56 VPWR.n3 0.122949
R113 VPWR.n57 VPWR.n56 0.122949
R114 VPWR.n58 VPWR.n57 0.122949
R115 VPWR.n58 VPWR.n0 0.122949
R116 a_1312_424.t0 a_1312_424.t1 63.3219
R117 VPB.t17 VPB.t10 1590.99
R118 VPB.t0 VPB.t5 543.952
R119 VPB.t1 VPB.t7 531.183
R120 VPB.t16 VPB.t18 500.538
R121 VPB.t9 VPB.t4 500.538
R122 VPB.t5 VPB.t3 303.899
R123 VPB.t12 VPB.t2 275.807
R124 VPB.t10 VPB.t15 268.146
R125 VPB.t18 VPB.t8 265.591
R126 VPB.t13 VPB.t9 260.485
R127 VPB.t14 VPB.t1 260.485
R128 VPB VPB.t6 252.823
R129 VPB.t8 VPB.t11 229.839
R130 VPB.t15 VPB.t16 229.839
R131 VPB.t6 VPB.t0 229.839
R132 VPB.t2 VPB.t17 214.517
R133 VPB.t4 VPB.t12 214.517
R134 VPB.t7 VPB.t13 214.517
R135 VPB.t3 VPB.t14 214.517
R136 a_601_119.n2 a_601_119.n1 679.027
R137 a_601_119.n3 a_601_119.n2 266.161
R138 a_601_119.n2 a_601_119.n0 243.743
R139 a_601_119.n0 a_601_119.t5 226.005
R140 a_601_119.n0 a_601_119.t4 163.898
R141 a_601_119.n1 a_601_119.t1 84.4291
R142 a_601_119.n1 a_601_119.t2 84.4291
R143 a_601_119.n3 a_601_119.t3 40.0005
R144 a_601_119.t0 a_601_119.n3 40.0005
R145 a_867_125.n0 a_867_125.t1 503.904
R146 a_867_125.n0 a_867_125.t2 45.8187
R147 a_867_125.t0 a_867_125.n0 30.546
R148 VNB.t5 VNB.t3 4619.42
R149 VNB.t16 VNB.t2 3083.46
R150 VNB.t12 VNB.t13 2436.75
R151 VNB.t18 VNB.t19 2321.26
R152 VNB.t9 VNB.t7 2286.61
R153 VNB.t7 VNB.t6 1512.86
R154 VNB.t17 VNB.t8 1316.54
R155 VNB.t13 VNB.t20 1247.24
R156 VNB.t1 VNB.t5 1154.86
R157 VNB.t15 VNB.t1 1154.86
R158 VNB VNB.t10 1143.31
R159 VNB.t19 VNB.t11 1097.11
R160 VNB.t14 VNB.t12 1085.56
R161 VNB.t11 VNB.t0 993.177
R162 VNB.t20 VNB.t18 993.177
R163 VNB.t8 VNB.t14 993.177
R164 VNB.t2 VNB.t15 993.177
R165 VNB.t4 VNB.t16 993.177
R166 VNB.t10 VNB.t9 993.177
R167 VNB.t3 VNB.t17 900.788
R168 VNB.t6 VNB.t4 831.496
R169 a_27_74.n1 a_27_74.n0 1365.67
R170 a_27_74.t6 a_27_74.n1 800.12
R171 a_27_74.n0 a_27_74.t5 782.332
R172 a_27_74.t2 a_27_74.t4 720.859
R173 a_27_74.t0 a_27_74.n3 284.483
R174 a_27_74.n2 a_27_74.t3 264.298
R175 a_27_74.n2 a_27_74.t6 204.048
R176 a_27_74.n3 a_27_74.t1 196.087
R177 a_27_74.n1 a_27_74.t2 176.733
R178 a_27_74.n3 a_27_74.n2 152
R179 a_529_119.t0 a_529_119.t1 60.0005
R180 SET_B.n2 SET_B.t0 258.673
R181 SET_B.n1 SET_B.t2 252.248
R182 SET_B.n1 SET_B.n0 236.983
R183 SET_B.n2 SET_B.t1 205.922
R184 SET_B SET_B.n1 180.885
R185 SET_B SET_B.n2 173.463
R186 VGND.n28 VGND.n27 361.13
R187 VGND.n17 VGND.t0 311.671
R188 VGND.n36 VGND.n11 224.429
R189 VGND.n7 VGND.n6 218.358
R190 VGND.n62 VGND.n61 209.243
R191 VGND.n2 VGND.n1 207.338
R192 VGND.n27 VGND.n26 185
R193 VGND.n16 VGND.t11 176.054
R194 VGND.n19 VGND.n18 119.867
R195 VGND.n11 VGND.t13 79.3832
R196 VGND.n15 VGND.t9 75.7148
R197 VGND.n1 VGND.t2 72.8576
R198 VGND.n1 VGND.t3 71.4291
R199 VGND.n6 VGND.t6 45.8187
R200 VGND.n27 VGND.n15 36.2908
R201 VGND.n30 VGND.n12 36.1417
R202 VGND.n34 VGND.n12 36.1417
R203 VGND.n35 VGND.n34 36.1417
R204 VGND.n37 VGND.n9 36.1417
R205 VGND.n41 VGND.n9 36.1417
R206 VGND.n42 VGND.n41 36.1417
R207 VGND.n43 VGND.n42 36.1417
R208 VGND.n48 VGND.n47 36.1417
R209 VGND.n49 VGND.n48 36.1417
R210 VGND.n49 VGND.n4 36.1417
R211 VGND.n53 VGND.n4 36.1417
R212 VGND.n54 VGND.n53 36.1417
R213 VGND.n55 VGND.n54 36.1417
R214 VGND.n60 VGND.n59 36.1417
R215 VGND.n37 VGND.n36 35.3887
R216 VGND.n18 VGND.t12 31.8755
R217 VGND.n6 VGND.t1 30.546
R218 VGND.n43 VGND.n7 30.4946
R219 VGND.n25 VGND.n16 29.7417
R220 VGND.n30 VGND.n29 28.9308
R221 VGND.n20 VGND.n19 28.2358
R222 VGND.n59 VGND.n2 27.4829
R223 VGND.n26 VGND.n25 26.9519
R224 VGND.n18 VGND.t8 25.4736
R225 VGND.n62 VGND.n60 24.4711
R226 VGND.n20 VGND.n16 23.7181
R227 VGND.n11 VGND.t5 22.7037
R228 VGND.n61 VGND.t4 22.7032
R229 VGND.n61 VGND.t7 22.7032
R230 VGND.n15 VGND.t10 20.2708
R231 VGND.n47 VGND.n7 16.9417
R232 VGND.n55 VGND.n2 15.0593
R233 VGND.n28 VGND.n14 9.84665
R234 VGND.n60 VGND.n0 9.3005
R235 VGND.n59 VGND.n58 9.3005
R236 VGND.n57 VGND.n2 9.3005
R237 VGND.n56 VGND.n55 9.3005
R238 VGND.n54 VGND.n3 9.3005
R239 VGND.n53 VGND.n52 9.3005
R240 VGND.n51 VGND.n4 9.3005
R241 VGND.n50 VGND.n49 9.3005
R242 VGND.n48 VGND.n5 9.3005
R243 VGND.n47 VGND.n46 9.3005
R244 VGND.n45 VGND.n7 9.3005
R245 VGND.n44 VGND.n43 9.3005
R246 VGND.n42 VGND.n8 9.3005
R247 VGND.n41 VGND.n40 9.3005
R248 VGND.n39 VGND.n9 9.3005
R249 VGND.n38 VGND.n37 9.3005
R250 VGND.n35 VGND.n10 9.3005
R251 VGND.n34 VGND.n33 9.3005
R252 VGND.n32 VGND.n12 9.3005
R253 VGND.n31 VGND.n30 9.3005
R254 VGND.n29 VGND.n13 9.3005
R255 VGND.n23 VGND.n14 9.3005
R256 VGND.n25 VGND.n24 9.3005
R257 VGND.n22 VGND.n16 9.3005
R258 VGND.n21 VGND.n20 9.3005
R259 VGND.n63 VGND.n62 7.19894
R260 VGND.n19 VGND.n17 6.60325
R261 VGND.n36 VGND.n35 0.753441
R262 VGND.n29 VGND.n28 0.65691
R263 VGND.n21 VGND.n17 0.655275
R264 VGND VGND.n63 0.156997
R265 VGND.n63 VGND.n0 0.150766
R266 VGND.n22 VGND.n21 0.122949
R267 VGND.n24 VGND.n22 0.122949
R268 VGND.n24 VGND.n23 0.122949
R269 VGND.n23 VGND.n13 0.122949
R270 VGND.n31 VGND.n13 0.122949
R271 VGND.n32 VGND.n31 0.122949
R272 VGND.n33 VGND.n32 0.122949
R273 VGND.n33 VGND.n10 0.122949
R274 VGND.n38 VGND.n10 0.122949
R275 VGND.n39 VGND.n38 0.122949
R276 VGND.n40 VGND.n39 0.122949
R277 VGND.n40 VGND.n8 0.122949
R278 VGND.n44 VGND.n8 0.122949
R279 VGND.n45 VGND.n44 0.122949
R280 VGND.n46 VGND.n45 0.122949
R281 VGND.n46 VGND.n5 0.122949
R282 VGND.n50 VGND.n5 0.122949
R283 VGND.n51 VGND.n50 0.122949
R284 VGND.n52 VGND.n51 0.122949
R285 VGND.n52 VGND.n3 0.122949
R286 VGND.n56 VGND.n3 0.122949
R287 VGND.n57 VGND.n56 0.122949
R288 VGND.n58 VGND.n57 0.122949
R289 VGND.n58 VGND.n0 0.122949
R290 VGND.n26 VGND.n14 0.109902
R291 a_1335_112.t2 a_1335_112.n2 418.055
R292 a_1335_112.n2 a_1335_112.n1 349.118
R293 a_1335_112.n1 a_1335_112.t3 258.673
R294 a_1335_112.n1 a_1335_112.n0 231.629
R295 a_1335_112.n2 a_1335_112.t0 205.155
R296 a_1335_112.t2 a_1335_112.t1 113.599
R297 a_1832_74.n0 a_1832_74.t1 556.125
R298 a_1832_74.n0 a_1832_74.t2 22.7032
R299 a_1832_74.t0 a_1832_74.n0 22.7032
R300 a_975_322.t1 a_975_322.n4 711.361
R301 a_975_322.n3 a_975_322.n0 587.611
R302 a_975_322.n2 a_975_322.n1 298.572
R303 a_975_322.n4 a_975_322.t0 252.482
R304 a_975_322.n0 a_975_322.t4 252.248
R305 a_975_322.n0 a_975_322.t3 211.278
R306 a_975_322.n2 a_975_322.t2 178.34
R307 a_975_322.n3 a_975_322.n2 152
R308 a_975_322.n4 a_975_322.n3 61.1351
R309 a_930_424.t0 a_930_424.t1 63.3219
R310 D.n0 D.t1 358.486
R311 D.n1 D.n0 152
R312 D.n0 D.t0 138.373
R313 D.n1 D 16.8732
R314 D D.n1 1.74595
R315 a_311_119.n0 a_311_119.t0 856.856
R316 a_311_119.n1 a_311_119.t1 817.038
R317 a_311_119.n0 a_311_119.t3 258.81
R318 a_311_119.t2 a_311_119.n1 231.912
R319 a_311_119.n1 a_311_119.n0 164.089
R320 a_200_74.n0 a_200_74.t5 388.765
R321 a_200_74.n0 a_200_74.t2 351.704
R322 a_200_74.n2 a_200_74.t3 311.524
R323 a_200_74.n1 a_200_74.t4 289.012
R324 a_200_74.n3 a_200_74.t1 217.465
R325 a_200_74.t0 a_200_74.n3 216.137
R326 a_200_74.n3 a_200_74.n2 211.18
R327 a_200_74.n1 a_200_74.n0 21.9278
R328 a_200_74.n2 a_200_74.n1 17.5456
R329 CLK_N.n0 CLK_N.t1 259.132
R330 CLK_N.n0 CLK_N.t0 198.882
R331 CLK_N CLK_N.n0 156.667
R332 RESET_B.n0 RESET_B.t0 173.788
R333 RESET_B RESET_B.n0 158.995
R334 RESET_B.n0 RESET_B.t1 126.927
R335 a_1640_138.t0 a_1640_138.t1 68.5719
R336 a_536_503.t0 a_536_503.t1 126.644
R337 a_2516_368.n1 a_2516_368.t5 253.343
R338 a_2516_368.t0 a_2516_368.n3 250.364
R339 a_2516_368.n0 a_2516_368.t4 248.231
R340 a_2516_368.n3 a_2516_368.n2 181.868
R341 a_2516_368.n0 a_2516_368.t3 172.499
R342 a_2516_368.n1 a_2516_368.t2 170.308
R343 a_2516_368.n3 a_2516_368.t1 155.846
R344 a_2516_368.n2 a_2516_368.n0 54.7732
R345 a_2516_368.n2 a_2516_368.n1 5.84292
R346 Q.n2 Q 589.85
R347 Q.n2 Q.n0 585
R348 Q.n3 Q.n2 585
R349 Q Q.n1 169.084
R350 Q.n2 Q.t1 26.3844
R351 Q.n2 Q.t0 26.3844
R352 Q.n1 Q.t2 22.7032
R353 Q.n1 Q.t3 22.7032
R354 Q Q.n3 12.9944
R355 Q Q.n0 11.249
R356 Q Q.n0 3.10353
R357 Q.n3 Q 1.35808
R358 a_1504_508.t0 a_1504_508.t1 126.644
R359 Q_N.n1 Q_N.n0 280.01
R360 Q_N.n2 Q_N.n1 185
R361 Q_N.n3 Q_N.n2 185
R362 Q_N.n0 Q_N.t1 26.3844
R363 Q_N.n0 Q_N.t0 26.3844
R364 Q_N.n2 Q_N.t2 22.7032
R365 Q_N.n2 Q_N.t3 22.7032
R366 Q_N Q_N.n3 7.03149
R367 Q_N Q_N.n1 6.31036
R368 Q_N.n3 Q_N 6.31036
R369 a_1240_125.n0 a_1240_125.t0 58.2266
C0 Q_N a_1555_410# 0.213875f
C1 VPB SET_B 0.1333f
C2 VPWR D 0.005151f
C3 Q a_1555_410# 0.002437f
C4 VPWR a_1931_392# 0.002476f
C5 VPB VGND 0.025156f
C6 VPWR SET_B 0.162483f
C7 VPB RESET_B 0.044984f
C8 CLK_N SET_B 1.13e-20
C9 VPWR VGND 0.152967f
C10 D SET_B 2.05e-20
C11 VPWR RESET_B 0.005604f
C12 VPB Q_N 0.007219f
C13 CLK_N VGND 0.017214f
C14 VPB a_1555_410# 0.337971f
C15 SET_B a_1931_392# 4.85e-19
C16 VPB Q 0.0089f
C17 D VGND 0.011675f
C18 VPWR Q_N 0.118365f
C19 VPWR a_1555_410# 0.38687f
C20 VGND a_1931_392# 7.13e-19
C21 SET_B VGND 0.06728f
C22 VPWR Q 0.200926f
C23 SET_B RESET_B 2.09e-19
C24 VGND RESET_B 0.006023f
C25 SET_B Q_N 2.22e-19
C26 a_1555_410# a_1931_392# 0.009561f
C27 SET_B a_1555_410# 0.097856f
C28 VPB VPWR 0.414842f
C29 SET_B Q 6.02e-20
C30 VGND Q_N 0.108641f
C31 VGND a_1555_410# 0.171636f
C32 VPB CLK_N 0.039657f
C33 RESET_B Q_N 0.001182f
C34 VGND Q 0.132764f
C35 RESET_B a_1555_410# 0.111543f
C36 VPWR CLK_N 0.01506f
C37 VPB D 0.100032f
C38 RESET_B Q 9.33e-20
C39 Q VNB 0.057529f
C40 Q_N VNB 0.012295f
C41 RESET_B VNB 0.110096f
C42 VGND VNB 1.61643f
C43 SET_B VNB 0.208552f
C44 D VNB 0.142698f
C45 CLK_N VNB 0.161399f
C46 VPWR VNB 1.30819f
C47 VPB VNB 3.2989f
C48 a_1555_410# VNB 0.505581f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfbbn_1 VNB VPB VPWR SET_B VGND Q D RESET_B CLK_N Q_N
X0 a_933_424.t0 a_595_119.t4 a_474_405.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1008 pd=1.08 as=0.2352 ps=2.24 w=0.84 l=0.15
X1 a_595_119.t1 a_27_74.t2 a_523_119.t0 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_1349_114# a_27_74.t3 a_1254_119.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.314125 pd=1.71 as=0.09155 ps=0.9 w=0.55 l=0.15
X3 a_1818_76.t2 SET_B.t0 VGND.t9 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.14955 ps=1.235 w=0.74 l=0.15
X4 a_1818_76.t1 a_1349_114# a_1534_446.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.296 pd=2.52 as=0.1184 ps=1.06 w=0.74 l=0.15
X5 VGND.t2 D.t0 a_311_119.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.137925 pd=1.13 as=0.1197 ps=1.41 w=0.42 l=0.15
X6 VGND.t8 SET_B.t1 a_867_119.t2 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.09625 ps=0.9 w=0.55 l=0.15
X7 a_200_74.t1 a_27_74.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VGND.t0 CLK_N.t0 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_523_119.t1 a_474_405.t4 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.137925 ps=1.13 w=0.42 l=0.15
X10 a_311_119.t1 a_200_74.t2 a_595_119.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.40005 pd=2.58 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_1297_424# a_474_405.t5 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1008 pd=1.08 as=0.2352 ps=2.24 w=0.84 l=0.15
X12 VPWR.t7 D.t1 a_311_119.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0945 pd=0.87 as=0.17805 ps=1.75 w=0.42 l=0.15
X13 a_1534_446.t2 a_1349_114# a_1917_392.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X14 Q_N.t0 a_1534_446.t4 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.1884 ps=1.495 w=1.12 l=0.15
X15 Q_N.t1 a_1534_446.t5 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.172025 ps=1.385 w=0.74 l=0.15
X16 Q.t1 a_2412_410.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.11565 ps=1.085 w=0.74 l=0.15
X17 a_867_119.t0 a_978_357.t2 a_474_405.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.09625 ps=0.9 w=0.55 l=0.15
X18 a_595_119.t2 a_200_74.t3 a_537_503.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1917_392.t0 a_978_357.t3 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.269075 ps=1.705 w=1 l=0.15
X20 a_311_119.t0 a_27_74.t5 a_595_119.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1704 pd=1.72 as=0.0756 ps=0.78 w=0.42 l=0.15
X21 VGND.t4 RESET_B.t0 a_978_357.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.172025 pd=1.385 as=0.1134 ps=1.38 w=0.42 l=0.15
X22 VPWR.t12 a_978_357.t4 a_933_424.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1008 ps=1.08 w=0.84 l=0.15
X23 VPWR.t6 CLK_N.t1 a_27_74.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X24 a_474_405.t0 SET_B.t2 VPWR.t9 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=2.24 as=0.126 ps=1.14 w=0.84 l=0.15
X25 VPWR.t8 SET_B.t3 a_1534_446.t3 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.269075 pd=1.705 as=0.295 ps=2.59 w=1 l=0.15
X26 a_200_74.t0 a_27_74.t6 VGND.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 VGND.t7 a_1534_446.t6 a_2412_410.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.11565 pd=1.085 as=0.1134 ps=1.38 w=0.42 l=0.15
X28 a_474_405.t3 a_595_119.t5 a_867_119.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.15675 ps=1.67 w=0.55 l=0.15
X29 a_1534_446.t0 a_978_357.t5 a_1818_76.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X30 VPWR.t4 a_1534_446.t7 a_2412_410.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1974 pd=1.495 as=0.2394 ps=2.25 w=0.84 l=0.15
X31 VPWR.t0 RESET_B.t1 a_978_357.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1884 pd=1.495 as=0.1792 ps=1.84 w=0.64 l=0.15
X32 VGND.t5 a_1534_446.t8 a_1611_140.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.14955 pd=1.235 as=0.0504 ps=0.66 w=0.42 l=0.15
X33 a_537_503.t1 a_474_405.t6 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X34 a_1254_119.t1 a_474_405.t7 VGND.t11 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.09155 pd=0.9 as=0.09625 ps=0.9 w=0.55 l=0.15
X35 Q.t0 a_2412_410.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1974 ps=1.495 w=1.12 l=0.15
R0 a_200_74.n2 a_200_74.n1 375.502
R1 a_200_74.n2 a_200_74.n0 312.223
R2 a_200_74.n4 a_200_74.t3 310.728
R3 a_200_74.n3 a_200_74.t2 287.849
R4 a_200_74.n5 a_200_74.t0 219.405
R5 a_200_74.t1 a_200_74.n5 215.762
R6 a_200_74.n5 a_200_74.n4 214.659
R7 a_200_74.n3 a_200_74.n2 21.9278
R8 a_200_74.n4 a_200_74.n3 15.7974
R9 VNB.t17 VNB.t5 3926.51
R10 VNB.t12 VNB.t11 3152.76
R11 VNB.t13 VNB.t4 2367.45
R12 VNB.t9 VNB.t1 2286.61
R13 VNB.t6 VNB.t8 2217.32
R14 VNB.t5 VNB.t10 1489.76
R15 VNB.t1 VNB.t14 1443.57
R16 VNB.t4 VNB.t6 1304.99
R17 VNB.t15 VNB.t18 1154.86
R18 VNB.t2 VNB.t15 1154.86
R19 VNB.t11 VNB.t2 1154.86
R20 VNB.t8 VNB.t3 1143.31
R21 VNB VNB.t0 1143.31
R22 VNB.t18 VNB.t17 1097.11
R23 VNB.t7 VNB.t13 1085.56
R24 VNB.t10 VNB.t7 993.177
R25 VNB.t16 VNB.t12 993.177
R26 VNB.t0 VNB.t9 993.177
R27 VNB.t14 VNB.t16 831.496
R28 a_27_74.n1 a_27_74.t3 1401.01
R29 a_27_74.t6 a_27_74.n1 790.481
R30 a_27_74.t2 a_27_74.t5 744.154
R31 a_27_74.t3 a_27_74.n0 738.799
R32 a_27_74.t1 a_27_74.n3 284.834
R33 a_27_74.n2 a_27_74.t4 264.298
R34 a_27_74.n2 a_27_74.t6 204.048
R35 a_27_74.n3 a_27_74.t0 196.438
R36 a_27_74.n1 a_27_74.t2 176.733
R37 a_27_74.n3 a_27_74.n2 152
R38 VPB.t13 VPB.t15 1266.67
R39 VPB.t2 VPB.t9 543.952
R40 VPB.t1 VPB.t10 536.29
R41 VPB.t7 VPB.t8 503.091
R42 VPB.t12 VPB.t0 500.538
R43 VPB.t4 VPB.t13 500.538
R44 VPB.t15 VPB.t5 316.668
R45 VPB.t9 VPB.t14 306.452
R46 VPB.t8 VPB.t3 268.146
R47 VPB.t0 VPB.t7 268.146
R48 VPB.t11 VPB.t1 260.485
R49 VPB VPB.t6 252.823
R50 VPB.t16 VPB.t4 229.839
R51 VPB.t6 VPB.t2 229.839
R52 VPB.t5 VPB.t12 214.517
R53 VPB.t14 VPB.t11 214.517
R54 VPB.t10 VPB.t16 199.195
R55 a_595_119.n2 a_595_119.n1 672.049
R56 a_595_119.n2 a_595_119.n0 328.861
R57 a_595_119.n0 a_595_119.t4 292.95
R58 a_595_119.n3 a_595_119.n2 257.125
R59 a_595_119.n0 a_595_119.t5 202.44
R60 a_595_119.n1 a_595_119.t0 84.4291
R61 a_595_119.n1 a_595_119.t2 84.4291
R62 a_595_119.n3 a_595_119.t3 40.0005
R63 a_595_119.t1 a_595_119.n3 40.0005
R64 a_474_405.n2 a_474_405.t4 416.127
R65 a_474_405.t0 a_474_405.n5 332.834
R66 a_474_405.n3 a_474_405.n2 326.844
R67 a_474_405.n3 a_474_405.t2 323.712
R68 a_474_405.n4 a_474_405.n1 284.993
R69 a_474_405.n0 a_474_405.t7 265.142
R70 a_474_405.n0 a_474_405.t5 202.75
R71 a_474_405.n5 a_474_405.n0 198.25
R72 a_474_405.n2 a_474_405.t6 138.441
R73 a_474_405.n5 a_474_405.n4 62.7286
R74 a_474_405.n1 a_474_405.t3 45.8187
R75 a_474_405.n1 a_474_405.t1 30.546
R76 a_474_405.n4 a_474_405.n3 21.8738
R77 a_933_424.t0 a_933_424.t1 56.2862
R78 a_523_119.t0 a_523_119.t1 60.0005
R79 a_1254_119.n0 a_1254_119.t1 40.2203
R80 a_1254_119.n0 a_1254_119.t0 23.0774
R81 a_1254_119.n1 a_1254_119.n0 7.2005
R82 SET_B.n0 SET_B.t3 290.539
R83 SET_B.n1 SET_B.t1 268.313
R84 SET_B.n1 SET_B.t2 207.138
R85 SET_B SET_B.n0 185.395
R86 SET_B.n0 SET_B.t0 184.745
R87 SET_B SET_B.n1 174.042
R88 VGND.n17 VGND.n16 251.679
R89 VGND.n2 VGND.n1 235.94
R90 VGND.n25 VGND.n11 221.793
R91 VGND.n15 VGND.n14 221.008
R92 VGND.n7 VGND.n6 218.745
R93 VGND.n51 VGND.n50 209.243
R94 VGND.n11 VGND.t5 100.811
R95 VGND.n16 VGND.t4 70.0005
R96 VGND.n1 VGND.t10 68.5719
R97 VGND.n1 VGND.t2 67.1434
R98 VGND.n14 VGND.t7 58.5719
R99 VGND.n6 VGND.t8 45.8187
R100 VGND.n19 VGND.n18 36.1417
R101 VGND.n19 VGND.n12 36.1417
R102 VGND.n23 VGND.n12 36.1417
R103 VGND.n24 VGND.n23 36.1417
R104 VGND.n26 VGND.n9 36.1417
R105 VGND.n30 VGND.n9 36.1417
R106 VGND.n31 VGND.n30 36.1417
R107 VGND.n32 VGND.n31 36.1417
R108 VGND.n37 VGND.n36 36.1417
R109 VGND.n38 VGND.n37 36.1417
R110 VGND.n38 VGND.n4 36.1417
R111 VGND.n42 VGND.n4 36.1417
R112 VGND.n43 VGND.n42 36.1417
R113 VGND.n44 VGND.n43 36.1417
R114 VGND.n49 VGND.n48 36.1417
R115 VGND.n6 VGND.t11 30.546
R116 VGND.n26 VGND.n25 30.1181
R117 VGND.n16 VGND.t6 27.5681
R118 VGND.n48 VGND.n2 27.4829
R119 VGND.n32 VGND.n7 25.224
R120 VGND.n51 VGND.n49 24.4711
R121 VGND.n14 VGND.t3 23.321
R122 VGND.n11 VGND.t9 22.7037
R123 VGND.n50 VGND.t1 22.7032
R124 VGND.n50 VGND.t0 22.7032
R125 VGND.n36 VGND.n7 22.2123
R126 VGND.n18 VGND.n17 19.2005
R127 VGND.n44 VGND.n2 17.3181
R128 VGND.n49 VGND.n0 9.3005
R129 VGND.n48 VGND.n47 9.3005
R130 VGND.n46 VGND.n2 9.3005
R131 VGND.n45 VGND.n44 9.3005
R132 VGND.n43 VGND.n3 9.3005
R133 VGND.n42 VGND.n41 9.3005
R134 VGND.n40 VGND.n4 9.3005
R135 VGND.n39 VGND.n38 9.3005
R136 VGND.n37 VGND.n5 9.3005
R137 VGND.n36 VGND.n35 9.3005
R138 VGND.n34 VGND.n7 9.3005
R139 VGND.n18 VGND.n13 9.3005
R140 VGND.n20 VGND.n19 9.3005
R141 VGND.n21 VGND.n12 9.3005
R142 VGND.n23 VGND.n22 9.3005
R143 VGND.n24 VGND.n10 9.3005
R144 VGND.n27 VGND.n26 9.3005
R145 VGND.n28 VGND.n9 9.3005
R146 VGND.n30 VGND.n29 9.3005
R147 VGND.n31 VGND.n8 9.3005
R148 VGND.n33 VGND.n32 9.3005
R149 VGND.n17 VGND.n15 7.30311
R150 VGND.n52 VGND.n51 7.19894
R151 VGND.n25 VGND.n24 6.02403
R152 VGND.n15 VGND.n13 0.212973
R153 VGND VGND.n52 0.156997
R154 VGND.n52 VGND.n0 0.150766
R155 VGND.n20 VGND.n13 0.122949
R156 VGND.n21 VGND.n20 0.122949
R157 VGND.n22 VGND.n21 0.122949
R158 VGND.n22 VGND.n10 0.122949
R159 VGND.n27 VGND.n10 0.122949
R160 VGND.n28 VGND.n27 0.122949
R161 VGND.n29 VGND.n28 0.122949
R162 VGND.n29 VGND.n8 0.122949
R163 VGND.n33 VGND.n8 0.122949
R164 VGND.n34 VGND.n33 0.122949
R165 VGND.n35 VGND.n34 0.122949
R166 VGND.n35 VGND.n5 0.122949
R167 VGND.n39 VGND.n5 0.122949
R168 VGND.n40 VGND.n39 0.122949
R169 VGND.n41 VGND.n40 0.122949
R170 VGND.n41 VGND.n3 0.122949
R171 VGND.n45 VGND.n3 0.122949
R172 VGND.n46 VGND.n45 0.122949
R173 VGND.n47 VGND.n46 0.122949
R174 VGND.n47 VGND.n0 0.122949
R175 a_1818_76.n0 a_1818_76.t1 598.523
R176 a_1818_76.t0 a_1818_76.n0 22.7032
R177 a_1818_76.n0 a_1818_76.t2 22.7032
R178 a_1534_446.n6 a_1534_446.t3 815.39
R179 a_1534_446.n5 a_1534_446.t8 412.329
R180 a_1534_446.n3 a_1534_446.n1 354.474
R181 a_1534_446.t2 a_1534_446.n7 320.517
R182 a_1534_446.n2 a_1534_446.t7 294.021
R183 a_1534_446.n2 a_1534_446.t6 277.954
R184 a_1534_446.n0 a_1534_446.t4 258.942
R185 a_1534_446.n6 a_1534_446.n5 198.512
R186 a_1534_446.n0 a_1534_446.t5 191.339
R187 a_1534_446.n5 a_1534_446.n4 171.379
R188 a_1534_446.n3 a_1534_446.n0 152
R189 a_1534_446.n7 a_1534_446.n3 135.772
R190 a_1534_446.n7 a_1534_446.n6 98.3925
R191 a_1534_446.n0 a_1534_446.n2 94.0357
R192 a_1534_446.n1 a_1534_446.t1 25.9464
R193 a_1534_446.n1 a_1534_446.t0 25.9464
R194 D.n0 D.t1 359.777
R195 D.n1 D.n0 152
R196 D.n0 D.t0 139.665
R197 D.n1 D 18.0369
R198 D D.n1 0.582318
R199 a_311_119.n1 a_311_119.t0 868.184
R200 a_311_119.n0 a_311_119.t3 814.707
R201 a_311_119.t1 a_311_119.n1 261.668
R202 a_311_119.n0 a_311_119.t2 231.172
R203 a_311_119.n1 a_311_119.n0 162.363
R204 a_867_119.n0 a_867_119.t1 487.065
R205 a_867_119.t0 a_867_119.n0 45.8187
R206 a_867_119.n0 a_867_119.t2 30.546
R207 VPWR.n32 VPWR.t11 775.191
R208 VPWR.n24 VPWR.n23 649.534
R209 VPWR.n46 VPWR.n45 623.024
R210 VPWR.n16 VPWR.n15 607.417
R211 VPWR.n38 VPWR.n6 606.333
R212 VPWR.n53 VPWR.n1 331.5
R213 VPWR.n14 VPWR.n13 243.151
R214 VPWR.n45 VPWR.t7 138.369
R215 VPWR.n45 VPWR.t10 72.7029
R216 VPWR.n15 VPWR.t0 70.7974
R217 VPWR.n13 VPWR.t4 53.1234
R218 VPWR.n23 VPWR.t3 46.2955
R219 VPWR.n23 VPWR.t8 46.2955
R220 VPWR.n39 VPWR.n38 36.1417
R221 VPWR.n39 VPWR.n4 36.1417
R222 VPWR.n43 VPWR.n4 36.1417
R223 VPWR.n44 VPWR.n43 36.1417
R224 VPWR.n47 VPWR.n44 36.1417
R225 VPWR.n51 VPWR.n2 36.1417
R226 VPWR.n52 VPWR.n51 36.1417
R227 VPWR.n53 VPWR.n52 36.1417
R228 VPWR.n37 VPWR.n7 36.1417
R229 VPWR.n31 VPWR.n30 36.1417
R230 VPWR.n33 VPWR.n31 36.1417
R231 VPWR.n26 VPWR.n25 36.1417
R232 VPWR.n18 VPWR.n17 36.1417
R233 VPWR.n18 VPWR.n11 36.1417
R234 VPWR.n22 VPWR.n11 35.909
R235 VPWR.n30 VPWR.n9 35.4437
R236 VPWR.n6 VPWR.t9 35.1791
R237 VPWR.n6 VPWR.t12 35.1791
R238 VPWR.n13 VPWR.t2 28.2205
R239 VPWR.n1 VPWR.t1 26.3844
R240 VPWR.n1 VPWR.t6 26.3844
R241 VPWR.n15 VPWR.t5 25.505
R242 VPWR.n26 VPWR.n9 19.8562
R243 VPWR.n47 VPWR.n46 19.577
R244 VPWR.n17 VPWR.n16 18.4476
R245 VPWR.n46 VPWR.n2 16.5652
R246 VPWR.n25 VPWR.n24 16.4172
R247 VPWR.n38 VPWR.n37 11.2946
R248 VPWR.n33 VPWR.n32 9.78874
R249 VPWR.n17 VPWR.n12 9.3005
R250 VPWR.n19 VPWR.n18 9.3005
R251 VPWR.n20 VPWR.n11 9.3005
R252 VPWR.n22 VPWR.n21 9.3005
R253 VPWR.n25 VPWR.n10 9.3005
R254 VPWR.n27 VPWR.n26 9.3005
R255 VPWR.n28 VPWR.n9 9.3005
R256 VPWR.n30 VPWR.n29 9.3005
R257 VPWR.n31 VPWR.n8 9.3005
R258 VPWR.n34 VPWR.n33 9.3005
R259 VPWR.n35 VPWR.n7 9.3005
R260 VPWR.n37 VPWR.n36 9.3005
R261 VPWR.n38 VPWR.n5 9.3005
R262 VPWR.n40 VPWR.n39 9.3005
R263 VPWR.n41 VPWR.n4 9.3005
R264 VPWR.n43 VPWR.n42 9.3005
R265 VPWR.n44 VPWR.n3 9.3005
R266 VPWR.n48 VPWR.n47 9.3005
R267 VPWR.n49 VPWR.n2 9.3005
R268 VPWR.n51 VPWR.n50 9.3005
R269 VPWR.n52 VPWR.n0 9.3005
R270 VPWR.n54 VPWR.n53 7.70379
R271 VPWR.n16 VPWR.n14 7.33232
R272 VPWR.n24 VPWR.n22 4.60275
R273 VPWR.n32 VPWR.n7 1.50638
R274 VPWR.n14 VPWR.n12 0.214838
R275 VPWR VPWR.n54 0.163644
R276 VPWR.n54 VPWR.n0 0.144205
R277 VPWR.n19 VPWR.n12 0.122949
R278 VPWR.n20 VPWR.n19 0.122949
R279 VPWR.n21 VPWR.n20 0.122949
R280 VPWR.n21 VPWR.n10 0.122949
R281 VPWR.n27 VPWR.n10 0.122949
R282 VPWR.n28 VPWR.n27 0.122949
R283 VPWR.n29 VPWR.n28 0.122949
R284 VPWR.n29 VPWR.n8 0.122949
R285 VPWR.n34 VPWR.n8 0.122949
R286 VPWR.n35 VPWR.n34 0.122949
R287 VPWR.n36 VPWR.n35 0.122949
R288 VPWR.n36 VPWR.n5 0.122949
R289 VPWR.n40 VPWR.n5 0.122949
R290 VPWR.n41 VPWR.n40 0.122949
R291 VPWR.n42 VPWR.n41 0.122949
R292 VPWR.n42 VPWR.n3 0.122949
R293 VPWR.n48 VPWR.n3 0.122949
R294 VPWR.n49 VPWR.n48 0.122949
R295 VPWR.n50 VPWR.n49 0.122949
R296 VPWR.n50 VPWR.n0 0.122949
R297 CLK_N.n0 CLK_N.t1 259.132
R298 CLK_N.n0 CLK_N.t0 198.882
R299 CLK_N CLK_N.n0 156.667
R300 a_1917_392.t0 a_1917_392.t1 53.1905
R301 Q_N.n1 Q_N 589.572
R302 Q_N.n1 Q_N.n0 585
R303 Q_N.n2 Q_N.n1 585
R304 Q_N Q_N.t1 202.718
R305 Q_N.n1 Q_N.t0 26.3844
R306 Q_N Q_N.n2 12.2519
R307 Q_N Q_N.n0 10.6062
R308 Q_N Q_N.n0 2.92621
R309 Q_N.n2 Q_N 1.2805
R310 a_2412_410.t0 a_2412_410.n1 425.692
R311 a_2412_410.n0 a_2412_410.t3 267.252
R312 a_2412_410.n1 a_2412_410.t1 259.56
R313 a_2412_410.n0 a_2412_410.t2 180.493
R314 a_2412_410.n1 a_2412_410.n0 168.874
R315 Q.n3 Q 589.777
R316 Q.n3 Q.n0 585
R317 Q.n4 Q.n3 585
R318 Q.n2 Q.t1 285
R319 Q.t1 Q.n1 285
R320 Q.n3 Q.t0 26.3844
R321 Q Q.n4 12.8005
R322 Q.n1 Q 12.4184
R323 Q Q.n0 11.0811
R324 Q Q.n2 9.36169
R325 Q.n2 Q 4.77662
R326 Q Q.n0 3.05722
R327 Q.n1 Q 1.7199
R328 Q.n4 Q 1.33781
R329 a_978_357.t0 a_978_357.n3 713.995
R330 a_978_357.n2 a_978_357.n0 554.585
R331 a_978_357.n1 a_978_357.t3 295.894
R332 a_978_357.n0 a_978_357.t4 281.301
R333 a_978_357.n3 a_978_357.t1 247.213
R334 a_978_357.n1 a_978_357.t5 178.34
R335 a_978_357.n0 a_978_357.t2 173.52
R336 a_978_357.n2 a_978_357.n1 166.546
R337 a_978_357.n3 a_978_357.n2 60.2358
R338 a_537_503.t0 a_537_503.t1 126.644
R339 RESET_B.n0 RESET_B.t1 173.788
R340 RESET_B RESET_B.n0 156.019
R341 RESET_B.n0 RESET_B.t0 151.028
C0 D SET_B 2.05e-20
C1 CLK_N VGND 0.017214f
C2 a_1349_114# RESET_B 0.017129f
C3 VPWR CLK_N 0.01506f
C4 VPB D 0.098607f
C5 a_1349_114# a_1483_508# 0.005327f
C6 D VGND 0.011449f
C7 a_1349_114# Q_N 2.94e-19
C8 VPB SET_B 0.150066f
C9 VPWR D 0.005088f
C10 SET_B VGND 0.06745f
C11 a_1297_424# SET_B 0.003506f
C12 VPB VGND 0.021815f
C13 VPWR SET_B 0.161304f
C14 VPB VPWR 0.373583f
C15 SET_B RESET_B 2.2e-19
C16 a_1483_508# SET_B 0.001757f
C17 VPWR VGND 0.120309f
C18 VPB RESET_B 0.044732f
C19 a_1297_424# VPWR 0.007961f
C20 SET_B Q_N 2.47e-19
C21 VGND RESET_B 0.004539f
C22 VPWR RESET_B 0.004679f
C23 VPB Q_N 0.016039f
C24 a_1483_508# VPWR 0.003589f
C25 VGND Q_N 0.04076f
C26 SET_B Q 7.36e-20
C27 VPWR Q_N 0.07198f
C28 VPB Q 0.014088f
C29 VGND Q 0.07861f
C30 RESET_B Q_N 0.001428f
C31 VPWR Q 0.127503f
C32 RESET_B Q 1.49e-19
C33 a_1349_114# SET_B 0.206713f
C34 a_1349_114# VPB 0.094218f
C35 CLK_N SET_B 1.13e-20
C36 a_1349_114# VGND 0.028769f
C37 VPB CLK_N 0.039657f
C38 a_1349_114# a_1297_424# 0.005799f
C39 a_1349_114# VPWR 0.113979f
C40 Q VNB 0.111529f
C41 Q_N VNB 0.014842f
C42 RESET_B VNB 0.115003f
C43 VGND VNB 1.48812f
C44 SET_B VNB 0.221839f
C45 D VNB 0.139776f
C46 CLK_N VNB 0.161399f
C47 VPWR VNB 1.19507f
C48 VPB VNB 3.08462f
C49 a_1349_114# VNB 0.13507f
.ends

* NGSPICE file created from sky130_fd_sc_hs__decap_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__decap_8 VNB VPB VPWR VGND
X0 VPWR.t2 VGND.t3 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1375 pd=1.275 as=0 ps=0 w=1 l=1
X1 VPWR.t1 VGND.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2 VGND.t1 VPWR.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3 VGND.t2 VPWR.t4 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=1
R0 VGND.n6 VGND.t4 271.815
R1 VGND.n2 VGND.t3 268.562
R2 VGND.t2 VGND.n2 225
R3 VGND.n6 VGND.t1 225
R4 VGND.n4 VGND.n3 209.825
R5 VGND.n3 VGND.t2 40.0005
R6 VGND.n3 VGND.t0 40.0005
R7 VGND.n7 VGND.n5 34.6358
R8 VGND.n5 VGND.n4 18.824
R9 VGND.n2 VGND.n1 15.8334
R10 VGND.n7 VGND.n6 14.3724
R11 VGND.n5 VGND.n0 9.3005
R12 VGND.n4 VGND.n1 6.96404
R13 VGND.n8 VGND.n7 4.62059
R14 VGND.n1 VGND.n0 0.512494
R15 VGND.n8 VGND.n0 0.184273
R16 VGND VGND.n8 0.123049
R17 VPWR.t2 VPWR.n1 255.988
R18 VPWR.n7 VPWR.t1 252.012
R19 VPWR.n4 VPWR.n3 192.861
R20 VPWR.n2 VPWR.t4 101.233
R21 VPWR.n2 VPWR.t3 100.415
R22 VPWR.n4 VPWR.n2 75.2651
R23 VPWR.n6 VPWR.n5 32.0005
R24 VPWR.n3 VPWR.t0 27.5805
R25 VPWR.n3 VPWR.t2 26.5955
R26 VPWR.n7 VPWR.n6 22.2123
R27 VPWR.n5 VPWR.n4 11.8714
R28 VPWR.n6 VPWR.n0 9.3005
R29 VPWR.n8 VPWR.n7 9.3005
R30 VPWR.n5 VPWR.n1 3.15412
R31 VPWR.n1 VPWR.n0 0.495413
R32 VPWR.n8 VPWR.n0 0.122949
R33 VPWR VPWR.n8 0.0617245
R34 VPB.t0 VPB.t1 651.211
R35 VPB VPB.t0 464.786
R36 VNB.t1 VNB.t0 2956.43
R37 VNB VNB.t1 2251.97
C0 VGND VPWR 0.878569f
C1 VPB VPWR 0.180477f
C2 VPB VGND 0.213851f
C3 VPWR VNB 1.11129f
C4 VGND VNB 1.0624f
C5 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__decap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__decap_4 VNB VPB VPWR VGND
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
R0 VGND.n0 VGND.t2 271.815
R1 VGND.n1 VGND.t0 256.68
R2 VGND.n0 VGND.t1 225
R3 VGND.n1 VGND.n0 18.2828
R4 VGND VGND.n1 0.374088
R5 VPWR.n0 VPWR.t2 278.632
R6 VPWR.n1 VPWR.t1 258.839
R7 VPWR.n0 VPWR.t0 219.089
R8 VPWR.n1 VPWR.n0 23.567
R9 VPWR VPWR.n1 0.322181
R10 VPB VPB.t0 464.786
R11 VNB VNB.t0 2251.97
C0 VGND VPB 0.106687f
C1 VPWR VPB 0.09177f
C2 VGND VPWR 0.425061f
C3 VPWR VNB 0.685621f
C4 VGND VNB 0.609974f
C5 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__conb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__conb_1 VNB VPB VPWR VGND LO HI
X0 VPWR.t0 HI.t0 sky130_fd_pr__res_generic_po w=0.51 l=0.045
X1 LO.t0 VGND.t0 sky130_fd_pr__res_generic_po w=0.51 l=0.045
R0 VPWR VPWR.t0 214.004
R1 HI.n0 HI.t0 155.44
R2 HI.n1 HI 15.0715
R3 HI HI.n0 6.10389
R4 HI.n0 HI 2.75926
R5 HI HI.n1 0.206952
R6 HI.n1 HI 0.121255
R7 LO.n0 LO.t0 188.905
R8 LO.n1 LO 7.0405
R9 LO LO.n1 3.98541
R10 LO.n1 LO.n0 3.80527
R11 LO.n0 LO 1.13544
R12 VGND VGND.t0 181.356
C0 VPWR HI 0.068326f
C1 VPB HI 0.007052f
C2 VPB VPWR 0.189101f
C3 HI VGND 0.224519f
C4 HI LO 0.051631f
C5 VPWR VGND 0.028636f
C6 VPWR LO 0.258375f
C7 VPB VGND 0.005087f
C8 VPB LO 0.159645f
C9 LO VGND 0.052542f
C10 VGND VNB 0.459009f
C11 LO VNB 0.203197f
C12 HI VNB 0.30832f
C13 VPWR VNB 0.321691f
C14 VPB VNB 0.406224f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkinv_16 VNB VPB VPWR VGND A Y
X0 Y.t39 A.t0 VPWR.t23 VPB.t23 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t22 A.t1 Y.t38 VPB.t22 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t21 A.t2 Y.t37 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VGND.t15 A.t3 Y.t15 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y.t14 A.t4 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0882 ps=0.84 w=0.42 l=0.15
X5 VGND.t13 A.t5 Y.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND.t12 A.t6 Y.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 Y.t36 A.t7 VPWR.t20 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Y.t11 A.t8 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VPWR.t19 A.t9 Y.t35 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t34 A.t10 VPWR.t18 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t33 A.t11 VPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VGND.t10 A.t12 Y.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR.t16 A.t13 Y.t32 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR.t15 A.t14 Y.t31 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 Y.t30 A.t15 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.196 ps=1.47 w=1.12 l=0.15
X16 Y.t29 A.t16 VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 Y.t28 A.t17 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VPWR.t11 A.t18 Y.t27 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VPWR.t10 A.t19 Y.t26 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2016 ps=1.48 w=1.12 l=0.15
X20 Y.t9 A.t20 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 Y.t25 A.t21 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X22 VPWR.t8 A.t22 Y.t24 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 VPWR.t7 A.t23 Y.t23 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X24 Y.t22 A.t24 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 Y.t8 A.t25 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X26 VPWR.t5 A.t26 Y.t21 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 Y.t20 A.t27 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 Y.t7 A.t28 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X29 VPWR.t3 A.t29 Y.t19 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X30 Y.t6 A.t30 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X31 Y.t18 A.t31 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X32 VGND.t5 A.t32 Y.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 Y.t4 A.t33 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 VGND.t3 A.t34 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 Y.t2 A.t35 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 VPWR.t1 A.t36 Y.t17 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X37 VGND.t1 A.t37 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 Y.t16 A.t38 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X39 VGND.t0 A.t39 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.71835 pd=5.57 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A.n16 A.t23 262.288
R1 A.n82 A.t28 229.486
R2 A.n83 A.t3 228.148
R3 A.n81 A.t8 228.148
R4 A.n79 A.t37 228.148
R5 A.n76 A.t30 228.148
R6 A.n74 A.t34 228.148
R7 A.n66 A.t25 228.148
R8 A.n67 A.t12 228.148
R9 A.n64 A.t4 228.148
R10 A.n62 A.t32 228.148
R11 A.n59 A.t20 228.148
R12 A.n57 A.t6 228.148
R13 A.n50 A.t35 228.148
R14 A.n52 A.t5 228.148
R15 A.n48 A.t33 228.148
R16 A.n47 A.t39 228.148
R17 A.n15 A.t27 226.809
R18 A.n20 A.t36 226.809
R19 A.n11 A.t7 226.809
R20 A.n30 A.t9 226.809
R21 A.n31 A.t11 226.809
R22 A.n41 A.t13 226.809
R23 A.n5 A.t17 226.809
R24 A.n46 A.t19 226.809
R25 A.n49 A.t15 226.809
R26 A.n51 A.t29 226.809
R27 A.n3 A.t31 226.809
R28 A.n58 A.t2 226.809
R29 A.n60 A.t38 226.809
R30 A.n63 A.t1 226.809
R31 A.n65 A.t10 226.809
R32 A.n68 A.t14 226.809
R33 A.n1 A.t16 226.809
R34 A.n73 A.t18 226.809
R35 A.n75 A.t21 226.809
R36 A.n78 A.t22 226.809
R37 A.n80 A.t24 226.809
R38 A.n84 A.t26 226.809
R39 A.n82 A.t0 204.048
R40 A.n86 A.n85 168.9
R41 A.n77 A.n0 168.671
R42 A.n72 A.n71 168.671
R43 A.n70 A.n69 168.671
R44 A.n61 A.n2 168.671
R45 A.n56 A.n55 168.671
R46 A.n54 A.n53 168.671
R47 A.n45 A.n44 155.584
R48 A.n17 A.n16 153.024
R49 A.n19 A.n18 152
R50 A.n23 A.n22 152
R51 A.n21 A.n12 152
R52 A.n29 A.n28 152
R53 A.n33 A.n32 152
R54 A.n8 A.n7 152
R55 A.n40 A.n39 152
R56 A.n43 A.n42 152
R57 A.n48 A.n47 57.5727
R58 A.n67 A.n66 57.5727
R59 A.n83 A.n82 56.2338
R60 A.n75 A.n74 54.8949
R61 A.n80 A.n79 50.8783
R62 A.n22 A.n21 45.5227
R63 A.n40 A.n7 45.5227
R64 A.n64 A.n63 45.5227
R65 A.n51 A.n50 44.1838
R66 A.n20 A.n19 39.4977
R67 A.n32 A.n31 38.1588
R68 A.n42 A.n41 38.1588
R69 A.n29 A.n11 36.8199
R70 A.n46 A.n45 36.8199
R71 A.n62 A.n61 36.8199
R72 A.n69 A.n68 36.8199
R73 A.n77 A.n76 34.1422
R74 A.n73 A.n72 32.8033
R75 A.n59 A.n58 32.1338
R76 A.n85 A.n81 30.1255
R77 A.n60 A.n59 28.1172
R78 A.n53 A.n52 27.4477
R79 A.n72 A.n1 27.4477
R80 A.n53 A.n49 26.1088
R81 A.n56 A.n3 26.1088
R82 A.n58 A.n57 25.4394
R83 A.n16 A.n15 24.7699
R84 A.n30 A.n29 23.4311
R85 A.n45 A.n5 23.4311
R86 A.n69 A.n65 23.4311
R87 A.n78 A.n77 23.4311
R88 A.n85 A.n84 23.4311
R89 A.n32 A.n30 22.0922
R90 A.n42 A.n5 22.0922
R91 A.n19 A.n15 20.7533
R92 A.n50 A.n3 16.0672
R93 A.n57 A.n56 15.3977
R94 A.n65 A.n64 14.7283
R95 A.n52 A.n51 13.3894
R96 A.n63 A.n62 12.0505
R97 A.n61 A.n60 11.3811
R98 A.n17 A.n13 9.49615
R99 A.n79 A.n78 9.37272
R100 A.n44 A.n4 9.3005
R101 A.n36 A.n6 9.3005
R102 A.n38 A.n37 9.3005
R103 A.n35 A.n34 9.3005
R104 A.n10 A.n9 9.3005
R105 A.n27 A.n26 9.3005
R106 A.n25 A.n24 9.3005
R107 A.n14 A.n13 9.3005
R108 A.n21 A.n11 8.70328
R109 A.n18 A.n17 7.6805
R110 A.n31 A.n7 7.36439
R111 A.n41 A.n40 7.36439
R112 A.n23 A.n14 7.1685
R113 A.n47 A.n46 6.69494
R114 A.n81 A.n80 6.69494
R115 A.n24 A.n12 6.6565
R116 A.n28 A.n27 6.1445
R117 A.n22 A.n20 6.0255
R118 A.n33 A.n10 5.6325
R119 A.n74 A.n73 5.35606
R120 A.n34 A.n8 5.1205
R121 A.n44 A.n43 5.1205
R122 A.n39 A.n38 4.6085
R123 A.n39 A.n6 4.6085
R124 A.n38 A.n8 4.0965
R125 A.n43 A.n6 4.0965
R126 A.n49 A.n48 4.01717
R127 A.n84 A.n83 4.01717
R128 A.n34 A.n33 3.5845
R129 A.n28 A.n10 3.0725
R130 A.n76 A.n75 2.67828
R131 A.n27 A.n12 2.5605
R132 A.n24 A.n23 2.0485
R133 A.n18 A.n14 1.5365
R134 A.n68 A.n67 1.33939
R135 A.n66 A.n1 1.33939
R136 A.n54 A.n4 0.609196
R137 A.n70 A.n2 0.538543
R138 A.n71 A.n0 0.527674
R139 A.n55 A.n54 0.516804
R140 A.n71 A.n70 0.505935
R141 A.n86 A.n0 0.48963
R142 A.n55 A.n2 0.457022
R143 A.n25 A.n13 0.196152
R144 A.n26 A.n25 0.196152
R145 A.n26 A.n9 0.196152
R146 A.n35 A.n9 0.196152
R147 A.n37 A.n35 0.196152
R148 A.n37 A.n36 0.196152
R149 A.n36 A.n4 0.196152
R150 A A.n86 0.0793043
R151 VPWR.n18 VPWR.t7 256.671
R152 VPWR.n60 VPWR.t23 250.081
R153 VPWR.n4 VPWR.n3 243.916
R154 VPWR.n52 VPWR.n6 243.916
R155 VPWR.n46 VPWR.n45 243.916
R156 VPWR.n43 VPWR.n9 243.916
R157 VPWR.n58 VPWR.n2 232.787
R158 VPWR.n37 VPWR.n36 232.787
R159 VPWR.n26 VPWR.n15 232.787
R160 VPWR.n34 VPWR.n12 228.188
R161 VPWR.n28 VPWR.n27 223.696
R162 VPWR.n17 VPWR.n16 223.696
R163 VPWR.n20 VPWR.n19 223.696
R164 VPWR.n42 VPWR.n10 36.1417
R165 VPWR.n47 VPWR.n44 36.1417
R166 VPWR.n51 VPWR.n7 36.1417
R167 VPWR.n54 VPWR.n53 36.1417
R168 VPWR.n38 VPWR.n35 36.1417
R169 VPWR.n33 VPWR.n13 36.1417
R170 VPWR.n36 VPWR.t2 35.1791
R171 VPWR.n12 VPWR.t14 35.1791
R172 VPWR.n29 VPWR.n26 34.2593
R173 VPWR.n58 VPWR.n57 31.2476
R174 VPWR.n57 VPWR.n4 30.1181
R175 VPWR.n25 VPWR.n17 29.7417
R176 VPWR.n2 VPWR.t6 26.3844
R177 VPWR.n2 VPWR.t5 26.3844
R178 VPWR.n3 VPWR.t9 26.3844
R179 VPWR.n3 VPWR.t8 26.3844
R180 VPWR.n6 VPWR.t13 26.3844
R181 VPWR.n6 VPWR.t11 26.3844
R182 VPWR.n45 VPWR.t18 26.3844
R183 VPWR.n45 VPWR.t15 26.3844
R184 VPWR.n9 VPWR.t0 26.3844
R185 VPWR.n9 VPWR.t22 26.3844
R186 VPWR.n36 VPWR.t21 26.3844
R187 VPWR.n12 VPWR.t3 26.3844
R188 VPWR.n27 VPWR.t12 26.3844
R189 VPWR.n27 VPWR.t10 26.3844
R190 VPWR.n15 VPWR.t17 26.3844
R191 VPWR.n15 VPWR.t16 26.3844
R192 VPWR.n16 VPWR.t20 26.3844
R193 VPWR.n16 VPWR.t19 26.3844
R194 VPWR.n19 VPWR.t4 26.3844
R195 VPWR.n19 VPWR.t1 26.3844
R196 VPWR.n53 VPWR.n52 25.6005
R197 VPWR.n21 VPWR.n20 25.224
R198 VPWR.n59 VPWR.n58 22.2123
R199 VPWR.n46 VPWR.n7 21.0829
R200 VPWR.n60 VPWR.n59 20.7064
R201 VPWR.n43 VPWR.n42 19.577
R202 VPWR.n26 VPWR.n25 19.2005
R203 VPWR.n21 VPWR.n17 17.6946
R204 VPWR.n44 VPWR.n43 16.5652
R205 VPWR.n47 VPWR.n46 15.0593
R206 VPWR.n34 VPWR.n33 12.424
R207 VPWR.n38 VPWR.n37 11.6711
R208 VPWR.n52 VPWR.n51 10.5417
R209 VPWR.n22 VPWR.n21 9.3005
R210 VPWR.n23 VPWR.n17 9.3005
R211 VPWR.n25 VPWR.n24 9.3005
R212 VPWR.n26 VPWR.n14 9.3005
R213 VPWR.n30 VPWR.n29 9.3005
R214 VPWR.n31 VPWR.n13 9.3005
R215 VPWR.n33 VPWR.n32 9.3005
R216 VPWR.n35 VPWR.n11 9.3005
R217 VPWR.n39 VPWR.n38 9.3005
R218 VPWR.n40 VPWR.n10 9.3005
R219 VPWR.n42 VPWR.n41 9.3005
R220 VPWR.n44 VPWR.n8 9.3005
R221 VPWR.n48 VPWR.n47 9.3005
R222 VPWR.n49 VPWR.n7 9.3005
R223 VPWR.n51 VPWR.n50 9.3005
R224 VPWR.n53 VPWR.n5 9.3005
R225 VPWR.n55 VPWR.n54 9.3005
R226 VPWR.n57 VPWR.n56 9.3005
R227 VPWR.n58 VPWR.n1 9.3005
R228 VPWR.n59 VPWR.n0 9.3005
R229 VPWR.n61 VPWR.n60 9.3005
R230 VPWR.n29 VPWR.n28 8.65932
R231 VPWR.n20 VPWR.n18 6.50549
R232 VPWR.n54 VPWR.n4 6.02403
R233 VPWR.n37 VPWR.n10 5.64756
R234 VPWR.n28 VPWR.n13 2.63579
R235 VPWR.n35 VPWR.n34 2.25932
R236 VPWR.n22 VPWR.n18 0.686474
R237 VPWR.n23 VPWR.n22 0.122949
R238 VPWR.n24 VPWR.n23 0.122949
R239 VPWR.n24 VPWR.n14 0.122949
R240 VPWR.n30 VPWR.n14 0.122949
R241 VPWR.n31 VPWR.n30 0.122949
R242 VPWR.n32 VPWR.n31 0.122949
R243 VPWR.n32 VPWR.n11 0.122949
R244 VPWR.n39 VPWR.n11 0.122949
R245 VPWR.n40 VPWR.n39 0.122949
R246 VPWR.n41 VPWR.n40 0.122949
R247 VPWR.n41 VPWR.n8 0.122949
R248 VPWR.n48 VPWR.n8 0.122949
R249 VPWR.n49 VPWR.n48 0.122949
R250 VPWR.n50 VPWR.n49 0.122949
R251 VPWR.n50 VPWR.n5 0.122949
R252 VPWR.n55 VPWR.n5 0.122949
R253 VPWR.n56 VPWR.n55 0.122949
R254 VPWR.n56 VPWR.n1 0.122949
R255 VPWR.n1 VPWR.n0 0.122949
R256 VPWR.n61 VPWR.n0 0.122949
R257 VPWR VPWR.n61 0.0617245
R258 Y.n37 Y.n36 283.704
R259 Y.n17 Y.n15 279.776
R260 Y.n21 Y.n19 267.248
R261 Y.n13 Y.n11 261.435
R262 Y.n33 Y.n31 260.041
R263 Y.n9 Y.n7 258.527
R264 Y.n25 Y.n23 253.325
R265 Y.n29 Y.n27 244.208
R266 Y.n2 Y.n0 220.27
R267 Y.n6 Y.n5 219.78
R268 Y.n4 Y.n3 219.78
R269 Y.n2 Y.n1 219.78
R270 Y.n37 Y.n35 207.712
R271 Y.n9 Y.n8 204.954
R272 Y.n25 Y.n24 204.399
R273 Y.n13 Y.n12 202.802
R274 Y.n17 Y.n16 202.475
R275 Y.n33 Y.n32 202.457
R276 Y.n29 Y.n28 202.457
R277 Y.n21 Y.n20 202.457
R278 Y.n36 Y.t15 40.0005
R279 Y.n36 Y.t7 40.0005
R280 Y.n31 Y.t1 40.0005
R281 Y.n31 Y.t11 40.0005
R282 Y.n27 Y.t3 40.0005
R283 Y.n27 Y.t6 40.0005
R284 Y.n23 Y.t10 40.0005
R285 Y.n23 Y.t8 40.0005
R286 Y.n19 Y.t5 40.0005
R287 Y.n19 Y.t14 40.0005
R288 Y.n15 Y.t12 40.0005
R289 Y.n15 Y.t9 40.0005
R290 Y.n11 Y.t13 40.0005
R291 Y.n11 Y.t2 40.0005
R292 Y.n7 Y.t0 40.0005
R293 Y.n7 Y.t4 40.0005
R294 Y.n8 Y.t26 31.6612
R295 Y.n8 Y.t30 31.6612
R296 Y.n35 Y.t21 26.3844
R297 Y.n35 Y.t39 26.3844
R298 Y.n32 Y.t24 26.3844
R299 Y.n32 Y.t22 26.3844
R300 Y.n28 Y.t27 26.3844
R301 Y.n28 Y.t25 26.3844
R302 Y.n24 Y.t31 26.3844
R303 Y.n24 Y.t29 26.3844
R304 Y.n20 Y.t38 26.3844
R305 Y.n20 Y.t34 26.3844
R306 Y.n16 Y.t37 26.3844
R307 Y.n16 Y.t16 26.3844
R308 Y.n12 Y.t19 26.3844
R309 Y.n12 Y.t18 26.3844
R310 Y.n5 Y.t32 26.3844
R311 Y.n5 Y.t28 26.3844
R312 Y.n3 Y.t35 26.3844
R313 Y.n3 Y.t33 26.3844
R314 Y.n1 Y.t17 26.3844
R315 Y.n1 Y.t36 26.3844
R316 Y.n0 Y.t23 26.3844
R317 Y.n0 Y.t20 26.3844
R318 Y.n38 Y.n37 10.497
R319 Y.n10 Y.n9 10.2162
R320 Y.n26 Y.n25 10.1611
R321 Y.n14 Y.n13 10.0053
R322 Y.n34 Y.n33 9.97218
R323 Y.n30 Y.n29 9.97218
R324 Y.n22 Y.n21 9.97218
R325 Y.n18 Y.n17 9.94427
R326 Y.n14 Y.n10 0.533109
R327 Y.n18 Y.n14 0.516804
R328 Y.n10 Y.n6 0.505935
R329 Y.n30 Y.n26 0.505935
R330 Y.n38 Y.n34 0.495065
R331 Y.n4 Y.n2 0.48963
R332 Y.n6 Y.n4 0.48963
R333 Y.n22 Y.n18 0.48963
R334 Y.n34 Y.n30 0.48963
R335 Y.n26 Y.n22 0.473326
R336 Y Y.n38 0.0793043
R337 VPB.t14 VPB.t10 260.485
R338 VPB VPB.t23 257.93
R339 VPB.t3 VPB.t14 255.376
R340 VPB.t21 VPB.t2 255.376
R341 VPB.t4 VPB.t7 229.839
R342 VPB.t1 VPB.t4 229.839
R343 VPB.t20 VPB.t1 229.839
R344 VPB.t19 VPB.t20 229.839
R345 VPB.t17 VPB.t19 229.839
R346 VPB.t16 VPB.t17 229.839
R347 VPB.t12 VPB.t16 229.839
R348 VPB.t10 VPB.t12 229.839
R349 VPB.t2 VPB.t3 229.839
R350 VPB.t0 VPB.t21 229.839
R351 VPB.t22 VPB.t0 229.839
R352 VPB.t18 VPB.t22 229.839
R353 VPB.t15 VPB.t18 229.839
R354 VPB.t13 VPB.t15 229.839
R355 VPB.t11 VPB.t13 229.839
R356 VPB.t9 VPB.t11 229.839
R357 VPB.t8 VPB.t9 229.839
R358 VPB.t6 VPB.t8 229.839
R359 VPB.t5 VPB.t6 229.839
R360 VPB.t23 VPB.t5 229.839
R361 VGND.n37 VGND.t7 248.661
R362 VGND.n28 VGND.n27 216.232
R363 VGND.n31 VGND.n30 212.887
R364 VGND.n14 VGND.n13 212.397
R365 VGND.n35 VGND.n2 212.397
R366 VGND.n11 VGND.n10 209.4
R367 VGND.n19 VGND.n7 209.4
R368 VGND.n22 VGND.n21 208.661
R369 VGND.n9 VGND.t0 184.867
R370 VGND.n7 VGND.t9 60.0005
R371 VGND.n7 VGND.t5 60.0005
R372 VGND.n21 VGND.t14 60.0005
R373 VGND.n21 VGND.t10 60.0005
R374 VGND.n27 VGND.t8 60.0005
R375 VGND.n30 VGND.t6 60.0005
R376 VGND.n10 VGND.t4 40.0005
R377 VGND.n10 VGND.t13 40.0005
R378 VGND.n13 VGND.t2 40.0005
R379 VGND.n13 VGND.t12 40.0005
R380 VGND.n27 VGND.t3 40.0005
R381 VGND.n30 VGND.t1 40.0005
R382 VGND.n2 VGND.t11 40.0005
R383 VGND.n2 VGND.t15 40.0005
R384 VGND.n15 VGND.n12 36.1417
R385 VGND.n26 VGND.n4 36.1417
R386 VGND.n31 VGND.n29 35.7652
R387 VGND.n22 VGND.n20 35.0123
R388 VGND.n19 VGND.n6 32.7534
R389 VGND.n35 VGND.n1 31.624
R390 VGND.n37 VGND.n36 20.7064
R391 VGND.n36 VGND.n35 19.2005
R392 VGND.n20 VGND.n19 15.4358
R393 VGND.n29 VGND.n28 15.4358
R394 VGND.n31 VGND.n1 15.4358
R395 VGND.n11 VGND.n9 13.5087
R396 VGND.n14 VGND.n6 13.177
R397 VGND.n22 VGND.n4 12.424
R398 VGND.n38 VGND.n37 9.3005
R399 VGND.n12 VGND.n8 9.3005
R400 VGND.n16 VGND.n15 9.3005
R401 VGND.n17 VGND.n6 9.3005
R402 VGND.n19 VGND.n18 9.3005
R403 VGND.n20 VGND.n5 9.3005
R404 VGND.n23 VGND.n22 9.3005
R405 VGND.n24 VGND.n4 9.3005
R406 VGND.n26 VGND.n25 9.3005
R407 VGND.n29 VGND.n3 9.3005
R408 VGND.n32 VGND.n31 9.3005
R409 VGND.n33 VGND.n1 9.3005
R410 VGND.n35 VGND.n34 9.3005
R411 VGND.n36 VGND.n0 9.3005
R412 VGND.n12 VGND.n11 5.64756
R413 VGND.n28 VGND.n26 1.88285
R414 VGND.n15 VGND.n14 1.50638
R415 VGND.n9 VGND.n8 0.634035
R416 VGND.n16 VGND.n8 0.122949
R417 VGND.n17 VGND.n16 0.122949
R418 VGND.n18 VGND.n17 0.122949
R419 VGND.n18 VGND.n5 0.122949
R420 VGND.n23 VGND.n5 0.122949
R421 VGND.n24 VGND.n23 0.122949
R422 VGND.n25 VGND.n24 0.122949
R423 VGND.n25 VGND.n3 0.122949
R424 VGND.n32 VGND.n3 0.122949
R425 VGND.n33 VGND.n32 0.122949
R426 VGND.n34 VGND.n33 0.122949
R427 VGND.n34 VGND.n0 0.122949
R428 VGND.n38 VGND.n0 0.122949
R429 VGND VGND.n38 0.0617245
R430 VNB.t5 VNB.t9 1316.54
R431 VNB.t10 VNB.t14 1316.54
R432 VNB.t3 VNB.t8 1154.86
R433 VNB.t1 VNB.t6 1154.86
R434 VNB VNB.t7 1143.31
R435 VNB.t4 VNB.t0 993.177
R436 VNB.t13 VNB.t4 993.177
R437 VNB.t2 VNB.t13 993.177
R438 VNB.t12 VNB.t2 993.177
R439 VNB.t9 VNB.t12 993.177
R440 VNB.t14 VNB.t5 993.177
R441 VNB.t8 VNB.t10 993.177
R442 VNB.t6 VNB.t3 993.177
R443 VNB.t11 VNB.t1 993.177
R444 VNB.t15 VNB.t11 993.177
R445 VNB.t7 VNB.t15 993.177
C0 VPB A 0.871924f
C1 VPB VPWR 0.319568f
C2 VPB Y 0.067344f
C3 A VPWR 0.76022f
C4 A Y 2.38127f
C5 VPB VGND 0.007236f
C6 A VGND 0.949899f
C7 VPWR Y 3.11059f
C8 VPWR VGND 0.054447f
C9 Y VGND 0.803793f
C10 VGND VNB 1.44736f
C11 Y VNB 0.144682f
C12 VPWR VNB 1.154254f
C13 A VNB 2.616634f
C14 VPB VNB 2.65608f
C15 Y.t23 VNB 0.033776f
C16 Y.t20 VNB 0.033776f
C17 Y.n0 VNB 0.076585f
C18 Y.t17 VNB 0.033776f
C19 Y.t36 VNB 0.033776f
C20 Y.n1 VNB 0.076307f
C21 Y.n2 VNB 0.279056f
C22 Y.t35 VNB 0.033776f
C23 Y.t33 VNB 0.033776f
C24 Y.n3 VNB 0.076307f
C25 Y.n4 VNB 0.153771f
C26 Y.t32 VNB 0.033776f
C27 Y.t28 VNB 0.033776f
C28 Y.n5 VNB 0.076307f
C29 Y.n6 VNB 0.155158f
C30 Y.t0 VNB 0.011821f
C31 Y.t4 VNB 0.011821f
C32 Y.n7 VNB 0.049807f
C33 Y.t26 VNB 0.040531f
C34 Y.t30 VNB 0.040531f
C35 Y.n8 VNB 0.086814f
C36 Y.n9 VNB 0.216139f
C37 Y.n10 VNB 0.096368f
C38 Y.t13 VNB 0.011821f
C39 Y.t2 VNB 0.011821f
C40 Y.n11 VNB 0.047022f
C41 Y.t19 VNB 0.033776f
C42 Y.t18 VNB 0.033776f
C43 Y.n12 VNB 0.073408f
C44 Y.n13 VNB 0.241886f
C45 Y.n14 VNB 0.097486f
C46 Y.t12 VNB 0.011821f
C47 Y.t9 VNB 0.011821f
C48 Y.n15 VNB 0.050396f
C49 Y.t37 VNB 0.033776f
C50 Y.t16 VNB 0.033776f
C51 Y.n16 VNB 0.073426f
C52 Y.n17 VNB 0.227656f
C53 Y.n18 VNB 0.093498f
C54 Y.t5 VNB 0.011821f
C55 Y.t14 VNB 0.011821f
C56 Y.n19 VNB 0.056599f
C57 Y.t38 VNB 0.033776f
C58 Y.t34 VNB 0.033776f
C59 Y.n20 VNB 0.073426f
C60 Y.n21 VNB 0.257119f
C61 Y.n22 VNB 0.09012f
C62 Y.t10 VNB 0.011821f
C63 Y.t8 VNB 0.011821f
C64 Y.n23 VNB 0.051687f
C65 Y.t31 VNB 0.033776f
C66 Y.t29 VNB 0.033776f
C67 Y.n24 VNB 0.073331f
C68 Y.n25 VNB 0.23544f
C69 Y.n26 VNB 0.091332f
C70 Y.t3 VNB 0.011821f
C71 Y.t6 VNB 0.011821f
C72 Y.n27 VNB 0.051478f
C73 Y.t27 VNB 0.033776f
C74 Y.t25 VNB 0.033776f
C75 Y.n28 VNB 0.073426f
C76 Y.n29 VNB 0.287229f
C77 Y.n30 VNB 0.092894f
C78 Y.t1 VNB 0.011821f
C79 Y.t11 VNB 0.011821f
C80 Y.n31 VNB 0.049693f
C81 Y.t24 VNB 0.033776f
C82 Y.t22 VNB 0.033776f
C83 Y.n32 VNB 0.073426f
C84 Y.n33 VNB 0.249046f
C85 Y.n34 VNB 0.091969f
C86 Y.t21 VNB 0.033776f
C87 Y.t39 VNB 0.033776f
C88 Y.n35 VNB 0.073173f
C89 Y.t15 VNB 0.011821f
C90 Y.t7 VNB 0.011821f
C91 Y.n36 VNB 0.047697f
C92 Y.n37 VNB 0.156949f
C93 Y.n38 VNB 0.05659f
C94 VPWR.n0 VNB 0.043497f
C95 VPWR.t23 VNB 0.064192f
C96 VPWR.n1 VNB 0.043497f
C97 VPWR.t6 VNB 0.015535f
C98 VPWR.t5 VNB 0.015535f
C99 VPWR.n2 VNB 0.040279f
C100 VPWR.t9 VNB 0.015535f
C101 VPWR.t8 VNB 0.015535f
C102 VPWR.n3 VNB 0.03861f
C103 VPWR.n4 VNB 0.044806f
C104 VPWR.n5 VNB 0.043497f
C105 VPWR.t13 VNB 0.015535f
C106 VPWR.t11 VNB 0.015535f
C107 VPWR.n6 VNB 0.03861f
C108 VPWR.n7 VNB 0.011947f
C109 VPWR.n8 VNB 0.043497f
C110 VPWR.t0 VNB 0.015535f
C111 VPWR.t22 VNB 0.015535f
C112 VPWR.n9 VNB 0.03861f
C113 VPWR.n10 VNB 0.008724f
C114 VPWR.n11 VNB 0.043497f
C115 VPWR.t14 VNB 0.020713f
C116 VPWR.t3 VNB 0.015535f
C117 VPWR.n12 VNB 0.045652f
C118 VPWR.n13 VNB 0.008096f
C119 VPWR.n14 VNB 0.043497f
C120 VPWR.t17 VNB 0.015535f
C121 VPWR.t16 VNB 0.015535f
C122 VPWR.n15 VNB 0.040279f
C123 VPWR.t20 VNB 0.015535f
C124 VPWR.t19 VNB 0.015535f
C125 VPWR.n16 VNB 0.040675f
C126 VPWR.n17 VNB 0.097639f
C127 VPWR.t7 VNB 0.067399f
C128 VPWR.n18 VNB 0.126563f
C129 VPWR.t4 VNB 0.015535f
C130 VPWR.t1 VNB 0.015535f
C131 VPWR.n19 VNB 0.040675f
C132 VPWR.n20 VNB 0.099254f
C133 VPWR.n21 VNB 0.00896f
C134 VPWR.n22 VNB 0.146524f
C135 VPWR.n23 VNB 0.043497f
C136 VPWR.n24 VNB 0.043497f
C137 VPWR.n25 VNB 0.010218f
C138 VPWR.n26 VNB 0.075695f
C139 VPWR.t12 VNB 0.015535f
C140 VPWR.t10 VNB 0.015535f
C141 VPWR.n27 VNB 0.040675f
C142 VPWR.n28 VNB 0.090094f
C143 VPWR.n29 VNB 0.00896f
C144 VPWR.n30 VNB 0.043497f
C145 VPWR.n31 VNB 0.043497f
C146 VPWR.n32 VNB 0.043497f
C147 VPWR.n33 VNB 0.010139f
C148 VPWR.n34 VNB 0.077715f
C149 VPWR.n35 VNB 0.008017f
C150 VPWR.t2 VNB 0.020713f
C151 VPWR.t21 VNB 0.015535f
C152 VPWR.n36 VNB 0.045457f
C153 VPWR.n37 VNB 0.068149f
C154 VPWR.n38 VNB 0.009982f
C155 VPWR.n39 VNB 0.043497f
C156 VPWR.n40 VNB 0.043497f
C157 VPWR.n41 VNB 0.043497f
C158 VPWR.n42 VNB 0.011632f
C159 VPWR.n43 VNB 0.044806f
C160 VPWR.n44 VNB 0.011004f
C161 VPWR.t18 VNB 0.015535f
C162 VPWR.t15 VNB 0.015535f
C163 VPWR.n45 VNB 0.03861f
C164 VPWR.n46 VNB 0.044806f
C165 VPWR.n47 VNB 0.010689f
C166 VPWR.n48 VNB 0.043497f
C167 VPWR.n49 VNB 0.043497f
C168 VPWR.n50 VNB 0.043497f
C169 VPWR.n51 VNB 0.009746f
C170 VPWR.n52 VNB 0.044806f
C171 VPWR.n53 VNB 0.01289f
C172 VPWR.n54 VNB 0.008803f
C173 VPWR.n55 VNB 0.043497f
C174 VPWR.n56 VNB 0.043497f
C175 VPWR.n57 VNB 0.012811f
C176 VPWR.n58 VNB 0.075695f
C177 VPWR.n59 VNB 0.00896f
C178 VPWR.n60 VNB 0.090078f
C179 VPWR.n61 VNB 0.032623f
C180 A.n0 VNB 0.058448f
C181 A.t8 VNB 0.010386f
C182 A.t24 VNB 0.01873f
C183 A.t37 VNB 0.010386f
C184 A.t22 VNB 0.01873f
C185 A.t30 VNB 0.010386f
C186 A.t21 VNB 0.01873f
C187 A.t34 VNB 0.010386f
C188 A.t18 VNB 0.01873f
C189 A.t16 VNB 0.01873f
C190 A.n1 VNB 0.015293f
C191 A.n2 VNB 0.057716f
C192 A.t10 VNB 0.01873f
C193 A.t4 VNB 0.010386f
C194 A.t1 VNB 0.01873f
C195 A.t32 VNB 0.010386f
C196 A.t38 VNB 0.01873f
C197 A.t20 VNB 0.010386f
C198 A.t2 VNB 0.01873f
C199 A.t6 VNB 0.010386f
C200 A.t31 VNB 0.01873f
C201 A.n3 VNB 0.018158f
C202 A.n4 VNB 0.027091f
C203 A.t15 VNB 0.01873f
C204 A.t33 VNB 0.010386f
C205 A.t39 VNB 0.010386f
C206 A.t19 VNB 0.01873f
C207 A.t17 VNB 0.01873f
C208 A.n5 VNB 0.018874f
C209 A.n6 VNB 0.013529f
C210 A.t13 VNB 0.01873f
C211 A.n7 VNB 0.011317f
C212 A.n8 VNB 0.014325f
C213 A.n9 VNB 0.013179f
C214 A.n10 VNB 0.013529f
C215 A.t9 VNB 0.01873f
C216 A.t7 VNB 0.01873f
C217 A.n11 VNB 0.018874f
C218 A.n12 VNB 0.014325f
C219 A.n13 VNB 0.027701f
C220 A.n14 VNB 0.013529f
C221 A.t36 VNB 0.01873f
C222 A.t27 VNB 0.01873f
C223 A.n15 VNB 0.018874f
C224 A.t23 VNB 0.02169f
C225 A.n16 VNB 0.031914f
C226 A.n17 VNB 0.02846f
C227 A.n18 VNB 0.014325f
C228 A.n19 VNB 0.012893f
C229 A.n20 VNB 0.018874f
C230 A.n21 VNB 0.011603f
C231 A.n22 VNB 0.011031f
C232 A.n23 VNB 0.014325f
C233 A.n24 VNB 0.013529f
C234 A.n25 VNB 0.013179f
C235 A.n26 VNB 0.013179f
C236 A.n27 VNB 0.013529f
C237 A.n28 VNB 0.014325f
C238 A.n29 VNB 0.012893f
C239 A.n30 VNB 0.018874f
C240 A.t11 VNB 0.01873f
C241 A.n31 VNB 0.018874f
C242 A.n32 VNB 0.012893f
C243 A.n33 VNB 0.014325f
C244 A.n34 VNB 0.013529f
C245 A.n35 VNB 0.013179f
C246 A.n36 VNB 0.013179f
C247 A.n37 VNB 0.013179f
C248 A.n38 VNB 0.013529f
C249 A.n39 VNB 0.014325f
C250 A.n40 VNB 0.011317f
C251 A.n41 VNB 0.018874f
C252 A.n42 VNB 0.012893f
C253 A.n43 VNB 0.014325f
C254 A.n44 VNB 0.031801f
C255 A.n45 VNB 0.013324f
C256 A.n46 VNB 0.018444f
C257 A.n47 VNB 0.022228f
C258 A.n48 VNB 0.021655f
C259 A.n49 VNB 0.015579f
C260 A.t5 VNB 0.010386f
C261 A.t29 VNB 0.01873f
C262 A.t35 VNB 0.010386f
C263 A.n50 VNB 0.021369f
C264 A.n51 VNB 0.021453f
C265 A.n52 VNB 0.017214f
C266 A.n53 VNB 0.013505f
C267 A.n54 VNB 0.062109f
C268 A.n55 VNB 0.056984f
C269 A.n56 VNB 0.010926f
C270 A.n57 VNB 0.017214f
C271 A.n58 VNB 0.021453f
C272 A.n59 VNB 0.021369f
C273 A.n60 VNB 0.017585f
C274 A.n61 VNB 0.012359f
C275 A.n62 VNB 0.018933f
C276 A.n63 VNB 0.021453f
C277 A.n64 VNB 0.021369f
C278 A.n65 VNB 0.017298f
C279 A.t14 VNB 0.01873f
C280 A.t12 VNB 0.010386f
C281 A.t25 VNB 0.010386f
C282 A.n66 VNB 0.021082f
C283 A.n67 VNB 0.021082f
C284 A.n68 VNB 0.017298f
C285 A.n69 VNB 0.014938f
C286 A.n70 VNB 0.059363f
C287 A.n71 VNB 0.058997f
C288 A.n72 VNB 0.014938f
C289 A.n73 VNB 0.017298f
C290 A.n74 VNB 0.021369f
C291 A.n75 VNB 0.021453f
C292 A.n76 VNB 0.016355f
C293 A.n77 VNB 0.014365f
C294 A.n78 VNB 0.016152f
C295 A.n79 VNB 0.021369f
C296 A.n80 VNB 0.021453f
C297 A.n81 VNB 0.016355f
C298 A.t26 VNB 0.01873f
C299 A.t3 VNB 0.010386f
C300 A.t0 VNB 0.017847f
C301 A.t28 VNB 0.010463f
C302 A.n82 VNB 0.035458f
C303 A.n83 VNB 0.021369f
C304 A.n84 VNB 0.015006f
C305 A.n85 VNB 0.013458f
C306 A.n86 VNB 0.042597f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkinv_8 VNB VPB VPWR VGND A Y
X0 VPWR.t11 A.t0 Y.t9 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t10 A.t1 Y.t18 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t7 A.t2 Y.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.4221 ps=2.43 w=0.42 l=0.15
X3 VGND.t6 A.t3 Y.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y.t17 A.t4 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5 Y.t16 A.t5 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6 Y.t12 A.t6 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0882 ps=0.84 w=0.42 l=0.15
X7 VPWR.t7 A.t7 Y.t15 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t6 A.t8 Y.t14 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t11 A.t9 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.4221 pd=2.43 as=0.1281 ps=1.45 w=0.42 l=0.15
X10 Y.t13 A.t10 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X11 VGND.t3 A.t11 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 VGND.t2 A.t12 Y.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR.t4 A.t13 Y.t8 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X14 Y.t19 A.t14 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0882 ps=0.84 w=0.42 l=0.15
X15 Y.t7 A.t15 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X16 VPWR.t2 A.t16 Y.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X17 Y.t5 A.t17 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3584 ps=2.88 w=1.12 l=0.15
X18 Y.t4 A.t18 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X19 Y.t10 A.t19 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0882 ps=0.84 w=0.42 l=0.15
R0 A.n22 A.t9 239.978
R1 A.n3 A.t11 239.978
R2 A.n18 A.t2 237.787
R3 A.n17 A.t19 237.787
R4 A.n42 A.t12 237.787
R5 A.n14 A.t6 237.787
R6 A.n1 A.t3 237.787
R7 A.n6 A.t14 237.787
R8 A.n3 A.t16 226.809
R9 A.n5 A.t18 226.809
R10 A.n8 A.t0 226.809
R11 A.n13 A.t4 226.809
R12 A.n43 A.t7 226.809
R13 A.n16 A.t10 226.809
R14 A.n37 A.t13 226.809
R15 A.n32 A.t15 226.809
R16 A.n30 A.t1 226.809
R17 A.n20 A.t5 226.809
R18 A.n24 A.t8 226.809
R19 A.n22 A.t17 226.809
R20 A.n4 A.n2 162.121
R21 A.n23 A 161.674
R22 A.n7 A.n2 152
R23 A.n10 A.n9 152
R24 A.n12 A.n11 152
R25 A.n15 A.n0 152
R26 A.n45 A.n44 152
R27 A.n41 A.n40 152
R28 A.n39 A.n38 152
R29 A.n36 A.n35 152
R30 A.n34 A.n33 152
R31 A.n31 A.n19 152
R32 A.n29 A.n28 152
R33 A.n27 A.n26 152
R34 A.n25 A.n21 152
R35 A.n9 A.n7 49.6611
R36 A.n44 A.n15 49.6611
R37 A.n26 A.n25 49.6611
R38 A.n29 A.n20 48.2005
R39 A.n38 A.n37 42.3581
R40 A.n32 A.n31 40.8975
R41 A.n5 A.n4 39.4369
R42 A.n23 A.n22 37.9763
R43 A.n31 A.n30 32.1338
R44 A.n13 A.n12 29.2126
R45 A.n24 A.n23 27.752
R46 A.n33 A.n18 27.0217
R47 A.n4 A.n3 26.2914
R48 A.n42 A.n41 24.1005
R49 A.n43 A.n42 22.6399
R50 A.n36 A.n18 22.6399
R51 A.n25 A.n24 21.9096
R52 A.n12 A.n1 21.1793
R53 A.n17 A.n16 19.7187
R54 A.n41 A.n16 18.9884
R55 A.n30 A.n29 17.5278
R56 A.n8 A.n1 15.3369
R57 A.n9 A.n8 13.146
R58 A.n14 A.n13 12.4157
R59 A.n38 A.n17 10.955
R60 A.n10 A.n2 10.1214
R61 A.n11 A.n10 10.1214
R62 A.n11 A.n0 10.1214
R63 A.n40 A.n39 10.1214
R64 A.n34 A.n19 10.1214
R65 A.n27 A.n21 10.1214
R66 A.n45 A 9.97259
R67 A.n33 A.n32 8.76414
R68 A.n35 A 8.18655
R69 A.n15 A.n14 8.03383
R70 A.n28 A 7.88887
R71 A.n37 A.n36 7.30353
R72 A.n28 A 6.4005
R73 A.n35 A 6.10283
R74 A A.n0 5.80515
R75 A.n6 A.n5 5.11262
R76 A.n7 A.n6 5.11262
R77 A A.n45 4.31678
R78 A.n39 A 4.0191
R79 A A.n27 3.72143
R80 A.n44 A.n43 2.92171
R81 A A.n19 2.23306
R82 A A.n34 1.93538
R83 A.n26 A.n20 1.46111
R84 A A.n21 0.447012
R85 A.n40 A 0.149337
R86 Y.n27 Y.n2 203.812
R87 Y.n26 Y.n3 203.812
R88 Y.n25 Y.n4 203.812
R89 Y.n15 Y.n8 203.394
R90 Y.n14 Y.n9 203.394
R91 Y.n13 Y.n10 203.394
R92 Y.n12 Y.n11 203.394
R93 Y.n1 Y.n0 203.394
R94 Y.n16 Y.n7 203.394
R95 Y.n18 Y.n17 185
R96 Y.n19 Y.n6 185
R97 Y.n21 Y.n20 185
R98 Y.n22 Y.n5 185
R99 Y.n24 Y.n23 185
R100 Y.n23 Y.n22 120.001
R101 Y.n22 Y.n21 120.001
R102 Y.n21 Y.n6 120.001
R103 Y.n17 Y.n6 120.001
R104 Y.n18 Y.n16 95.9221
R105 Y Y.n1 62.1018
R106 Y.n2 Y.t3 60.0005
R107 Y.n17 Y.t11 54.2862
R108 Y.n25 Y.n24 53.3809
R109 Y.n27 Y.n26 50.4476
R110 Y.n26 Y.n25 50.4476
R111 Y.n16 Y.n15 46.6829
R112 Y.n15 Y.n14 46.6829
R113 Y.n14 Y.n13 46.6829
R114 Y.n13 Y.n12 46.6829
R115 Y.n12 Y.n1 46.6829
R116 Y.n23 Y.t2 40.0005
R117 Y.n2 Y.t19 40.0005
R118 Y.n3 Y.t1 40.0005
R119 Y.n3 Y.t12 40.0005
R120 Y.n4 Y.t0 40.0005
R121 Y.n4 Y.t10 40.0005
R122 Y.n7 Y.t14 26.3844
R123 Y.n7 Y.t5 26.3844
R124 Y.n8 Y.t18 26.3844
R125 Y.n8 Y.t16 26.3844
R126 Y.n9 Y.t8 26.3844
R127 Y.n9 Y.t7 26.3844
R128 Y.n10 Y.t15 26.3844
R129 Y.n10 Y.t13 26.3844
R130 Y.n11 Y.t9 26.3844
R131 Y.n11 Y.t17 26.3844
R132 Y.n0 Y.t6 26.3844
R133 Y.n0 Y.t4 26.3844
R134 Y Y.n27 25.977
R135 Y.n24 Y.n5 7.46717
R136 Y.n20 Y.n5 7.46717
R137 Y.n20 Y.n19 7.46717
R138 Y.n19 Y.n18 7.46717
R139 VPWR.n9 VPWR.t2 356.822
R140 VPWR.n25 VPWR.t1 349.623
R141 VPWR.n23 VPWR.n2 323.406
R142 VPWR.n4 VPWR.n3 323.406
R143 VPWR.n17 VPWR.n6 323.406
R144 VPWR.n8 VPWR.n7 323.406
R145 VPWR.n11 VPWR.n10 323.406
R146 VPWR.n2 VPWR.t8 35.1791
R147 VPWR.n3 VPWR.t3 35.1791
R148 VPWR.n6 VPWR.t5 35.1791
R149 VPWR.n7 VPWR.t9 35.1791
R150 VPWR.n10 VPWR.t0 35.1791
R151 VPWR.n24 VPWR.n23 30.1181
R152 VPWR.n22 VPWR.n4 29.3652
R153 VPWR.n18 VPWR.n17 28.6123
R154 VPWR.n16 VPWR.n8 27.8593
R155 VPWR.n12 VPWR.n11 27.1064
R156 VPWR.n2 VPWR.t6 26.3844
R157 VPWR.n3 VPWR.t10 26.3844
R158 VPWR.n6 VPWR.t4 26.3844
R159 VPWR.n7 VPWR.t7 26.3844
R160 VPWR.n10 VPWR.t11 26.3844
R161 VPWR.n12 VPWR.n8 25.6005
R162 VPWR.n25 VPWR.n24 24.8476
R163 VPWR.n17 VPWR.n16 24.8476
R164 VPWR.n18 VPWR.n4 24.0946
R165 VPWR.n23 VPWR.n22 23.3417
R166 VPWR.n13 VPWR.n12 9.3005
R167 VPWR.n14 VPWR.n8 9.3005
R168 VPWR.n16 VPWR.n15 9.3005
R169 VPWR.n17 VPWR.n5 9.3005
R170 VPWR.n19 VPWR.n18 9.3005
R171 VPWR.n20 VPWR.n4 9.3005
R172 VPWR.n22 VPWR.n21 9.3005
R173 VPWR.n23 VPWR.n1 9.3005
R174 VPWR.n24 VPWR.n0 9.3005
R175 VPWR.n26 VPWR.n25 9.3005
R176 VPWR.n11 VPWR.n9 6.85153
R177 VPWR.n13 VPWR.n9 0.568865
R178 VPWR.n14 VPWR.n13 0.122949
R179 VPWR.n15 VPWR.n14 0.122949
R180 VPWR.n15 VPWR.n5 0.122949
R181 VPWR.n19 VPWR.n5 0.122949
R182 VPWR.n20 VPWR.n19 0.122949
R183 VPWR.n21 VPWR.n20 0.122949
R184 VPWR.n21 VPWR.n1 0.122949
R185 VPWR.n1 VPWR.n0 0.122949
R186 VPWR.n26 VPWR.n0 0.122949
R187 VPWR VPWR.n26 0.0617245
R188 VPB VPB.t1 270.7
R189 VPB.t11 VPB.t0 255.376
R190 VPB.t7 VPB.t9 255.376
R191 VPB.t4 VPB.t5 255.376
R192 VPB.t10 VPB.t3 255.376
R193 VPB.t6 VPB.t8 255.376
R194 VPB.t0 VPB.t2 229.839
R195 VPB.t9 VPB.t11 229.839
R196 VPB.t5 VPB.t7 229.839
R197 VPB.t3 VPB.t4 229.839
R198 VPB.t8 VPB.t10 229.839
R199 VPB.t1 VPB.t6 229.839
R200 VGND.n6 VGND.t3 255.365
R201 VGND.n23 VGND.t4 254.375
R202 VGND.n8 VGND.n7 208.661
R203 VGND.n11 VGND.n10 208.661
R204 VGND.n15 VGND.n4 208.661
R205 VGND.n7 VGND.t1 60.0005
R206 VGND.n7 VGND.t6 60.0005
R207 VGND.n10 VGND.t5 60.0005
R208 VGND.n10 VGND.t2 60.0005
R209 VGND.n4 VGND.t0 60.0005
R210 VGND.n4 VGND.t7 60.0005
R211 VGND.n17 VGND.n16 36.1417
R212 VGND.n17 VGND.n1 36.1417
R213 VGND.n21 VGND.n1 36.1417
R214 VGND.n22 VGND.n21 36.1417
R215 VGND.n15 VGND.n3 35.7652
R216 VGND.n11 VGND.n9 32.7534
R217 VGND.n23 VGND.n22 20.7064
R218 VGND.n9 VGND.n8 17.6946
R219 VGND.n11 VGND.n3 14.6829
R220 VGND.n16 VGND.n15 11.6711
R221 VGND.n24 VGND.n23 9.3005
R222 VGND.n9 VGND.n5 9.3005
R223 VGND.n12 VGND.n11 9.3005
R224 VGND.n13 VGND.n3 9.3005
R225 VGND.n15 VGND.n14 9.3005
R226 VGND.n16 VGND.n2 9.3005
R227 VGND.n18 VGND.n17 9.3005
R228 VGND.n19 VGND.n1 9.3005
R229 VGND.n21 VGND.n20 9.3005
R230 VGND.n22 VGND.n0 9.3005
R231 VGND.n8 VGND.n6 6.96039
R232 VGND.n6 VGND.n5 0.594857
R233 VGND.n12 VGND.n5 0.122949
R234 VGND.n13 VGND.n12 0.122949
R235 VGND.n14 VGND.n13 0.122949
R236 VGND.n14 VGND.n2 0.122949
R237 VGND.n18 VGND.n2 0.122949
R238 VGND.n19 VGND.n18 0.122949
R239 VGND.n20 VGND.n19 0.122949
R240 VGND.n20 VGND.n0 0.122949
R241 VGND.n24 VGND.n0 0.122949
R242 VGND VGND.n24 0.0617245
R243 VNB.t4 VNB.t7 4988.98
R244 VNB.t6 VNB.t1 1316.54
R245 VNB.t2 VNB.t5 1316.54
R246 VNB.t7 VNB.t0 1316.54
R247 VNB VNB.t4 1189.5
R248 VNB.t1 VNB.t3 1154.86
R249 VNB.t5 VNB.t6 993.177
R250 VNB.t0 VNB.t2 993.177
C0 VPB Y 0.033179f
C1 A VPWR 0.214922f
C2 A Y 1.38961f
C3 VPB VGND 0.007817f
C4 A VGND 0.140983f
C5 VPWR Y 1.14616f
C6 VPWR VGND 0.108113f
C7 Y VGND 0.642053f
C8 VPB A 0.451292f
C9 VPB VPWR 0.178075f
C10 VGND VNB 0.809477f
C11 Y VNB 0.230081f
C12 VPWR VNB 0.63369f
C13 A VNB 1.35264f
C14 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxbp_1 VNB VPB VPWR VGND D CLK Q Q_N
X0 a_701_463.t2 a_543_447.t4 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2541 pd=1.445 as=0.232575 ps=1.715 w=0.84 l=0.15
X1 a_420_503.t2 D.t0 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.368725 ps=2.64 w=0.42 l=0.15
X2 a_543_447.t1 a_27_74.t2 a_420_503.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.075675 pd=0.83 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR.t2 a_1191_120# a_1158_482.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4 VGND.t5 CLK.t0 a_27_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2017 pd=1.35 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 a_1005_120.t1 a_205_368.t2 a_701_463.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.12965 pd=1.09 as=0.11825 ps=1.13 w=0.55 l=0.15
X6 a_205_368.t0 a_27_74.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.3252 pd=2.59 as=0.2017 ps=1.35 w=0.74 l=0.15
X7 Q.t1 a_1191_120# VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1934 ps=1.475 w=1.12 l=0.15
X8 VPWR.t3 a_1191_120# a_1644_94.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2394 ps=2.25 w=0.84 l=0.15
X9 a_543_447.t2 a_205_368.t3 a_420_503.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.107525 pd=1.11 as=0.146375 ps=1.335 w=0.42 l=0.15
X10 a_1158_482.t0 a_205_368.t4 a_1005_120.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.14085 ps=1.225 w=0.42 l=0.15
X11 a_205_368.t1 a_27_74.t4 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VPWR.t1 a_701_463.t4 a_650_508.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.232575 pd=1.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_701_463.t3 a_543_447.t5 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.11825 pd=1.13 as=0.145125 ps=1.19 w=0.55 l=0.15
X14 a_650_508.t1 a_27_74.t5 a_543_447.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.107525 ps=1.11 w=0.42 l=0.15
X15 VGND.t0 a_701_463.t5 a_713_102.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.145125 pd=1.19 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 Q.t0 a_1191_120# VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1469 ps=1.16 w=0.74 l=0.15
X17 VPWR.t0 CLK.t1 a_27_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
X18 a_713_102.t1 a_205_368.t5 a_543_447.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.075675 ps=0.83 w=0.42 l=0.15
X19 Q_N.t0 a_1644_94.t1 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.12945 ps=1.1 w=0.74 l=0.15
X20 a_420_503.t3 D.t1 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.146375 pd=1.335 as=0.2282 ps=2.1 w=0.42 l=0.15
X21 a_1005_120.t0 a_27_74.t6 a_701_463.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.14085 pd=1.225 as=0.2541 ps=1.445 w=0.84 l=0.15
X22 VGND.t3 a_1191_120# a_1143_146# VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_543_447.n2 a_543_447.n1 588.23
R1 a_543_447.n0 a_543_447.t5 329.368
R2 a_543_447.n3 a_543_447.n2 287.25
R3 a_543_447.n2 a_543_447.n0 265.303
R4 a_543_447.n1 a_543_447.t3 243.191
R5 a_543_447.n0 a_543_447.t4 197.888
R6 a_543_447.n1 a_543_447.t2 68.0124
R7 a_543_447.n3 a_543_447.t1 41.0879
R8 a_543_447.n4 a_543_447.t0 25.6415
R9 a_543_447.n5 a_543_447.n4 21.6005
R10 a_543_447.n4 a_543_447.n3 21.493
R11 VPWR.n2 VPWR.t5 773.793
R12 VPWR.n12 VPWR.t2 682.896
R13 VPWR.n20 VPWR.n19 613.144
R14 VPWR.n9 VPWR.t3 410.954
R15 VPWR.n8 VPWR.t4 369.661
R16 VPWR.n32 VPWR.n1 326.231
R17 VPWR.n19 VPWR.t7 162.994
R18 VPWR.n19 VPWR.t1 124.299
R19 VPWR.n25 VPWR.n4 36.1417
R20 VPWR.n26 VPWR.n25 36.1417
R21 VPWR.n27 VPWR.n26 36.1417
R22 VPWR.n13 VPWR.n6 36.1417
R23 VPWR.n17 VPWR.n6 36.1417
R24 VPWR.n18 VPWR.n17 36.1417
R25 VPWR.n12 VPWR.n11 35.0123
R26 VPWR.n21 VPWR.n18 33.6831
R27 VPWR.n31 VPWR.n30 29.7488
R28 VPWR.n32 VPWR.n31 29.3652
R29 VPWR.n1 VPWR.t6 26.3844
R30 VPWR.n1 VPWR.t0 26.3844
R31 VPWR.n27 VPWR.n2 24.6913
R32 VPWR.n11 VPWR.n8 21.0829
R33 VPWR.n20 VPWR.n4 15.6356
R34 VPWR.n13 VPWR.n12 12.424
R35 VPWR.n11 VPWR.n10 9.3005
R36 VPWR.n12 VPWR.n7 9.3005
R37 VPWR.n14 VPWR.n13 9.3005
R38 VPWR.n15 VPWR.n6 9.3005
R39 VPWR.n17 VPWR.n16 9.3005
R40 VPWR.n18 VPWR.n5 9.3005
R41 VPWR.n22 VPWR.n21 9.3005
R42 VPWR.n23 VPWR.n4 9.3005
R43 VPWR.n25 VPWR.n24 9.3005
R44 VPWR.n26 VPWR.n3 9.3005
R45 VPWR.n28 VPWR.n27 9.3005
R46 VPWR.n30 VPWR.n29 9.3005
R47 VPWR.n31 VPWR.n0 9.3005
R48 VPWR.n9 VPWR.n8 7.45966
R49 VPWR.n33 VPWR.n32 7.25439
R50 VPWR.n21 VPWR.n20 3.78826
R51 VPWR.n30 VPWR.n2 0.966538
R52 VPWR.n10 VPWR.n9 0.215804
R53 VPWR VPWR.n33 0.157727
R54 VPWR.n33 VPWR.n0 0.150046
R55 VPWR.n10 VPWR.n7 0.122949
R56 VPWR.n14 VPWR.n7 0.122949
R57 VPWR.n15 VPWR.n14 0.122949
R58 VPWR.n16 VPWR.n15 0.122949
R59 VPWR.n16 VPWR.n5 0.122949
R60 VPWR.n22 VPWR.n5 0.122949
R61 VPWR.n23 VPWR.n22 0.122949
R62 VPWR.n24 VPWR.n23 0.122949
R63 VPWR.n24 VPWR.n3 0.122949
R64 VPWR.n28 VPWR.n3 0.122949
R65 VPWR.n29 VPWR.n28 0.122949
R66 VPWR.n29 VPWR.n0 0.122949
R67 a_701_463.n3 a_701_463.n2 665.566
R68 a_701_463.n1 a_701_463.t4 485.031
R69 a_701_463.n2 a_701_463.n0 192.606
R70 a_701_463.n2 a_701_463.n1 171.651
R71 a_701_463.n1 a_701_463.t5 123.757
R72 a_701_463.t1 a_701_463.n3 89.1195
R73 a_701_463.n0 a_701_463.t3 61.0919
R74 a_701_463.n3 a_701_463.t2 52.7684
R75 a_701_463.n0 a_701_463.t0 30.5465
R76 VPB.t6 VPB.t5 766.13
R77 VPB.t8 VPB.t7 549.059
R78 VPB.t5 VPB.t4 505.646
R79 VPB.t0 VPB.t11 423.925
R80 VPB.t11 VPB.t10 385.618
R81 VPB.t7 VPB.t1 314.113
R82 VPB.t10 VPB.t2 273.253
R83 VPB.t1 VPB.t9 273.253
R84 VPB VPB.t3 255.376
R85 VPB.t3 VPB.t8 229.839
R86 VPB.t9 VPB.t0 214.517
R87 VPB.t2 VPB.t6 199.195
R88 D.n0 D.t0 357.654
R89 D D.t1 316.622
R90 D.n0 D 10.3116
R91 D D.n0 2.84494
R92 VGND.n1 VGND.t2 366.918
R93 VGND.n8 VGND.t4 269.262
R94 VGND.n10 VGND.t3 258.94
R95 VGND.n18 VGND.n17 240.066
R96 VGND.n32 VGND.n31 198.305
R97 VGND.n7 VGND.t6 160.272
R98 VGND.n17 VGND.t0 72.8576
R99 VGND.n17 VGND.t7 40.3641
R100 VGND.n31 VGND.t1 39.7302
R101 VGND.n31 VGND.t5 39.7302
R102 VGND.n11 VGND.n9 36.1417
R103 VGND.n15 VGND.n5 36.1417
R104 VGND.n16 VGND.n15 36.1417
R105 VGND.n19 VGND.n16 36.1417
R106 VGND.n24 VGND.n23 36.1417
R107 VGND.n25 VGND.n24 36.1417
R108 VGND.n30 VGND.n29 36.1417
R109 VGND.n25 VGND.n1 32.7534
R110 VGND.n23 VGND.n3 31.1981
R111 VGND.n19 VGND.n18 23.0907
R112 VGND.n32 VGND.n30 14.6829
R113 VGND.n9 VGND.n8 13.5534
R114 VGND.n29 VGND.n1 13.177
R115 VGND.n30 VGND.n0 9.3005
R116 VGND.n29 VGND.n28 9.3005
R117 VGND.n27 VGND.n1 9.3005
R118 VGND.n26 VGND.n25 9.3005
R119 VGND.n24 VGND.n2 9.3005
R120 VGND.n23 VGND.n22 9.3005
R121 VGND.n21 VGND.n3 9.3005
R122 VGND.n20 VGND.n19 9.3005
R123 VGND.n16 VGND.n4 9.3005
R124 VGND.n15 VGND.n14 9.3005
R125 VGND.n13 VGND.n5 9.3005
R126 VGND.n12 VGND.n11 9.3005
R127 VGND.n9 VGND.n6 9.3005
R128 VGND.n8 VGND.n7 7.52071
R129 VGND.n33 VGND.n32 7.46433
R130 VGND.n10 VGND.n5 6.02403
R131 VGND.n11 VGND.n10 5.27109
R132 VGND.n18 VGND.n3 1.68131
R133 VGND.n7 VGND.n6 0.206693
R134 VGND VGND.n33 0.160491
R135 VGND.n33 VGND.n0 0.147317
R136 VGND.n12 VGND.n6 0.122949
R137 VGND.n13 VGND.n12 0.122949
R138 VGND.n14 VGND.n13 0.122949
R139 VGND.n14 VGND.n4 0.122949
R140 VGND.n20 VGND.n4 0.122949
R141 VGND.n21 VGND.n20 0.122949
R142 VGND.n22 VGND.n21 0.122949
R143 VGND.n22 VGND.n2 0.122949
R144 VGND.n26 VGND.n2 0.122949
R145 VGND.n27 VGND.n26 0.122949
R146 VGND.n28 VGND.n27 0.122949
R147 VGND.n28 VGND.n0 0.122949
R148 a_420_503.n1 a_420_503.n0 926.83
R149 a_420_503.n0 a_420_503.t3 265.012
R150 a_420_503.n0 a_420_503.t1 89.1196
R151 a_420_503.t0 a_420_503.n1 40.0005
R152 a_420_503.n1 a_420_503.t2 40.0005
R153 VNB.t5 VNB.t6 3603.15
R154 VNB.t6 VNB.t9 3464.57
R155 VNB.t3 VNB.t4 3349.08
R156 VNB.t8 VNB.t5 2494.49
R157 VNB.t7 VNB.t3 1478.22
R158 VNB.t0 VNB.t10 1362.73
R159 VNB.t10 VNB.t8 1177.95
R160 VNB VNB.t7 1143.31
R161 VNB.t2 VNB.t1 1097.11
R162 VNB.t4 VNB.t2 993.177
R163 VNB.t1 VNB.t0 831.496
R164 a_27_74.n1 a_27_74.t6 565.548
R165 a_27_74.n2 a_27_74.n1 398.166
R166 a_27_74.n0 a_27_74.t2 317.647
R167 a_27_74.t0 a_27_74.n5 289.589
R168 a_27_74.n4 a_27_74.t4 281.017
R169 a_27_74.n2 a_27_74.n0 238.519
R170 a_27_74.n3 a_27_74.t1 227.845
R171 a_27_74.n3 a_27_74.n2 221.365
R172 a_27_74.n0 a_27_74.t5 211.607
R173 a_27_74.n4 a_27_74.t3 173.638
R174 a_27_74.n5 a_27_74.n4 152
R175 a_27_74.n5 a_27_74.n3 17.3719
R176 a_1158_482.t0 a_1158_482.t1 112.572
R177 a_1644_94.t0 a_1644_94.n1 602.271
R178 a_1644_94.n1 a_1644_94.n0 264.298
R179 a_1644_94.n1 a_1644_94.t1 204.048
R180 Q_N.n1 Q_N.n0 1214.44
R181 Q_N Q_N.t0 205.88
R182 Q_N Q_N.n1 12.0794
R183 Q_N Q_N.n0 7.05556
R184 Q_N.n0 Q_N 6.21275
R185 Q_N.n1 Q_N 1.26247
R186 CLK.n0 CLK.t1 280.555
R187 CLK.n0 CLK.t0 173.177
R188 CLK CLK.n0 158.227
R189 a_205_368.n0 a_205_368.t5 1135.91
R190 a_205_368.n2 a_205_368.t4 509.288
R191 a_205_368.n0 a_205_368.t3 458.192
R192 a_205_368.n2 a_205_368.t2 421.082
R193 a_205_368.n1 a_205_368.t0 342.512
R194 a_205_368.n3 a_205_368.n2 260.286
R195 a_205_368.t1 a_205_368.n3 217.857
R196 a_205_368.n1 a_205_368.n0 152
R197 a_205_368.n3 a_205_368.n1 19.9957
R198 a_1005_120.n4 a_1005_120.n3 666.388
R199 a_1005_120.n2 a_1005_120.n0 272.464
R200 a_1005_120.n3 a_1005_120.t1 263.3
R201 a_1005_120.n3 a_1005_120.n2 249.506
R202 a_1005_120.n2 a_1005_120.n1 182.758
R203 a_1005_120.n4 a_1005_120.t2 110.227
R204 a_1005_120.n6 a_1005_120.n5 50.5066
R205 a_1005_120.n5 a_1005_120.t0 30.5882
R206 a_1005_120.n5 a_1005_120.n4 6.87376
R207 Q.t1 Q 875.811
R208 Q.n0 Q.t1 726.702
R209 Q.n0 Q.t0 221.031
R210 Q Q.n0 3.95112
R211 a_650_508.t0 a_650_508.t1 126.644
R212 a_713_102.t0 a_713_102.t1 60.0005
C0 a_1191_120# Q 0.152712f
C1 a_1143_146# VPWR 6.06e-19
C2 VGND Q_N 0.104726f
C3 a_1191_120# Q_N 0.002408f
C4 VPB VPWR 0.28133f
C5 VPB CLK 0.036196f
C6 a_1143_146# VGND 0.005069f
C7 a_1191_120# a_1143_146# 2.28e-19
C8 VPB D 0.101066f
C9 VPWR CLK 0.021816f
C10 VPWR D 0.014471f
C11 VPB VGND 0.020709f
C12 a_1191_120# VPB 0.250077f
C13 VPB Q 0.015185f
C14 VPWR VGND 0.153212f
C15 a_1191_120# VPWR 0.25605f
C16 VPB Q_N 0.01462f
C17 VPWR Q 0.134561f
C18 CLK VGND 0.013627f
C19 D VGND 0.008405f
C20 VPWR Q_N 0.135113f
C21 a_1191_120# VGND 0.190805f
C22 VGND Q 0.086306f
C23 Q_N VNB 0.112924f
C24 Q VNB 0.013942f
C25 VGND VNB 1.11695f
C26 D VNB 0.133991f
C27 CLK VNB 0.161665f
C28 VPWR VNB 0.871044f
C29 VPB VNB 2.22754f
C30 a_1191_120# VNB 0.431206f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfstp_4 VNB VPB VPWR SET_B VGND CLK D Q
X0 a_1321_392.t1 a_225_74.t2 a_1220_347.t1 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.21665 pd=1.645 as=0.197175 ps=1.58 w=1 l=0.15
X1 a_612_74.t1 a_398_74.t2 a_27_74.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X2 a_1321_392.t3 a_398_74.t3 a_1225_74.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.105725 pd=1 as=0.1264 ps=1.035 w=0.64 l=0.15
X3 a_1225_74.t1 a_612_74.t4 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1264 pd=1.035 as=0.11745 ps=1.05 w=0.64 l=0.15
X4 VGND.t6 D.t0 a_27_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X5 Q.t6 a_1940_74.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1946 ps=1.49 w=1.12 l=0.15
X6 a_398_74.t0 a_225_74.t3 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_1321_392.t0 SET_B.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.39 as=0.063 ps=0.72 w=0.42 l=0.15
X8 VGND.t8 a_767_402.t3 a_732_74.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.147 pd=1.54 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 a_1514_88.t0 a_1484_62.t2 a_1436_88.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X10 a_1220_347.t0 a_612_74.t5 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.197175 pd=1.58 as=0.1955 ps=1.565 w=1 l=0.15
X11 VPWR.t3 a_1484_62.t3 a_1480_508.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR.t13 CLK.t0 a_225_74.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X13 a_1480_508.t1 a_398_74.t4 a_1321_392.t4 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.21665 ps=1.645 w=0.42 l=0.15
X14 VGND.t11 SET_B.t1 a_1035_118.t0 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.11745 pd=1.05 as=0.0504 ps=0.66 w=0.42 l=0.15
X15 VGND.t10 CLK.t1 a_225_74.t0 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X16 a_1484_62.t0 a_1321_392.t5 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.21735 ps=1.455 w=0.42 l=0.15
X17 Q.t3 a_1940_74.t4 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 VGND.t4 a_1940_74.t5 Q.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.12025 ps=1.065 w=0.74 l=0.15
X19 VPWR.t4 a_767_402.t4 a_716_463.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.16485 pd=1.205 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_398_74.t1 a_225_74.t4 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 Q.t1 a_1940_74.t6 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.2627 ps=1.45 w=0.74 l=0.15
X22 a_612_74.t2 a_225_74.t5 a_27_74.t3 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0945 pd=0.87 as=0.18665 ps=1.8 w=0.42 l=0.15
X23 VGND.t12 SET_B.t2 a_1514_88.t1 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.21735 pd=1.455 as=0.0504 ps=0.66 w=0.42 l=0.15
X24 a_716_463.t1 a_225_74.t6 a_612_74.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0735 ps=0.77 w=0.42 l=0.15
X25 a_732_74.t1 a_398_74.t5 a_612_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0945 ps=0.87 w=0.42 l=0.15
X26 a_1436_88.t1 a_225_74.t7 a_1321_392.t2 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.105725 ps=1 w=0.42 l=0.15
X27 VGND.t2 a_1940_74.t7 Q.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=1.45 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 VPWR.t8 D.t1 a_27_74.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1239 ps=1.43 w=0.42 l=0.15
X29 a_767_402.t1 a_612_74.t6 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.16485 ps=1.205 w=0.42 l=0.15
X30 a_1484_62.t1 a_1321_392.t6 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.39 as=0.1176 ps=1.4 w=0.42 l=0.15
X31 a_1035_118.t1 a_612_74.t7 a_767_402.t2 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1491 ps=1.55 w=0.42 l=0.15
X32 VPWR.t11 a_1321_392.t7 a_1940_74.t0 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1946 pd=1.49 as=0.126 ps=1.14 w=0.84 l=0.15
X33 VGND.t1 a_1321_392.t8 a_1940_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X34 VPWR.t1 a_1940_74.t8 Q.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X35 VPWR.t14 SET_B.t3 a_767_402.t0 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.1955 pd=1.565 as=0.063 ps=0.72 w=0.42 l=0.15
X36 a_1940_74.t2 a_1321_392.t9 VPWR.t12 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2352 ps=2.24 w=0.84 l=0.15
X37 Q.t4 a_1940_74.t9 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 a_1940_74.n13 a_1940_74.n12 310.733
R1 a_1940_74.n8 a_1940_74.t4 278.426
R2 a_1940_74.n2 a_1940_74.t8 244.524
R3 a_1940_74.n6 a_1940_74.n1 234.841
R4 a_1940_74.n9 a_1940_74.t3 234.841
R5 a_1940_74.n3 a_1940_74.t9 232.466
R6 a_1940_74.n2 a_1940_74.t5 186.374
R7 a_1940_74.n12 a_1940_74.t1 172.901
R8 a_1940_74.n5 a_1940_74.n0 165.189
R9 a_1940_74.n8 a_1940_74.t7 155.847
R10 a_1940_74.n4 a_1940_74.t6 155.847
R11 a_1940_74.n11 a_1940_74.n10 152
R12 a_1940_74.n7 a_1940_74.n0 152
R13 a_1940_74.n3 a_1940_74.n2 54.3023
R14 a_1940_74.n10 a_1940_74.n7 38.5605
R15 a_1940_74.t0 a_1940_74.n13 35.1791
R16 a_1940_74.n13 a_1940_74.t2 35.1791
R17 a_1940_74.n12 a_1940_74.n11 30.255
R18 a_1940_74.n6 a_1940_74.n5 30.0546
R19 a_1940_74.n11 a_1940_74.n0 13.1884
R20 a_1940_74.n4 a_1940_74.n3 10.6823
R21 a_1940_74.n5 a_1940_74.n4 10.2076
R22 a_1940_74.n7 a_1940_74.n6 8.50638
R23 a_1940_74.n9 a_1940_74.n8 6.23815
R24 a_1940_74.n10 a_1940_74.n9 3.96991
R25 Q.n1 Q.t6 270.442
R26 Q.n1 Q.n0 203.242
R27 Q.n4 Q.n2 176.218
R28 Q.n4 Q.n3 100.547
R29 Q.n3 Q.t1 30.0005
R30 Q Q.n4 27.6465
R31 Q.n0 Q.t5 26.3844
R32 Q.n0 Q.t4 26.3844
R33 Q.n2 Q.t0 22.7032
R34 Q.n2 Q.t3 22.7032
R35 Q.n3 Q.t2 22.7032
R36 Q Q.n1 15.3217
R37 VPWR.n27 VPWR.t10 681.726
R38 VPWR.n54 VPWR.t8 678.63
R39 VPWR.n45 VPWR.n5 627.761
R40 VPWR.n38 VPWR.n8 620.938
R41 VPWR.n12 VPWR.n11 617.378
R42 VPWR.n52 VPWR.n2 607.885
R43 VPWR.n14 VPWR.t12 436.861
R44 VPWR.n18 VPWR.t1 349.418
R45 VPWR.n17 VPWR.t0 343.442
R46 VPWR.n5 VPWR.t7 290.81
R47 VPWR.n21 VPWR.n16 239.084
R48 VPWR.n8 VPWR.t14 180.583
R49 VPWR.n5 VPWR.t4 77.3934
R50 VPWR.n11 VPWR.t5 70.3576
R51 VPWR.n11 VPWR.t3 70.3576
R52 VPWR.n16 VPWR.t11 52.3396
R53 VPWR.n8 VPWR.t6 47.7026
R54 VPWR.n40 VPWR.n39 36.1417
R55 VPWR.n40 VPWR.n6 36.1417
R56 VPWR.n44 VPWR.n6 36.1417
R57 VPWR.n47 VPWR.n46 36.1417
R58 VPWR.n47 VPWR.n3 36.1417
R59 VPWR.n51 VPWR.n3 36.1417
R60 VPWR.n32 VPWR.n31 36.1417
R61 VPWR.n33 VPWR.n32 36.1417
R62 VPWR.n33 VPWR.n9 36.1417
R63 VPWR.n37 VPWR.n9 36.1417
R64 VPWR.n46 VPWR.n45 35.3887
R65 VPWR.n28 VPWR.n12 32.377
R66 VPWR.n22 VPWR.n21 30.4946
R67 VPWR.n26 VPWR.n14 29.7417
R68 VPWR.n16 VPWR.t2 29.7402
R69 VPWR.n28 VPWR.n27 28.6123
R70 VPWR.n53 VPWR.n52 28.2358
R71 VPWR.n2 VPWR.t9 26.3844
R72 VPWR.n2 VPWR.t13 26.3844
R73 VPWR.n20 VPWR.n17 25.977
R74 VPWR.n27 VPWR.n26 24.8476
R75 VPWR.n22 VPWR.n14 23.7181
R76 VPWR.n54 VPWR.n53 22.9652
R77 VPWR.n21 VPWR.n20 20.7064
R78 VPWR.n52 VPWR.n51 19.2005
R79 VPWR.n39 VPWR.n38 12.0476
R80 VPWR.n20 VPWR.n19 9.3005
R81 VPWR.n21 VPWR.n15 9.3005
R82 VPWR.n23 VPWR.n22 9.3005
R83 VPWR.n24 VPWR.n14 9.3005
R84 VPWR.n26 VPWR.n25 9.3005
R85 VPWR.n27 VPWR.n13 9.3005
R86 VPWR.n29 VPWR.n28 9.3005
R87 VPWR.n31 VPWR.n30 9.3005
R88 VPWR.n32 VPWR.n10 9.3005
R89 VPWR.n34 VPWR.n33 9.3005
R90 VPWR.n35 VPWR.n9 9.3005
R91 VPWR.n37 VPWR.n36 9.3005
R92 VPWR.n39 VPWR.n7 9.3005
R93 VPWR.n41 VPWR.n40 9.3005
R94 VPWR.n42 VPWR.n6 9.3005
R95 VPWR.n44 VPWR.n43 9.3005
R96 VPWR.n46 VPWR.n4 9.3005
R97 VPWR.n48 VPWR.n47 9.3005
R98 VPWR.n49 VPWR.n3 9.3005
R99 VPWR.n51 VPWR.n50 9.3005
R100 VPWR.n52 VPWR.n1 9.3005
R101 VPWR.n53 VPWR.n0 9.3005
R102 VPWR.n55 VPWR.n54 7.27223
R103 VPWR.n18 VPWR.n17 6.46335
R104 VPWR.n38 VPWR.n37 4.51815
R105 VPWR.n31 VPWR.n12 3.76521
R106 VPWR.n45 VPWR.n44 0.753441
R107 VPWR.n19 VPWR.n18 0.686829
R108 VPWR VPWR.n55 0.157962
R109 VPWR.n55 VPWR.n0 0.149814
R110 VPWR.n19 VPWR.n15 0.122949
R111 VPWR.n23 VPWR.n15 0.122949
R112 VPWR.n24 VPWR.n23 0.122949
R113 VPWR.n25 VPWR.n24 0.122949
R114 VPWR.n25 VPWR.n13 0.122949
R115 VPWR.n29 VPWR.n13 0.122949
R116 VPWR.n30 VPWR.n29 0.122949
R117 VPWR.n30 VPWR.n10 0.122949
R118 VPWR.n34 VPWR.n10 0.122949
R119 VPWR.n35 VPWR.n34 0.122949
R120 VPWR.n36 VPWR.n35 0.122949
R121 VPWR.n36 VPWR.n7 0.122949
R122 VPWR.n41 VPWR.n7 0.122949
R123 VPWR.n42 VPWR.n41 0.122949
R124 VPWR.n43 VPWR.n42 0.122949
R125 VPWR.n43 VPWR.n4 0.122949
R126 VPWR.n48 VPWR.n4 0.122949
R127 VPWR.n49 VPWR.n48 0.122949
R128 VPWR.n50 VPWR.n49 0.122949
R129 VPWR.n50 VPWR.n1 0.122949
R130 VPWR.n1 VPWR.n0 0.122949
R131 VPB.t9 VPB.t15 531.183
R132 VPB.t8 VPB.t14 515.861
R133 VPB.t11 VPB.t13 497.985
R134 VPB.t5 VPB.t11 497.985
R135 VPB.t4 VPB.t7 477.555
R136 VPB.t2 VPB.t0 459.678
R137 VPB.t17 VPB.t16 406.048
R138 VPB.t18 VPB.t6 365.188
R139 VPB.t12 VPB.t2 265.591
R140 VPB.t6 VPB.t17 257.93
R141 VPB VPB.t8 257.93
R142 VPB.t15 VPB.t10 255.376
R143 VPB.t0 VPB.t1 229.839
R144 VPB.t13 VPB.t12 229.839
R145 VPB.t3 VPB.t5 229.839
R146 VPB.t7 VPB.t18 229.839
R147 VPB.t14 VPB.t9 229.839
R148 VPB.t16 VPB.t3 214.517
R149 VPB.t10 VPB.t4 214.517
R150 a_225_74.n0 a_225_74.t2 1129.75
R151 a_225_74.t1 a_225_74.n4 862.136
R152 a_225_74.n1 a_225_74.n0 747.101
R153 a_225_74.t2 a_225_74.t7 705.327
R154 a_225_74.n1 a_225_74.t5 359.894
R155 a_225_74.n2 a_225_74.t3 226.809
R156 a_225_74.n4 a_225_74.n3 206.178
R157 a_225_74.n2 a_225_74.t4 203.316
R158 a_225_74.n4 a_225_74.t0 198.974
R159 a_225_74.n0 a_225_74.t6 182.625
R160 a_225_74.n3 a_225_74.n1 54.7732
R161 a_225_74.n3 a_225_74.n2 21.1793
R162 a_1220_347.t0 a_1220_347.t1 80.7086
R163 a_1321_392.t1 a_1321_392.n0 813.662
R164 a_1321_392.n9 a_1321_392.t0 669.128
R165 a_1321_392.n2 a_1321_392.n1 286.337
R166 a_1321_392.n10 a_1321_392.n4 585
R167 a_1321_392.n5 a_1321_392.t7 303.661
R168 a_1321_392.n0 a_1321_392.n3 283.404
R169 a_1321_392.n7 a_1321_392.t5 243.411
R170 a_1321_392.n6 a_1321_392.t8 202.44
R171 a_1321_392.n7 a_1321_392.n6 171.16
R172 a_1321_392.n2 a_1321_392.n4 176.076
R173 a_1321_392.n5 a_1321_392.t9 159.06
R174 a_1321_392.n8 a_1321_392.t6 156.946
R175 a_1321_392.n10 a_1321_392.n9 78.7657
R176 a_1321_392.n4 a_1321_392.t4 70.3576
R177 a_1321_392.n9 a_1321_392.n8 66.7249
R178 a_1321_392.n3 a_1321_392.t2 62.8576
R179 a_1321_392.n8 a_1321_392.n7 35.0731
R180 a_1321_392.n1 a_1321_392.n0 25.6005
R181 a_1321_392.n3 a_1321_392.t3 22.0228
R182 a_1321_392.n1 a_1321_392.n10 9.20897
R183 a_1321_392.t1 a_1321_392.n2 20.0333
R184 a_1321_392.n6 a_1321_392.n5 4.8205
R185 a_398_74.t0 a_398_74.n3 884.077
R186 a_398_74.n2 a_398_74.t4 547.874
R187 a_398_74.n0 a_398_74.t1 380.079
R188 a_398_74.n3 a_398_74.n2 346.875
R189 a_398_74.n2 a_398_74.t3 314.274
R190 a_398_74.n1 a_398_74.t5 285.988
R191 a_398_74.n3 a_398_74.n1 210.163
R192 a_398_74.n0 a_398_74.t2 157.81
R193 a_398_74.n1 a_398_74.n0 103.18
R194 a_27_74.n1 a_27_74.t2 676.093
R195 a_27_74.n0 a_27_74.t1 666.771
R196 a_27_74.t0 a_27_74.n1 348.8
R197 a_27_74.n0 a_27_74.t3 340.469
R198 a_27_74.n1 a_27_74.n0 163.012
R199 a_612_74.n4 a_612_74.n3 671.212
R200 a_612_74.n1 a_612_74.t6 322.762
R201 a_612_74.n0 a_612_74.t5 243.679
R202 a_612_74.n2 a_612_74.n0 220.572
R203 a_612_74.n5 a_612_74.n4 213.161
R204 a_612_74.n0 a_612_74.t4 187.981
R205 a_612_74.n2 a_612_74.n1 152
R206 a_612_74.n1 a_612_74.t7 122.465
R207 a_612_74.n4 a_612_74.n2 114.624
R208 a_612_74.n3 a_612_74.t1 93.81
R209 a_612_74.n5 a_612_74.t2 88.5719
R210 a_612_74.n3 a_612_74.t3 70.3576
R211 a_612_74.t0 a_612_74.n5 40.0005
R212 a_1225_74.t0 a_1225_74.t1 74.063
R213 VNB.n0 VNB 15117.1
R214 VNB VNB.t17 13420
R215 VNB.t18 VNB.t2 2737.01
R216 VNB.t10 VNB.t12 2598.43
R217 VNB.t14 VNB.t15 2471.39
R218 VNB.t2 VNB.t1 2448.29
R219 VNB.t16 VNB.t7 2286.61
R220 VNB.t3 VNB.t4 1986.35
R221 VNB.t8 VNB.t14 1385.83
R222 VNB.t17 VNB.t11 1350.04
R223 VNB.t11 VNB.n0 1210
R224 VNB.t9 VNB.t13 1177.95
R225 VNB.t1 VNB.t6 1154.86
R226 VNB.t7 VNB 1143.31
R227 VNB.t4 VNB.t5 1097.11
R228 VNB.t6 VNB.t3 993.177
R229 VNB.t15 VNB.t16 993.177
R230 VNB.t0 VNB.t18 900.788
R231 VNB.t13 VNB.t0 900.788
R232 VNB.t17 VNB.t10 900.788
R233 VNB.t12 VNB.t8 900.788
R234 VNB.n0 VNB.t9 59.3797
R235 VGND.n58 VGND.t6 254.696
R236 VGND.n16 VGND.t4 250.792
R237 VGND.n4 VGND.t8 250.261
R238 VGND.n20 VGND.n19 185
R239 VGND.n18 VGND.n17 185
R240 VGND.n33 VGND.n32 185
R241 VGND.n31 VGND.n11 185
R242 VGND.n30 VGND.n29 185
R243 VGND.n7 VGND.n6 123.576
R244 VGND.n56 VGND.n2 122.118
R245 VGND.n23 VGND.n22 116.644
R246 VGND.n31 VGND.n30 98.5719
R247 VGND.n32 VGND.n31 97.1434
R248 VGND.n6 VGND.t11 76.0899
R249 VGND.n19 VGND.n18 69.7302
R250 VGND.n30 VGND.t0 60.0005
R251 VGND.n32 VGND.t12 40.0005
R252 VGND.n27 VGND.n12 36.1417
R253 VGND.n38 VGND.n9 36.1417
R254 VGND.n39 VGND.n38 36.1417
R255 VGND.n40 VGND.n39 36.1417
R256 VGND.n40 VGND.n7 36.1417
R257 VGND.n45 VGND.n44 36.1417
R258 VGND.n46 VGND.n45 36.1417
R259 VGND.n51 VGND.n50 36.1417
R260 VGND.n52 VGND.n51 36.1417
R261 VGND.n52 VGND.n1 36.1417
R262 VGND.n22 VGND.t5 34.0546
R263 VGND.n28 VGND.n27 32.0578
R264 VGND.n50 VGND.n4 32.0005
R265 VGND.n57 VGND.n56 31.2476
R266 VGND.n58 VGND.n57 30.4946
R267 VGND.n21 VGND.n20 29.9863
R268 VGND.n23 VGND.n12 25.6005
R269 VGND.n18 VGND.t3 22.7032
R270 VGND.n19 VGND.t2 22.7032
R271 VGND.n22 VGND.t1 22.7032
R272 VGND.n2 VGND.t9 22.7032
R273 VGND.n2 VGND.t10 22.7032
R274 VGND.n56 VGND.n1 22.2123
R275 VGND.n23 VGND.n21 21.8358
R276 VGND.n6 VGND.t7 20.5082
R277 VGND.n44 VGND.n7 11.2946
R278 VGND.n46 VGND.n4 10.5417
R279 VGND.n57 VGND.n0 9.3005
R280 VGND.n56 VGND.n55 9.3005
R281 VGND.n54 VGND.n1 9.3005
R282 VGND.n53 VGND.n52 9.3005
R283 VGND.n51 VGND.n3 9.3005
R284 VGND.n50 VGND.n49 9.3005
R285 VGND.n48 VGND.n4 9.3005
R286 VGND.n47 VGND.n46 9.3005
R287 VGND.n45 VGND.n5 9.3005
R288 VGND.n44 VGND.n43 9.3005
R289 VGND.n42 VGND.n7 9.3005
R290 VGND.n41 VGND.n40 9.3005
R291 VGND.n39 VGND.n8 9.3005
R292 VGND.n38 VGND.n37 9.3005
R293 VGND.n36 VGND.n9 9.3005
R294 VGND.n35 VGND.n34 9.3005
R295 VGND.n28 VGND.n10 9.3005
R296 VGND.n27 VGND.n26 9.3005
R297 VGND.n25 VGND.n12 9.3005
R298 VGND.n24 VGND.n23 9.3005
R299 VGND.n15 VGND.n14 9.3005
R300 VGND.n21 VGND.n13 9.3005
R301 VGND.n17 VGND.n16 7.81645
R302 VGND.n59 VGND.n58 7.19894
R303 VGND.n17 VGND.n14 6.14739
R304 VGND.n29 VGND.n11 5.84951
R305 VGND.n34 VGND.n33 5.08659
R306 VGND.n33 VGND.n9 3.92726
R307 VGND.n29 VGND.n28 1.6111
R308 VGND.n34 VGND.n11 0.678646
R309 VGND.n16 VGND.n15 0.582656
R310 VGND VGND.n59 0.156997
R311 VGND.n59 VGND.n0 0.150766
R312 VGND.n15 VGND.n13 0.122949
R313 VGND.n24 VGND.n13 0.122949
R314 VGND.n25 VGND.n24 0.122949
R315 VGND.n26 VGND.n25 0.122949
R316 VGND.n26 VGND.n10 0.122949
R317 VGND.n35 VGND.n10 0.122949
R318 VGND.n36 VGND.n35 0.122949
R319 VGND.n37 VGND.n36 0.122949
R320 VGND.n37 VGND.n8 0.122949
R321 VGND.n41 VGND.n8 0.122949
R322 VGND.n42 VGND.n41 0.122949
R323 VGND.n43 VGND.n42 0.122949
R324 VGND.n43 VGND.n5 0.122949
R325 VGND.n47 VGND.n5 0.122949
R326 VGND.n48 VGND.n47 0.122949
R327 VGND.n49 VGND.n48 0.122949
R328 VGND.n49 VGND.n3 0.122949
R329 VGND.n53 VGND.n3 0.122949
R330 VGND.n54 VGND.n53 0.122949
R331 VGND.n55 VGND.n54 0.122949
R332 VGND.n55 VGND.n0 0.122949
R333 VGND.n20 VGND.n14 0.0728164
R334 D.n0 D.t1 233.811
R335 D D.n0 161.504
R336 D.n1 D 154.522
R337 D.n3 D.n2 152
R338 D.n1 D.t0 148.927
R339 D.n2 D.n0 42.021
R340 D.n2 D.n1 42.021
R341 D.n3 D 10.6672
R342 D D.n3 3.68535
R343 SET_B.n1 SET_B.t1 297.841
R344 SET_B.n0 SET_B.t0 292.76
R345 SET_B.n0 SET_B.t2 251.285
R346 SET_B.n1 SET_B.t3 180.019
R347 SET_B SET_B.n1 169.185
R348 SET_B SET_B.n0 79.675
R349 a_767_402.n1 a_767_402.n0 801.658
R350 a_767_402.t2 a_767_402.n2 406.067
R351 a_767_402.n2 a_767_402.n1 199.227
R352 a_767_402.n2 a_767_402.t3 197.912
R353 a_767_402.n1 a_767_402.t4 197.352
R354 a_767_402.n0 a_767_402.t0 70.3576
R355 a_767_402.n0 a_767_402.t1 70.3576
R356 a_732_74.t0 a_732_74.t1 68.5719
R357 a_1484_62.n1 a_1484_62.t1 788.537
R358 a_1484_62.n0 a_1484_62.t3 325.959
R359 a_1484_62.n1 a_1484_62.n0 267.656
R360 a_1484_62.t0 a_1484_62.n1 235.667
R361 a_1484_62.n0 a_1484_62.t2 234.38
R362 a_1436_88.t0 a_1436_88.t1 68.5719
R363 a_1514_88.t0 a_1514_88.t1 68.5719
R364 a_1480_508.t0 a_1480_508.t1 126.644
R365 CLK.n0 CLK.t0 285.719
R366 CLK.n0 CLK.t1 178.34
R367 CLK CLK.n0 156.87
R368 a_1035_118.t0 a_1035_118.t1 68.5719
R369 a_716_463.t0 a_716_463.t1 126.644
C0 VPB VGND 0.025938f
C1 VGND Q 0.373059f
C2 D VGND 0.045351f
C3 VPB Q 0.0163f
C4 VPB D 0.11717f
C5 CLK VGND 0.034532f
C6 VPB CLK 0.033597f
C7 VPWR VGND 0.157985f
C8 D CLK 0.025591f
C9 VPB VPWR 0.371429f
C10 VPWR Q 0.418261f
C11 SET_B VGND 0.1259f
C12 D VPWR 0.017924f
C13 VPB SET_B 0.200379f
C14 SET_B Q 7.11e-20
C15 D SET_B 7.37e-20
C16 CLK VPWR 0.01799f
C17 CLK SET_B 6.29e-20
C18 VPWR SET_B 0.113433f
C19 Q VNB 0.075526f
C20 VGND VNB 1.53393f
C21 SET_B VNB 0.289225f
C22 VPWR VNB 1.17278f
C23 CLK VNB 0.115192f
C24 D VNB 0.214526f
C25 VPB VNB 2.99059f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfstp_2 VNB VPB VPWR SET_B VGND CLK D Q
X0 a_1596_118.t0 a_1566_92# a_1489_118.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.08085 ps=0.805 w=0.42 l=0.15
X1 VPWR.t5 a_767_384.t3 a_716_456.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.246825 pd=1.575 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND.t8 a_1356_74# a_2022_94.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 a_1489_118.t1 a_225_74.t2 a_1356_74# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.08085 pd=0.805 as=0.13565 ps=1.155 w=0.42 l=0.15
X4 VGND.t3 SET_B.t0 a_1596_118.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.17955 pd=1.275 as=0.0882 ps=0.84 w=0.42 l=0.15
X5 a_716_456.t0 a_225_74.t3 a_612_74.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR.t1 D.t0 a_27_74.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1239 ps=1.43 w=0.42 l=0.15
X7 VGND.t0 D.t1 a_27_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 a_1566_92# a_1356_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1239 ps=1.43 w=0.42 l=0.15
X9 a_1356_74# a_398_74.t2 a_1278_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.13565 pd=1.155 as=0.0768 ps=0.88 w=0.64 l=0.15
X10 a_612_74.t0 a_398_74.t3 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X11 a_767_384.t2 a_612_74.t4 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.246825 ps=1.575 w=0.42 l=0.15
X12 VPWR.t3 SET_B.t1 a_767_384.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2447 pd=1.88 as=0.063 ps=0.72 w=0.42 l=0.15
X13 VGND.t4 CLK.t0 a_225_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 VPWR.t0 a_1566_92# a_1521_508.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VPWR.t6 a_2022_94.t2 Q.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_1521_508.t1 a_398_74.t4 a_1356_74# VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.21575 ps=1.62 w=0.42 l=0.15
X17 a_1356_74# SET_B.t2 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.0819 ps=0.81 w=0.42 l=0.15
X18 VGND.t6 a_2022_94.t3 Q.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2294 pd=2.1 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_398_74.t1 a_225_74.t4 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_1266_341.t0 a_612_74.t5 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1998 pd=1.61 as=0.2447 ps=1.88 w=1 l=0.15
X21 VPWR.t10 a_1356_74# a_2022_94.t0 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.295 ps=2.59 w=1 l=0.15
X22 VGND.t7 a_767_384.t4 a_781_74.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 VPWR.t9 CLK.t1 a_225_74.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X24 a_398_74.t0 a_225_74.t5 VGND.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 a_1057_118.t0 a_612_74.t6 a_767_384.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X26 a_1566_92# a_1356_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.17955 ps=1.275 w=0.42 l=0.15
X27 a_781_74.t0 a_398_74.t5 a_612_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.14595 ps=1.115 w=0.42 l=0.15
X28 a_612_74.t3 a_225_74.t6 a_27_74.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.14595 pd=1.115 as=0.18665 ps=1.8 w=0.42 l=0.15
X29 Q.t0 a_2022_94.t4 VGND.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.15535 ps=1.17 w=0.74 l=0.15
X30 a_1278_74.t0 a_612_74.t7 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1522 ps=1.205 w=0.64 l=0.15
R0 a_1489_118.t0 a_1489_118.t1 110.001
R1 a_1596_118.t0 a_1596_118.t1 120.001
R2 VNB.t1 VNB 15486.6
R3 VNB VNB.n0 14256.5
R4 VNB.t10 VNB.t14 4607.87
R5 VNB.t9 VNB.t8 2538.01
R6 VNB.t4 VNB.t12 2348.25
R7 VNB.t11 VNB.t0 2348.25
R8 VNB.t3 VNB.t9 2004.31
R9 VNB.t1 VNB.t7 1458.09
R10 VNB.n0 VNB.t5 1441.81
R11 VNB.t14 VNB.t13 1339.63
R12 VNB.t2 VNB.t10 1316.54
R13 VNB.n0 VNB.t4 1245.28
R14 VNB.t7 VNB.t2 1235.7
R15 VNB.t0 VNB 1174.12
R16 VNB.t8 VNB.t11 1019.95
R17 VNB.t13 VNB.t6 993.177
R18 VNB.t5 VNB.t1 969.492
R19 VNB.t12 VNB.t3 925.067
R20 a_767_384.n1 a_767_384.n0 795.544
R21 a_767_384.t0 a_767_384.n2 390.132
R22 a_767_384.n1 a_767_384.t3 241
R23 a_767_384.n2 a_767_384.n1 201.125
R24 a_767_384.n2 a_767_384.t4 177.025
R25 a_767_384.n0 a_767_384.t1 70.3576
R26 a_767_384.n0 a_767_384.t2 70.3576
R27 a_716_456.t0 a_716_456.t1 126.644
R28 VPWR.n9 VPWR.n8 694.966
R29 VPWR.n47 VPWR.t1 677.66
R30 VPWR.n6 VPWR.n5 616.624
R31 VPWR.n45 VPWR.n2 608.274
R32 VPWR.n23 VPWR.n13 605.17
R33 VPWR.n16 VPWR.t10 362.695
R34 VPWR.n5 VPWR.t7 268.204
R35 VPWR.n17 VPWR.t6 266.168
R36 VPWR.n8 VPWR.t3 199.345
R37 VPWR.n5 VPWR.t5 116.493
R38 VPWR.n13 VPWR.t0 112.572
R39 VPWR.n13 VPWR.t4 70.3576
R40 VPWR.n8 VPWR.t8 43.6029
R41 VPWR.n34 VPWR.n33 36.1417
R42 VPWR.n35 VPWR.n34 36.1417
R43 VPWR.n39 VPWR.n38 36.1417
R44 VPWR.n40 VPWR.n39 36.1417
R45 VPWR.n40 VPWR.n3 36.1417
R46 VPWR.n44 VPWR.n3 36.1417
R47 VPWR.n27 VPWR.n11 36.1417
R48 VPWR.n28 VPWR.n27 36.1417
R49 VPWR.n29 VPWR.n28 36.1417
R50 VPWR.n20 VPWR.n15 36.1417
R51 VPWR.n23 VPWR.n22 33.8829
R52 VPWR.n35 VPWR.n6 30.4946
R53 VPWR.n21 VPWR.n20 30.1181
R54 VPWR.n46 VPWR.n45 28.2358
R55 VPWR.n29 VPWR.n9 27.8593
R56 VPWR.n2 VPWR.t2 26.3844
R57 VPWR.n2 VPWR.t9 26.3844
R58 VPWR.n33 VPWR.n9 25.6005
R59 VPWR.n16 VPWR.n15 25.224
R60 VPWR.n47 VPWR.n46 22.9652
R61 VPWR.n45 VPWR.n44 19.2005
R62 VPWR.n22 VPWR.n21 17.3181
R63 VPWR.n23 VPWR.n11 13.5534
R64 VPWR.n18 VPWR.n15 9.3005
R65 VPWR.n20 VPWR.n19 9.3005
R66 VPWR.n21 VPWR.n14 9.3005
R67 VPWR.n22 VPWR.n12 9.3005
R68 VPWR.n24 VPWR.n23 9.3005
R69 VPWR.n25 VPWR.n11 9.3005
R70 VPWR.n27 VPWR.n26 9.3005
R71 VPWR.n28 VPWR.n10 9.3005
R72 VPWR.n30 VPWR.n29 9.3005
R73 VPWR.n31 VPWR.n9 9.3005
R74 VPWR.n33 VPWR.n32 9.3005
R75 VPWR.n34 VPWR.n7 9.3005
R76 VPWR.n36 VPWR.n35 9.3005
R77 VPWR.n38 VPWR.n37 9.3005
R78 VPWR.n39 VPWR.n4 9.3005
R79 VPWR.n41 VPWR.n40 9.3005
R80 VPWR.n42 VPWR.n3 9.3005
R81 VPWR.n44 VPWR.n43 9.3005
R82 VPWR.n45 VPWR.n1 9.3005
R83 VPWR.n46 VPWR.n0 9.3005
R84 VPWR.n48 VPWR.n47 7.27223
R85 VPWR.n17 VPWR.n16 6.59649
R86 VPWR.n38 VPWR.n6 5.64756
R87 VPWR.n18 VPWR.n17 0.612104
R88 VPWR VPWR.n48 0.157962
R89 VPWR.n48 VPWR.n0 0.149814
R90 VPWR.n19 VPWR.n18 0.122949
R91 VPWR.n19 VPWR.n14 0.122949
R92 VPWR.n14 VPWR.n12 0.122949
R93 VPWR.n24 VPWR.n12 0.122949
R94 VPWR.n25 VPWR.n24 0.122949
R95 VPWR.n26 VPWR.n25 0.122949
R96 VPWR.n26 VPWR.n10 0.122949
R97 VPWR.n30 VPWR.n10 0.122949
R98 VPWR.n31 VPWR.n30 0.122949
R99 VPWR.n32 VPWR.n31 0.122949
R100 VPWR.n32 VPWR.n7 0.122949
R101 VPWR.n36 VPWR.n7 0.122949
R102 VPWR.n37 VPWR.n36 0.122949
R103 VPWR.n37 VPWR.n4 0.122949
R104 VPWR.n41 VPWR.n4 0.122949
R105 VPWR.n42 VPWR.n41 0.122949
R106 VPWR.n43 VPWR.n42 0.122949
R107 VPWR.n43 VPWR.n1 0.122949
R108 VPWR.n1 VPWR.n0 0.122949
R109 VPB.n0 VPB 3460.35
R110 VPB.t7 VPB.t13 1031.72
R111 VPB.t8 VPB.t10 554.582
R112 VPB.t5 VPB.t0 517.279
R113 VPB.t13 VPB.t9 503.091
R114 VPB VPB.n1 479.974
R115 VPB.n0 VPB.t3 385.618
R116 VPB.t6 VPB.t11 380.498
R117 VPB.t1 VPB.t7 275.807
R118 VPB.n1 VPB.t12 273.56
R119 VPB.t11 VPB.n0 258.639
R120 VPB.t2 VPB 257.93
R121 VPB.t0 VPB.t4 248.691
R122 VPB.n1 VPB.t2 234.946
R123 VPB.t10 VPB.t6 223.822
R124 VPB.t12 VPB.t5 223.822
R125 VPB.t3 VPB.t1 214.517
R126 VPB.t4 VPB.t8 208.901
R127 a_2022_94.t0 a_2022_94.n3 249.915
R128 a_2022_94.n2 a_2022_94.t2 242.388
R129 a_2022_94.n0 a_2022_94.n1 240.197
R130 a_2022_94.n3 a_2022_94.n0 182.589
R131 a_2022_94.n0 a_2022_94.t4 179.947
R132 a_2022_94.n2 a_2022_94.t3 179.947
R133 a_2022_94.n3 a_2022_94.t1 151.512
R134 a_2022_94.n0 a_2022_94.n2 63.5369
R135 VGND.n21 VGND.n20 329.286
R136 VGND.n47 VGND.t0 254.696
R137 VGND.n35 VGND.t7 245.559
R138 VGND.n22 VGND.n21 185
R139 VGND.n12 VGND.t6 174.998
R140 VGND.n6 VGND.t1 150.822
R141 VGND.n45 VGND.n2 122.118
R142 VGND.n14 VGND.n13 116.644
R143 VGND.n13 VGND.t8 41.2505
R144 VGND.n21 VGND.t3 40.0005
R145 VGND.n15 VGND.n11 36.1417
R146 VGND.n19 VGND.n11 36.1417
R147 VGND.n23 VGND.n8 36.1417
R148 VGND.n27 VGND.n8 36.1417
R149 VGND.n28 VGND.n27 36.1417
R150 VGND.n29 VGND.n28 36.1417
R151 VGND.n34 VGND.n33 36.1417
R152 VGND.n39 VGND.n4 36.1417
R153 VGND.n40 VGND.n39 36.1417
R154 VGND.n41 VGND.n40 36.1417
R155 VGND.n41 VGND.n1 36.1417
R156 VGND.n35 VGND.n34 33.1299
R157 VGND.n46 VGND.n45 31.2476
R158 VGND.n47 VGND.n46 30.4946
R159 VGND.n13 VGND.t5 30.2643
R160 VGND.n2 VGND.t2 22.7032
R161 VGND.n2 VGND.t4 22.7032
R162 VGND.n45 VGND.n1 22.2123
R163 VGND.n15 VGND.n14 21.0829
R164 VGND.n29 VGND.n6 17.6946
R165 VGND.n35 VGND.n4 14.3064
R166 VGND.n23 VGND.n22 11.5564
R167 VGND.n33 VGND.n6 9.78874
R168 VGND.n46 VGND.n0 9.3005
R169 VGND.n45 VGND.n44 9.3005
R170 VGND.n43 VGND.n1 9.3005
R171 VGND.n42 VGND.n41 9.3005
R172 VGND.n40 VGND.n3 9.3005
R173 VGND.n39 VGND.n38 9.3005
R174 VGND.n37 VGND.n4 9.3005
R175 VGND.n36 VGND.n35 9.3005
R176 VGND.n34 VGND.n5 9.3005
R177 VGND.n33 VGND.n32 9.3005
R178 VGND.n31 VGND.n6 9.3005
R179 VGND.n30 VGND.n29 9.3005
R180 VGND.n28 VGND.n7 9.3005
R181 VGND.n27 VGND.n26 9.3005
R182 VGND.n25 VGND.n8 9.3005
R183 VGND.n24 VGND.n23 9.3005
R184 VGND.n10 VGND.n9 9.3005
R185 VGND.n19 VGND.n18 9.3005
R186 VGND.n17 VGND.n11 9.3005
R187 VGND.n16 VGND.n15 9.3005
R188 VGND.n48 VGND.n47 7.19894
R189 VGND.n14 VGND.n12 6.8559
R190 VGND.n20 VGND.n10 4.0939
R191 VGND.n22 VGND.n10 2.46954
R192 VGND.n20 VGND.n19 2.14466
R193 VGND.n16 VGND.n12 0.565232
R194 VGND VGND.n48 0.156997
R195 VGND.n48 VGND.n0 0.150766
R196 VGND.n17 VGND.n16 0.122949
R197 VGND.n18 VGND.n17 0.122949
R198 VGND.n18 VGND.n9 0.122949
R199 VGND.n24 VGND.n9 0.122949
R200 VGND.n25 VGND.n24 0.122949
R201 VGND.n26 VGND.n25 0.122949
R202 VGND.n26 VGND.n7 0.122949
R203 VGND.n30 VGND.n7 0.122949
R204 VGND.n31 VGND.n30 0.122949
R205 VGND.n32 VGND.n31 0.122949
R206 VGND.n32 VGND.n5 0.122949
R207 VGND.n36 VGND.n5 0.122949
R208 VGND.n37 VGND.n36 0.122949
R209 VGND.n38 VGND.n37 0.122949
R210 VGND.n38 VGND.n3 0.122949
R211 VGND.n42 VGND.n3 0.122949
R212 VGND.n43 VGND.n42 0.122949
R213 VGND.n44 VGND.n43 0.122949
R214 VGND.n44 VGND.n0 0.122949
R215 a_225_74.n1 a_225_74.n0 1203.66
R216 a_225_74.t1 a_225_74.n5 862.136
R217 a_225_74.n2 a_225_74.n1 763.168
R218 a_225_74.n0 a_225_74.t2 668.374
R219 a_225_74.n2 a_225_74.t6 343.827
R220 a_225_74.n3 a_225_74.t4 226.809
R221 a_225_74.n5 a_225_74.n4 209.123
R222 a_225_74.n5 a_225_74.t0 202.351
R223 a_225_74.n1 a_225_74.t3 191.998
R224 a_225_74.n3 a_225_74.t5 187.25
R225 a_225_74.n4 a_225_74.n2 54.7732
R226 a_225_74.n4 a_225_74.n3 21.1793
R227 SET_B.n2 SET_B.n1 340.524
R228 SET_B.n0 SET_B.t0 264.767
R229 SET_B.n0 SET_B.t2 220.761
R230 SET_B SET_B.n2 177.874
R231 SET_B.n2 SET_B.t1 136.744
R232 SET_B SET_B.n0 78.7135
R233 a_612_74.n4 a_612_74.n3 676.015
R234 a_612_74.n1 a_612_74.t4 290.716
R235 a_612_74.n0 a_612_74.t5 224.272
R236 a_612_74.n5 a_612_74.n4 205.946
R237 a_612_74.n2 a_612_74.n0 187.292
R238 a_612_74.n0 a_612_74.t7 185.444
R239 a_612_74.n1 a_612_74.t6 158.701
R240 a_612_74.n2 a_612_74.n1 152
R241 a_612_74.n4 a_612_74.n2 120.859
R242 a_612_74.n5 a_612_74.t3 111.43
R243 a_612_74.n3 a_612_74.t0 93.81
R244 a_612_74.t1 a_612_74.n5 87.1434
R245 a_612_74.n3 a_612_74.t2 70.3576
R246 D.n0 D.t0 239.167
R247 D D.n0 161.504
R248 D.n1 D 154.522
R249 D.n3 D.n2 152
R250 D.n1 D.t1 148.927
R251 D.n2 D.n0 42.021
R252 D.n2 D.n1 42.021
R253 D.n3 D 10.6672
R254 D D.n3 3.68535
R255 a_27_74.n1 a_27_74.t2 679.678
R256 a_27_74.n0 a_27_74.t0 664.573
R257 a_27_74.t1 a_27_74.n1 346.118
R258 a_27_74.n0 a_27_74.t3 339.716
R259 a_27_74.n1 a_27_74.n0 157.465
R260 a_1266_341.n0 a_1266_341.t0 69.3667
R261 a_398_74.t1 a_398_74.n3 966.638
R262 a_398_74.n0 a_398_74.t4 549.559
R263 a_398_74.n1 a_398_74.t0 373.961
R264 a_398_74.n3 a_398_74.n0 330.276
R265 a_398_74.n0 a_398_74.t2 314.274
R266 a_398_74.n2 a_398_74.t5 265.83
R267 a_398_74.n3 a_398_74.n2 186.429
R268 a_398_74.n1 a_398_74.t3 169.506
R269 a_398_74.n2 a_398_74.n1 131.107
R270 a_1278_74.t0 a_1278_74.t1 45.0005
R271 CLK.n0 CLK.t1 272.33
R272 CLK.n0 CLK.t0 178.34
R273 CLK CLK.n0 156.87
R274 a_1521_508.t0 a_1521_508.t1 126.644
R275 Q.n1 Q.t2 227.394
R276 Q.n1 Q.n0 157.274
R277 Q.n0 Q.t1 22.7032
R278 Q.n0 Q.t0 22.7032
R279 Q Q.n1 3.9258
R280 a_781_74.t0 a_781_74.t1 68.5719
C0 a_1356_74# VGND 0.044435f
C1 VPB D 0.120753f
C2 a_1566_92# a_1356_74# 0.207845f
C3 a_1356_74# Q 0.00637f
C4 VPB VPWR 0.328837f
C5 VPB CLK 0.034679f
C6 D VPWR 0.019449f
C7 D CLK 0.023743f
C8 VPB SET_B 0.202273f
C9 VPWR CLK 0.0175f
C10 VPB VGND 0.030663f
C11 D SET_B 5.06e-20
C12 a_1566_92# VPB 0.108376f
C13 VPB Q 0.008184f
C14 VPWR SET_B 0.131547f
C15 D VGND 0.042139f
C16 a_1356_74# VPB 0.259859f
C17 CLK SET_B 5.46e-20
C18 VPWR VGND 0.159513f
C19 a_1566_92# VPWR 0.070472f
C20 CLK VGND 0.034572f
C21 VPWR Q 0.227948f
C22 a_1356_74# VPWR 0.305798f
C23 SET_B VGND 0.091486f
C24 a_1566_92# SET_B 0.232617f
C25 SET_B Q 4.62e-19
C26 a_1356_74# SET_B 0.183363f
C27 a_1566_92# VGND 0.152923f
C28 VGND Q 0.172216f
C29 Q VNB 0.031262f
C30 VGND VNB 1.47264f
C31 SET_B VNB 0.224742f
C32 CLK VNB 0.110888f
C33 VPWR VNB 1.11319f
C34 D VNB 0.213977f
C35 VPB VNB 2.80868f
C36 a_1356_74# VNB 0.328164f
C37 a_1566_92# VNB 0.165118f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfstp_1 VNB VPB VPWR SET_B VGND Q D CLK
X0 a_1298_392.t3 a_224_350.t2 a_1197_341.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.21665 pd=1.645 as=0.1998 ps=1.61 w=1 l=0.15
X1 VGND.t3 a_760_395.t3 a_740_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1449 pd=1.53 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 VGND.t4 SET_B.t0 a_1027_118.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.12165 pd=1.07 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 a_740_74.t0 a_398_74.t2 a_604_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1113 ps=0.95 w=0.42 l=0.15
X4 a_1027_118.t1 a_604_74.t4 a_760_395.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1176 ps=1.4 w=0.42 l=0.15
X5 a_1298_392.t0 a_398_74.t3 a_1215_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10695 pd=1 as=0.12 ps=1.015 w=0.64 l=0.15
X6 VGND.t5 SET_B.t1 a_1500_74.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.19215 pd=1.335 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 VGND.t0 D.t0 a_27_74.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X8 a_1500_74.t1 a_1470_48# a_1422_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 VGND.t6 a_1298_392.t4 a_1902_74.t0 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X10 VPWR.t7 a_1470_48# a_1457_508.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1197_341.t1 a_604_74.t5 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1998 pd=1.61 as=0.23615 ps=1.86 w=1 l=0.15
X12 a_1457_508.t0 a_398_74.t4 a_1298_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.21665 ps=1.645 w=0.42 l=0.15
X13 VPWR.t2 a_760_395.t4 a_709_463.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.14175 pd=1.095 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VGND.t1 CLK.t0 a_224_350.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 a_604_74.t2 a_224_350.t3 a_27_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.17595 ps=1.76 w=0.42 l=0.15
X16 VPWR.t8 a_1298_392.t5 a_1902_74.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1946 pd=1.49 as=0.231 ps=2.23 w=0.84 l=0.15
X17 a_1470_48# a_1298_392.t6 VPWR.t9 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.39 as=0.1176 ps=1.4 w=0.42 l=0.15
X18 a_709_463.t0 a_224_350.t4 a_604_74.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0735 ps=0.77 w=0.42 l=0.15
X19 a_398_74.t1 a_224_350.t5 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_398_74.t0 a_224_350.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VPWR.t0 CLK.t1 a_224_350.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X22 a_1422_74.t0 a_224_350.t7 a_1298_392.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.10695 ps=1 w=0.42 l=0.15
X23 Q.t0 a_1902_74.t2 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X24 a_760_395.t2 a_604_74.t6 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.14175 ps=1.095 w=0.42 l=0.15
X25 VPWR.t4 D.t1 a_27_74.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.1197 ps=1.41 w=0.42 l=0.15
X26 VPWR.t3 SET_B.t2 a_760_395.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.23615 pd=1.86 as=0.063 ps=0.72 w=0.42 l=0.15
X27 Q.t1 a_1902_74.t3 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1946 ps=1.49 w=1.12 l=0.15
X28 a_604_74.t0 a_398_74.t5 a_27_74.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
R0 a_224_350.n0 a_224_350.t2 1104.05
R1 a_224_350.t0 a_224_350.n4 871.861
R2 a_224_350.n1 a_224_350.n0 776.02
R3 a_224_350.t2 a_224_350.t7 742.28
R4 a_224_350.n1 a_224_350.t3 329.368
R5 a_224_350.n2 a_224_350.t5 226.809
R6 a_224_350.n4 a_224_350.n3 215.493
R7 a_224_350.n4 a_224_350.t1 198.404
R8 a_224_350.n0 a_224_350.t4 182.625
R9 a_224_350.n2 a_224_350.t6 169.285
R10 a_224_350.n3 a_224_350.n1 43.8187
R11 a_224_350.n3 a_224_350.n2 32.1338
R12 a_1197_341.t0 a_1197_341.t1 82.5648
R13 a_1298_392.t3 a_1298_392.n3 799.59
R14 a_1298_392.n13 a_1298_392.n4 591.394
R15 a_1298_392.n10 a_1298_392.n5 585
R16 a_1298_392.n12 a_1298_392.n11 585
R17 a_1298_392.n6 a_1298_392.t4 367.928
R18 a_1298_392.n3 a_1298_392.n2 272.269
R19 a_1298_392.n1 a_1298_392.n6 242.607
R20 a_1298_392.n6 a_1298_392.t5 208.868
R21 a_1298_392.n12 a_1298_392.n5 161.821
R22 a_1298_392.n9 a_1298_392.n8 152
R23 a_1298_392.n1 a_1298_392.n0 20.052
R24 a_1298_392.n8 a_1298_392.t6 137.454
R25 a_1298_392.n10 a_1298_392.n9 107.034
R26 a_1298_392.n5 a_1298_392.t1 70.3576
R27 a_1298_392.n2 a_1298_392.t2 62.8576
R28 a_1298_392.n8 a_1298_392.n1 48.2005
R29 a_1298_392.n0 a_1298_392.n7 299.036
R30 a_1298_392.n2 a_1298_392.t0 26.2505
R31 a_1298_392.n13 a_1298_392.n12 21.7396
R32 a_1298_392.t3 a_1298_392.n13 13.2606
R33 a_1298_392.n9 a_1298_392.n0 81.9064
R34 a_1298_392.n4 a_1298_392.n3 12.9915
R35 a_1298_392.n11 a_1298_392.n10 12.4399
R36 a_1298_392.n11 a_1298_392.n4 4.96766
R37 VPB.t3 VPB.t2 506.668
R38 VPB VPB.n0 457.95
R39 VPB.t6 VPB.t10 401.923
R40 VPB.t8 VPB.t9 362.95
R41 VPB.n0 VPB.t0 263.077
R42 VPB.t7 VPB 252.823
R43 VPB.t9 VPB.t5 246.026
R44 VPB.t2 VPB.t4 243.59
R45 VPB.n0 VPB.t7 227.286
R46 VPB.t10 VPB.t8 219.232
R47 VPB.t0 VPB.t3 219.232
R48 VPB.t4 VPB.t6 204.615
R49 VPB.t1 VPB 66.3026
R50 VPB.t5 VPB.t1 37.3584
R51 VPB.t11 VPB.t12 6.92758
R52 VPB.t5 VPB.t11 4.94842
R53 a_760_395.n1 a_760_395.n0 819.014
R54 a_760_395.t1 a_760_395.n2 391.046
R55 a_760_395.n1 a_760_395.t4 217.971
R56 a_760_395.n2 a_760_395.t3 185.571
R57 a_760_395.n2 a_760_395.n1 168.445
R58 a_760_395.n0 a_760_395.t0 70.3576
R59 a_760_395.n0 a_760_395.t2 70.3576
R60 a_740_74.t0 a_740_74.t1 68.5719
R61 VGND.n14 VGND.n13 345
R62 VGND.n40 VGND.t0 254.696
R63 VGND.n29 VGND.t3 250.475
R64 VGND.n22 VGND.t4 205.387
R65 VGND.n15 VGND.n14 185
R66 VGND.n2 VGND.n1 129.522
R67 VGND.n12 VGND.n11 123.999
R68 VGND.n11 VGND.t6 50.9375
R69 VGND.n14 VGND.t5 41.4291
R70 VGND.n20 VGND.n8 36.1417
R71 VGND.n21 VGND.n20 36.1417
R72 VGND.n23 VGND.n21 36.1417
R73 VGND.n27 VGND.n6 36.1417
R74 VGND.n28 VGND.n27 36.1417
R75 VGND.n33 VGND.n4 36.1417
R76 VGND.n34 VGND.n33 36.1417
R77 VGND.n35 VGND.n34 36.1417
R78 VGND.n39 VGND.n38 36.1417
R79 VGND.n29 VGND.n4 35.0123
R80 VGND.n35 VGND.n2 34.6358
R81 VGND.n16 VGND.n8 33.3113
R82 VGND.n11 VGND.t7 32.6953
R83 VGND.n40 VGND.n39 30.4946
R84 VGND.n1 VGND.t2 22.7032
R85 VGND.n1 VGND.t1 22.7032
R86 VGND.n13 VGND.n12 19.6902
R87 VGND.n39 VGND.n0 9.3005
R88 VGND.n38 VGND.n37 9.3005
R89 VGND.n36 VGND.n35 9.3005
R90 VGND.n34 VGND.n3 9.3005
R91 VGND.n33 VGND.n32 9.3005
R92 VGND.n31 VGND.n4 9.3005
R93 VGND.n30 VGND.n29 9.3005
R94 VGND.n28 VGND.n5 9.3005
R95 VGND.n27 VGND.n26 9.3005
R96 VGND.n25 VGND.n6 9.3005
R97 VGND.n10 VGND.n9 9.3005
R98 VGND.n17 VGND.n16 9.3005
R99 VGND.n18 VGND.n8 9.3005
R100 VGND.n20 VGND.n19 9.3005
R101 VGND.n21 VGND.n7 9.3005
R102 VGND.n24 VGND.n23 9.3005
R103 VGND.n29 VGND.n28 7.90638
R104 VGND.n22 VGND.n6 7.52991
R105 VGND.n41 VGND.n40 7.19894
R106 VGND.n15 VGND.n10 6.82094
R107 VGND.n23 VGND.n22 3.76521
R108 VGND.n13 VGND.n10 3.6443
R109 VGND.n16 VGND.n15 2.14941
R110 VGND.n38 VGND.n2 1.50638
R111 VGND.n12 VGND.n9 0.226933
R112 VGND VGND.n41 0.156997
R113 VGND.n41 VGND.n0 0.150766
R114 VGND.n17 VGND.n9 0.122949
R115 VGND.n18 VGND.n17 0.122949
R116 VGND.n19 VGND.n18 0.122949
R117 VGND.n19 VGND.n7 0.122949
R118 VGND.n24 VGND.n7 0.122949
R119 VGND.n25 VGND.n24 0.122949
R120 VGND.n26 VGND.n25 0.122949
R121 VGND.n26 VGND.n5 0.122949
R122 VGND.n30 VGND.n5 0.122949
R123 VGND.n31 VGND.n30 0.122949
R124 VGND.n32 VGND.n31 0.122949
R125 VGND.n32 VGND.n3 0.122949
R126 VGND.n36 VGND.n3 0.122949
R127 VGND.n37 VGND.n36 0.122949
R128 VGND.n37 VGND.n0 0.122949
R129 VNB.n0 VNB 14851.4
R130 VNB.t10 VNB.t12 4746.46
R131 VNB VNB.n0 2707.69
R132 VNB.t11 VNB.t7 2533.33
R133 VNB.t5 VNB.t4 2496.97
R134 VNB.t1 VNB.t0 2400
R135 VNB.t6 VNB.t5 1648.48
R136 VNB.t12 VNB.t13 1339.63
R137 VNB.t0 VNB 1200
R138 VNB.t2 VNB.t3 1177.95
R139 VNB.t4 VNB.t1 1042.42
R140 VNB.t7 VNB.t6 945.456
R141 VNB.t8 VNB.t10 900.788
R142 VNB.t3 VNB.t8 900.788
R143 VNB.n0 VNB.t11 800
R144 VNB.n0 VNB.t2 219.423
R145 VNB.n0 VNB.t9 65.6721
R146 SET_B.n2 SET_B.t0 346.697
R147 SET_B.n1 SET_B.t1 264.356
R148 SET_B.n1 SET_B.n0 220.054
R149 SET_B SET_B.n2 174.392
R150 SET_B.n2 SET_B.t2 134.617
R151 SET_B SET_B.n1 57.0418
R152 a_1027_118.t0 a_1027_118.t1 60.0005
R153 a_604_74.n5 a_604_74.n4 692.703
R154 a_604_74.n2 a_604_74.t6 309.454
R155 a_604_74.n1 a_604_74.t5 230.919
R156 a_604_74.n6 a_604_74.n5 198.77
R157 a_604_74.n1 a_604_74.n0 192.091
R158 a_604_74.n3 a_604_74.n1 188.073
R159 a_604_74.n2 a_604_74.t4 157.453
R160 a_604_74.n3 a_604_74.n2 152
R161 a_604_74.n5 a_604_74.n3 123.483
R162 a_604_74.t2 a_604_74.n6 111.43
R163 a_604_74.n4 a_604_74.t0 93.81
R164 a_604_74.n4 a_604_74.t1 70.3576
R165 a_604_74.n6 a_604_74.t3 40.0005
R166 a_398_74.t1 a_398_74.n3 976.965
R167 a_398_74.n2 a_398_74.t4 547.314
R168 a_398_74.n0 a_398_74.t0 356.149
R169 a_398_74.n3 a_398_74.n2 337.575
R170 a_398_74.n2 a_398_74.t3 314.274
R171 a_398_74.n1 a_398_74.t2 274.74
R172 a_398_74.n3 a_398_74.n1 195.09
R173 a_398_74.n1 a_398_74.n0 176.316
R174 a_398_74.n0 a_398_74.t5 174.529
R175 a_1500_74.t0 a_1500_74.t1 68.5719
R176 D.n0 D.t1 238.657
R177 D D.n0 161.504
R178 D.n1 D 154.522
R179 D.n3 D.n2 152
R180 D.n1 D.t0 148.417
R181 D.n2 D.n0 40.9705
R182 D.n2 D.n1 40.9705
R183 D.n3 D 10.6672
R184 D D.n3 3.68535
R185 a_27_74.n0 a_27_74.t3 677.63
R186 a_27_74.n1 a_27_74.t1 673.173
R187 a_27_74.n0 a_27_74.t2 347.594
R188 a_27_74.t0 a_27_74.n1 345.539
R189 a_27_74.n1 a_27_74.n0 160.376
R190 a_1422_74.t0 a_1422_74.t1 68.5719
R191 VPWR.n25 VPWR.n9 1464.52
R192 VPWR.n18 VPWR.t7 687.735
R193 VPWR.n12 VPWR.t9 681.726
R194 VPWR.n40 VPWR.t4 676.885
R195 VPWR.n31 VPWR.n6 618.83
R196 VPWR.n38 VPWR.n2 609.824
R197 VPWR.n6 VPWR.t5 239.214
R198 VPWR.n14 VPWR.n13 231.458
R199 VPWR.n9 VPWR.t6 132.673
R200 VPWR.n9 VPWR.t3 117.263
R201 VPWR.n6 VPWR.t2 77.3934
R202 VPWR.n13 VPWR.t8 52.3309
R203 VPWR.n33 VPWR.n32 36.1417
R204 VPWR.n33 VPWR.n3 36.1417
R205 VPWR.n37 VPWR.n3 36.1417
R206 VPWR.n26 VPWR.n7 36.1417
R207 VPWR.n30 VPWR.n7 36.1417
R208 VPWR.n17 VPWR.n16 36.1417
R209 VPWR.n19 VPWR.n10 36.1417
R210 VPWR.n23 VPWR.n10 36.1417
R211 VPWR.n24 VPWR.n23 36.1417
R212 VPWR.n19 VPWR.n18 31.2476
R213 VPWR.n13 VPWR.t10 28.4351
R214 VPWR.n2 VPWR.t1 26.3844
R215 VPWR.n2 VPWR.t0 26.3844
R216 VPWR.n32 VPWR.n31 26.3534
R217 VPWR.n39 VPWR.n38 25.6005
R218 VPWR.n31 VPWR.n30 24.8476
R219 VPWR.n40 VPWR.n39 23.7181
R220 VPWR.n38 VPWR.n37 21.8358
R221 VPWR.n16 VPWR.n12 19.9534
R222 VPWR.n25 VPWR.n24 16.1887
R223 VPWR.n16 VPWR.n15 9.3005
R224 VPWR.n17 VPWR.n11 9.3005
R225 VPWR.n20 VPWR.n19 9.3005
R226 VPWR.n21 VPWR.n10 9.3005
R227 VPWR.n23 VPWR.n22 9.3005
R228 VPWR.n24 VPWR.n8 9.3005
R229 VPWR.n27 VPWR.n26 9.3005
R230 VPWR.n28 VPWR.n7 9.3005
R231 VPWR.n30 VPWR.n29 9.3005
R232 VPWR.n31 VPWR.n5 9.3005
R233 VPWR.n32 VPWR.n4 9.3005
R234 VPWR.n34 VPWR.n33 9.3005
R235 VPWR.n35 VPWR.n3 9.3005
R236 VPWR.n37 VPWR.n36 9.3005
R237 VPWR.n38 VPWR.n1 9.3005
R238 VPWR.n39 VPWR.n0 9.3005
R239 VPWR.n14 VPWR.n12 7.50963
R240 VPWR.n41 VPWR.n40 7.23624
R241 VPWR.n18 VPWR.n17 4.89462
R242 VPWR.n26 VPWR.n25 1.12991
R243 VPWR.n15 VPWR.n14 0.205157
R244 VPWR VPWR.n41 0.157488
R245 VPWR.n41 VPWR.n0 0.150282
R246 VPWR.n15 VPWR.n11 0.122949
R247 VPWR.n20 VPWR.n11 0.122949
R248 VPWR.n21 VPWR.n20 0.122949
R249 VPWR.n22 VPWR.n21 0.122949
R250 VPWR.n22 VPWR.n8 0.122949
R251 VPWR.n27 VPWR.n8 0.122949
R252 VPWR.n28 VPWR.n27 0.122949
R253 VPWR.n29 VPWR.n28 0.122949
R254 VPWR.n29 VPWR.n5 0.122949
R255 VPWR.n5 VPWR.n4 0.122949
R256 VPWR.n34 VPWR.n4 0.122949
R257 VPWR.n35 VPWR.n34 0.122949
R258 VPWR.n36 VPWR.n35 0.122949
R259 VPWR.n36 VPWR.n1 0.122949
R260 VPWR.n1 VPWR.n0 0.122949
R261 a_1902_74.t1 a_1902_74.n1 419.923
R262 a_1902_74.n0 a_1902_74.t3 279.293
R263 a_1902_74.n1 a_1902_74.t0 253.255
R264 a_1902_74.n1 a_1902_74.n0 173.333
R265 a_1902_74.n0 a_1902_74.t2 171.913
R266 a_1457_508.t0 a_1457_508.t1 126.644
R267 a_709_463.t0 a_709_463.t1 126.644
R268 CLK.n0 CLK.t1 261.62
R269 CLK.n0 CLK.t0 178.34
R270 CLK CLK.n0 156.667
R271 Q.n3 Q 591.4
R272 Q.n3 Q.n0 585
R273 Q.n4 Q.n3 585
R274 Q.t0 Q.n1 279.738
R275 Q.n2 Q.t0 246.054
R276 Q.n3 Q.t1 26.3844
R277 Q Q.n4 17.1525
R278 Q Q.n0 14.8485
R279 Q Q.n2 13.0477
R280 Q.n1 Q 9.56372
R281 Q Q.n0 4.0965
R282 Q.n4 Q 1.7925
R283 Q.n2 Q 1.32464
R284 Q.n1 Q 1.32464
C0 VPB Q 0.01354f
C1 D VGND 0.045523f
C2 VPWR SET_B 0.144502f
C3 CLK SET_B 6.57e-20
C4 VPWR VGND 0.123412f
C5 VPB a_1470_48# 0.100267f
C6 CLK VGND 0.035713f
C7 VPWR Q 0.122539f
C8 SET_B VGND 0.110738f
C9 VPWR a_1470_48# 0.073304f
C10 SET_B Q 2.97e-19
C11 VGND Q 0.105495f
C12 SET_B a_1470_48# 0.220182f
C13 VPB D 0.123048f
C14 VGND a_1470_48# 0.175264f
C15 VPB VPWR 0.295302f
C16 D VPWR 0.018907f
C17 VPB CLK 0.035618f
C18 VPB SET_B 0.235994f
C19 D CLK 0.022292f
C20 D SET_B 6.15e-20
C21 VPWR CLK 0.016075f
C22 VPB VGND 0.02579f
C23 Q VNB 0.115862f
C24 VGND VNB 1.30574f
C25 SET_B VNB 0.285238f
C26 CLK VNB 0.10776f
C27 VPWR VNB 0.990004f
C28 D VNB 0.214578f
C29 VPB VNB 2.61385f
C30 a_1470_48# VNB 0.177497f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfsbp_2 VNB VPB VPWR SET_B VGND CLK D Q_N Q
X0 VPWR.t10 a_757_401.t3 a_706_463.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1961 pd=1.425 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_1261_74# a_595_97.t4 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1934 ps=1.43 w=0.64 l=0.15
X2 a_706_463.t0 a_225_74.t2 a_595_97.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X3 VPWR.t5 SET_B.t0 a_757_401.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2543 pd=1.885 as=0.07665 ps=0.785 w=0.42 l=0.15
X4 a_595_97.t0 a_398_74.t2 a_27_74.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X5 VGND.t2 a_1339_74# Q_N.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 Q_N.t0 a_1339_74# VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 VGND.t3 a_1339_74# a_2221_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1469 pd=1.16 as=0.1824 ps=1.85 w=0.64 l=0.15
X8 VPWR.t8 D.t0 a_27_74.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1239 ps=1.43 w=0.42 l=0.15
X9 VGND.t8 D.t1 a_27_74.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X10 a_1258_341# a_595_97.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1998 pd=1.61 as=0.2543 ps=1.885 w=1 l=0.15
X11 a_731_97.t0 a_398_74.t3 a_595_97.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1113 ps=0.95 w=0.42 l=0.15
X12 VPWR.t1 a_1339_74# Q_N.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t10 SET_B.t1 a_1531_118.t0 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.260625 pd=1.505 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 VGND.t9 a_757_401.t4 a_731_97.t1 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_1339_74# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.063 ps=0.72 w=0.42 l=0.15
X16 Q.t1 a_2221_74.t2 VGND.t12 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1469 ps=1.16 w=0.74 l=0.15
X17 VGND.t6 CLK.t0 a_225_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X18 VPWR.t9 a_1501_92.t2 a_1521_508.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 Q_N a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1841 ps=1.505 w=1.12 l=0.15
X20 VPWR.t7 a_2221_74.t3 Q.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_1001_74.t0 a_595_97.t6 a_757_401.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X22 a_1521_508.t0 a_398_74.t4 a_1339_74# VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.22415 ps=1.66 w=0.42 l=0.15
X23 VPWR.t0 a_1339_74# a_1501_92.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1841 pd=1.505 as=0.2544 ps=2.27 w=0.42 l=0.15
X24 a_398_74.t1 a_225_74.t3 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X25 VGND.t11 SET_B.t2 a_1001_74.t1 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1934 pd=1.43 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 VGND.t5 a_2221_74.t4 Q.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 VPWR.t11 CLK.t1 a_225_74.t1 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X28 a_398_74.t0 a_225_74.t4 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 a_595_97.t3 a_225_74.t5 a_27_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1197 ps=1.41 w=0.42 l=0.15
X30 a_757_401.t0 a_595_97.t7 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.1961 ps=1.425 w=0.42 l=0.15
X31 VPWR.t2 a_1339_74# a_2221_74.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2074 pd=1.5 as=0.295 ps=2.59 w=1 l=0.15
X32 a_1453_118.t0 a_225_74.t6 a_1339_74# VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1157 ps=1.06 w=0.42 l=0.15
X33 a_1501_92.t0 a_1339_74# VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1533 pd=1.57 as=0.260625 ps=1.505 w=0.42 l=0.15
R0 a_757_401.n1 a_757_401.n0 792.278
R1 a_757_401.t1 a_757_401.n2 398.233
R2 a_757_401.n2 a_757_401.t4 229.85
R3 a_757_401.n1 a_757_401.t3 203.804
R4 a_757_401.n2 a_757_401.n1 202.081
R5 a_757_401.n0 a_757_401.t2 100.846
R6 a_757_401.n0 a_757_401.t0 70.3576
R7 a_706_463.t0 a_706_463.t1 126.644
R8 VPWR.n22 VPWR.t0 1079.54
R9 VPWR.n28 VPWR.t9 687.735
R10 VPWR.n50 VPWR.t8 677.66
R11 VPWR.n41 VPWR.n6 662.524
R12 VPWR.n48 VPWR.n2 608.274
R13 VPWR.n35 VPWR.n9 606.968
R14 VPWR.n16 VPWR.t2 282.637
R15 VPWR.n15 VPWR.t7 266.248
R16 VPWR.n14 VPWR.t1 258.81
R17 VPWR.n6 VPWR.t3 253.286
R18 VPWR.n9 VPWR.t5 238.132
R19 VPWR.n6 VPWR.t10 110.227
R20 VPWR.n9 VPWR.t4 87.2109
R21 VPWR.n43 VPWR.n42 36.1417
R22 VPWR.n43 VPWR.n3 36.1417
R23 VPWR.n47 VPWR.n3 36.1417
R24 VPWR.n36 VPWR.n7 36.1417
R25 VPWR.n40 VPWR.n7 36.1417
R26 VPWR.n23 VPWR.n12 36.1417
R27 VPWR.n27 VPWR.n12 36.1417
R28 VPWR.n30 VPWR.n29 36.1417
R29 VPWR.n30 VPWR.n10 36.1417
R30 VPWR.n34 VPWR.n10 36.1417
R31 VPWR.n42 VPWR.n41 31.624
R32 VPWR.n17 VPWR.n14 31.624
R33 VPWR.n35 VPWR.n34 30.8711
R34 VPWR.n49 VPWR.n48 28.2358
R35 VPWR.n22 VPWR.n21 27.1064
R36 VPWR.n2 VPWR.t6 26.3844
R37 VPWR.n2 VPWR.t11 26.3844
R38 VPWR.n17 VPWR.n16 25.224
R39 VPWR.n50 VPWR.n49 22.9652
R40 VPWR.n21 VPWR.n14 21.4593
R41 VPWR.n23 VPWR.n22 20.3299
R42 VPWR.n48 VPWR.n47 19.2005
R43 VPWR.n29 VPWR.n28 19.2005
R44 VPWR.n28 VPWR.n27 16.9417
R45 VPWR.n41 VPWR.n40 15.8123
R46 VPWR.n36 VPWR.n35 13.5534
R47 VPWR.n18 VPWR.n17 9.3005
R48 VPWR.n19 VPWR.n14 9.3005
R49 VPWR.n21 VPWR.n20 9.3005
R50 VPWR.n22 VPWR.n13 9.3005
R51 VPWR.n24 VPWR.n23 9.3005
R52 VPWR.n25 VPWR.n12 9.3005
R53 VPWR.n27 VPWR.n26 9.3005
R54 VPWR.n29 VPWR.n11 9.3005
R55 VPWR.n31 VPWR.n30 9.3005
R56 VPWR.n32 VPWR.n10 9.3005
R57 VPWR.n34 VPWR.n33 9.3005
R58 VPWR.n35 VPWR.n8 9.3005
R59 VPWR.n37 VPWR.n36 9.3005
R60 VPWR.n38 VPWR.n7 9.3005
R61 VPWR.n40 VPWR.n39 9.3005
R62 VPWR.n41 VPWR.n5 9.3005
R63 VPWR.n42 VPWR.n4 9.3005
R64 VPWR.n44 VPWR.n43 9.3005
R65 VPWR.n45 VPWR.n3 9.3005
R66 VPWR.n47 VPWR.n46 9.3005
R67 VPWR.n48 VPWR.n1 9.3005
R68 VPWR.n49 VPWR.n0 9.3005
R69 VPWR.n51 VPWR.n50 7.27223
R70 VPWR.n16 VPWR.n15 6.95806
R71 VPWR.n18 VPWR.n15 0.546775
R72 VPWR VPWR.n51 0.157962
R73 VPWR.n51 VPWR.n0 0.149814
R74 VPWR.n19 VPWR.n18 0.122949
R75 VPWR.n20 VPWR.n19 0.122949
R76 VPWR.n20 VPWR.n13 0.122949
R77 VPWR.n24 VPWR.n13 0.122949
R78 VPWR.n25 VPWR.n24 0.122949
R79 VPWR.n26 VPWR.n25 0.122949
R80 VPWR.n26 VPWR.n11 0.122949
R81 VPWR.n31 VPWR.n11 0.122949
R82 VPWR.n32 VPWR.n31 0.122949
R83 VPWR.n33 VPWR.n32 0.122949
R84 VPWR.n33 VPWR.n8 0.122949
R85 VPWR.n37 VPWR.n8 0.122949
R86 VPWR.n38 VPWR.n37 0.122949
R87 VPWR.n39 VPWR.n38 0.122949
R88 VPWR.n39 VPWR.n5 0.122949
R89 VPWR.n5 VPWR.n4 0.122949
R90 VPWR.n44 VPWR.n4 0.122949
R91 VPWR.n45 VPWR.n44 0.122949
R92 VPWR.n46 VPWR.n45 0.122949
R93 VPWR.n46 VPWR.n1 0.122949
R94 VPWR.n1 VPWR.n0 0.122949
R95 VPB.n0 VPB 3439.92
R96 VPB.t12 VPB.t1 784.005
R97 VPB.t9 VPB.t6 517.279
R98 VPB.t2 VPB.t0 513.307
R99 VPB.t1 VPB.t2 503.091
R100 VPB.t0 VPB.t10 500.538
R101 VPB VPB.n1 479.974
R102 VPB.t13 VPB.t3 460.079
R103 VPB.t5 VPB.t4 447.644
R104 VPB.n0 VPB.t7 406.048
R105 VPB.n1 VPB.t14 273.56
R106 VPB.t4 VPB.n0 258.639
R107 VPB.t11 VPB 257.93
R108 VPB.t3 VPB.t5 256.152
R109 VPB.n1 VPB.t11 234.946
R110 VPB.t6 VPB.t8 223.822
R111 VPB.t14 VPB.t9 223.822
R112 VPB.t7 VPB.t12 214.517
R113 VPB.t8 VPB.t13 208.901
R114 a_595_97.n4 a_595_97.n3 674.215
R115 a_595_97.n0 a_595_97.t6 337.401
R116 a_595_97.n2 a_595_97.n1 307.063
R117 a_595_97.n1 a_595_97.t5 301.25
R118 a_595_97.n0 a_595_97.t7 210.742
R119 a_595_97.n5 a_595_97.n4 210.099
R120 a_595_97.n1 a_595_97.t4 158.257
R121 a_595_97.n2 a_595_97.n0 157.797
R122 a_595_97.n5 a_595_97.t3 111.43
R123 a_595_97.n4 a_595_97.n2 110.683
R124 a_595_97.n3 a_595_97.t2 70.3576
R125 a_595_97.n3 a_595_97.t0 70.3576
R126 a_595_97.t1 a_595_97.n5 40.0005
R127 VGND.n4 VGND.t9 258.536
R128 VGND.n56 VGND.t8 254.696
R129 VGND.n11 VGND.t1 233.886
R130 VGND.n25 VGND.n9 185
R131 VGND.n27 VGND.n26 185
R132 VGND.n42 VGND.n41 185
R133 VGND.n40 VGND.n39 185
R134 VGND.n15 VGND.t5 178.799
R135 VGND.n18 VGND.t2 171.77
R136 VGND.n41 VGND.n40 140
R137 VGND.n54 VGND.n2 121.365
R138 VGND.n14 VGND.n13 115.751
R139 VGND.n26 VGND.n25 76.6159
R140 VGND.n25 VGND.t10 48.1983
R141 VGND.n26 VGND.t0 48.1983
R142 VGND.n41 VGND.t11 40.0005
R143 VGND.n13 VGND.t3 39.3755
R144 VGND.n24 VGND.n23 36.1417
R145 VGND.n32 VGND.n31 36.1417
R146 VGND.n33 VGND.n32 36.1417
R147 VGND.n33 VGND.n7 36.1417
R148 VGND.n44 VGND.n43 36.1417
R149 VGND.n49 VGND.n48 36.1417
R150 VGND.n50 VGND.n49 36.1417
R151 VGND.n50 VGND.n1 36.1417
R152 VGND.n13 VGND.t12 35.7861
R153 VGND.n40 VGND.t7 33.438
R154 VGND.n18 VGND.n17 32.0005
R155 VGND.n55 VGND.n54 30.4946
R156 VGND.n56 VGND.n55 30.4946
R157 VGND.n48 VGND.n4 29.3652
R158 VGND.n38 VGND.n7 26.7717
R159 VGND.n43 VGND.n42 25.3495
R160 VGND.n19 VGND.n11 24.4711
R161 VGND.n44 VGND.n4 24.0946
R162 VGND.n17 VGND.n14 22.9652
R163 VGND.n23 VGND.n11 22.9652
R164 VGND.n2 VGND.t4 22.7032
R165 VGND.n2 VGND.t6 22.7032
R166 VGND.n54 VGND.n1 22.2123
R167 VGND.n19 VGND.n18 21.4593
R168 VGND.n31 VGND.n9 16.3508
R169 VGND.n55 VGND.n0 9.3005
R170 VGND.n54 VGND.n53 9.3005
R171 VGND.n52 VGND.n1 9.3005
R172 VGND.n51 VGND.n50 9.3005
R173 VGND.n49 VGND.n3 9.3005
R174 VGND.n48 VGND.n47 9.3005
R175 VGND.n46 VGND.n4 9.3005
R176 VGND.n45 VGND.n44 9.3005
R177 VGND.n43 VGND.n5 9.3005
R178 VGND.n36 VGND.n6 9.3005
R179 VGND.n38 VGND.n37 9.3005
R180 VGND.n35 VGND.n7 9.3005
R181 VGND.n34 VGND.n33 9.3005
R182 VGND.n32 VGND.n8 9.3005
R183 VGND.n31 VGND.n30 9.3005
R184 VGND.n29 VGND.n28 9.3005
R185 VGND.n24 VGND.n10 9.3005
R186 VGND.n23 VGND.n22 9.3005
R187 VGND.n21 VGND.n11 9.3005
R188 VGND.n20 VGND.n19 9.3005
R189 VGND.n17 VGND.n16 9.3005
R190 VGND.n18 VGND.n12 9.3005
R191 VGND.n39 VGND.n6 7.94821
R192 VGND.n57 VGND.n56 7.19894
R193 VGND.n15 VGND.n14 6.74444
R194 VGND.n27 VGND.n24 5.43315
R195 VGND.n28 VGND.n27 4.74752
R196 VGND.n28 VGND.n9 2.28924
R197 VGND.n16 VGND.n15 0.585372
R198 VGND.n42 VGND.n6 0.25148
R199 VGND VGND.n57 0.156997
R200 VGND.n57 VGND.n0 0.150766
R201 VGND.n16 VGND.n12 0.122949
R202 VGND.n20 VGND.n12 0.122949
R203 VGND.n21 VGND.n20 0.122949
R204 VGND.n22 VGND.n21 0.122949
R205 VGND.n22 VGND.n10 0.122949
R206 VGND.n29 VGND.n10 0.122949
R207 VGND.n30 VGND.n29 0.122949
R208 VGND.n30 VGND.n8 0.122949
R209 VGND.n34 VGND.n8 0.122949
R210 VGND.n35 VGND.n34 0.122949
R211 VGND.n37 VGND.n35 0.122949
R212 VGND.n37 VGND.n36 0.122949
R213 VGND.n36 VGND.n5 0.122949
R214 VGND.n45 VGND.n5 0.122949
R215 VGND.n46 VGND.n45 0.122949
R216 VGND.n47 VGND.n46 0.122949
R217 VGND.n47 VGND.n3 0.122949
R218 VGND.n51 VGND.n3 0.122949
R219 VGND.n52 VGND.n51 0.122949
R220 VGND.n53 VGND.n52 0.122949
R221 VGND.n53 VGND.n0 0.122949
R222 VGND.n39 VGND.n38 0.0841601
R223 VNB.n0 VNB 15555.9
R224 VNB VNB.n1 14157.1
R225 VNB.t0 VNB.t2 2471.39
R226 VNB.t8 VNB.t13 2348.25
R227 VNB.t7 VNB.t10 2348.25
R228 VNB.t11 VNB.t5 2336.39
R229 VNB.t14 VNB.t0 2321.26
R230 VNB.t3 VNB.t1 2286.61
R231 VNB.t12 VNB.t14 1801.57
R232 VNB.t4 VNB.t11 1612.94
R233 VNB.n1 VNB.t9 1329.94
R234 VNB.t1 VNB.t16 1316.54
R235 VNB.t9 VNB.n0 1255.37
R236 VNB.t10 VNB 1174.12
R237 VNB.n0 VNB.t12 1050.92
R238 VNB.t5 VNB.t7 1019.95
R239 VNB.t16 VNB.t6 993.177
R240 VNB.t2 VNB.t3 993.177
R241 VNB.n1 VNB.t15 960.648
R242 VNB.t15 VNB.t8 853.909
R243 VNB.t13 VNB.t4 853.909
R244 a_225_74.n1 a_225_74.n0 1206.87
R245 a_225_74.t1 a_225_74.n5 862.136
R246 a_225_74.n2 a_225_74.n1 747.101
R247 a_225_74.n0 a_225_74.t6 623.388
R248 a_225_74.n2 a_225_74.t5 279.56
R249 a_225_74.n3 a_225_74.t3 226.809
R250 a_225_74.n5 a_225_74.n4 209.123
R251 a_225_74.n5 a_225_74.t0 200.375
R252 a_225_74.n3 a_225_74.t4 187.25
R253 a_225_74.n1 a_225_74.t2 182.625
R254 a_225_74.n4 a_225_74.n2 54.7732
R255 a_225_74.n4 a_225_74.n3 21.1793
R256 SET_B.n2 SET_B.t2 377.767
R257 SET_B.n1 SET_B.n0 371.409
R258 SET_B.n1 SET_B.t1 228.732
R259 SET_B.n2 SET_B.t0 174.591
R260 SET_B SET_B.n1 172.885
R261 SET_B SET_B.n2 169.656
R262 a_398_74.t1 a_398_74.n4 951.146
R263 a_398_74.n1 a_398_74.t4 554.239
R264 a_398_74.n2 a_398_74.t0 378.575
R265 a_398_74.n4 a_398_74.n1 319.735
R266 a_398_74.n1 a_398_74.n0 314.274
R267 a_398_74.n3 a_398_74.t3 237.787
R268 a_398_74.n4 a_398_74.n3 225.839
R269 a_398_74.n2 a_398_74.t2 164.149
R270 a_398_74.n3 a_398_74.n2 103.355
R271 a_27_74.n0 a_27_74.t2 679.678
R272 a_27_74.n1 a_27_74.t1 667.524
R273 a_27_74.n0 a_27_74.t3 345.034
R274 a_27_74.t0 a_27_74.n1 316.957
R275 a_27_74.n1 a_27_74.n0 157.465
R276 Q_N Q_N.t2 232.159
R277 Q_N.n1 Q_N.n0 185
R278 Q_N.n2 Q_N.n1 185
R279 Q_N.n1 Q_N.t1 22.7032
R280 Q_N.n1 Q_N.t0 22.7032
R281 Q_N.n2 Q_N 16.0005
R282 Q_N.n0 Q_N 12.062
R283 Q_N.n0 Q_N 6.15435
R284 Q_N Q_N.n2 2.21588
R285 a_2221_74.t1 a_2221_74.n4 245.808
R286 a_2221_74.n1 a_2221_74.t3 240.197
R287 a_2221_74.n3 a_2221_74.n0 240.197
R288 a_2221_74.n4 a_2221_74.n3 188.258
R289 a_2221_74.n1 a_2221_74.t4 181.407
R290 a_2221_74.n2 a_2221_74.t2 179.947
R291 a_2221_74.n4 a_2221_74.t0 149.524
R292 a_2221_74.n2 a_2221_74.n1 61.346
R293 a_2221_74.n3 a_2221_74.n2 4.38232
R294 D.n0 D.t0 239.167
R295 D D.n0 161.504
R296 D.n1 D 154.522
R297 D.n3 D.n2 152
R298 D.n1 D.t1 148.927
R299 D.n2 D.n0 42.021
R300 D.n2 D.n1 42.021
R301 D.n3 D 10.6672
R302 D D.n3 3.68535
R303 a_731_97.t0 a_731_97.t1 60.0005
R304 Q.n0 Q.t2 293.426
R305 Q.n1 Q.n0 185
R306 Q.n2 Q.n1 185
R307 Q.n1 Q.t0 22.7032
R308 Q.n1 Q.t1 22.7032
R309 Q.n2 Q 12.2358
R310 Q.n0 Q 4.70638
R311 Q Q.n2 1.69462
R312 CLK.n0 CLK.t1 272.33
R313 CLK.n0 CLK.t0 178.34
R314 CLK CLK.n0 156.87
R315 a_1501_92.n2 a_1501_92.t1 989.374
R316 a_1501_92.n1 a_1501_92.t2 299.108
R317 a_1501_92.n1 a_1501_92.n0 268.606
R318 a_1501_92.n2 a_1501_92.n1 261.699
R319 a_1501_92.t0 a_1501_92.n2 247.857
R320 a_1521_508.t0 a_1521_508.t1 126.644
R321 a_1001_74.t0 a_1001_74.t1 60.0005
C0 CLK SET_B 6.26e-20
C1 VPWR VGND 0.181418f
C2 a_1339_74# Q 0.002268f
C3 D SET_B 7.37e-20
C4 VPB VGND 0.030612f
C5 VPWR Q_N 0.16233f
C6 CLK VGND 0.037727f
C7 a_1258_341# SET_B 0.00454f
C8 D VGND 0.045364f
C9 VPB Q_N 0.005899f
C10 VPWR Q 0.227139f
C11 SET_B VGND 0.128646f
C12 a_1258_341# VGND 1.17e-19
C13 VPB Q 0.00698f
C14 a_1339_74# a_1261_74# 5.14e-19
C15 SET_B Q_N 8.58e-19
C16 VGND Q_N 0.138113f
C17 SET_B Q 2.14e-19
C18 VGND Q 0.160567f
C19 a_1339_74# VPWR 0.296488f
C20 a_1261_74# SET_B 5.63e-19
C21 a_1339_74# VPB 0.276702f
C22 a_1261_74# VGND 0.001266f
C23 a_1339_74# SET_B 0.20218f
C24 VPB VPWR 0.372482f
C25 a_1339_74# a_1258_341# 0.007436f
C26 VPWR CLK 0.0175f
C27 a_1339_74# VGND 0.092551f
C28 D VPWR 0.019443f
C29 VPB CLK 0.034679f
C30 VPB D 0.120753f
C31 VPWR SET_B 0.113148f
C32 a_1258_341# VPWR 0.009892f
C33 a_1339_74# Q_N 0.078127f
C34 D CLK 0.023743f
C35 VPB SET_B 0.216742f
C36 Q VNB 0.031218f
C37 Q_N VNB 0.009534f
C38 VGND VNB 1.56213f
C39 SET_B VNB 0.293694f
C40 CLK VNB 0.110851f
C41 VPWR VNB 1.19716f
C42 D VNB 0.21434f
C43 VPB VNB 3.02272f
C44 a_1339_74# VNB 0.576289f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfsbp_1 VNB VPB VPWR SET_B VGND Q Q_N D CLK
X0 VGND.t7 a_779_380.t3 a_748_81.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 a_1262_74.t1 a_596_81.t4 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1088 pd=0.98 as=0.129 ps=1.105 w=0.64 l=0.15
X2 VPWR.t7 SET_B.t0 a_779_380.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.222525 pd=1.715 as=0.0756 ps=0.78 w=0.42 l=0.15
X3 Q_N a_1355_377# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1673 ps=1.475 w=1.12 l=0.15
X4 VPWR.t4 D.t0 a_27_80.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1239 ps=1.43 w=0.42 l=0.15
X5 a_596_81.t0 a_398_74.t2 a_27_80.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.1239 ps=1.43 w=0.42 l=0.15
X6 a_1510_48.t1 a_1355_377# VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1491 ps=1.13 w=0.42 l=0.15
X7 Q.t1 a_2113_74.t1 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X8 a_748_81.t0 a_398_74.t3 a_596_81.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_1462_74.t1 a_225_74.t2 a_1355_377# VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.10695 ps=1 w=0.42 l=0.15
X10 VPWR.t2 a_1355_377# a_1510_48.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1673 pd=1.475 as=0.1596 ps=1.6 w=0.42 l=0.15
X11 VPWR.t3 a_1355_377# a_2113_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X12 VGND.t0 CLK.t0 a_225_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 a_1061_74.t0 a_596_81.t5 a_779_380.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1113 ps=1.37 w=0.42 l=0.15
X14 Q.t0 a_2113_74.t2 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X15 a_1254_341.t0 a_596_81.t6 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.19325 pd=1.535 as=0.222525 ps=1.715 w=1 l=0.15
X16 VGND.t1 D.t1 a_27_80.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1197 ps=1.41 w=0.42 l=0.15
X17 a_398_74.t1 a_225_74.t3 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VPWR.t5 CLK.t1 a_225_74.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X19 a_398_74.t0 a_225_74.t4 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_1355_377# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X21 VPWR.t8 a_779_380.t4 a_728_463.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15855 pd=1.175 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 VPWR.t6 a_1510_48.t2 a_1517_508.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_1355_377# a_398_74.t4 a_1262_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.10695 pd=1 as=0.1088 ps=0.98 w=0.64 l=0.15
X24 a_779_380.t0 a_596_81.t7 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.0756 pd=0.78 as=0.15855 ps=1.175 w=0.42 l=0.15
X25 VGND.t6 SET_B.t1 a_1540_74.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1491 pd=1.13 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 Q_N.t0 a_1355_377# VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X27 a_728_463.t0 a_225_74.t5 a_596_81.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0735 ps=0.77 w=0.42 l=0.15
X28 a_1517_508.t0 a_398_74.t5 a_1355_377# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.2204 ps=1.735 w=0.42 l=0.15
X29 a_596_81.t2 a_225_74.t6 a_27_80.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1281 pd=1.03 as=0.1197 ps=1.41 w=0.42 l=0.15
X30 a_1540_74.t0 a_1510_48.t3 a_1462_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_779_380.n1 a_779_380.n0 801.548
R1 a_779_380.t1 a_779_380.n2 394.844
R2 a_779_380.n1 a_779_380.t4 236.448
R3 a_779_380.n2 a_779_380.t3 230.046
R4 a_779_380.n2 a_779_380.n1 183.452
R5 a_779_380.n0 a_779_380.t2 98.5005
R6 a_779_380.n0 a_779_380.t0 70.3576
R7 a_748_81.t0 a_748_81.t1 68.5719
R8 VGND.n44 VGND.t1 256.233
R9 VGND.n31 VGND.t7 246.333
R10 VGND.n10 VGND.t4 240.387
R11 VGND.n18 VGND.n17 185
R12 VGND.n16 VGND.n15 185
R13 VGND.n11 VGND.t8 156.681
R14 VGND.n6 VGND.t2 139.144
R15 VGND.n42 VGND.n2 121.365
R16 VGND.n17 VGND.n16 102.858
R17 VGND.n16 VGND.t3 60.0005
R18 VGND.n17 VGND.t6 40.0005
R19 VGND.n14 VGND.n13 36.1417
R20 VGND.n23 VGND.n8 36.1417
R21 VGND.n24 VGND.n23 36.1417
R22 VGND.n25 VGND.n24 36.1417
R23 VGND.n30 VGND.n29 36.1417
R24 VGND.n32 VGND.n30 36.1417
R25 VGND.n36 VGND.n4 36.1417
R26 VGND.n37 VGND.n36 36.1417
R27 VGND.n38 VGND.n37 36.1417
R28 VGND.n38 VGND.n1 36.1417
R29 VGND.n43 VGND.n42 30.4946
R30 VGND.n44 VGND.n43 30.4946
R31 VGND.n29 VGND.n6 25.224
R32 VGND.n2 VGND.t5 22.7032
R33 VGND.n2 VGND.t0 22.7032
R34 VGND.n25 VGND.n6 22.2123
R35 VGND.n42 VGND.n1 22.2123
R36 VGND.n18 VGND.n8 13.7155
R37 VGND.n15 VGND.n14 12.2096
R38 VGND.n11 VGND.n10 9.47227
R39 VGND.n13 VGND.n10 9.41227
R40 VGND.n32 VGND.n31 9.41227
R41 VGND.n43 VGND.n0 9.3005
R42 VGND.n42 VGND.n41 9.3005
R43 VGND.n13 VGND.n12 9.3005
R44 VGND.n14 VGND.n9 9.3005
R45 VGND.n20 VGND.n19 9.3005
R46 VGND.n21 VGND.n8 9.3005
R47 VGND.n23 VGND.n22 9.3005
R48 VGND.n24 VGND.n7 9.3005
R49 VGND.n26 VGND.n25 9.3005
R50 VGND.n27 VGND.n6 9.3005
R51 VGND.n29 VGND.n28 9.3005
R52 VGND.n30 VGND.n5 9.3005
R53 VGND.n33 VGND.n32 9.3005
R54 VGND.n34 VGND.n4 9.3005
R55 VGND.n36 VGND.n35 9.3005
R56 VGND.n37 VGND.n3 9.3005
R57 VGND.n39 VGND.n38 9.3005
R58 VGND.n40 VGND.n1 9.3005
R59 VGND.n45 VGND.n44 7.19894
R60 VGND.n19 VGND.n15 3.22169
R61 VGND.n19 VGND.n18 2.88262
R62 VGND.n31 VGND.n4 1.88285
R63 VGND.n12 VGND.n11 0.20927
R64 VGND VGND.n45 0.156997
R65 VGND.n45 VGND.n0 0.150766
R66 VGND.n12 VGND.n9 0.122949
R67 VGND.n20 VGND.n9 0.122949
R68 VGND.n21 VGND.n20 0.122949
R69 VGND.n22 VGND.n21 0.122949
R70 VGND.n22 VGND.n7 0.122949
R71 VGND.n26 VGND.n7 0.122949
R72 VGND.n27 VGND.n26 0.122949
R73 VGND.n28 VGND.n27 0.122949
R74 VGND.n28 VGND.n5 0.122949
R75 VGND.n33 VGND.n5 0.122949
R76 VGND.n34 VGND.n33 0.122949
R77 VGND.n35 VGND.n34 0.122949
R78 VGND.n35 VGND.n3 0.122949
R79 VGND.n39 VGND.n3 0.122949
R80 VGND.n40 VGND.n39 0.122949
R81 VGND.n41 VGND.n40 0.122949
R82 VGND.n41 VGND.n0 0.122949
R83 VNB.n0 VNB 15509.7
R84 VNB VNB.n1 14107.3
R85 VNB.t7 VNB.t13 3626.25
R86 VNB.t3 VNB.t12 2787.06
R87 VNB.t8 VNB.t7 2448.29
R88 VNB.t9 VNB.t10 2348.25
R89 VNB.t0 VNB.t1 2348.25
R90 VNB.t11 VNB.t8 1986.35
R91 VNB.t4 VNB.t9 1802.7
R92 VNB.n1 VNB.t2 1392.09
R93 VNB.t2 VNB.n0 1193.22
R94 VNB.t5 VNB.t14 1177.95
R95 VNB.t1 VNB 1174.12
R96 VNB.n1 VNB.t3 1055.53
R97 VNB.t10 VNB.t0 1019.95
R98 VNB.t12 VNB.t4 925.067
R99 VNB.t6 VNB.t11 900.788
R100 VNB.t14 VNB.t6 900.788
R101 VNB.n0 VNB.t5 11.9733
R102 a_596_81.n4 a_596_81.n3 690.539
R103 a_596_81.n1 a_596_81.t7 336.774
R104 a_596_81.n0 a_596_81.t6 254.175
R105 a_596_81.n2 a_596_81.n0 211.78
R106 a_596_81.n5 a_596_81.n4 203.177
R107 a_596_81.n1 a_596_81.t5 175.036
R108 a_596_81.n0 a_596_81.t4 159.381
R109 a_596_81.n2 a_596_81.n1 152
R110 a_596_81.n4 a_596_81.n2 142.603
R111 a_596_81.n5 a_596_81.t2 134.286
R112 a_596_81.n3 a_596_81.t0 93.81
R113 a_596_81.n3 a_596_81.t3 70.3576
R114 a_596_81.t1 a_596_81.n5 40.0005
R115 a_1262_74.t0 a_1262_74.t1 63.7505
R116 SET_B.n1 SET_B.n0 387.474
R117 SET_B.n3 SET_B.n2 356.452
R118 SET_B.n1 SET_B.t1 324.839
R119 SET_B.n3 SET_B.t0 188.554
R120 SET_B SET_B.n1 170.489
R121 SET_B SET_B.n3 169.242
R122 VPWR.n15 VPWR.t2 690.609
R123 VPWR.n21 VPWR.t6 687.735
R124 VPWR.n43 VPWR.t4 677.66
R125 VPWR.n28 VPWR.n9 611.354
R126 VPWR.n41 VPWR.n2 609.63
R127 VPWR.n34 VPWR.n6 608.981
R128 VPWR.n14 VPWR.n13 327.83
R129 VPWR.n6 VPWR.t1 269.702
R130 VPWR.n9 VPWR.t7 174.451
R131 VPWR.n9 VPWR.t0 99.8391
R132 VPWR.n6 VPWR.t8 84.4291
R133 VPWR.n13 VPWR.t9 42.7085
R134 VPWR.n36 VPWR.n35 36.1417
R135 VPWR.n36 VPWR.n3 36.1417
R136 VPWR.n40 VPWR.n3 36.1417
R137 VPWR.n29 VPWR.n7 36.1417
R138 VPWR.n33 VPWR.n7 36.1417
R139 VPWR.n16 VPWR.n12 36.1417
R140 VPWR.n20 VPWR.n12 36.1417
R141 VPWR.n23 VPWR.n22 36.1417
R142 VPWR.n23 VPWR.n10 36.1417
R143 VPWR.n27 VPWR.n10 36.1417
R144 VPWR.n13 VPWR.t3 35.1791
R145 VPWR.n35 VPWR.n34 33.5064
R146 VPWR.n28 VPWR.n27 32.377
R147 VPWR.n42 VPWR.n41 28.2358
R148 VPWR.n2 VPWR.t10 26.3844
R149 VPWR.n2 VPWR.t5 26.3844
R150 VPWR.n43 VPWR.n42 22.9652
R151 VPWR.n41 VPWR.n40 19.2005
R152 VPWR.n21 VPWR.n20 18.4476
R153 VPWR.n22 VPWR.n21 17.6946
R154 VPWR.n16 VPWR.n15 15.0593
R155 VPWR.n29 VPWR.n28 14.3064
R156 VPWR.n17 VPWR.n16 9.3005
R157 VPWR.n18 VPWR.n12 9.3005
R158 VPWR.n20 VPWR.n19 9.3005
R159 VPWR.n22 VPWR.n11 9.3005
R160 VPWR.n24 VPWR.n23 9.3005
R161 VPWR.n25 VPWR.n10 9.3005
R162 VPWR.n27 VPWR.n26 9.3005
R163 VPWR.n28 VPWR.n8 9.3005
R164 VPWR.n30 VPWR.n29 9.3005
R165 VPWR.n31 VPWR.n7 9.3005
R166 VPWR.n33 VPWR.n32 9.3005
R167 VPWR.n34 VPWR.n5 9.3005
R168 VPWR.n35 VPWR.n4 9.3005
R169 VPWR.n37 VPWR.n36 9.3005
R170 VPWR.n38 VPWR.n3 9.3005
R171 VPWR.n40 VPWR.n39 9.3005
R172 VPWR.n41 VPWR.n1 9.3005
R173 VPWR.n42 VPWR.n0 9.3005
R174 VPWR.n34 VPWR.n33 9.03579
R175 VPWR.n15 VPWR.n14 7.40095
R176 VPWR.n44 VPWR.n43 7.27223
R177 VPWR.n17 VPWR.n14 0.219551
R178 VPWR VPWR.n44 0.157962
R179 VPWR.n44 VPWR.n0 0.149814
R180 VPWR.n18 VPWR.n17 0.122949
R181 VPWR.n19 VPWR.n18 0.122949
R182 VPWR.n19 VPWR.n11 0.122949
R183 VPWR.n24 VPWR.n11 0.122949
R184 VPWR.n25 VPWR.n24 0.122949
R185 VPWR.n26 VPWR.n25 0.122949
R186 VPWR.n26 VPWR.n8 0.122949
R187 VPWR.n30 VPWR.n8 0.122949
R188 VPWR.n31 VPWR.n30 0.122949
R189 VPWR.n32 VPWR.n31 0.122949
R190 VPWR.n32 VPWR.n5 0.122949
R191 VPWR.n5 VPWR.n4 0.122949
R192 VPWR.n37 VPWR.n4 0.122949
R193 VPWR.n38 VPWR.n37 0.122949
R194 VPWR.n39 VPWR.n38 0.122949
R195 VPWR.n39 VPWR.n1 0.122949
R196 VPWR.n1 VPWR.n0 0.122949
R197 VPB.n0 VPB 3429.7
R198 VPB.t8 VPB.t4 789.114
R199 VPB.t4 VPB.t3 773.79
R200 VPB.t13 VPB.t0 547.12
R201 VPB VPB.n1 479.974
R202 VPB.t11 VPB.t1 450.132
R203 VPB.n0 VPB.t5 406.048
R204 VPB.t9 VPB.t2 395.42
R205 VPB.n1 VPB.t7 273.56
R206 VPB.t2 VPB.n0 258.639
R207 VPB.t3 VPB.t12 257.93
R208 VPB.t6 VPB 257.93
R209 VPB.t1 VPB.t9 253.666
R210 VPB.t0 VPB.t10 248.691
R211 VPB.n1 VPB.t6 234.946
R212 VPB.t7 VPB.t13 223.822
R213 VPB.t5 VPB.t8 214.517
R214 VPB.t10 VPB.t11 208.901
R215 Q_N.n1 Q_N.n0 1208.67
R216 Q_N Q_N.t0 155.002
R217 Q_N Q_N.n1 13.6132
R218 Q_N Q_N.n0 7.96062
R219 Q_N.n0 Q_N 6.98145
R220 Q_N.n1 Q_N 1.42272
R221 D.n0 D.t0 231.133
R222 D D.n0 162.667
R223 D.n1 D 153.358
R224 D.n3 D.n2 152
R225 D.n1 D.t1 148.927
R226 D.n2 D.n0 42.021
R227 D.n2 D.n1 42.021
R228 D.n3 D 11.8308
R229 D D.n3 2.52171
R230 a_27_80.n0 a_27_80.t2 679.678
R231 a_27_80.n1 a_27_80.t0 666.942
R232 a_27_80.n0 a_27_80.t3 342.776
R233 a_27_80.t1 a_27_80.n1 322.882
R234 a_27_80.n1 a_27_80.n0 163.489
R235 a_398_74.t1 a_398_74.n3 905.835
R236 a_398_74.n0 a_398_74.t5 551.582
R237 a_398_74.n1 a_398_74.t0 366.618
R238 a_398_74.n3 a_398_74.n0 325.5
R239 a_398_74.n0 a_398_74.t4 314.274
R240 a_398_74.n2 a_398_74.t3 239.393
R241 a_398_74.n3 a_398_74.n2 214.036
R242 a_398_74.n1 a_398_74.t2 174.192
R243 a_398_74.n2 a_398_74.n1 112.037
R244 a_1510_48.n1 a_1510_48.t0 863.635
R245 a_1510_48.n0 a_1510_48.t3 382.68
R246 a_1510_48.n0 a_1510_48.t2 262.959
R247 a_1510_48.n1 a_1510_48.n0 246.119
R248 a_1510_48.t1 a_1510_48.n1 238.382
R249 a_2113_74.t0 a_2113_74.n0 617.74
R250 a_2113_74.n0 a_2113_74.t2 285.719
R251 a_2113_74.n0 a_2113_74.t1 178.34
R252 Q.n1 Q 589.85
R253 Q.n1 Q.n0 585
R254 Q.n2 Q.n1 585
R255 Q Q.t1 203.387
R256 Q.n1 Q.t0 26.3844
R257 Q Q.n2 12.9944
R258 Q Q.n0 11.249
R259 Q Q.n0 3.10353
R260 Q.n2 Q 1.35808
R261 a_225_74.n1 a_225_74.n0 1185.18
R262 a_225_74.t1 a_225_74.n5 862.136
R263 a_225_74.n2 a_225_74.n1 782.447
R264 a_225_74.n0 a_225_74.t2 703.721
R265 a_225_74.n2 a_225_74.t6 306.873
R266 a_225_74.n3 a_225_74.t3 226.809
R267 a_225_74.n5 a_225_74.n4 215.147
R268 a_225_74.n5 a_225_74.t0 201.371
R269 a_225_74.n3 a_225_74.t4 188.728
R270 a_225_74.n1 a_225_74.t5 182.625
R271 a_225_74.n4 a_225_74.n2 43.0884
R272 a_225_74.n4 a_225_74.n3 32.8641
R273 a_1462_74.t0 a_1462_74.t1 68.5719
R274 CLK.n0 CLK.t1 272.33
R275 CLK.n0 CLK.t0 178.34
R276 CLK CLK.n0 156.667
R277 a_1254_341.n0 a_1254_341.t0 49.9442
R278 a_728_463.t0 a_728_463.t1 126.644
R279 a_1517_508.t0 a_1517_508.t1 126.644
R280 a_1540_74.t0 a_1540_74.t1 68.5719
C0 VPB VPWR 0.319901f
C1 SET_B Q 6.16e-20
C2 VGND a_1355_377# 0.064294f
C3 VPB CLK 0.034761f
C4 D VPWR 0.018852f
C5 Q_N a_1355_377# 0.067498f
C6 D CLK 0.023171f
C7 Q a_1355_377# 0.004685f
C8 VGND VPB 0.025985f
C9 SET_B a_1355_377# 0.191264f
C10 VPWR CLK 0.017323f
C11 VGND D 0.044811f
C12 Q_N VPB 0.014147f
C13 VGND VPWR 0.142591f
C14 Q VPB 0.014139f
C15 SET_B VPB 0.206662f
C16 VGND CLK 0.039539f
C17 Q_N VPWR 0.065567f
C18 SET_B D 7.37e-20
C19 Q VPWR 0.119134f
C20 SET_B VPWR 0.106724f
C21 a_1355_377# VPB 0.328083f
C22 VGND Q_N 0.069964f
C23 SET_B CLK 6.26e-20
C24 VGND Q 0.087399f
C25 a_1355_377# VPWR 0.264848f
C26 SET_B VGND 0.128283f
C27 VPB D 0.1214f
C28 SET_B Q_N 3.82e-19
C29 Q VNB 0.110954f
C30 Q_N VNB 0.015214f
C31 VGND VNB 1.40416f
C32 SET_B VNB 0.304227f
C33 CLK VNB 0.11198f
C34 VPWR VNB 1.07921f
C35 D VNB 0.20988f
C36 VPB VNB 2.80832f
C37 a_1355_377# VNB 0.528644f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfrtp_4 VNB VPB VPWR RESET_B VGND D CLK Q
X0 VPWR.t0 CLK.t0 a_313_74.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3248 ps=2.82 w=1.12 l=0.15
X1 VGND.t5 RESET_B.t0 a_124_78.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 a_494_366.t0 a_313_74.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X3 a_37_78.t3 D.t0 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X4 a_834_355.t0 a_699_463.t5 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.47175 pd=2.015 as=0.30625 ps=1.74 w=0.74 l=0.15
X5 VPWR.t10 a_2010_409.t3 Q.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.434 pd=1.895 as=0.1932 ps=1.465 w=1.12 l=0.15
X6 VPWR.t12 a_1350_392.t2 a_1678_395.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.195 as=0.063 ps=0.72 w=0.42 l=0.15
X7 VGND.t1 CLK.t1 a_313_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VGND.t4 RESET_B.t1 a_890_138.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.30625 pd=1.74 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 a_699_463.t2 RESET_B.t2 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1295 ps=1.115 w=0.42 l=0.15
X10 a_1827_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X11 a_1350_392.t0 a_313_74.t3 a_834_355.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3362 pd=2.235 as=0.15 ps=1.3 w=1 l=0.15
X12 a_890_138.t1 a_834_355.t4 a_812_138.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X13 a_834_355.t1 a_699_463.t6 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2845 ps=2.68 w=1 l=0.15
X14 a_812_138.t1 a_494_366.t2 a_699_463.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X15 Q.t2 a_2010_409.t4 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.13875 pd=1.115 as=0.2109 ps=2.05 w=0.74 l=0.15
X16 VGND.t7 a_2010_409.t5 Q.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VPWR.t13 a_1350_392.t3 a_2010_409.t2 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.126 ps=1.14 w=0.84 l=0.15
X18 Q.t5 a_2010_409.t6 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.1862 ps=1.475 w=1.12 l=0.15
X19 VGND.t8 a_2010_409.t7 Q.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.13875 ps=1.115 w=0.74 l=0.15
X20 VGND.t0 a_1678_395.t2 a_1647_81.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X21 VPWR.t3 RESET_B.t3 a_37_78.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X22 VPWR.t5 a_834_355.t5 a_789_463.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1295 pd=1.115 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 a_1678_395.t1 a_1350_392.t4 a_1827_81# VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X24 a_1350_392.t1 a_494_366.t3 a_834_355.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.47175 ps=2.015 w=0.74 l=0.15
X25 a_124_78.t1 D.t1 a_37_78.t4 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X26 a_699_463.t0 a_313_74.t4 a_37_78.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X27 a_789_463.t0 a_313_74.t5 a_699_463.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X28 a_2010_409.t0 a_1350_392.t5 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1302 ps=1.195 w=0.84 l=0.15
X29 VPWR.t7 a_2010_409.t8 Q.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_699_463.t3 a_494_366.t4 a_37_78.t2 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X31 Q.t3 a_2010_409.t9 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.434 ps=1.895 w=1.12 l=0.15
X32 a_494_366.t1 a_313_74.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X33 a_2010_409.t1 a_1350_392.t6 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
R0 CLK.n0 CLK.t0 258.942
R1 CLK.n0 CLK.t1 207.261
R2 CLK CLK.n0 157.625
R3 a_313_74.n2 a_313_74.n1 1169.7
R4 a_313_74.t1 a_313_74.n6 926.933
R5 a_313_74.n3 a_313_74.n2 767.987
R6 a_313_74.n1 a_313_74.n0 740.673
R7 a_313_74.n4 a_313_74.t4 408.094
R8 a_313_74.n1 a_313_74.t3 239.996
R9 a_313_74.n3 a_313_74.t6 216.671
R10 a_313_74.n6 a_313_74.n5 213.284
R11 a_313_74.n2 a_313_74.t5 182.625
R12 a_313_74.n4 a_313_74.t2 154.24
R13 a_313_74.n6 a_313_74.t0 145.959
R14 a_313_74.n5 a_313_74.n3 32.1338
R15 a_313_74.n5 a_313_74.n4 4.01717
R16 VPWR.n8 VPWR.t2 879.162
R17 VPWR.n53 VPWR.t9 685.053
R18 VPWR.n51 VPWR.t3 681.726
R19 VPWR.n40 VPWR.n7 667.909
R20 VPWR.n13 VPWR.n12 618.537
R21 VPWR.n3 VPWR.n2 606.139
R22 VPWR.n21 VPWR.n15 320.625
R23 VPWR.n18 VPWR.t7 264.014
R24 VPWR.n17 VPWR.n16 139.94
R25 VPWR.n7 VPWR.t11 107.882
R26 VPWR.n7 VPWR.t5 107.882
R27 VPWR.n12 VPWR.t12 89.1195
R28 VPWR.n16 VPWR.t10 63.1443
R29 VPWR.n16 VPWR.t8 63.1439
R30 VPWR.n15 VPWR.t13 46.9053
R31 VPWR.n12 VPWR.t4 45.7326
R32 VPWR.n44 VPWR.n5 36.1417
R33 VPWR.n45 VPWR.n44 36.1417
R34 VPWR.n46 VPWR.n45 36.1417
R35 VPWR.n39 VPWR.n38 36.1417
R36 VPWR.n28 VPWR.n10 36.1417
R37 VPWR.n32 VPWR.n10 36.1417
R38 VPWR.n33 VPWR.n32 36.1417
R39 VPWR.n34 VPWR.n33 36.1417
R40 VPWR.n27 VPWR.n26 33.8829
R41 VPWR.n22 VPWR.n13 31.624
R42 VPWR.n21 VPWR.n20 31.2476
R43 VPWR.n15 VPWR.t6 30.9049
R44 VPWR.n52 VPWR.n51 27.8593
R45 VPWR.n53 VPWR.n52 27.1064
R46 VPWR.n2 VPWR.t1 26.3844
R47 VPWR.n2 VPWR.t0 26.3844
R48 VPWR.n51 VPWR.n50 25.6005
R49 VPWR.n50 VPWR.n3 24.4711
R50 VPWR.n40 VPWR.n5 24.0946
R51 VPWR.n34 VPWR.n8 23.7181
R52 VPWR.n38 VPWR.n8 23.3417
R53 VPWR.n40 VPWR.n39 23.3417
R54 VPWR.n46 VPWR.n3 22.9652
R55 VPWR.n26 VPWR.n13 21.8358
R56 VPWR.n20 VPWR.n17 19.2005
R57 VPWR.n22 VPWR.n21 16.1887
R58 VPWR.n28 VPWR.n27 13.5534
R59 VPWR.n20 VPWR.n19 9.3005
R60 VPWR.n21 VPWR.n14 9.3005
R61 VPWR.n23 VPWR.n22 9.3005
R62 VPWR.n24 VPWR.n13 9.3005
R63 VPWR.n26 VPWR.n25 9.3005
R64 VPWR.n27 VPWR.n11 9.3005
R65 VPWR.n29 VPWR.n28 9.3005
R66 VPWR.n30 VPWR.n10 9.3005
R67 VPWR.n32 VPWR.n31 9.3005
R68 VPWR.n33 VPWR.n9 9.3005
R69 VPWR.n35 VPWR.n34 9.3005
R70 VPWR.n36 VPWR.n8 9.3005
R71 VPWR.n38 VPWR.n37 9.3005
R72 VPWR.n39 VPWR.n6 9.3005
R73 VPWR.n41 VPWR.n40 9.3005
R74 VPWR.n42 VPWR.n5 9.3005
R75 VPWR.n44 VPWR.n43 9.3005
R76 VPWR.n45 VPWR.n4 9.3005
R77 VPWR.n47 VPWR.n46 9.3005
R78 VPWR.n48 VPWR.n3 9.3005
R79 VPWR.n50 VPWR.n49 9.3005
R80 VPWR.n51 VPWR.n1 9.3005
R81 VPWR.n52 VPWR.n0 9.3005
R82 VPWR.n54 VPWR.n53 9.3005
R83 VPWR.n18 VPWR.n17 3.89738
R84 VPWR.n19 VPWR.n18 0.459696
R85 VPWR.n19 VPWR.n14 0.122949
R86 VPWR.n23 VPWR.n14 0.122949
R87 VPWR.n24 VPWR.n23 0.122949
R88 VPWR.n25 VPWR.n24 0.122949
R89 VPWR.n25 VPWR.n11 0.122949
R90 VPWR.n29 VPWR.n11 0.122949
R91 VPWR.n30 VPWR.n29 0.122949
R92 VPWR.n31 VPWR.n30 0.122949
R93 VPWR.n31 VPWR.n9 0.122949
R94 VPWR.n35 VPWR.n9 0.122949
R95 VPWR.n36 VPWR.n35 0.122949
R96 VPWR.n37 VPWR.n36 0.122949
R97 VPWR.n37 VPWR.n6 0.122949
R98 VPWR.n41 VPWR.n6 0.122949
R99 VPWR.n42 VPWR.n41 0.122949
R100 VPWR.n43 VPWR.n42 0.122949
R101 VPWR.n43 VPWR.n4 0.122949
R102 VPWR.n47 VPWR.n4 0.122949
R103 VPWR.n48 VPWR.n47 0.122949
R104 VPWR.n49 VPWR.n48 0.122949
R105 VPWR.n49 VPWR.n1 0.122949
R106 VPWR.n1 VPWR.n0 0.122949
R107 VPWR.n54 VPWR.n0 0.122949
R108 VPWR VPWR.n54 0.0617245
R109 VPB.t3 VPB.t15 1427.55
R110 VPB.t14 VPB.t4 692.071
R111 VPB.t1 VPB.t12 523.521
R112 VPB.t5 VPB.t0 508.2
R113 VPB.t13 VPB.t10 472.447
R114 VPB.t7 VPB.t14 311.56
R115 VPB.t16 VPB.t8 257.93
R116 VPB.t15 VPB.t6 257.93
R117 VPB VPB.t11 255.376
R118 VPB.t8 VPB.t13 252.823
R119 VPB.t0 VPB.t1 229.839
R120 VPB.t10 VPB.t9 229.839
R121 VPB.t6 VPB.t16 229.839
R122 VPB.t4 VPB.t3 229.839
R123 VPB.t12 VPB.t2 229.839
R124 VPB.t11 VPB.t5 229.839
R125 VPB.t2 VPB.t7 199.195
R126 RESET_B.n2 RESET_B.n1 451.474
R127 RESET_B.n3 RESET_B.t1 226.005
R128 RESET_B.n5 RESET_B.t3 222.395
R129 RESET_B.n4 RESET_B.n3 222.292
R130 RESET_B.n5 RESET_B.t0 219.93
R131 RESET_B.n4 RESET_B.n2 167.625
R132 RESET_B.n3 RESET_B.t2 158.038
R133 RESET_B.n2 RESET_B.n0 146.475
R134 RESET_B.n6 RESET_B.n5 58.5071
R135 RESET_B.n6 RESET_B.n4 3.75632
R136 RESET_B RESET_B.n6 0.0466957
R137 a_124_78.t0 a_124_78.t1 68.5719
R138 VGND.n13 VGND.t8 277.875
R139 VGND.n0 VGND.t5 263.776
R140 VGND.n24 VGND.t0 255.998
R141 VGND.n37 VGND.n36 220.173
R142 VGND.n48 VGND.n3 207.304
R143 VGND.n14 VGND.t7 169.036
R144 VGND.n17 VGND.t9 166.2
R145 VGND.n11 VGND.t6 159.535
R146 VGND.n36 VGND.t3 89.1897
R147 VGND.n36 VGND.t4 44.9426
R148 VGND.n52 VGND.n0 40.0803
R149 VGND.n23 VGND.n22 36.1417
R150 VGND.n28 VGND.n9 36.1417
R151 VGND.n29 VGND.n28 36.1417
R152 VGND.n30 VGND.n29 36.1417
R153 VGND.n30 VGND.n7 36.1417
R154 VGND.n34 VGND.n7 36.1417
R155 VGND.n35 VGND.n34 36.1417
R156 VGND.n42 VGND.n5 36.1417
R157 VGND.n43 VGND.n42 36.1417
R158 VGND.n44 VGND.n43 36.1417
R159 VGND.n44 VGND.n2 36.1417
R160 VGND.n50 VGND.n49 36.1417
R161 VGND.n3 VGND.t2 34.0546
R162 VGND.n3 VGND.t1 34.0546
R163 VGND.n18 VGND.n11 30.8711
R164 VGND.n24 VGND.n23 30.4946
R165 VGND.n38 VGND.n5 29.3032
R166 VGND.n49 VGND.n48 27.4829
R167 VGND.n37 VGND.n35 26.854
R168 VGND.n17 VGND.n16 26.3534
R169 VGND.n16 VGND.n13 24.0946
R170 VGND.n18 VGND.n17 24.0946
R171 VGND.n22 VGND.n11 20.7064
R172 VGND.n48 VGND.n2 19.9534
R173 VGND.n24 VGND.n9 16.9417
R174 VGND.n51 VGND.n50 9.3005
R175 VGND.n49 VGND.n1 9.3005
R176 VGND.n48 VGND.n47 9.3005
R177 VGND.n46 VGND.n2 9.3005
R178 VGND.n45 VGND.n44 9.3005
R179 VGND.n43 VGND.n4 9.3005
R180 VGND.n42 VGND.n41 9.3005
R181 VGND.n40 VGND.n5 9.3005
R182 VGND.n39 VGND.n38 9.3005
R183 VGND.n35 VGND.n6 9.3005
R184 VGND.n34 VGND.n33 9.3005
R185 VGND.n32 VGND.n7 9.3005
R186 VGND.n31 VGND.n30 9.3005
R187 VGND.n29 VGND.n8 9.3005
R188 VGND.n28 VGND.n27 9.3005
R189 VGND.n26 VGND.n9 9.3005
R190 VGND.n25 VGND.n24 9.3005
R191 VGND.n23 VGND.n10 9.3005
R192 VGND.n22 VGND.n21 9.3005
R193 VGND.n16 VGND.n15 9.3005
R194 VGND.n17 VGND.n12 9.3005
R195 VGND.n19 VGND.n18 9.3005
R196 VGND.n20 VGND.n11 9.3005
R197 VGND.n14 VGND.n13 6.62245
R198 VGND.n50 VGND.n0 3.76521
R199 VGND.n15 VGND.n14 0.655242
R200 VGND.n38 VGND.n37 0.563137
R201 VGND VGND.n52 0.163644
R202 VGND.n52 VGND.n51 0.144205
R203 VGND.n15 VGND.n12 0.122949
R204 VGND.n19 VGND.n12 0.122949
R205 VGND.n20 VGND.n19 0.122949
R206 VGND.n21 VGND.n20 0.122949
R207 VGND.n21 VGND.n10 0.122949
R208 VGND.n25 VGND.n10 0.122949
R209 VGND.n26 VGND.n25 0.122949
R210 VGND.n27 VGND.n26 0.122949
R211 VGND.n27 VGND.n8 0.122949
R212 VGND.n31 VGND.n8 0.122949
R213 VGND.n32 VGND.n31 0.122949
R214 VGND.n33 VGND.n32 0.122949
R215 VGND.n33 VGND.n6 0.122949
R216 VGND.n39 VGND.n6 0.122949
R217 VGND.n40 VGND.n39 0.122949
R218 VGND.n41 VGND.n40 0.122949
R219 VGND.n41 VGND.n4 0.122949
R220 VGND.n45 VGND.n4 0.122949
R221 VGND.n46 VGND.n45 0.122949
R222 VGND.n47 VGND.n46 0.122949
R223 VGND.n47 VGND.n1 0.122949
R224 VGND.n51 VGND.n1 0.122949
R225 VNB VNB.n0 6779
R226 VNB.t13 VNB.t0 3325.98
R227 VNB.t4 VNB.t13 3291.34
R228 VNB.t5 VNB.t8 2448.29
R229 VNB.t1 VNB.t7 2298.68
R230 VNB.t8 VNB.t15 2286.61
R231 VNB.t11 VNB.t10 2148.03
R232 VNB.t6 VNB.t4 2124.93
R233 VNB.t0 VNB.t5 2078.74
R234 VNB.t3 VNB.t1 1323.48
R235 VNB.n0 VNB.t2 1270.34
R236 VNB.t14 VNB 1265.44
R237 VNB.t15 VNB.t11 1212.6
R238 VNB.t2 VNB.t12 1154.86
R239 VNB.n0 VNB.t3 1021.64
R240 VNB.t7 VNB.t14 905.542
R241 VNB.t9 VNB.t6 900.788
R242 VNB.t12 VNB.t9 900.788
R243 a_494_366.t1 a_494_366.n4 874.292
R244 a_494_366.n1 a_494_366.t3 469.651
R245 a_494_366.n2 a_494_366.n1 461.154
R246 a_494_366.n3 a_494_366.t2 324.166
R247 a_494_366.n1 a_494_366.n0 316.575
R248 a_494_366.n2 a_494_366.t0 254.475
R249 a_494_366.n3 a_494_366.t4 209.403
R250 a_494_366.n4 a_494_366.n3 177.976
R251 a_494_366.n4 a_494_366.n2 75.3987
R252 D.n3 D.t0 220.296
R253 D D.n0 153.477
R254 D.n2 D.n1 152
R255 D.n4 D.n3 152
R256 D.n0 D.t1 148.417
R257 D.n3 D.n2 40.9705
R258 D.n2 D.n0 40.9705
R259 D.n1 D 9.68255
R260 D.n4 D 8.69794
R261 D D.n4 3.44665
R262 D.n1 D 2.46204
R263 a_37_78.n2 a_37_78.t2 659.236
R264 a_37_78.n1 a_37_78.n0 601.726
R265 a_37_78.n1 a_37_78.t4 367.041
R266 a_37_78.t0 a_37_78.n2 354.103
R267 a_37_78.n2 a_37_78.n1 159.209
R268 a_37_78.n0 a_37_78.t1 70.3576
R269 a_37_78.n0 a_37_78.t3 70.3576
R270 a_699_463.n1 a_699_463.t2 667.692
R271 a_699_463.n3 a_699_463.n2 609.02
R272 a_699_463.n0 a_699_463.t6 341.077
R273 a_699_463.n4 a_699_463.n3 300.865
R274 a_699_463.n1 a_699_463.n0 257.116
R275 a_699_463.n0 a_699_463.t5 174.903
R276 a_699_463.n2 a_699_463.t1 70.3576
R277 a_699_463.n2 a_699_463.t3 70.3576
R278 a_699_463.t0 a_699_463.n4 60.0005
R279 a_699_463.n3 a_699_463.n1 56.2863
R280 a_699_463.n4 a_699_463.t4 40.0005
R281 a_834_355.n5 a_834_355.n4 661.125
R282 a_834_355.n1 a_834_355.t4 301.05
R283 a_834_355.n3 a_834_355.n1 293.212
R284 a_834_355.n3 a_834_355.n2 185
R285 a_834_355.n1 a_834_355.t5 147.613
R286 a_834_355.n2 a_834_355.n0 104.697
R287 a_834_355.n4 a_834_355.n0 85.705
R288 a_834_355.n0 a_834_355.t3 67.0906
R289 a_834_355.n5 a_834_355.t2 29.5505
R290 a_834_355.t1 a_834_355.n5 29.5505
R291 a_834_355.n2 a_834_355.t0 22.7032
R292 a_834_355.n4 a_834_355.n3 13.1884
R293 a_2010_409.n13 a_2010_409.n12 353.483
R294 a_2010_409.n10 a_2010_409.t6 351.861
R295 a_2010_409.n2 a_2010_409.t5 287.594
R296 a_2010_409.n4 a_2010_409.t9 260.281
R297 a_2010_409.n2 a_2010_409.t8 240.197
R298 a_2010_409.n9 a_2010_409.t3 240.197
R299 a_2010_409.n3 a_2010_409.n1 237.787
R300 a_2010_409.n8 a_2010_409.t4 179.947
R301 a_2010_409.n6 a_2010_409.t7 179.947
R302 a_2010_409.n5 a_2010_409.n0 165.189
R303 a_2010_409.n12 a_2010_409.t1 157.095
R304 a_2010_409.n11 a_2010_409.n10 152
R305 a_2010_409.n7 a_2010_409.n0 152
R306 a_2010_409.n3 a_2010_409.n2 88.3672
R307 a_2010_409.n7 a_2010_409.n6 42.3581
R308 a_2010_409.n13 a_2010_409.t2 35.1791
R309 a_2010_409.t0 a_2010_409.n13 35.1791
R310 a_2010_409.n8 a_2010_409.n7 34.3247
R311 a_2010_409.n5 a_2010_409.n4 30.5272
R312 a_2010_409.n4 a_2010_409.n3 27.3138
R313 a_2010_409.n12 a_2010_409.n11 25.9884
R314 a_2010_409.n11 a_2010_409.n0 13.1884
R315 a_2010_409.n9 a_2010_409.n8 10.955
R316 a_2010_409.n6 a_2010_409.n5 7.30353
R317 a_2010_409.n10 a_2010_409.n9 4.38232
R318 Q.n2 Q.n0 286.283
R319 Q.n2 Q.n1 207.6
R320 Q.n4 Q.t1 145.78
R321 Q.n4 Q.n3 138.792
R322 Q.n0 Q.t5 34.2996
R323 Q.n5 Q.n2 31.9321
R324 Q.n3 Q.t0 30.8113
R325 Q.n3 Q.t2 30.0005
R326 Q.n1 Q.t4 26.3844
R327 Q.n1 Q.t3 26.3844
R328 Q.n0 Q.t6 26.3844
R329 Q.n5 Q.n4 16.392
R330 Q Q.n5 12.8005
R331 Q.n5 Q 6.4005
R332 a_1350_392.n5 a_1350_392.n4 514.227
R333 a_1350_392.n4 a_1350_392.n3 325.603
R334 a_1350_392.n2 a_1350_392.t2 285.962
R335 a_1350_392.n4 a_1350_392.t1 278.187
R336 a_1350_392.n3 a_1350_392.t4 268.313
R337 a_1350_392.n0 a_1350_392.t6 266.635
R338 a_1350_392.n0 a_1350_392.t3 250.105
R339 a_1350_392.n1 a_1350_392.t5 250.105
R340 a_1350_392.n1 a_1350_392.n0 86.7605
R341 a_1350_392.n2 a_1350_392.n1 67.4805
R342 a_1350_392.n6 a_1350_392.n5 26.0194
R343 a_1350_392.n5 a_1350_392.t0 25.4563
R344 a_1350_392.n3 a_1350_392.n2 13.146
R345 a_1678_395.n2 a_1678_395.t0 792.976
R346 a_1678_395.n1 a_1678_395.n0 417.923
R347 a_1678_395.t1 a_1678_395.n2 241.292
R348 a_1678_395.n2 a_1678_395.n1 225.412
R349 a_1678_395.n1 a_1678_395.t2 159.06
R350 a_890_138.t0 a_890_138.t1 68.5719
R351 a_812_138.t0 a_812_138.t1 68.5719
R352 a_789_463.t0 a_789_463.t1 112.572
C0 a_1627_493# VPWR 0.001485f
C1 RESET_B VGND 0.240838f
C2 VPWR CLK 0.017555f
C3 RESET_B Q 5.2e-19
C4 VPWR VGND 0.093874f
C5 CLK VGND 0.016048f
C6 VPWR Q 0.501463f
C7 VGND Q 0.328645f
C8 VPB D 0.09933f
C9 a_1827_81# VPWR 4.97e-19
C10 VPB RESET_B 0.348382f
C11 VPB VPWR 0.401044f
C12 D RESET_B 0.131724f
C13 a_1827_81# VGND 0.005927f
C14 D VPWR 0.036254f
C15 VPB CLK 0.036124f
C16 VPB VGND 0.018309f
C17 RESET_B VPWR 0.374762f
C18 a_1627_493# RESET_B 3.38e-19
C19 RESET_B CLK 0.045086f
C20 VPB Q 0.020233f
C21 D VGND 0.014594f
C22 Q VNB 0.055007f
C23 VGND VNB 1.5805f
C24 CLK VNB 0.112382f
C25 VPWR VNB 1.23129f
C26 RESET_B VNB 0.420822f
C27 D VNB 0.241627f
C28 VPB VNB 3.08647f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfrtp_2 VNB VPB RESET_B VPWR VGND D CLK Q
X0 a_786_457.t0 a_306_74.t2 a_696_457.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X1 a_696_457.t1 a_490_362.t2 a_30_78.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X2 a_1478_493.t0 a_490_362.t3 a_1271_74.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.22695 ps=1.83 w=0.42 l=0.15
X3 a_1921_409.t0 a_1271_74.t3 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1638 ps=1.275 w=0.84 l=0.15
X4 a_1525_212.t0 a_1271_74.t4 a_1663_81.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1176 pd=1.4 as=0.0504 ps=0.66 w=0.42 l=0.15
X5 VGND.t5 a_1921_409.t2 Q.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VGND.t6 RESET_B.t0 a_895_138.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.353275 pd=1.84 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_837_359.t1 a_696_457.t5 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.18405 pd=1.43 as=0.295 ps=2.59 w=1 l=0.15
X8 a_895_138.t0 a_837_359.t3 a_817_138.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X9 a_837_359.t2 a_696_457.t6 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.353275 ps=1.84 w=0.74 l=0.15
X10 Q.t2 a_1921_409.t3 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 a_817_138.t0 a_490_362.t4 a_696_457.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 VPWR.t9 RESET_B.t1 a_30_78.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X13 a_1921_409.t1 a_1271_74.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2072 ps=2.04 w=0.74 l=0.15
X14 a_117_78.t0 D.t0 a_30_78.t3 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X15 VPWR.t0 a_1921_409.t4 Q.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_1481_81.t0 a_306_74.t3 a_1271_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X17 a_1525_212.t2 RESET_B.t2 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=0.98 as=0.0735 ps=0.77 w=0.42 l=0.15
X18 Q.t0 a_1921_409.t5 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3584 ps=2.88 w=1.12 l=0.15
X19 VPWR.t3 a_1271_74.t6 a_1525_212.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.275 as=0.1176 ps=0.98 w=0.42 l=0.15
X20 a_490_362.t0 a_306_74.t4 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X21 a_696_457.t3 a_306_74.t5 a_30_78.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X22 VGND.t7 RESET_B.t3 a_117_78.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 a_696_457.t0 RESET_B.t4 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1393 ps=1.17 w=0.42 l=0.15
X24 a_1271_74.t0 a_306_74.t6 a_837_359.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.22695 pd=1.83 as=0.18405 ps=1.43 w=1 l=0.15
X25 a_490_362.t1 a_306_74.t7 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X26 VPWR.t8 a_837_359.t4 a_786_457.t1 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1393 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X27 a_30_78.t4 D.t1 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X28 VPWR.t7 CLK.t0 a_306_74.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X29 VPWR.t11 a_1525_212.t3 a_1478_493.t1 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.0567 ps=0.69 w=0.42 l=0.15
X30 VGND.t3 CLK.t1 a_306_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
R0 a_306_74.n0 a_306_74.t6 1018.89
R1 a_306_74.t1 a_306_74.n4 914.299
R2 a_306_74.t6 a_306_74.t3 792.087
R3 a_306_74.n1 a_306_74.n0 764.774
R4 a_306_74.n2 a_306_74.t5 340.613
R5 a_306_74.n1 a_306_74.t7 214.758
R6 a_306_74.n4 a_306_74.n3 213.617
R7 a_306_74.n0 a_306_74.t2 190.659
R8 a_306_74.n2 a_306_74.t4 151.028
R9 a_306_74.n4 a_306_74.t0 146.838
R10 a_306_74.n3 a_306_74.n1 28.3849
R11 a_306_74.n3 a_306_74.n2 13.3894
R12 a_696_457.n1 a_696_457.t0 675.644
R13 a_696_457.n3 a_696_457.n2 608.379
R14 a_696_457.n4 a_696_457.n3 293.776
R15 a_696_457.n1 a_696_457.n0 287.207
R16 a_696_457.n0 a_696_457.t5 221.738
R17 a_696_457.n0 a_696_457.t6 162.274
R18 a_696_457.n2 a_696_457.t4 70.3576
R19 a_696_457.n2 a_696_457.t1 70.3576
R20 a_696_457.n4 a_696_457.t3 60.0005
R21 a_696_457.n3 a_696_457.n1 49.2826
R22 a_696_457.t2 a_696_457.n4 40.0005
R23 a_786_457.t0 a_786_457.t1 126.644
R24 VPB.n0 VPB 3539.52
R25 VPB VPB.n1 672.01
R26 VPB.t0 VPB.t2 528.63
R27 VPB.t6 VPB.t4 497.964
R28 VPB.t3 VPB.t9 488.296
R29 VPB.t14 VPB.t11 362.635
R30 VPB.t12 VPB.t3 299.747
R31 VPB.t11 VPB.t0 298.791
R32 VPB.n1 VPB.t10 258.651
R33 VPB.t15 VPB.t14 255.376
R34 VPB.t16 VPB 252.823
R35 VPB.t7 VPB.n0 251.399
R36 VPB.t9 VPB.t7 244.149
R37 VPB.t2 VPB.t1 229.839
R38 VPB.t13 VPB.t16 229.839
R39 VPB.n1 VPB.t13 227.286
R40 VPB.t4 VPB.t8 217.558
R41 VPB.t10 VPB.t6 217.558
R42 VPB.t5 VPB.t15 214.517
R43 VPB.t8 VPB.t12 203.054
R44 VPB.n0 VPB.t5 196.641
R45 a_490_362.t1 a_490_362.n4 889.256
R46 a_490_362.n1 a_490_362.n0 471.397
R47 a_490_362.n2 a_490_362.n1 408.06
R48 a_490_362.n3 a_490_362.t4 339.793
R49 a_490_362.n1 a_490_362.t3 325.659
R50 a_490_362.n2 a_490_362.t0 207.703
R51 a_490_362.n3 a_490_362.t2 197.352
R52 a_490_362.n4 a_490_362.n3 166.546
R53 a_490_362.n4 a_490_362.n2 62.1892
R54 a_30_78.n2 a_30_78.t1 660.477
R55 a_30_78.n1 a_30_78.n0 601.98
R56 a_30_78.n1 a_30_78.t3 363.615
R57 a_30_78.t0 a_30_78.n2 359.687
R58 a_30_78.n2 a_30_78.n1 170.542
R59 a_30_78.n0 a_30_78.t2 70.3576
R60 a_30_78.n0 a_30_78.t4 70.3576
R61 a_1271_74.n4 a_1271_74.n0 585
R62 a_1271_74.n6 a_1271_74.n5 585
R63 a_1271_74.n3 a_1271_74.t4 349.894
R64 a_1271_74.n5 a_1271_74.t1 334.647
R65 a_1271_74.n4 a_1271_74.n3 319.666
R66 a_1271_74.n1 a_1271_74.t5 287.594
R67 a_1271_74.n6 a_1271_74.n0 234.117
R68 a_1271_74.n1 a_1271_74.t3 230.022
R69 a_1271_74.n2 a_1271_74.t6 225.47
R70 a_1271_74.n2 a_1271_74.n1 172.01
R71 a_1271_74.t0 a_1271_74.n6 82.2634
R72 a_1271_74.n0 a_1271_74.t2 71.8871
R73 a_1271_74.n5 a_1271_74.n4 15.9035
R74 a_1271_74.n3 a_1271_74.n2 10.7915
R75 a_1478_493.t0 a_1478_493.t1 126.644
R76 VPWR.n33 VPWR.n7 695.713
R77 VPWR.n46 VPWR.t12 677.855
R78 VPWR.n44 VPWR.t9 676.691
R79 VPWR.n24 VPWR.n12 610.407
R80 VPWR.n19 VPWR.n15 610.407
R81 VPWR.n3 VPWR.n2 606.915
R82 VPWR.n16 VPWR.t0 266.195
R83 VPWR.n31 VPWR.t6 260.43
R84 VPWR.n17 VPWR.t1 254.477
R85 VPWR.n7 VPWR.t4 110.227
R86 VPWR.n7 VPWR.t8 110.227
R87 VPWR.n15 VPWR.t3 110.227
R88 VPWR.n12 VPWR.t10 93.81
R89 VPWR.n12 VPWR.t11 70.3576
R90 VPWR.n15 VPWR.t2 52.7684
R91 VPWR.n37 VPWR.n5 36.1417
R92 VPWR.n38 VPWR.n37 36.1417
R93 VPWR.n39 VPWR.n38 36.1417
R94 VPWR.n26 VPWR.n25 36.1417
R95 VPWR.n26 VPWR.n9 36.1417
R96 VPWR.n30 VPWR.n9 36.1417
R97 VPWR.n23 VPWR.n13 36.1417
R98 VPWR.n32 VPWR.n31 35.7652
R99 VPWR.n19 VPWR.n18 31.624
R100 VPWR.n25 VPWR.n24 26.7299
R101 VPWR.n2 VPWR.t5 26.3844
R102 VPWR.n2 VPWR.t7 26.3844
R103 VPWR.n44 VPWR.n43 25.977
R104 VPWR.n33 VPWR.n5 25.6005
R105 VPWR.n39 VPWR.n3 24.4711
R106 VPWR.n18 VPWR.n17 23.3417
R107 VPWR.n43 VPWR.n3 22.9652
R108 VPWR.n33 VPWR.n32 21.8358
R109 VPWR.n45 VPWR.n44 21.4593
R110 VPWR.n46 VPWR.n45 21.4593
R111 VPWR.n24 VPWR.n23 20.7064
R112 VPWR.n19 VPWR.n13 15.8123
R113 VPWR.n31 VPWR.n30 11.6711
R114 VPWR.n18 VPWR.n14 9.3005
R115 VPWR.n20 VPWR.n19 9.3005
R116 VPWR.n21 VPWR.n13 9.3005
R117 VPWR.n23 VPWR.n22 9.3005
R118 VPWR.n24 VPWR.n11 9.3005
R119 VPWR.n25 VPWR.n10 9.3005
R120 VPWR.n27 VPWR.n26 9.3005
R121 VPWR.n28 VPWR.n9 9.3005
R122 VPWR.n30 VPWR.n29 9.3005
R123 VPWR.n31 VPWR.n8 9.3005
R124 VPWR.n32 VPWR.n6 9.3005
R125 VPWR.n34 VPWR.n33 9.3005
R126 VPWR.n35 VPWR.n5 9.3005
R127 VPWR.n37 VPWR.n36 9.3005
R128 VPWR.n38 VPWR.n4 9.3005
R129 VPWR.n40 VPWR.n39 9.3005
R130 VPWR.n41 VPWR.n3 9.3005
R131 VPWR.n43 VPWR.n42 9.3005
R132 VPWR.n44 VPWR.n1 9.3005
R133 VPWR.n45 VPWR.n0 9.3005
R134 VPWR.n47 VPWR.n46 9.3005
R135 VPWR.n17 VPWR.n16 6.72092
R136 VPWR.n16 VPWR.n14 0.589622
R137 VPWR.n20 VPWR.n14 0.122949
R138 VPWR.n21 VPWR.n20 0.122949
R139 VPWR.n22 VPWR.n21 0.122949
R140 VPWR.n22 VPWR.n11 0.122949
R141 VPWR.n11 VPWR.n10 0.122949
R142 VPWR.n27 VPWR.n10 0.122949
R143 VPWR.n28 VPWR.n27 0.122949
R144 VPWR.n29 VPWR.n28 0.122949
R145 VPWR.n29 VPWR.n8 0.122949
R146 VPWR.n8 VPWR.n6 0.122949
R147 VPWR.n34 VPWR.n6 0.122949
R148 VPWR.n35 VPWR.n34 0.122949
R149 VPWR.n36 VPWR.n35 0.122949
R150 VPWR.n36 VPWR.n4 0.122949
R151 VPWR.n40 VPWR.n4 0.122949
R152 VPWR.n41 VPWR.n40 0.122949
R153 VPWR.n42 VPWR.n41 0.122949
R154 VPWR.n42 VPWR.n1 0.122949
R155 VPWR.n1 VPWR.n0 0.122949
R156 VPWR.n47 VPWR.n0 0.122949
R157 VPWR VPWR.n47 0.0617245
R158 a_1921_409.t0 a_1921_409.n3 418.755
R159 a_1921_409.n0 a_1921_409.t4 308.481
R160 a_1921_409.n2 a_1921_409.t5 288.397
R161 a_1921_409.n3 a_1921_409.n2 275.714
R162 a_1921_409.n0 a_1921_409.t2 200.03
R163 a_1921_409.n1 a_1921_409.t3 179.947
R164 a_1921_409.n3 a_1921_409.t1 160.668
R165 a_1921_409.n1 a_1921_409.n0 104.433
R166 a_1921_409.n2 a_1921_409.n1 11.2472
R167 a_1525_212.n3 a_1525_212.n2 717.758
R168 a_1525_212.n1 a_1525_212.t3 414.788
R169 a_1525_212.t0 a_1525_212.n3 251.764
R170 a_1525_212.n3 a_1525_212.n1 212.988
R171 a_1525_212.n1 a_1525_212.n0 167.094
R172 a_1525_212.n2 a_1525_212.t1 131.333
R173 a_1525_212.n2 a_1525_212.t2 131.333
R174 VNB VNB.n0 16006.3
R175 VNB.t4 VNB.t1 3002.62
R176 VNB.n0 VNB.t5 2750
R177 VNB.t2 VNB.t3 2566.67
R178 VNB.t5 VNB.t11 2481.11
R179 VNB.t6 VNB.t12 2420
R180 VNB.t0 VNB.t8 2286.61
R181 VNB.t1 VNB.t0 2263.52
R182 VNB.t3 VNB.t6 1393.33
R183 VNB.t13 VNB 1246.67
R184 VNB.t7 VNB.t2 1222.22
R185 VNB.t8 VNB.t9 993.177
R186 VNB.t11 VNB.t10 953.333
R187 VNB.t10 VNB.t7 953.333
R188 VNB.t12 VNB.t13 953.333
R189 VNB.n0 VNB.t4 923.885
R190 Q.n4 Q 589.85
R191 Q.n4 Q.n0 585
R192 Q.n5 Q.n4 585
R193 Q.n3 Q.n2 185
R194 Q.n2 Q.n1 185
R195 Q.n4 Q.t1 26.3844
R196 Q.n4 Q.t0 26.3844
R197 Q.n2 Q.t3 22.7032
R198 Q.n2 Q.t2 22.7032
R199 Q Q.n5 12.9944
R200 Q.n1 Q 12.6066
R201 Q Q.n0 11.249
R202 Q Q.n3 9.50353
R203 Q.n3 Q 4.84898
R204 Q Q.n0 3.10353
R205 Q.n1 Q 1.74595
R206 Q.n5 Q 1.35808
R207 VGND.n41 VGND.t7 255.464
R208 VGND.n28 VGND.n27 213.053
R209 VGND.n39 VGND.n2 209.048
R210 VGND.n11 VGND.t5 179.673
R211 VGND.n10 VGND.t4 171.77
R212 VGND.n14 VGND.t0 163.141
R213 VGND.n27 VGND.t2 97.2978
R214 VGND.n27 VGND.t6 52.2399
R215 VGND.n15 VGND.n8 36.1417
R216 VGND.n21 VGND.n20 36.1417
R217 VGND.n21 VGND.n6 36.1417
R218 VGND.n25 VGND.n6 36.1417
R219 VGND.n26 VGND.n25 36.1417
R220 VGND.n33 VGND.n4 36.1417
R221 VGND.n34 VGND.n33 36.1417
R222 VGND.n35 VGND.n34 36.1417
R223 VGND.n35 VGND.n1 36.1417
R224 VGND.n2 VGND.t1 34.0546
R225 VGND.n2 VGND.t3 34.0546
R226 VGND.n41 VGND.n40 30.1181
R227 VGND.n29 VGND.n4 30.0045
R228 VGND.n13 VGND.n10 28.6123
R229 VGND.n14 VGND.n13 27.1064
R230 VGND.n15 VGND.n14 26.3534
R231 VGND.n20 VGND.n19 24.8476
R232 VGND.n40 VGND.n39 24.8476
R233 VGND.n39 VGND.n1 22.5887
R234 VGND.n28 VGND.n26 18.3694
R235 VGND.n19 VGND.n8 15.8123
R236 VGND.n40 VGND.n0 9.3005
R237 VGND.n39 VGND.n38 9.3005
R238 VGND.n37 VGND.n1 9.3005
R239 VGND.n36 VGND.n35 9.3005
R240 VGND.n34 VGND.n3 9.3005
R241 VGND.n33 VGND.n32 9.3005
R242 VGND.n31 VGND.n4 9.3005
R243 VGND.n30 VGND.n29 9.3005
R244 VGND.n26 VGND.n5 9.3005
R245 VGND.n25 VGND.n24 9.3005
R246 VGND.n23 VGND.n6 9.3005
R247 VGND.n22 VGND.n21 9.3005
R248 VGND.n20 VGND.n7 9.3005
R249 VGND.n19 VGND.n18 9.3005
R250 VGND.n17 VGND.n8 9.3005
R251 VGND.n16 VGND.n15 9.3005
R252 VGND.n14 VGND.n9 9.3005
R253 VGND.n13 VGND.n12 9.3005
R254 VGND.n42 VGND.n41 7.13181
R255 VGND.n11 VGND.n10 6.77202
R256 VGND.n29 VGND.n28 2.17408
R257 VGND.n12 VGND.n11 0.577493
R258 VGND VGND.n42 0.27433
R259 VGND.n42 VGND.n0 0.156458
R260 VGND.n12 VGND.n9 0.122949
R261 VGND.n16 VGND.n9 0.122949
R262 VGND.n17 VGND.n16 0.122949
R263 VGND.n18 VGND.n17 0.122949
R264 VGND.n18 VGND.n7 0.122949
R265 VGND.n22 VGND.n7 0.122949
R266 VGND.n23 VGND.n22 0.122949
R267 VGND.n24 VGND.n23 0.122949
R268 VGND.n24 VGND.n5 0.122949
R269 VGND.n30 VGND.n5 0.122949
R270 VGND.n31 VGND.n30 0.122949
R271 VGND.n32 VGND.n31 0.122949
R272 VGND.n32 VGND.n3 0.122949
R273 VGND.n36 VGND.n3 0.122949
R274 VGND.n37 VGND.n36 0.122949
R275 VGND.n38 VGND.n37 0.122949
R276 VGND.n38 VGND.n0 0.122949
R277 RESET_B.n1 RESET_B.n0 451.474
R278 RESET_B.n2 RESET_B.t0 286.087
R279 RESET_B.n4 RESET_B.t3 222.916
R280 RESET_B.n4 RESET_B.t1 219.874
R281 RESET_B.n3 RESET_B.n1 174.948
R282 RESET_B.n3 RESET_B.n2 164.185
R283 RESET_B.n1 RESET_B.t2 146.475
R284 RESET_B.n2 RESET_B.t4 130.911
R285 RESET_B.n5 RESET_B.n4 57.2968
R286 RESET_B.n5 RESET_B.n3 3.32775
R287 RESET_B RESET_B.n5 0.0466957
R288 a_895_138.t0 a_895_138.t1 68.5719
R289 a_837_359.n2 a_837_359.n1 362.404
R290 a_837_359.n1 a_837_359.n0 325.457
R291 a_837_359.n0 a_837_359.t3 310.985
R292 a_837_359.n1 a_837_359.t2 214.685
R293 a_837_359.n0 a_837_359.t4 137.732
R294 a_837_359.n2 a_837_359.t1 40.3644
R295 a_837_359.t0 a_837_359.n2 30.6131
R296 a_817_138.t0 a_817_138.t1 68.5719
R297 D.n3 D.t1 235.208
R298 D D.n0 153.558
R299 D.n2 D.n1 152
R300 D.n4 D.n3 152
R301 D.n0 D.t0 150.322
R302 D.n3 D.n2 44.8991
R303 D.n2 D.n0 44.8991
R304 D.n1 D 10.2059
R305 D.n4 D 9.16807
R306 D D.n4 3.63293
R307 D.n1 D 2.59509
R308 a_117_78.t0 a_117_78.t1 68.5719
R309 CLK.n0 CLK.t0 250.909
R310 CLK.n0 CLK.t1 210.474
R311 CLK CLK.n0 158.4
C0 VPB D 0.095356f
C1 VPB RESET_B 0.361111f
C2 VPB VPWR 0.375711f
C3 D RESET_B 0.130002f
C4 D VPWR 0.040378f
C5 VPB CLK 0.043085f
C6 RESET_B VPWR 0.403245f
C7 VPB VGND 0.021676f
C8 RESET_B CLK 0.043105f
C9 D VGND 0.013088f
C10 VPB Q 0.006935f
C11 RESET_B VGND 0.221429f
C12 VPWR CLK 0.017721f
C13 VPWR VGND 0.097462f
C14 RESET_B Q 1.86e-19
C15 CLK VGND 0.016443f
C16 VPWR Q 0.230314f
C17 VGND Q 0.164633f
C18 Q VNB 0.033274f
C19 VGND VNB 1.38669f
C20 CLK VNB 0.104552f
C21 VPWR VNB 1.08691f
C22 RESET_B VNB 0.387751f
C23 D VNB 0.236178f
C24 VPB VNB 2.72588f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfrtp_1 VNB VPB VPWR RESET_B VGND Q CLK D
X0 a_894_138.t0 a_830_359# a_816_138.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 VPWR.t2 a_1518_203.t2 a_1468_493.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1864_409.t0 a_1266_74.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3 a_816_138.t1 a_490_366.t2 a_695_457.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4 a_830_359# a_695_457.t5 VGND.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.211225 ps=1.45 w=0.74 l=0.15
X5 a_1476_81.t1 a_306_74.t2 a_1266_74.t3 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X6 VGND.t6 a_1864_409.t2 Q.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 a_490_366.t1 a_306_74.t3 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t5 CLK.t0 a_306_74.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X9 a_1468_493.t1 a_490_366.t3 a_1266_74.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X10 a_1266_74.t2 a_306_74.t4 a_830_359# VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.190625 ps=1.505 w=1 l=0.15
X11 a_1656_81.t0 RESET_B.t0 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X12 VPWR.t3 a_1864_409.t3 Q.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X13 a_1864_409.t1 a_1266_74.t5 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X14 VPWR.t1 a_1266_74.t6 a_1518_203.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X15 VPWR.t6 RESET_B.t1 a_30_78.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X16 a_117_78.t1 D.t0 a_30_78.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X17 a_695_457.t4 a_306_74.t5 a_30_78.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X18 a_1518_203.t1 a_1266_74.t7 a_1656_81.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 a_695_457.t2 RESET_B.t2 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.137125 ps=1.155 w=0.42 l=0.15
X20 a_490_366.t0 a_306_74.t6 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X21 VPWR.t4 a_830_359# a_785_457.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.137125 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 VGND.t0 a_1518_203.t3 a_1476_81.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 VGND.t7 RESET_B.t3 a_117_78.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X24 a_785_457.t1 a_306_74.t7 a_695_457.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X25 a_695_457.t1 a_490_366.t4 a_30_78.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X26 a_1266_74.t1 a_490_366.t5 a_830_359# VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X27 a_30_78.t3 D.t1 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X28 VGND.t1 CLK.t1 a_306_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X29 VGND.t8 RESET_B.t4 a_894_138.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.211225 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_816_138.t0 a_816_138.t1 68.5719
R1 a_894_138.t0 a_894_138.t1 68.5719
R2 VNB.n0 VNB 14782.2
R3 VNB VNB.n1 13004.4
R4 VNB.t12 VNB.t11 2588.92
R5 VNB.t6 VNB.t13 2298.68
R6 VNB.t1 VNB.t4 2286.61
R7 VNB.t2 VNB.t1 2286.61
R8 VNB.n0 VNB.t15 2090.29
R9 VNB.t0 VNB.t3 1992.22
R10 VNB.n1 VNB.t14 1242.22
R11 VNB.t5 VNB 1184.17
R12 VNB.t9 VNB.t8 1177.95
R13 VNB.t10 VNB.t12 1160.95
R14 VNB.t11 VNB.t6 1160.95
R15 VNB.t14 VNB.t7 905.542
R16 VNB.t7 VNB.t10 905.542
R17 VNB.t13 VNB.t5 905.542
R18 VNB.t15 VNB.t9 900.788
R19 VNB.t8 VNB.t2 831.496
R20 VNB.t3 VNB.n0 354.445
R21 VNB.n1 VNB.t0 293.334
R22 a_1518_203.n1 a_1518_203.t0 795.564
R23 a_1518_203.n0 a_1518_203.t2 416.93
R24 a_1518_203.t1 a_1518_203.n1 243.812
R25 a_1518_203.n1 a_1518_203.n0 210.73
R26 a_1518_203.n0 a_1518_203.t3 152.633
R27 a_1468_493.t0 a_1468_493.t1 126.644
R28 VPWR.n17 VPWR.t2 708.907
R29 VPWR.n26 VPWR.n7 686.106
R30 VPWR.n39 VPWR.t8 685.053
R31 VPWR.n37 VPWR.t6 681.726
R32 VPWR.n3 VPWR.n2 606.139
R33 VPWR.n13 VPWR.n12 319.026
R34 VPWR.n14 VPWR.t3 258.324
R35 VPWR.n7 VPWR.t7 110.227
R36 VPWR.n7 VPWR.t4 110.227
R37 VPWR.n12 VPWR.t1 110.227
R38 VPWR.n30 VPWR.n5 36.1417
R39 VPWR.n31 VPWR.n30 36.1417
R40 VPWR.n32 VPWR.n31 36.1417
R41 VPWR.n19 VPWR.n18 36.1417
R42 VPWR.n19 VPWR.n9 36.1417
R43 VPWR.n23 VPWR.n9 36.1417
R44 VPWR.n12 VPWR.t0 35.1791
R45 VPWR.n16 VPWR.n13 34.2593
R46 VPWR.n25 VPWR.n24 33.1299
R47 VPWR.n38 VPWR.n37 27.4829
R48 VPWR.n39 VPWR.n38 27.4829
R49 VPWR.n18 VPWR.n17 27.4829
R50 VPWR.n2 VPWR.t9 26.3844
R51 VPWR.n2 VPWR.t5 26.3844
R52 VPWR.n37 VPWR.n36 25.977
R53 VPWR.n32 VPWR.n3 24.4711
R54 VPWR.n26 VPWR.n25 24.4711
R55 VPWR.n36 VPWR.n3 22.9652
R56 VPWR.n26 VPWR.n5 22.9652
R57 VPWR.n17 VPWR.n16 19.9534
R58 VPWR.n24 VPWR.n23 14.3064
R59 VPWR.n16 VPWR.n15 9.3005
R60 VPWR.n17 VPWR.n11 9.3005
R61 VPWR.n18 VPWR.n10 9.3005
R62 VPWR.n20 VPWR.n19 9.3005
R63 VPWR.n21 VPWR.n9 9.3005
R64 VPWR.n23 VPWR.n22 9.3005
R65 VPWR.n24 VPWR.n8 9.3005
R66 VPWR.n25 VPWR.n6 9.3005
R67 VPWR.n27 VPWR.n26 9.3005
R68 VPWR.n28 VPWR.n5 9.3005
R69 VPWR.n30 VPWR.n29 9.3005
R70 VPWR.n31 VPWR.n4 9.3005
R71 VPWR.n33 VPWR.n32 9.3005
R72 VPWR.n34 VPWR.n3 9.3005
R73 VPWR.n36 VPWR.n35 9.3005
R74 VPWR.n37 VPWR.n1 9.3005
R75 VPWR.n38 VPWR.n0 9.3005
R76 VPWR.n40 VPWR.n39 9.3005
R77 VPWR.n14 VPWR.n13 6.37758
R78 VPWR.n15 VPWR.n14 0.190046
R79 VPWR.n15 VPWR.n11 0.122949
R80 VPWR.n11 VPWR.n10 0.122949
R81 VPWR.n20 VPWR.n10 0.122949
R82 VPWR.n21 VPWR.n20 0.122949
R83 VPWR.n22 VPWR.n21 0.122949
R84 VPWR.n22 VPWR.n8 0.122949
R85 VPWR.n8 VPWR.n6 0.122949
R86 VPWR.n27 VPWR.n6 0.122949
R87 VPWR.n28 VPWR.n27 0.122949
R88 VPWR.n29 VPWR.n28 0.122949
R89 VPWR.n29 VPWR.n4 0.122949
R90 VPWR.n33 VPWR.n4 0.122949
R91 VPWR.n34 VPWR.n33 0.122949
R92 VPWR.n35 VPWR.n34 0.122949
R93 VPWR.n35 VPWR.n1 0.122949
R94 VPWR.n1 VPWR.n0 0.122949
R95 VPWR.n40 VPWR.n0 0.122949
R96 VPWR VPWR.n40 0.0617245
R97 VPB.t13 VPB 3261.16
R98 VPB.t9 VPB.t13 774.734
R99 VPB VPB.n0 706.15
R100 VPB.t0 VPB.t5 656.317
R101 VPB.t2 VPB.t1 523.521
R102 VPB.t12 VPB.t4 520.722
R103 VPB.t13 VPB.t3 445.622
R104 VPB.t6 VPB.t9 314.974
R105 VPB.t1 VPB.t0 273.253
R106 VPB.n0 VPB.t7 271.791
R107 VPB.t10 VPB 252.823
R108 VPB.t8 VPB.t10 229.839
R109 VPB.t4 VPB.t11 228.611
R110 VPB.t7 VPB.t12 228.611
R111 VPB.n0 VPB.t8 227.286
R112 VPB.t3 VPB.t2 214.517
R113 VPB.t11 VPB.t6 198.129
R114 a_1266_74.n4 a_1266_74.n0 585
R115 a_1266_74.n7 a_1266_74.n6 585
R116 a_1266_74.n4 a_1266_74.n3 310.7
R117 a_1266_74.n1 a_1266_74.t5 284.38
R118 a_1266_74.n2 a_1266_74.t6 280.363
R119 a_1266_74.n3 a_1266_74.t7 257.284
R120 a_1266_74.n1 a_1266_74.t4 237.569
R121 a_1266_74.n6 a_1266_74.n5 198.107
R122 a_1266_74.n7 a_1266_74.n0 185.274
R123 a_1266_74.n5 a_1266_74.t3 139.399
R124 a_1266_74.n2 a_1266_74.n1 75.952
R125 a_1266_74.n5 a_1266_74.t1 71.5068
R126 a_1266_74.n0 a_1266_74.t0 70.3576
R127 a_1266_74.t2 a_1266_74.n7 51.4081
R128 a_1266_74.n6 a_1266_74.n4 15.3217
R129 a_1266_74.n3 a_1266_74.n2 3.65202
R130 a_1864_409.t0 a_1864_409.n1 434.01
R131 a_1864_409.n1 a_1864_409.n0 263.007
R132 a_1864_409.n1 a_1864_409.t1 248.089
R133 a_1864_409.n0 a_1864_409.t3 217.436
R134 a_1864_409.n0 a_1864_409.t2 209.452
R135 a_490_366.t1 a_490_366.n3 886.727
R136 a_490_366.n0 a_490_366.t5 472.753
R137 a_490_366.n1 a_490_366.n0 395.476
R138 a_490_366.n2 a_490_366.t2 320.851
R139 a_490_366.n0 a_490_366.t3 317.57
R140 a_490_366.n1 a_490_366.t0 219.054
R141 a_490_366.n2 a_490_366.t4 201.369
R142 a_490_366.n3 a_490_366.n2 166.739
R143 a_490_366.n3 a_490_366.n1 62.7097
R144 a_695_457.n2 a_695_457.t2 675.069
R145 a_695_457.n4 a_695_457.n3 608.063
R146 a_695_457.n5 a_695_457.n4 294.058
R147 a_695_457.n1 a_695_457.n0 285.743
R148 a_695_457.n2 a_695_457.n1 238.543
R149 a_695_457.n1 a_695_457.t5 186.374
R150 a_695_457.n3 a_695_457.t3 70.3576
R151 a_695_457.n3 a_695_457.t1 70.3576
R152 a_695_457.n5 a_695_457.t4 60.0005
R153 a_695_457.n4 a_695_457.n2 49.9054
R154 a_695_457.t0 a_695_457.n5 40.0005
R155 VGND.n38 VGND.t7 255.72
R156 VGND.n11 VGND.t2 246.01
R157 VGND.n16 VGND.n9 208.856
R158 VGND.n36 VGND.n2 207.304
R159 VGND.n25 VGND.n24 205.282
R160 VGND.n10 VGND.t6 179.31
R161 VGND.n9 VGND.t3 62.8576
R162 VGND.n24 VGND.t8 49.8075
R163 VGND.n24 VGND.t4 41.3519
R164 VGND.n9 VGND.t0 40.0005
R165 VGND.n12 VGND.n8 36.1417
R166 VGND.n18 VGND.n17 36.1417
R167 VGND.n18 VGND.n6 36.1417
R168 VGND.n22 VGND.n6 36.1417
R169 VGND.n23 VGND.n22 36.1417
R170 VGND.n30 VGND.n4 36.1417
R171 VGND.n31 VGND.n30 36.1417
R172 VGND.n32 VGND.n31 36.1417
R173 VGND.n32 VGND.n1 36.1417
R174 VGND.n2 VGND.t1 34.0546
R175 VGND.n38 VGND.n37 30.1181
R176 VGND.n26 VGND.n4 30.0632
R177 VGND.n37 VGND.n36 24.8476
R178 VGND.n16 VGND.n8 24.4711
R179 VGND.n17 VGND.n16 22.9652
R180 VGND.n2 VGND.t5 22.7032
R181 VGND.n36 VGND.n1 22.5887
R182 VGND.n12 VGND.n11 22.2123
R183 VGND.n25 VGND.n23 21.1456
R184 VGND.n37 VGND.n0 9.3005
R185 VGND.n36 VGND.n35 9.3005
R186 VGND.n34 VGND.n1 9.3005
R187 VGND.n33 VGND.n32 9.3005
R188 VGND.n31 VGND.n3 9.3005
R189 VGND.n30 VGND.n29 9.3005
R190 VGND.n28 VGND.n4 9.3005
R191 VGND.n27 VGND.n26 9.3005
R192 VGND.n23 VGND.n5 9.3005
R193 VGND.n22 VGND.n21 9.3005
R194 VGND.n20 VGND.n6 9.3005
R195 VGND.n19 VGND.n18 9.3005
R196 VGND.n17 VGND.n7 9.3005
R197 VGND.n16 VGND.n15 9.3005
R198 VGND.n14 VGND.n8 9.3005
R199 VGND.n13 VGND.n12 9.3005
R200 VGND.n11 VGND.n10 7.41876
R201 VGND.n39 VGND.n38 7.13181
R202 VGND.n26 VGND.n25 1.86717
R203 VGND VGND.n39 0.27433
R204 VGND.n13 VGND.n10 0.216393
R205 VGND.n39 VGND.n0 0.156458
R206 VGND.n14 VGND.n13 0.122949
R207 VGND.n15 VGND.n14 0.122949
R208 VGND.n15 VGND.n7 0.122949
R209 VGND.n19 VGND.n7 0.122949
R210 VGND.n20 VGND.n19 0.122949
R211 VGND.n21 VGND.n20 0.122949
R212 VGND.n21 VGND.n5 0.122949
R213 VGND.n27 VGND.n5 0.122949
R214 VGND.n28 VGND.n27 0.122949
R215 VGND.n29 VGND.n28 0.122949
R216 VGND.n29 VGND.n3 0.122949
R217 VGND.n33 VGND.n3 0.122949
R218 VGND.n34 VGND.n33 0.122949
R219 VGND.n35 VGND.n34 0.122949
R220 VGND.n35 VGND.n0 0.122949
R221 a_306_74.n0 a_306_74.t4 992.385
R222 a_306_74.t1 a_306_74.n4 935.407
R223 a_306_74.t4 a_306_74.t2 803.333
R224 a_306_74.n1 a_306_74.n0 772.808
R225 a_306_74.n1 a_306_74.t5 283.462
R226 a_306_74.n2 a_306_74.t3 261.007
R227 a_306_74.n4 a_306_74.n3 214.45
R228 a_306_74.n0 a_306_74.t7 190.659
R229 a_306_74.n2 a_306_74.t6 147.814
R230 a_306_74.n4 a_306_74.t0 146.505
R231 a_306_74.n3 a_306_74.n1 42.6919
R232 a_306_74.n3 a_306_74.n2 24.7891
R233 a_1476_81.t0 a_1476_81.t1 68.5719
R234 Q Q.n0 587.287
R235 Q.n2 Q.n0 585
R236 Q.n1 Q.n0 585
R237 Q Q.t1 188.859
R238 Q.n0 Q.t0 34.2996
R239 Q Q.n1 4.93764
R240 Q Q.n2 4.75479
R241 Q.n2 Q 2.01193
R242 Q.n1 Q 1.82907
R243 CLK.n0 CLK.t0 258.942
R244 CLK.n0 CLK.t1 207.261
R245 CLK CLK.n0 158.4
R246 RESET_B.n1 RESET_B.t0 444.688
R247 RESET_B.n2 RESET_B.t4 284.962
R248 RESET_B.n4 RESET_B.t1 219.607
R249 RESET_B.n4 RESET_B.t3 216.798
R250 RESET_B.n3 RESET_B.n1 173.704
R251 RESET_B.n3 RESET_B.n2 164.185
R252 RESET_B.n1 RESET_B.n0 151.47
R253 RESET_B.n2 RESET_B.t2 129.785
R254 RESET_B.n5 RESET_B.n4 59.2547
R255 RESET_B.n5 RESET_B.n3 3.32775
R256 RESET_B RESET_B.n5 0.0466957
R257 a_1656_81.t0 a_1656_81.t1 60.0005
R258 a_30_78.n0 a_30_78.t1 658.942
R259 a_30_78.n2 a_30_78.n1 601.922
R260 a_30_78.t2 a_30_78.n2 369.808
R261 a_30_78.n0 a_30_78.t4 357.579
R262 a_30_78.n2 a_30_78.n0 158.081
R263 a_30_78.n1 a_30_78.t0 70.3576
R264 a_30_78.n1 a_30_78.t3 70.3576
R265 D.n3 D.t1 235.208
R266 D D.n0 153.477
R267 D.n2 D.n1 152
R268 D.n4 D.n3 152
R269 D.n0 D.t0 150.322
R270 D.n3 D.n2 44.8991
R271 D.n2 D.n0 44.8991
R272 D.n1 D 9.68255
R273 D.n4 D 8.69794
R274 D D.n4 3.44665
R275 D.n1 D 2.46204
R276 a_117_78.t0 a_117_78.t1 68.5719
R277 a_785_457.t0 a_785_457.t1 112.572
C0 a_830_359# RESET_B 0.145411f
C1 VGND Q 0.105407f
C2 a_830_359# VPWR 0.120886f
C3 VPB D 0.0959f
C4 VPB RESET_B 0.343297f
C5 D RESET_B 0.129984f
C6 VPB VPWR 0.346367f
C7 VPB CLK 0.036397f
C8 D VPWR 0.035113f
C9 VGND a_830_359# 0.02944f
C10 VPB Q 0.028715f
C11 RESET_B VPWR 0.40365f
C12 RESET_B CLK 0.045935f
C13 VGND VPB 0.018485f
C14 RESET_B Q 7.03e-19
C15 VPWR CLK 0.017858f
C16 VGND D 0.013075f
C17 VPWR Q 0.178209f
C18 VGND RESET_B 0.219436f
C19 a_830_359# VPB 0.081281f
C20 VGND VPWR 0.077677f
C21 VGND CLK 0.016325f
C22 VGND VNB 1.33025f
C23 Q VNB 0.037352f
C24 CLK VNB 0.1118f
C25 VPWR VNB 1.04773f
C26 RESET_B VNB 0.401057f
C27 D VNB 0.236431f
C28 VPB VNB 2.56727f
C29 a_830_359# VNB 0.105931f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfrtn_1 VNB VPB VPWR RESET_B VGND CLK_N Q D
X0 a_714_127.t0 a_300_74.t2 a_33_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1 a_1266_119.t0 a_300_74.t3 a_856_304# VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.3067 pd=2.01 as=0.1073 ps=1.03 w=0.74 l=0.15
X2 a_33_74.t1 D.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X3 a_1266_119.t1 a_507_368.t2 a_856_304# VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.22385 pd=1.7 as=0.39 ps=1.78 w=1 l=0.15
X4 a_714_127.t3 a_507_368.t3 a_33_74.t4 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VPWR.t5 a_1266_119.t3 a_1598_93.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.39 as=0.063 ps=0.72 w=0.42 l=0.15
X6 VGND.t0 RESET_B.t0 a_120_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_507_368.t1 a_300_74.t4 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2596 pd=2.24 as=0.3593 ps=2.88 w=0.74 l=0.15
X8 a_300_74.t0 CLK_N.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.1673 ps=1.475 w=1.12 l=0.15
X9 a_1736_119.t0 RESET_B.t1 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 a_850_127.t0 a_300_74.t5 a_714_127.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1113 ps=0.95 w=0.42 l=0.15
X11 a_1550_119.t0 a_507_368.t4 a_1266_119.t2 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.3067 ps=2.01 w=0.42 l=0.15
X12 a_856_304# a_714_127.t5 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.240325 ps=1.715 w=0.74 l=0.15
X13 a_300_74.t1 CLK_N.t1 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1212 ps=1.1 w=0.74 l=0.15
X14 a_120_74.t1 D.t1 a_33_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X15 Q.t1 a_1934_94# VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.126075 ps=1.1 w=0.74 l=0.15
X16 VPWR.t7 RESET_B.t2 a_33_74.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1673 pd=1.475 as=0.063 ps=0.72 w=0.42 l=0.15
X17 VGND.t7 a_1266_119.t4 a_1934_94# VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X18 VGND.t2 RESET_B.t3 a_922_127.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.240325 pd=1.715 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 VPWR.t6 a_856_304# a_817_508.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X20 a_507_368.t0 a_300_74.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.4312 pd=3.01 as=0.3304 ps=2.83 w=1.12 l=0.15
X21 a_714_127.t2 RESET_B.t4 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.39 as=0.0756 ps=0.78 w=0.42 l=0.15
X22 Q.t0 a_1934_94# VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1862 ps=1.475 w=1.12 l=0.15
X23 a_1598_93.t1 a_1266_119.t5 a_1736_119.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X24 a_922_127.t1 a_856_304# a_850_127.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 a_817_508.t0 a_507_368.t5 a_714_127.t4 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X26 VGND.t6 a_1598_93.t2 a_1550_119.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_300_74.t5 a_300_74.t3 1086.11
R1 a_300_74.t0 a_300_74.n4 874.684
R2 a_300_74.t3 a_300_74.n0 642.616
R3 a_300_74.n1 a_300_74.t2 496.461
R4 a_300_74.n1 a_300_74.t5 483.608
R5 a_300_74.n3 a_300_74.t6 226.809
R6 a_300_74.n4 a_300_74.n3 207.504
R7 a_300_74.n4 a_300_74.t1 180.27
R8 a_300_74.n2 a_300_74.n1 178.048
R9 a_300_74.n2 a_300_74.t4 154.24
R10 a_300_74.n3 a_300_74.n2 2.19141
R11 a_33_74.n1 a_33_74.t0 729.749
R12 a_33_74.n2 a_33_74.n0 605.481
R13 a_33_74.n1 a_33_74.t4 395.825
R14 a_33_74.t2 a_33_74.n2 349.365
R15 a_33_74.n2 a_33_74.n1 118.947
R16 a_33_74.n0 a_33_74.t3 70.3576
R17 a_33_74.n0 a_33_74.t1 70.3576
R18 a_714_127.n3 a_714_127.t2 680.375
R19 a_714_127.n4 a_714_127.n0 616.615
R20 a_714_127.n5 a_714_127.n4 267.418
R21 a_714_127.n2 a_714_127.n1 217.023
R22 a_714_127.n3 a_714_127.n2 216.752
R23 a_714_127.n2 a_714_127.t5 162.274
R24 a_714_127.n5 a_714_127.t3 111.43
R25 a_714_127.n4 a_714_127.n3 75.2946
R26 a_714_127.n0 a_714_127.t4 70.3576
R27 a_714_127.n0 a_714_127.t0 70.3576
R28 a_714_127.t1 a_714_127.n5 40.0005
R29 VPB.n0 VPB 3534.41
R30 VPB VPB.n1 1660.57
R31 VPB.n0 VPB.t10 1098.12
R32 VPB.t4 VPB.t8 978.321
R33 VPB.t10 VPB.t5 753.361
R34 VPB.t1 VPB.t0 513.307
R35 VPB.n1 VPB.t1 390.726
R36 VPB.t6 VPB.t4 262.603
R37 VPB.t0 VPB.t7 257.93
R38 VPB.t3 VPB 255.376
R39 VPB.t2 VPB.t9 231.708
R40 VPB.t7 VPB.t3 229.839
R41 VPB.t9 VPB.t6 200.814
R42 VPB.n1 VPB.t2 172.494
R43 VPB.t8 VPB.n0 56.6401
R44 a_1266_119.n3 a_1266_119.n2 412.913
R45 a_1266_119.n6 a_1266_119.n5 412.283
R46 a_1266_119.n1 a_1266_119.t4 372.748
R47 a_1266_119.n3 a_1266_119.t3 217.436
R48 a_1266_119.n0 a_1266_119.t0 184.743
R49 a_1266_119.n5 a_1266_119.n4 155.357
R50 a_1266_119.n1 a_1266_119.t5 113.781
R51 a_1266_119.n0 a_1266_119.t2 100.29
R52 a_1266_119.n5 a_1266_119.n0 93.0189
R53 a_1266_119.n4 a_1266_119.n3 77.8012
R54 a_1266_119.n6 a_1266_119.t1 59.9403
R55 a_1266_119.n4 a_1266_119.n1 33.6491
R56 a_1266_119.n7 a_1266_119.n6 14.0719
R57 VNB.n0 VNB 15983.2
R58 VNB VNB.n1 7390.63
R59 VNB.t3 VNB.t1 2425.2
R60 VNB.t10 VNB.t11 2390.55
R61 VNB.t8 VNB.t13 2108.33
R62 VNB.n0 VNB.t15 1743.83
R63 VNB.n1 VNB.t3 1732.28
R64 VNB.t14 VNB.t2 1558.33
R65 VNB.t4 VNB.n0 1523.96
R66 VNB.t6 VNB.t0 1247.24
R67 VNB.t5 VNB 1212.6
R68 VNB.t11 VNB.t9 1177.95
R69 VNB.t1 VNB.t7 1177.95
R70 VNB.t13 VNB.t4 1008.33
R71 VNB.t0 VNB.t10 900.788
R72 VNB.t15 VNB.t6 900.788
R73 VNB.t7 VNB.t5 900.788
R74 VNB.t12 VNB.t8 825
R75 VNB.t2 VNB.t12 825
R76 VNB.n1 VNB.t14 618.75
R77 D.n1 D.t0 338.344
R78 D.n0 D.t1 164.173
R79 D.n0 D 156.107
R80 D.n2 D.n1 152
R81 D.n1 D.n0 49.6611
R82 D.n2 D 12.3175
R83 D D.n2 5.55522
R84 VPWR.n3 VPWR.t1 885.256
R85 VPWR.n13 VPWR.t5 685.053
R86 VPWR.n40 VPWR.t2 677.855
R87 VPWR.n27 VPWR.n7 607.497
R88 VPWR.n38 VPWR.n2 606.528
R89 VPWR.n12 VPWR.t4 363.771
R90 VPWR.n7 VPWR.t3 98.5005
R91 VPWR.n2 VPWR.t7 93.81
R92 VPWR.n7 VPWR.t6 70.3576
R93 VPWR.n2 VPWR.t0 48.7502
R94 VPWR.n31 VPWR.n5 36.1417
R95 VPWR.n32 VPWR.n31 36.1417
R96 VPWR.n33 VPWR.n32 36.1417
R97 VPWR.n19 VPWR.n18 36.1417
R98 VPWR.n20 VPWR.n19 36.1417
R99 VPWR.n20 VPWR.n9 36.1417
R100 VPWR.n24 VPWR.n9 36.1417
R101 VPWR.n26 VPWR.n25 33.8829
R102 VPWR.n14 VPWR.n11 30.8711
R103 VPWR.n37 VPWR.n3 29.3652
R104 VPWR.n27 VPWR.n5 28.6123
R105 VPWR.n39 VPWR.n38 25.6005
R106 VPWR.n14 VPWR.n13 24.8476
R107 VPWR.n38 VPWR.n37 21.8358
R108 VPWR.n40 VPWR.n39 21.0829
R109 VPWR.n27 VPWR.n26 18.824
R110 VPWR.n33 VPWR.n3 18.0711
R111 VPWR.n18 VPWR.n11 16.5652
R112 VPWR.n25 VPWR.n24 13.5534
R113 VPWR.n15 VPWR.n14 9.3005
R114 VPWR.n16 VPWR.n11 9.3005
R115 VPWR.n18 VPWR.n17 9.3005
R116 VPWR.n19 VPWR.n10 9.3005
R117 VPWR.n21 VPWR.n20 9.3005
R118 VPWR.n22 VPWR.n9 9.3005
R119 VPWR.n24 VPWR.n23 9.3005
R120 VPWR.n25 VPWR.n8 9.3005
R121 VPWR.n26 VPWR.n6 9.3005
R122 VPWR.n28 VPWR.n27 9.3005
R123 VPWR.n29 VPWR.n5 9.3005
R124 VPWR.n31 VPWR.n30 9.3005
R125 VPWR.n32 VPWR.n4 9.3005
R126 VPWR.n34 VPWR.n33 9.3005
R127 VPWR.n35 VPWR.n3 9.3005
R128 VPWR.n37 VPWR.n36 9.3005
R129 VPWR.n38 VPWR.n1 9.3005
R130 VPWR.n39 VPWR.n0 9.3005
R131 VPWR.n41 VPWR.n40 9.3005
R132 VPWR.n13 VPWR.n12 6.99826
R133 VPWR.n15 VPWR.n12 0.512215
R134 VPWR.n16 VPWR.n15 0.122949
R135 VPWR.n17 VPWR.n16 0.122949
R136 VPWR.n17 VPWR.n10 0.122949
R137 VPWR.n21 VPWR.n10 0.122949
R138 VPWR.n22 VPWR.n21 0.122949
R139 VPWR.n23 VPWR.n22 0.122949
R140 VPWR.n23 VPWR.n8 0.122949
R141 VPWR.n8 VPWR.n6 0.122949
R142 VPWR.n28 VPWR.n6 0.122949
R143 VPWR.n29 VPWR.n28 0.122949
R144 VPWR.n30 VPWR.n29 0.122949
R145 VPWR.n30 VPWR.n4 0.122949
R146 VPWR.n34 VPWR.n4 0.122949
R147 VPWR.n35 VPWR.n34 0.122949
R148 VPWR.n36 VPWR.n35 0.122949
R149 VPWR.n36 VPWR.n1 0.122949
R150 VPWR.n1 VPWR.n0 0.122949
R151 VPWR.n41 VPWR.n0 0.122949
R152 VPWR VPWR.n41 0.0617245
R153 a_507_368.t0 a_507_368.n3 801.462
R154 a_507_368.n3 a_507_368.t5 469.274
R155 a_507_368.n1 a_507_368.n0 404.274
R156 a_507_368.n0 a_507_368.t2 336.834
R157 a_507_368.n0 a_507_368.t4 231.23
R158 a_507_368.n2 a_507_368.t1 228.232
R159 a_507_368.n1 a_507_368.t3 199.113
R160 a_507_368.n2 a_507_368.n1 109.93
R161 a_507_368.n3 a_507_368.n2 21.4948
R162 a_1598_93.n2 a_1598_93.t0 671.455
R163 a_1598_93.n1 a_1598_93.t2 409.7
R164 a_1598_93.t1 a_1598_93.n2 349.065
R165 a_1598_93.n2 a_1598_93.n1 175.87
R166 a_1598_93.n1 a_1598_93.n0 150.492
R167 RESET_B.n4 RESET_B.t2 325.887
R168 RESET_B.n1 RESET_B.n0 295.091
R169 RESET_B.n2 RESET_B.t4 293.752
R170 RESET_B.n4 RESET_B.t0 271.527
R171 RESET_B.n1 RESET_B.t1 236.18
R172 RESET_B.n2 RESET_B.t3 224.934
R173 RESET_B.n3 RESET_B.n1 169.823
R174 RESET_B.n5 RESET_B.n4 167.999
R175 RESET_B.n3 RESET_B.n2 163.434
R176 RESET_B.n5 RESET_B.n3 3.32775
R177 RESET_B RESET_B.n5 0.0466957
R178 a_120_74.t0 a_120_74.t1 68.5719
R179 VGND.n1 VGND.t4 395.786
R180 VGND.n22 VGND.n21 230.579
R181 VGND.n35 VGND.n34 215.293
R182 VGND.n9 VGND.n8 206.528
R183 VGND.n11 VGND.n10 134.641
R184 VGND.n21 VGND.t8 131.141
R185 VGND.n34 VGND.t0 62.2404
R186 VGND.n21 VGND.t2 59.2552
R187 VGND.n8 VGND.t1 55.7148
R188 VGND.n8 VGND.t6 55.7148
R189 VGND.n10 VGND.t7 47.6797
R190 VGND.n14 VGND.n7 36.1417
R191 VGND.n15 VGND.n14 36.1417
R192 VGND.n16 VGND.n15 36.1417
R193 VGND.n16 VGND.n5 36.1417
R194 VGND.n20 VGND.n5 36.1417
R195 VGND.n23 VGND.n3 36.1417
R196 VGND.n27 VGND.n3 36.1417
R197 VGND.n28 VGND.n27 36.1417
R198 VGND.n29 VGND.n28 36.1417
R199 VGND.n23 VGND.n22 35.0123
R200 VGND.n35 VGND.n33 28.9887
R201 VGND.n33 VGND.n32 28.8587
R202 VGND.n29 VGND.n1 25.6758
R203 VGND.n34 VGND.t3 22.7037
R204 VGND.n10 VGND.t5 21.551
R205 VGND.n9 VGND.n7 14.6829
R206 VGND.n22 VGND.n20 12.424
R207 VGND.n33 VGND.n0 9.3005
R208 VGND.n32 VGND.n31 9.3005
R209 VGND.n30 VGND.n29 9.3005
R210 VGND.n28 VGND.n2 9.3005
R211 VGND.n27 VGND.n26 9.3005
R212 VGND.n25 VGND.n3 9.3005
R213 VGND.n24 VGND.n23 9.3005
R214 VGND.n22 VGND.n4 9.3005
R215 VGND.n20 VGND.n19 9.3005
R216 VGND.n18 VGND.n5 9.3005
R217 VGND.n17 VGND.n16 9.3005
R218 VGND.n15 VGND.n6 9.3005
R219 VGND.n14 VGND.n13 9.3005
R220 VGND.n12 VGND.n7 9.3005
R221 VGND.n36 VGND.n35 7.19068
R222 VGND.n11 VGND.n9 7.17529
R223 VGND.n32 VGND.n1 0.582318
R224 VGND VGND.n36 0.27524
R225 VGND.n12 VGND.n11 0.168522
R226 VGND.n36 VGND.n0 0.155562
R227 VGND.n13 VGND.n12 0.122949
R228 VGND.n13 VGND.n6 0.122949
R229 VGND.n17 VGND.n6 0.122949
R230 VGND.n18 VGND.n17 0.122949
R231 VGND.n19 VGND.n18 0.122949
R232 VGND.n19 VGND.n4 0.122949
R233 VGND.n24 VGND.n4 0.122949
R234 VGND.n25 VGND.n24 0.122949
R235 VGND.n26 VGND.n25 0.122949
R236 VGND.n26 VGND.n2 0.122949
R237 VGND.n30 VGND.n2 0.122949
R238 VGND.n31 VGND.n30 0.122949
R239 VGND.n31 VGND.n0 0.122949
R240 CLK_N.n0 CLK_N.t0 284.022
R241 CLK_N.n0 CLK_N.t1 176.643
R242 CLK_N CLK_N.n0 159.226
R243 a_1736_119.t0 a_1736_119.t1 68.5719
R244 a_850_127.t0 a_850_127.t1 60.0005
R245 a_1550_119.t0 a_1550_119.t1 68.5719
R246 Q.n1 Q 589.572
R247 Q.n1 Q.n0 585
R248 Q.n2 Q.n1 585
R249 Q Q.t1 194.948
R250 Q.n1 Q.t0 26.3844
R251 Q Q.n2 12.2519
R252 Q Q.n0 10.6062
R253 Q Q.n0 2.92621
R254 Q.n2 Q 1.2805
R255 a_922_127.t0 a_922_127.t1 60.0005
R256 a_817_508.t0 a_817_508.t1 112.572
C0 VPWR a_1934_94# 0.185841f
C1 VPWR D 0.035971f
C2 VGND VPB 0.011158f
C3 VGND a_1934_94# 0.118023f
C4 VPWR RESET_B 0.27413f
C5 VGND D 0.010616f
C6 Q VPB 0.015444f
C7 a_1547_508# RESET_B 0.001058f
C8 CLK_N VPWR 0.015318f
C9 Q a_1934_94# 0.076734f
C10 VGND RESET_B 0.275239f
C11 a_856_304# VPB 0.093787f
C12 CLK_N VGND 0.015894f
C13 Q RESET_B 1.2e-19
C14 VPWR a_1547_508# 0.004658f
C15 a_856_304# RESET_B 0.256952f
C16 VPWR VGND 0.057778f
C17 VPWR Q 0.108125f
C18 a_1934_94# VPB 0.054586f
C19 VPB D 0.102404f
C20 VGND Q 0.090062f
C21 VPWR a_856_304# 0.156998f
C22 a_856_304# a_1547_508# 3e-19
C23 VPB RESET_B 0.298499f
C24 CLK_N VPB 0.03608f
C25 VGND a_856_304# 0.022135f
C26 a_1934_94# RESET_B 0.001067f
C27 D RESET_B 0.107316f
C28 CLK_N RESET_B 0.094108f
C29 VPWR VPB 0.339811f
C30 Q VNB 0.10807f
C31 VGND VNB 1.29822f
C32 VPWR VNB 0.999716f
C33 CLK_N VNB 0.118448f
C34 RESET_B VNB 0.396022f
C35 D VNB 0.257672f
C36 VPB VNB 2.54229f
C37 a_1934_94# VNB 0.153078f
C38 a_856_304# VNB 0.121416f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxtp_1 VNB VPB VPWR VGND CLK Q D
X0 VPWR.t1 CLK.t0 a_27_74.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_668_503.t0 a_27_74.t2 a_561_463.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X2 Q.t0 a_1210_314.t2 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X3 a_454_503.t1 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X4 VPWR.t6 a_1011_424.t4 a_1210_314.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 VGND.t1 CLK.t1 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_1118_508# a_206_368.t2 a_1011_424.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X7 a_713_458.t0 a_561_463.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X8 VGND.t5 a_713_458.t4 a_731_101.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_561_463.t2 a_206_368.t3 a_454_503.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X10 a_206_368.t1 a_27_74.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_1011_424.t1 a_27_74.t4 a_713_458.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X12 a_1168_124.t0 a_27_74.t5 a_1011_424.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X13 Q.t1 a_1210_314.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X14 a_713_458.t1 a_561_463.t5 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X15 a_561_463.t0 a_27_74.t6 a_454_503.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.155625 ps=1.215 w=0.42 l=0.15
X16 VPWR.t4 a_713_458.t5 a_668_503.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X17 VGND.t6 a_1011_424.t5 a_1210_314.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X18 a_206_368.t0 a_27_74.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X19 a_731_101.t1 a_206_368.t4 a_561_463.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X20 a_1011_424.t3 a_206_368.t5 a_713_458.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X21 a_454_503.t2 D.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.155625 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
R0 CLK.n0 CLK.t0 259.132
R1 CLK.n0 CLK.t1 198.882
R2 CLK CLK.n0 156.934
R3 a_27_74.t5 a_27_74.t4 733.712
R4 a_27_74.n1 a_27_74.t5 449.469
R5 a_27_74.n0 a_27_74.t6 315.515
R6 a_27_74.n2 a_27_74.n1 303.166
R7 a_27_74.t1 a_27_74.n4 290.298
R8 a_27_74.n3 a_27_74.t3 282.276
R9 a_27_74.n1 a_27_74.n0 236.078
R10 a_27_74.n0 a_27_74.t2 209.476
R11 a_27_74.n3 a_27_74.t7 174.898
R12 a_27_74.n2 a_27_74.t0 172.839
R13 a_27_74.n4 a_27_74.n3 152
R14 a_27_74.n4 a_27_74.n2 9.46137
R15 VPWR.n2 VPWR.t0 840.035
R16 VPWR.n6 VPWR.n5 659.098
R17 VPWR.n8 VPWR.n7 333.757
R18 VPWR.n18 VPWR.n1 331.5
R19 VPWR.n5 VPWR.t4 131.333
R20 VPWR.n5 VPWR.t3 45.4599
R21 VPWR.n7 VPWR.t5 43.8979
R22 VPWR.n11 VPWR.n4 36.1417
R23 VPWR.n12 VPWR.n11 36.1417
R24 VPWR.n13 VPWR.n12 36.1417
R25 VPWR.n18 VPWR.n17 35.3887
R26 VPWR.n7 VPWR.t6 35.1791
R27 VPWR.n17 VPWR.n16 31.2225
R28 VPWR.n1 VPWR.t2 26.3844
R29 VPWR.n1 VPWR.t1 26.3844
R30 VPWR.n13 VPWR.n2 23.6596
R31 VPWR.n6 VPWR.n4 19.7527
R32 VPWR.n8 VPWR.n6 10.8455
R33 VPWR.n9 VPWR.n4 9.3005
R34 VPWR.n11 VPWR.n10 9.3005
R35 VPWR.n12 VPWR.n3 9.3005
R36 VPWR.n14 VPWR.n13 9.3005
R37 VPWR.n16 VPWR.n15 9.3005
R38 VPWR.n17 VPWR.n0 9.3005
R39 VPWR.n19 VPWR.n18 8.45673
R40 VPWR.n16 VPWR.n2 1.70717
R41 VPWR VPWR.n19 0.163644
R42 VPWR.n9 VPWR.n8 0.150798
R43 VPWR.n19 VPWR.n0 0.144205
R44 VPWR.n10 VPWR.n9 0.122949
R45 VPWR.n10 VPWR.n3 0.122949
R46 VPWR.n14 VPWR.n3 0.122949
R47 VPWR.n15 VPWR.n14 0.122949
R48 VPWR.n15 VPWR.n0 0.122949
R49 VPB.t7 VPB.t10 835.082
R50 VPB.t3 VPB.t0 633.333
R51 VPB.t6 VPB.t2 360.082
R52 VPB.t8 VPB.t6 316.668
R53 VPB.t2 VPB.t7 273.253
R54 VPB.t5 VPB.t4 273.253
R55 VPB.t0 VPB.t5 273.253
R56 VPB.t10 VPB.t9 257.93
R57 VPB VPB.t1 257.93
R58 VPB.t1 VPB.t3 229.839
R59 VPB.t4 VPB.t8 199.195
R60 a_561_463.n2 a_561_463.n1 589.926
R61 a_561_463.n0 a_561_463.t4 380.639
R62 a_561_463.n3 a_561_463.n2 300.101
R63 a_561_463.n2 a_561_463.n0 260.5
R64 a_561_463.n0 a_561_463.t5 203.294
R65 a_561_463.n1 a_561_463.t1 157.345
R66 a_561_463.n1 a_561_463.t2 68.0124
R67 a_561_463.n3 a_561_463.t3 57.7148
R68 a_561_463.n5 a_561_463.n4 28.8005
R69 a_561_463.n4 a_561_463.t0 23.1765
R70 a_561_463.n4 a_561_463.n3 8.0005
R71 a_668_503.t0 a_668_503.t1 112.572
R72 a_1210_314.t0 a_1210_314.n5 401.988
R73 a_1210_314.n4 a_1210_314.t1 288.435
R74 a_1210_314.n2 a_1210_314.n1 282.675
R75 a_1210_314.n3 a_1210_314.t2 250.909
R76 a_1210_314.n3 a_1210_314.t3 220.113
R77 a_1210_314.n2 a_1210_314.n0 198.083
R78 a_1210_314.n4 a_1210_314.n3 152
R79 a_1210_314.n5 a_1210_314.n2 97.1059
R80 a_1210_314.n5 a_1210_314.n4 36.7273
R81 Q.n0 Q.t0 305.339
R82 Q.t1 Q.n0 279.738
R83 Q.n1 Q.t1 279.738
R84 Q.n1 Q 11.5561
R85 Q.n0 Q 4.44494
R86 Q Q.n1 1.6005
R87 D D.t1 355.692
R88 D.n0 D.t0 291.063
R89 D.n0 D 3.42907
R90 D D.n0 2.52682
R91 a_454_503.n1 a_454_503.n0 918.856
R92 a_454_503.n0 a_454_503.t1 155
R93 a_454_503.t0 a_454_503.n1 72.8576
R94 a_454_503.n1 a_454_503.t2 71.2386
R95 a_454_503.n0 a_454_503.t3 70.3576
R96 a_1011_424.n3 a_1011_424.n2 695.769
R97 a_1011_424.n1 a_1011_424.t4 246.456
R98 a_1011_424.n2 a_1011_424.n1 244.236
R99 a_1011_424.n2 a_1011_424.n0 218.673
R100 a_1011_424.n1 a_1011_424.t5 182.481
R101 a_1011_424.n3 a_1011_424.t2 112.572
R102 a_1011_424.n0 a_1011_424.t0 70.0005
R103 a_1011_424.n0 a_1011_424.t3 56.4605
R104 a_1011_424.t1 a_1011_424.n3 34.0065
R105 VGND.n1 VGND.t3 315.938
R106 VGND.n17 VGND.n16 214.185
R107 VGND.n6 VGND.n5 212.548
R108 VGND.n4 VGND.n3 211.452
R109 VGND.n3 VGND.t0 67.6369
R110 VGND.n16 VGND.t2 53.514
R111 VGND.n3 VGND.t5 53.0654
R112 VGND.n9 VGND.n8 36.1417
R113 VGND.n10 VGND.n9 36.1417
R114 VGND.n15 VGND.n14 36.1417
R115 VGND.n8 VGND.n4 35.3887
R116 VGND.n5 VGND.t6 31.8755
R117 VGND.n17 VGND.n15 30.4946
R118 VGND.n5 VGND.t4 29.2236
R119 VGND.n10 VGND.n1 24.4711
R120 VGND.n14 VGND.n1 22.9652
R121 VGND.n16 VGND.t1 22.7032
R122 VGND.n15 VGND.n0 9.3005
R123 VGND.n14 VGND.n13 9.3005
R124 VGND.n12 VGND.n1 9.3005
R125 VGND.n11 VGND.n10 9.3005
R126 VGND.n9 VGND.n2 9.3005
R127 VGND.n8 VGND.n7 9.3005
R128 VGND.n18 VGND.n17 7.19894
R129 VGND.n6 VGND.n4 6.8022
R130 VGND.n7 VGND.n6 0.163018
R131 VGND VGND.n18 0.156997
R132 VGND.n18 VGND.n0 0.150766
R133 VGND.n7 VGND.n2 0.122949
R134 VGND.n11 VGND.n2 0.122949
R135 VGND.n12 VGND.n11 0.122949
R136 VGND.n13 VGND.n12 0.122949
R137 VGND.n13 VGND.n0 0.122949
R138 VNB.t4 VNB.t10 3245.14
R139 VNB.t2 VNB.t5 3071.92
R140 VNB.t8 VNB.t0 1570.6
R141 VNB.t5 VNB.t3 1524.41
R142 VNB.t9 VNB.t4 1466.67
R143 VNB.t1 VNB.t2 1432.02
R144 VNB.t0 VNB.t9 1177.95
R145 VNB.t10 VNB.t6 1143.31
R146 VNB VNB.t1 1143.31
R147 VNB.t3 VNB.t7 1097.11
R148 VNB.t7 VNB.t8 831.496
R149 a_206_368.n0 a_206_368.t4 1132.7
R150 a_206_368.n0 a_206_368.t3 541.106
R151 a_206_368.n2 a_206_368.t5 412.152
R152 a_206_368.n2 a_206_368.t2 372.413
R153 a_206_368.n3 a_206_368.n2 264.704
R154 a_206_368.n1 a_206_368.t0 258.969
R155 a_206_368.t1 a_206_368.n3 217.333
R156 a_206_368.n1 a_206_368.n0 152
R157 a_206_368.n3 a_206_368.n1 30.1502
R158 a_713_458.n3 a_713_458.n2 662.327
R159 a_713_458.n1 a_713_458.t5 478.647
R160 a_713_458.n2 a_713_458.n0 230.298
R161 a_713_458.n2 a_713_458.n1 177.44
R162 a_713_458.n1 a_713_458.t4 139.028
R163 a_713_458.n3 a_713_458.t2 92.6374
R164 a_713_458.n0 a_713_458.t0 49.4918
R165 a_713_458.t1 a_713_458.n3 37.5243
R166 a_713_458.n0 a_713_458.t3 24.2336
R167 a_731_101.t0 a_731_101.t1 60.0005
C0 VPWR VGND 0.127399f
C1 VGND Q 0.068667f
C2 CLK VGND 0.017148f
C3 D VGND 0.009382f
C4 a_1118_508# VPWR 0.005135f
C5 a_1118_508# VGND 4.56e-19
C6 VPB VPWR 0.240274f
C7 VPB Q 0.013643f
C8 VPB CLK 0.0398f
C9 VPWR Q 0.119773f
C10 VPWR CLK 0.015092f
C11 VPB D 0.098179f
C12 VPWR D 0.01058f
C13 VPB VGND 0.01901f
C14 Q VNB 0.111234f
C15 VGND VNB 0.949043f
C16 D VNB 0.129717f
C17 CLK VNB 0.163617f
C18 VPWR VNB 0.755441f
C19 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxtp_2 VNB VPB VPWR VGND Q CLK D
X0 a_431_508.t1 D.t0 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.318675 ps=2.49 w=0.42 l=0.15
X1 VPWR.t5 CLK.t0 a_27_74.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t4 a_1217_314# Q.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_1019_424.t2 a_27_74.t2 a_695_459.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1407 pd=1.22 as=0.2625 ps=1.465 w=0.84 l=0.15
X4 Q.t2 a_1217_314# VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1934 ps=1.475 w=1.12 l=0.15
X5 a_206_368.t0 a_27_74.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2775 pd=2.23 as=0.1628 ps=1.18 w=0.74 l=0.15
X6 a_644_504.t0 a_27_74.t4 a_538_429.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1126 ps=1.175 w=0.42 l=0.15
X7 VGND.t5 a_1217_314# a_1172_124.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X8 a_538_429.t3 a_27_74.t5 a_431_508.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.076125 pd=0.835 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND.t0 CLK.t1 a_27_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 a_1172_124.t1 a_27_74.t6 a_1019_424.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.122775 ps=1.175 w=0.42 l=0.15
X11 VGND.t2 a_695_459.t4 a_708_101.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2088 pd=1.405 as=0.0504 ps=0.66 w=0.42 l=0.15
X12 a_1125_508.t0 a_206_368.t2 a_1019_424.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1407 ps=1.22 w=0.42 l=0.15
X13 VGND.t4 a_1217_314# Q.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_1019_424.t0 a_206_368.t3 a_695_459.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.122775 pd=1.175 as=0.077 ps=0.83 w=0.55 l=0.15
X15 a_206_368.t1 a_27_74.t7 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_708_101.t0 a_206_368.t4 a_538_429.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.076125 ps=0.835 w=0.42 l=0.15
X17 a_695_459.t0 a_538_429.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2625 pd=1.465 as=0.209825 ps=1.605 w=0.84 l=0.15
X18 a_431_508.t2 D.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1154 pd=1.2 as=0.2474 ps=2.13 w=0.42 l=0.15
X19 a_538_429.t1 a_206_368.t5 a_431_508.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1126 pd=1.175 as=0.1154 ps=1.2 w=0.42 l=0.15
X20 VPWR.t0 a_695_459.t5 a_644_504.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.209825 pd=1.605 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR.t2 a_1217_314# a_1125_508.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.09975 ps=0.895 w=0.42 l=0.15
X22 Q.t0 a_1217_314# VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1405 ps=1.14 w=0.74 l=0.15
X23 VGND.t8 a_1019_424.t4 a_1217_314# VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1405 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X24 a_695_459.t3 a_538_429.t5 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.2088 ps=1.405 w=0.55 l=0.15
R0 D.n0 D.t0 360.868
R1 D.n0 D.t1 348.827
R2 D D.n0 3.44665
R3 VGND.n1 VGND.t6 377.608
R4 VGND.n12 VGND.t5 257.195
R5 VGND.n31 VGND.n30 214.185
R6 VGND.n4 VGND.n3 211.452
R7 VGND.n10 VGND.n9 207.346
R8 VGND.n8 VGND.t4 178.799
R9 VGND.n3 VGND.t7 102.546
R10 VGND.n3 VGND.t2 53.0654
R11 VGND.n30 VGND.t1 48.6491
R12 VGND.n9 VGND.t3 40.4736
R13 VGND.n16 VGND.n6 36.1417
R14 VGND.n17 VGND.n16 36.1417
R15 VGND.n18 VGND.n17 36.1417
R16 VGND.n23 VGND.n22 36.1417
R17 VGND.n24 VGND.n23 36.1417
R18 VGND.n29 VGND.n28 36.1417
R19 VGND.n24 VGND.n1 34.6358
R20 VGND.n9 VGND.t8 30.938
R21 VGND.n12 VGND.n11 30.4946
R22 VGND.n31 VGND.n29 30.4946
R23 VGND.n22 VGND.n4 28.9887
R24 VGND.n11 VGND.n10 25.6005
R25 VGND.n18 VGND.n4 24.4711
R26 VGND.n28 VGND.n1 22.9652
R27 VGND.n30 VGND.t0 22.7032
R28 VGND.n12 VGND.n6 16.9417
R29 VGND.n29 VGND.n0 9.3005
R30 VGND.n28 VGND.n27 9.3005
R31 VGND.n26 VGND.n1 9.3005
R32 VGND.n25 VGND.n24 9.3005
R33 VGND.n23 VGND.n2 9.3005
R34 VGND.n22 VGND.n21 9.3005
R35 VGND.n20 VGND.n4 9.3005
R36 VGND.n19 VGND.n18 9.3005
R37 VGND.n17 VGND.n5 9.3005
R38 VGND.n16 VGND.n15 9.3005
R39 VGND.n14 VGND.n6 9.3005
R40 VGND.n11 VGND.n7 9.3005
R41 VGND.n13 VGND.n12 9.3005
R42 VGND.n32 VGND.n31 7.19894
R43 VGND.n10 VGND.n8 6.74444
R44 VGND.n8 VGND.n7 0.585372
R45 VGND VGND.n32 0.156997
R46 VGND.n32 VGND.n0 0.150766
R47 VGND.n13 VGND.n7 0.122949
R48 VGND.n14 VGND.n13 0.122949
R49 VGND.n15 VGND.n14 0.122949
R50 VGND.n15 VGND.n5 0.122949
R51 VGND.n19 VGND.n5 0.122949
R52 VGND.n20 VGND.n19 0.122949
R53 VGND.n21 VGND.n20 0.122949
R54 VGND.n21 VGND.n2 0.122949
R55 VGND.n25 VGND.n2 0.122949
R56 VGND.n26 VGND.n25 0.122949
R57 VGND.n27 VGND.n26 0.122949
R58 VGND.n27 VGND.n0 0.122949
R59 a_431_508.n0 a_431_508.t2 948.65
R60 a_431_508.n1 a_431_508.n0 862.327
R61 a_431_508.n0 a_431_508.t3 70.3576
R62 a_431_508.t0 a_431_508.n1 40.0005
R63 a_431_508.n1 a_431_508.t1 40.0005
R64 VNB.t2 VNB.t9 3406.82
R65 VNB.t6 VNB.t11 2286.61
R66 VNB.t3 VNB.t10 1940.16
R67 VNB.t7 VNB.t12 1524.41
R68 VNB.t0 VNB.t2 1362.73
R69 VNB.t11 VNB.t4 1270.34
R70 VNB VNB.t0 1143.31
R71 VNB.t1 VNB.t8 1097.11
R72 VNB.t4 VNB.t5 993.177
R73 VNB.t10 VNB.t7 993.177
R74 VNB.t9 VNB.t1 993.177
R75 VNB.t12 VNB.t6 900.788
R76 VNB.t8 VNB.t3 900.788
R77 CLK.n0 CLK.t0 259.132
R78 CLK.n0 CLK.t1 198.882
R79 CLK CLK.n0 156.934
R80 a_27_74.t6 a_27_74.t2 733.842
R81 a_27_74.n1 a_27_74.t6 449.469
R82 a_27_74.n0 a_27_74.t5 393.769
R83 a_27_74.n2 a_27_74.n1 317.849
R84 a_27_74.t1 a_27_74.n4 290.298
R85 a_27_74.n3 a_27_74.t7 284.022
R86 a_27_74.n1 a_27_74.n0 235.953
R87 a_27_74.n0 a_27_74.t4 207.144
R88 a_27_74.n3 a_27_74.t3 176.643
R89 a_27_74.n2 a_27_74.t0 172.839
R90 a_27_74.n4 a_27_74.n3 152
R91 a_27_74.n4 a_27_74.n2 9.46137
R92 VPWR.n2 VPWR.t6 757.668
R93 VPWR.n12 VPWR.t2 677.855
R94 VPWR.n20 VPWR.n19 635.658
R95 VPWR.n8 VPWR.t3 360.286
R96 VPWR.n32 VPWR.n1 331.5
R97 VPWR.n9 VPWR.t4 266.226
R98 VPWR.n19 VPWR.t0 120.567
R99 VPWR.n19 VPWR.t1 89.8658
R100 VPWR.n25 VPWR.n4 36.1417
R101 VPWR.n26 VPWR.n25 36.1417
R102 VPWR.n27 VPWR.n26 36.1417
R103 VPWR.n13 VPWR.n6 36.1417
R104 VPWR.n17 VPWR.n6 36.1417
R105 VPWR.n18 VPWR.n17 36.1417
R106 VPWR.n32 VPWR.n31 35.3887
R107 VPWR.n21 VPWR.n18 35.2047
R108 VPWR.n31 VPWR.n30 31.2225
R109 VPWR.n12 VPWR.n11 29.7417
R110 VPWR.n1 VPWR.t7 26.3844
R111 VPWR.n1 VPWR.t5 26.3844
R112 VPWR.n27 VPWR.n2 22.0617
R113 VPWR.n11 VPWR.n8 21.0829
R114 VPWR.n13 VPWR.n12 17.6946
R115 VPWR.n20 VPWR.n4 13.8295
R116 VPWR.n11 VPWR.n10 9.3005
R117 VPWR.n12 VPWR.n7 9.3005
R118 VPWR.n14 VPWR.n13 9.3005
R119 VPWR.n15 VPWR.n6 9.3005
R120 VPWR.n17 VPWR.n16 9.3005
R121 VPWR.n18 VPWR.n5 9.3005
R122 VPWR.n22 VPWR.n21 9.3005
R123 VPWR.n23 VPWR.n4 9.3005
R124 VPWR.n25 VPWR.n24 9.3005
R125 VPWR.n26 VPWR.n3 9.3005
R126 VPWR.n28 VPWR.n27 9.3005
R127 VPWR.n30 VPWR.n29 9.3005
R128 VPWR.n31 VPWR.n0 9.3005
R129 VPWR.n33 VPWR.n32 8.45673
R130 VPWR.n9 VPWR.n8 6.8559
R131 VPWR.n21 VPWR.n20 4.97828
R132 VPWR.n30 VPWR.n2 2.13383
R133 VPWR.n10 VPWR.n9 0.565232
R134 VPWR VPWR.n33 0.163644
R135 VPWR.n33 VPWR.n0 0.144205
R136 VPWR.n10 VPWR.n7 0.122949
R137 VPWR.n14 VPWR.n7 0.122949
R138 VPWR.n15 VPWR.n14 0.122949
R139 VPWR.n16 VPWR.n15 0.122949
R140 VPWR.n16 VPWR.n5 0.122949
R141 VPWR.n22 VPWR.n5 0.122949
R142 VPWR.n23 VPWR.n22 0.122949
R143 VPWR.n24 VPWR.n23 0.122949
R144 VPWR.n24 VPWR.n3 0.122949
R145 VPWR.n28 VPWR.n3 0.122949
R146 VPWR.n29 VPWR.n28 0.122949
R147 VPWR.n29 VPWR.n0 0.122949
R148 VPB.t2 VPB.t3 771.237
R149 VPB.t8 VPB.t6 574.597
R150 VPB.t1 VPB.t10 395.834
R151 VPB.t0 VPB.t1 347.312
R152 VPB.t11 VPB.t2 319.221
R153 VPB.t6 VPB.t7 273.253
R154 VPB.t10 VPB.t11 270.7
R155 VPB.t7 VPB.t9 270.7
R156 VPB VPB.t5 257.93
R157 VPB.t3 VPB.t4 229.839
R158 VPB.t5 VPB.t8 229.839
R159 VPB.t9 VPB.t0 214.517
R160 Q Q.n0 589.444
R161 Q.n3 Q.n0 585
R162 Q.n2 Q.n0 585
R163 Q.n2 Q.n1 174.262
R164 Q.n0 Q.t3 26.3844
R165 Q.n0 Q.t2 26.3844
R166 Q.n1 Q.t1 22.7032
R167 Q.n1 Q.t0 22.7032
R168 Q Q.n3 7.64494
R169 Q Q.n2 6.57828
R170 Q.n3 Q 5.51161
R171 a_695_459.n3 a_695_459.n2 644.582
R172 a_695_459.n1 a_695_459.t5 518.953
R173 a_695_459.n2 a_695_459.n0 214.567
R174 a_695_459.n2 a_695_459.n1 187.876
R175 a_695_459.n1 a_695_459.t4 161.738
R176 a_695_459.n3 a_695_459.t2 110.227
R177 a_695_459.t0 a_695_459.n3 36.3517
R178 a_695_459.n0 a_695_459.t1 30.546
R179 a_695_459.n0 a_695_459.t3 30.546
R180 a_1019_424.n4 a_1019_424.n3 688.992
R181 a_1019_424.n2 a_1019_424.n1 272.464
R182 a_1019_424.n3 a_1019_424.n2 251.766
R183 a_1019_424.n3 a_1019_424.n0 215.675
R184 a_1019_424.n2 a_1019_424.t4 182.758
R185 a_1019_424.n4 a_1019_424.t3 110.227
R186 a_1019_424.n0 a_1019_424.t0 92.1913
R187 a_1019_424.n0 a_1019_424.t1 73.0918
R188 a_1019_424.t2 a_1019_424.n4 34.0065
R189 a_206_368.n0 a_206_368.t4 1093.74
R190 a_206_368.n0 a_206_368.t5 452.545
R191 a_206_368.n2 a_206_368.t3 435.118
R192 a_206_368.n2 a_206_368.t2 372.036
R193 a_206_368.n1 a_206_368.t0 264.344
R194 a_206_368.n3 a_206_368.n2 256.623
R195 a_206_368.t1 a_206_368.n3 217.333
R196 a_206_368.n1 a_206_368.n0 152
R197 a_206_368.n3 a_206_368.n1 24.1499
R198 a_538_429.n2 a_538_429.n1 588.587
R199 a_538_429.n1 a_538_429.t2 539.356
R200 a_538_429.n0 a_538_429.t5 338.861
R201 a_538_429.n3 a_538_429.n2 298.74
R202 a_538_429.n2 a_538_429.n0 269
R203 a_538_429.n0 a_538_429.t4 183.161
R204 a_538_429.n1 a_538_429.t1 68.0124
R205 a_538_429.n3 a_538_429.t3 48.4421
R206 a_538_429.n4 a_538_429.t0 25.4063
R207 a_538_429.n5 a_538_429.n4 21.6005
R208 a_538_429.n4 a_538_429.n3 14.546
R209 a_644_504.t0 a_644_504.t1 126.644
R210 a_1172_124.t0 a_1172_124.t1 68.5719
R211 a_708_101.t0 a_708_101.t1 68.5719
R212 a_1125_508.t0 a_1125_508.t1 222.798
C0 VGND Q 0.132986f
C1 VPB a_1217_314# 0.212825f
C2 VPB VPWR 0.256487f
C3 VPWR a_1217_314# 0.233601f
C4 VPB CLK 0.0398f
C5 VPB D 0.103618f
C6 VPWR CLK 0.015092f
C7 VPWR D 0.013266f
C8 VPB VGND 0.019699f
C9 VGND a_1217_314# 0.203521f
C10 VPB Q 0.005761f
C11 VPWR VGND 0.146695f
C12 Q a_1217_314# 0.161821f
C13 VPWR Q 0.217363f
C14 CLK VGND 0.017147f
C15 D VGND 0.007245f
C16 Q VNB 0.029895f
C17 VGND VNB 1.03587f
C18 D VNB 0.135431f
C19 CLK VNB 0.163339f
C20 VPWR VNB 0.839266f
C21 VPB VNB 2.01326f
C22 a_1217_314# VNB 0.374141f
.ends

* NGSPICE file created from sky130_fd_sc_hs__diode_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__diode_2 DIODE VNB VPB VPWR VGND
X0 VNB.t0 DIODE.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=3.24e+06 area=6.417e+11
R0 DIODE.n1 DIODE.t0 92.5005
R1 DIODE.t0 DIODE.n0 45.0815
R2 DIODE.n1 DIODE 4.73816
R3 DIODE.n0 DIODE 3.45585
R4 DIODE.n0 DIODE 2.55298
R5 DIODE DIODE.n1 1.41349
R6 VNB VNB.t0 2577.61
C0 DIODE VPB 0.057788f
C1 DIODE VPWR 0.107207f
C2 VPWR VPB 0.026311f
C3 DIODE VGND 0.107207f
C4 VPB VGND 0.003242f
C5 VPWR VGND 0.015199f
C6 VGND VNB 0.155443f
C7 VPWR VNB 0.132374f
C8 DIODE VNB 0.231428f
C9 VPB VNB 0.299088f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlclkp_1 VNB VPB VPWR VGND GCLK GATE CLK
X0 a_258_392.t0 GATE.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2959 ps=1.68 w=1 l=0.15
X1 VPWR.t2 a_83_260.t4 a_27_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2959 pd=1.68 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t3 a_27_74.t2 a_484_508.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.149975 pd=1.365 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_484_508.t1 a_315_54.t2 a_83_260.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.19445 ps=1.56 w=0.42 l=0.15
X4 GCLK.t1 a_987_393.t3 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5 VGND.t5 a_27_74.t3 a_477_124.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.141875 pd=1.23 as=0.0504 ps=0.66 w=0.42 l=0.15
X6 a_309_338.t0 a_315_54.t3 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.149975 ps=1.365 w=0.84 l=0.15
X7 VPWR.t4 CLK.t0 a_315_54.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.23 as=0.2478 ps=2.27 w=0.84 l=0.15
X8 a_987_393.t0 a_27_74.t4 a_984_125.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0768 ps=0.88 w=0.64 l=0.15
X9 VGND.t1 a_83_260.t5 a_27_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.219725 pd=1.415 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 a_83_260.t0 a_315_54.t4 a_267_80.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1346 pd=1.15 as=0.0768 ps=0.88 w=0.64 l=0.15
X11 a_477_124.t0 a_309_338.t2 a_83_260.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1346 ps=1.15 w=0.42 l=0.15
X12 VGND.t3 CLK.t1 a_315_54.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.2183 ps=2.07 w=0.74 l=0.15
X13 a_987_393.t2 CLK.t2 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.15 as=0.1638 ps=1.23 w=0.84 l=0.15
X14 a_984_125.t0 CLK.t3 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.12945 ps=1.1 w=0.64 l=0.15
X15 GCLK.t0 a_987_393.t4 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3318 ps=1.795 w=1.12 l=0.15
X16 VPWR.t1 a_27_74.t5 a_987_393.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3318 pd=1.795 as=0.1302 ps=1.15 w=0.84 l=0.15
X17 a_267_80.t1 GATE.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.219725 ps=1.415 w=0.64 l=0.15
X18 a_309_338.t1 a_315_54.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.141875 ps=1.23 w=0.74 l=0.15
X19 a_83_260.t2 a_309_338.t3 a_258_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.19445 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
R0 GATE.n0 GATE.t1 265.101
R1 GATE.n0 GATE.t0 231.629
R2 GATE GATE.n0 154.133
R3 VPWR.n13 VPWR.n4 604.976
R4 VPWR.n8 VPWR.n7 323.447
R5 VPWR.n20 VPWR.n1 315.736
R6 VPWR.n9 VPWR.n6 227.614
R7 VPWR.n6 VPWR.t1 113.403
R8 VPWR.n4 VPWR.t7 99.5923
R9 VPWR.n4 VPWR.t3 77.1507
R10 VPWR.n1 VPWR.t0 70.9205
R11 VPWR.n7 VPWR.t4 46.9053
R12 VPWR.n7 VPWR.t6 44.56
R13 VPWR.n1 VPWR.t2 37.541
R14 VPWR.n14 VPWR.n2 36.1417
R15 VPWR.n18 VPWR.n2 36.1417
R16 VPWR.n19 VPWR.n18 36.1417
R17 VPWR.n12 VPWR.n5 36.1417
R18 VPWR.n6 VPWR.t5 34.3894
R19 VPWR.n13 VPWR.n12 32.7534
R20 VPWR.n8 VPWR.n5 26.3534
R21 VPWR.n20 VPWR.n19 19.2005
R22 VPWR.n14 VPWR.n13 14.6829
R23 VPWR.n10 VPWR.n5 9.3005
R24 VPWR.n12 VPWR.n11 9.3005
R25 VPWR.n13 VPWR.n3 9.3005
R26 VPWR.n15 VPWR.n14 9.3005
R27 VPWR.n16 VPWR.n2 9.3005
R28 VPWR.n18 VPWR.n17 9.3005
R29 VPWR.n19 VPWR.n0 9.3005
R30 VPWR.n21 VPWR.n20 7.43488
R31 VPWR.n9 VPWR.n8 6.8968
R32 VPWR.n10 VPWR.n9 0.260241
R33 VPWR VPWR.n21 0.160103
R34 VPWR.n21 VPWR.n0 0.1477
R35 VPWR.n11 VPWR.n10 0.122949
R36 VPWR.n11 VPWR.n3 0.122949
R37 VPWR.n15 VPWR.n3 0.122949
R38 VPWR.n16 VPWR.n15 0.122949
R39 VPWR.n17 VPWR.n16 0.122949
R40 VPWR.n17 VPWR.n0 0.122949
R41 a_258_392.t0 a_258_392.t1 53.1905
R42 VPB.n0 VPB 2571.64
R43 VPB VPB.n1 1461.96
R44 VPB.t9 VPB.t5 553.027
R45 VPB.t1 VPB.t6 421.372
R46 VPB.t8 VPB.t3 362.635
R47 VPB.t0 VPB.t2 362.635
R48 VPB.t4 VPB.t9 298.416
R49 VPB.t5 VPB.t7 295.678
R50 VPB.t2 VPB 257.93
R51 VPB.t3 VPB.t0 214.517
R52 VPB.n1 VPB.t8 165.995
R53 VPB.n0 VPB.t1 145.565
R54 VPB.t7 VPB.n0 95.8218
R55 VPB.n1 VPB.t4 52.0178
R56 a_83_260.n3 a_83_260.n2 725.652
R57 a_83_260.n2 a_83_260.n0 280.087
R58 a_83_260.n1 a_83_260.t4 262.921
R59 a_83_260.n1 a_83_260.t5 202.671
R60 a_83_260.n2 a_83_260.n1 152
R61 a_83_260.n3 a_83_260.t3 131.333
R62 a_83_260.t2 a_83_260.n3 95.9676
R63 a_83_260.n0 a_83_260.t1 72.8576
R64 a_83_260.n0 a_83_260.t0 60.5809
R65 a_27_74.n0 a_27_74.t4 978.461
R66 a_27_74.t3 a_27_74.t2 567.616
R67 a_27_74.t4 a_27_74.t5 422.019
R68 a_27_74.n1 a_27_74.n0 353.58
R69 a_27_74.t0 a_27_74.n1 295.24
R70 a_27_74.n1 a_27_74.t1 142.268
R71 a_27_74.n0 a_27_74.t3 126.927
R72 a_484_508.t0 a_484_508.t1 126.644
R73 a_315_54.t1 a_315_54.n3 776.162
R74 a_315_54.t1 a_315_54.n4 768.644
R75 a_315_54.n1 a_315_54.t4 368.375
R76 a_315_54.n4 a_315_54.t0 318.923
R77 a_315_54.n1 a_315_54.t2 290.442
R78 a_315_54.n0 a_315_54.t3 205.922
R79 a_315_54.n0 a_315_54.t5 186.374
R80 a_315_54.n2 a_315_54.n0 173.78
R81 a_315_54.n3 a_315_54.n2 63.2476
R82 a_315_54.n2 a_315_54.n1 31.6126
R83 a_315_54.n4 a_315_54.n3 14.8322
R84 a_987_393.n2 a_987_393.n1 342.396
R85 a_987_393.n0 a_987_393.t4 240.197
R86 a_987_393.n1 a_987_393.n0 206.906
R87 a_987_393.n0 a_987_393.t3 194.304
R88 a_987_393.n1 a_987_393.t0 139.819
R89 a_987_393.n2 a_987_393.t2 37.5243
R90 a_987_393.t1 a_987_393.n2 35.1791
R91 VGND.n11 VGND.n3 240.161
R92 VGND.n20 VGND.n19 208.297
R93 VGND.n7 VGND.t4 178.06
R94 VGND.n6 VGND.n5 125.822
R95 VGND.n19 VGND.t2 74.063
R96 VGND.n3 VGND.t5 59.6881
R97 VGND.n3 VGND.t0 54.9696
R98 VGND.n5 VGND.t6 41.2505
R99 VGND.n10 VGND.n4 36.1417
R100 VGND.n13 VGND.n12 36.1417
R101 VGND.n13 VGND.n1 36.1417
R102 VGND.n17 VGND.n1 36.1417
R103 VGND.n18 VGND.n17 36.1417
R104 VGND.n19 VGND.t1 31.4443
R105 VGND.n11 VGND.n10 29.3652
R106 VGND.n20 VGND.n18 24.4711
R107 VGND.n6 VGND.n4 22.9652
R108 VGND.n5 VGND.t3 21.3263
R109 VGND.n18 VGND.n0 9.3005
R110 VGND.n17 VGND.n16 9.3005
R111 VGND.n15 VGND.n1 9.3005
R112 VGND.n14 VGND.n13 9.3005
R113 VGND.n12 VGND.n2 9.3005
R114 VGND.n10 VGND.n9 9.3005
R115 VGND.n8 VGND.n4 9.3005
R116 VGND.n21 VGND.n20 7.46433
R117 VGND.n7 VGND.n6 7.11986
R118 VGND.n12 VGND.n11 6.77697
R119 VGND.n8 VGND.n7 0.223262
R120 VGND VGND.n21 0.160491
R121 VGND.n21 VGND.n0 0.147317
R122 VGND.n9 VGND.n8 0.122949
R123 VGND.n9 VGND.n2 0.122949
R124 VGND.n14 VGND.n2 0.122949
R125 VGND.n15 VGND.n14 0.122949
R126 VGND.n16 VGND.n15 0.122949
R127 VGND.n16 VGND.n0 0.122949
R128 GCLK.n1 GCLK 589
R129 GCLK.n1 GCLK.n0 585
R130 GCLK.n2 GCLK.n1 585
R131 GCLK GCLK.t1 167.752
R132 GCLK.n1 GCLK.t0 26.3844
R133 GCLK GCLK.n2 10.7205
R134 GCLK GCLK.n0 9.2805
R135 GCLK GCLK.n0 2.5605
R136 GCLK.n2 GCLK 1.1205
R137 VNB.n0 VNB 11629.4
R138 VNB.t6 VNB.t5 2286.61
R139 VNB.t3 VNB.t2 1766.93
R140 VNB.t4 VNB.t1 1524.41
R141 VNB VNB.n0 1311.63
R142 VNB.t2 VNB 1143.31
R143 VNB.t1 VNB.t3 900.788
R144 VNB.n0 VNB.t4 831.496
R145 VNB.n0 VNB.t6 461.942
R146 VNB.t7 VNB.t8 213.953
R147 VNB.t8 VNB.t0 93.0238
R148 VNB.n0 VNB.t7 53.3856
R149 a_477_124.t0 a_477_124.t1 68.5719
R150 a_309_338.t0 a_309_338.n1 838.037
R151 a_309_338.n0 a_309_338.t3 384.286
R152 a_309_338.n0 a_309_338.t2 242.607
R153 a_309_338.n1 a_309_338.n0 238.702
R154 a_309_338.n1 a_309_338.t1 140.756
R155 CLK.n0 CLK.t2 179.825
R156 CLK.n0 CLK.t3 170.308
R157 CLK.n1 CLK.t0 163.524
R158 CLK.n1 CLK.t1 154.24
R159 CLK.n3 CLK.n2 152
R160 CLK.n2 CLK.n1 49.9857
R161 CLK.n3 CLK 10.8611
R162 CLK.n2 CLK.n0 10.7116
R163 CLK CLK.n3 7.75808
R164 a_984_125.t0 a_984_125.t1 45.0005
R165 a_267_80.t0 a_267_80.t1 45.0005
C0 VPB GATE 0.045531f
C1 VPB VPWR 0.208586f
C2 GATE VPWR 0.01339f
C3 VPB VGND 0.015333f
C4 GATE VGND 0.00606f
C5 VPB CLK 0.075428f
C6 VPB GCLK 0.018072f
C7 VPWR VGND 0.114725f
C8 VPWR CLK 0.075523f
C9 VGND CLK 0.070617f
C10 VPWR GCLK 0.132646f
C11 VGND GCLK 0.102728f
C12 GCLK VNB 0.110551f
C13 CLK VNB 0.184922f
C14 VGND VNB 0.823996f
C15 VPWR VNB 0.631769f
C16 GATE VNB 0.116158f
C17 VPB VNB 1.54924f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlclkp_2 VNB VPB VPWR VGND GATE CLK GCLK
X0 VGND.t3 CLK.t0 a_315_48.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VPWR.t0 a_83_244.t4 a_27_74.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3109 pd=1.71 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_264_392.t1 GATE.t0 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.3109 ps=1.71 w=1 l=0.15
X3 VPWR.t1 a_1041_387.t3 GCLK.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t1 a_1041_387.t4 GCLK.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 GCLK.t0 a_1041_387.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.50165 ps=2.09 w=1.12 l=0.15
X6 VPWR.t7 a_27_74.t2 a_508_508.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR.t4 CLK.t1 a_315_48.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1703 pd=1.355 as=0.2646 ps=2.31 w=0.84 l=0.15
X8 VGND.t5 a_83_244.t5 a_27_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2093 pd=1.355 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_508_508.t0 a_315_48.t2 a_83_244.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.21335 ps=1.65 w=0.42 l=0.15
X10 a_315_338.t1 a_315_48.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.17335 ps=1.375 w=0.74 l=0.15
X11 GCLK.t2 a_1041_387.t6 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.21835 ps=2.21 w=0.74 l=0.15
X12 a_1041_387.t1 a_27_74.t3 a_1044_119.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0777 ps=0.95 w=0.74 l=0.15
X13 VGND.t6 a_27_74.t4 a_494_118.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.17335 pd=1.375 as=0.077425 ps=0.85 w=0.42 l=0.15
X14 a_267_74.t1 GATE.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2093 ps=1.355 w=0.64 l=0.15
X15 VPWR.t6 a_27_74.t5 a_1041_387.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.50165 pd=2.09 as=0.1625 ps=1.325 w=1 l=0.15
X16 a_1041_387.t0 CLK.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.1703 ps=1.355 w=1 l=0.15
X17 a_315_338.t0 a_315_48.t4 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.17325 ps=1.4 w=0.84 l=0.15
X18 a_1044_119.t0 CLK.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1295 ps=1.09 w=0.74 l=0.15
X19 a_494_118.t1 a_315_338.t2 a_83_244.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.077425 pd=0.85 as=0.15245 ps=1.235 w=0.42 l=0.15
X20 a_83_244.t3 a_315_338.t3 a_264_392.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.21335 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X21 a_83_244.t2 a_315_48.t5 a_267_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.15245 pd=1.235 as=0.0768 ps=0.88 w=0.64 l=0.15
R0 CLK.n1 CLK.t1 227.588
R1 CLK.n0 CLK.t2 207.529
R2 CLK.n0 CLK.t3 156.431
R3 CLK.n1 CLK.t0 154.24
R4 CLK CLK.n2 68.4956
R5 CLK.n2 CLK.n0 32.0605
R6 CLK.n2 CLK.n1 32.0547
R7 a_315_48.t1 a_315_48.n3 409.772
R8 a_315_48.n0 a_315_48.t5 402.002
R9 a_315_48.n0 a_315_48.t2 290.442
R10 a_315_48.n3 a_315_48.n2 281.603
R11 a_315_48.n1 a_315_48.n0 266.776
R12 a_315_48.n1 a_315_48.t4 207.553
R13 a_315_48.n2 a_315_48.t3 176.2
R14 a_315_48.n3 a_315_48.t0 165.595
R15 a_315_48.n2 a_315_48.n1 12.6087
R16 VGND.n6 VGND.t7 263.909
R17 VGND.n28 VGND.n27 204.679
R18 VGND.n7 VGND.t1 183.407
R19 VGND.n19 VGND.n18 126.341
R20 VGND.n12 VGND.n11 124.657
R21 VGND.n27 VGND.t0 89.063
R22 VGND.n18 VGND.t6 82.0388
R23 VGND.n18 VGND.t4 62.0408
R24 VGND.n10 VGND.n5 36.1417
R25 VGND.n13 VGND.n3 36.1417
R26 VGND.n17 VGND.n3 36.1417
R27 VGND.n21 VGND.n20 36.1417
R28 VGND.n21 VGND.n1 36.1417
R29 VGND.n25 VGND.n1 36.1417
R30 VGND.n26 VGND.n25 36.1417
R31 VGND.n11 VGND.t3 34.0546
R32 VGND.n12 VGND.n10 32.0005
R33 VGND.n28 VGND.n26 24.0946
R34 VGND.n6 VGND.n5 22.9652
R35 VGND.n11 VGND.t2 22.7032
R36 VGND.n27 VGND.t5 22.6611
R37 VGND.n20 VGND.n19 16.5652
R38 VGND.n13 VGND.n12 15.4358
R39 VGND.n26 VGND.n0 9.3005
R40 VGND.n25 VGND.n24 9.3005
R41 VGND.n23 VGND.n1 9.3005
R42 VGND.n22 VGND.n21 9.3005
R43 VGND.n20 VGND.n2 9.3005
R44 VGND.n17 VGND.n16 9.3005
R45 VGND.n15 VGND.n3 9.3005
R46 VGND.n14 VGND.n13 9.3005
R47 VGND.n8 VGND.n5 9.3005
R48 VGND.n10 VGND.n9 9.3005
R49 VGND.n12 VGND.n4 9.3005
R50 VGND.n29 VGND.n28 7.19894
R51 VGND.n7 VGND.n6 6.74444
R52 VGND.n19 VGND.n17 4.89462
R53 VGND.n8 VGND.n7 0.585372
R54 VGND VGND.n29 0.156997
R55 VGND.n29 VGND.n0 0.150766
R56 VGND.n9 VGND.n8 0.122949
R57 VGND.n9 VGND.n4 0.122949
R58 VGND.n14 VGND.n4 0.122949
R59 VGND.n15 VGND.n14 0.122949
R60 VGND.n16 VGND.n15 0.122949
R61 VGND.n16 VGND.n2 0.122949
R62 VGND.n22 VGND.n2 0.122949
R63 VGND.n23 VGND.n22 0.122949
R64 VGND.n24 VGND.n23 0.122949
R65 VGND.n24 VGND.n0 0.122949
R66 VNB.n0 VNB 14331.8
R67 VNB.n1 VNB 9581
R68 VNB VNB.n2 2520.49
R69 VNB.t8 VNB.t6 1705.68
R70 VNB.t5 VNB.t0 1618.77
R71 VNB.t9 VNB.n0 1540
R72 VNB.n2 VNB.t7 1535.96
R73 VNB.t6 VNB.n1 1520.99
R74 VNB.n0 VNB.t10 1270.34
R75 VNB.t7 VNB 1143.31
R76 VNB.t4 VNB.t3 1100
R77 VNB.t0 VNB.t8 1032.1
R78 VNB.t10 VNB.t2 993.177
R79 VNB.t1 VNB.t5 847.408
R80 VNB.t3 VNB.t9 792
R81 VNB.n1 VNB.t4 638
R82 VNB.n2 VNB.t1 217.285
R83 a_83_244.n3 a_83_244.n2 408.091
R84 a_83_244.n1 a_83_244.t4 284.342
R85 a_83_244.n2 a_83_244.n0 275.731
R86 a_83_244.n1 a_83_244.t5 176.964
R87 a_83_244.n2 a_83_244.n1 152
R88 a_83_244.n3 a_83_244.t1 143.269
R89 a_83_244.t3 a_83_244.n3 106.251
R90 a_83_244.n0 a_83_244.t0 95.7148
R91 a_83_244.n0 a_83_244.t2 62.0094
R92 a_27_74.n0 a_27_74.t3 1013.37
R93 a_27_74.t4 a_27_74.t2 574.652
R94 a_27_74.t3 a_27_74.t5 435.377
R95 a_27_74.n1 a_27_74.n0 369.976
R96 a_27_74.t1 a_27_74.n1 305.942
R97 a_27_74.n1 a_27_74.t0 217.659
R98 a_27_74.n0 a_27_74.t4 124.617
R99 VPWR.n19 VPWR.n18 585
R100 VPWR.n12 VPWR.n6 318.685
R101 VPWR.n27 VPWR.n1 312.889
R102 VPWR.n9 VPWR.t1 266.438
R103 VPWR.n18 VPWR.t7 119.608
R104 VPWR.n18 VPWR.t5 111.4
R105 VPWR.n8 VPWR.n7 83.9007
R106 VPWR.n7 VPWR.t2 78.2803
R107 VPWR.n7 VPWR.t6 77.8946
R108 VPWR.n1 VPWR.t0 57.2409
R109 VPWR.n1 VPWR.t8 57.1305
R110 VPWR.n6 VPWR.t4 42.2148
R111 VPWR.n6 VPWR.t3 37.5177
R112 VPWR.n21 VPWR.n2 36.1417
R113 VPWR.n25 VPWR.n2 36.1417
R114 VPWR.n26 VPWR.n25 36.1417
R115 VPWR.n13 VPWR.n4 36.1417
R116 VPWR.n17 VPWR.n4 36.1417
R117 VPWR.n12 VPWR.n11 35.7652
R118 VPWR.n21 VPWR.n20 25.8933
R119 VPWR.n11 VPWR.n8 15.8123
R120 VPWR.n19 VPWR.n17 13.177
R121 VPWR.n13 VPWR.n12 11.6711
R122 VPWR.n27 VPWR.n26 9.41227
R123 VPWR.n11 VPWR.n10 9.3005
R124 VPWR.n12 VPWR.n5 9.3005
R125 VPWR.n14 VPWR.n13 9.3005
R126 VPWR.n15 VPWR.n4 9.3005
R127 VPWR.n17 VPWR.n16 9.3005
R128 VPWR.n20 VPWR.n3 9.3005
R129 VPWR.n22 VPWR.n21 9.3005
R130 VPWR.n23 VPWR.n2 9.3005
R131 VPWR.n25 VPWR.n24 9.3005
R132 VPWR.n26 VPWR.n0 9.3005
R133 VPWR.n28 VPWR.n27 7.6232
R134 VPWR.n9 VPWR.n8 3.77294
R135 VPWR.n20 VPWR.n19 1.59004
R136 VPWR.n10 VPWR.n9 0.450875
R137 VPWR VPWR.n28 0.162583
R138 VPWR.n28 VPWR.n0 0.145253
R139 VPWR.n10 VPWR.n5 0.122949
R140 VPWR.n14 VPWR.n5 0.122949
R141 VPWR.n15 VPWR.n14 0.122949
R142 VPWR.n16 VPWR.n15 0.122949
R143 VPWR.n16 VPWR.n3 0.122949
R144 VPWR.n22 VPWR.n3 0.122949
R145 VPWR.n23 VPWR.n22 0.122949
R146 VPWR.n24 VPWR.n23 0.122949
R147 VPWR.n24 VPWR.n0 0.122949
R148 VPB VPB.n0 2344.05
R149 VPB.t7 VPB.t2 602.833
R150 VPB.t4 VPB.t3 271.813
R151 VPB.t3 VPB.t7 255.667
R152 VPB.t2 VPB.t1 242.21
R153 VPB.n0 VPB.t4 145.327
R154 VPB.t6 VPB 70.0225
R155 VPB.n0 VPB.t5 22.9928
R156 VPB.n0 VPB.t6 20.9026
R157 VPB.t5 VPB.t8 16.7222
R158 VPB.t8 VPB.t0 12.5418
R159 GATE.n0 GATE.t1 268.313
R160 GATE.n0 GATE.t0 236.983
R161 GATE GATE.n0 154.133
R162 a_264_392.t0 a_264_392.t1 53.1905
R163 a_1041_387.n0 a_1041_387.t3 245.553
R164 a_1041_387.n2 a_1041_387.t5 245.553
R165 a_1041_387.n4 a_1041_387.n3 237.297
R166 a_1041_387.n3 a_1041_387.n2 176.702
R167 a_1041_387.n0 a_1041_387.t4 174.906
R168 a_1041_387.n1 a_1041_387.t6 173.52
R169 a_1041_387.n3 a_1041_387.t1 144.387
R170 a_1041_387.n1 a_1041_387.n0 84.3505
R171 a_1041_387.t0 a_1041_387.n4 34.4755
R172 a_1041_387.n4 a_1041_387.t2 29.5505
R173 a_1041_387.n2 a_1041_387.n1 6.0255
R174 GCLK.n4 GCLK 589.85
R175 GCLK.n4 GCLK.n0 585
R176 GCLK.n5 GCLK.n4 585
R177 GCLK.n3 GCLK.n2 185
R178 GCLK.n2 GCLK.n1 185
R179 GCLK.n4 GCLK.t1 26.3844
R180 GCLK.n4 GCLK.t0 26.3844
R181 GCLK.n2 GCLK.t3 22.7032
R182 GCLK.n2 GCLK.t2 22.7032
R183 GCLK GCLK.n5 12.9944
R184 GCLK GCLK.n0 11.249
R185 GCLK.n1 GCLK 9.11565
R186 GCLK.n3 GCLK 8.33989
R187 GCLK GCLK.n3 6.01262
R188 GCLK.n1 GCLK 5.23686
R189 GCLK GCLK.n0 3.10353
R190 GCLK.n5 GCLK 1.35808
R191 a_508_508.t0 a_508_508.t1 126.644
R192 a_315_338.t0 a_315_338.n1 449.82
R193 a_315_338.n0 a_315_338.t3 390.712
R194 a_315_338.n1 a_315_338.n0 253.511
R195 a_315_338.n0 a_315_338.t2 252.248
R196 a_315_338.n1 a_315_338.t1 153.845
R197 a_1044_119.t0 a_1044_119.t1 34.0546
R198 a_494_118.t0 a_494_118.t1 100.001
R199 a_267_74.t0 a_267_74.t1 45.0005
C0 VPB GCLK 0.008358f
C1 VPWR VGND 0.148602f
C2 VPWR CLK 0.069079f
C3 VPWR GCLK 0.218851f
C4 VGND CLK 0.067337f
C5 VGND GCLK 0.125441f
C6 CLK GCLK 8.35e-20
C7 VPB GATE 0.040145f
C8 VPB VPWR 0.228019f
C9 VPB VGND 0.017281f
C10 GATE VPWR 0.015886f
C11 VPB CLK 0.084452f
C12 GATE VGND 0.006343f
C13 GCLK VNB 0.030438f
C14 CLK VNB 0.169963f
C15 VGND VNB 0.974179f
C16 VPWR VNB 0.756363f
C17 GATE VNB 0.125644f
C18 VPB VNB 1.73189f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlclkp_4 VNB VPB VPWR VGND GATE CLK GCLK
X0 VPWR.t9 a_27_74.t2 a_524_508.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.52 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_1047_74.t1 CLK.t0 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t2 a_1044_368.t3 GCLK.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_524_508.t0 a_334_54.t2 a_84_48.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.2102 ps=1.635 w=0.42 l=0.15
X4 GCLK.t5 a_1044_368.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1876 ps=1.455 w=1.12 l=0.15
X5 VGND.t0 a_1044_368.t5 GCLK.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_1044_368.t2 CLK.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.2114 ps=1.52 w=1.12 l=0.15
X7 a_286_80.t1 GATE.t0 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.240975 ps=1.45 w=0.64 l=0.15
X8 VPWR.t6 a_84_48.t4 a_27_74.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3109 pd=1.71 as=0.3304 ps=2.83 w=1.12 l=0.15
X9 a_84_48.t0 a_334_338.t2 a_283_392.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.635 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t5 a_84_48.t5 a_27_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.240975 pd=1.45 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 a_283_392.t1 GATE.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.3109 ps=1.71 w=1 l=0.15
X12 VPWR.t8 a_27_74.t3 a_1044_368.t1 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.5348 pd=2.075 as=0.1876 ps=1.455 w=1.12 l=0.15
X13 GCLK.t4 a_1044_368.t6 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.5348 ps=2.075 w=1.12 l=0.15
X14 a_334_338.t1 a_334_54.t3 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1848 ps=1.52 w=0.84 l=0.15
X15 a_1044_368.t0 a_27_74.t4 a_1047_74.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X16 VPWR.t1 CLK.t2 a_334_54.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2114 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X17 VGND.t1 a_1044_368.t7 GCLK.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_84_48.t1 a_334_54.t4 a_286_80.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.12935 pd=1.125 as=0.0768 ps=0.88 w=0.64 l=0.15
X19 a_491_124.t0 a_334_338.t3 a_84_48.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.118875 pd=1.195 as=0.12935 ps=1.125 w=0.42 l=0.15
X20 a_334_338.t0 a_334_54.t5 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2675 pd=2.66 as=0.16425 ps=1.305 w=0.74 l=0.15
X21 VGND.t7 a_27_74.t5 a_491_124.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.16425 pd=1.305 as=0.118875 ps=1.195 w=0.42 l=0.15
X22 GCLK.t1 a_1044_368.t8 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X23 VGND.t9 CLK.t3 a_334_54.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2333 ps=2.19 w=0.74 l=0.15
X24 GCLK.t0 a_1044_368.t9 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2977 ps=2.9 w=0.74 l=0.15
R0 a_27_74.t5 a_27_74.t2 457.632
R1 a_27_74.n1 a_27_74.t5 372.113
R2 a_27_74.n1 a_27_74.n0 365.493
R3 a_27_74.t1 a_27_74.n2 277.678
R4 a_27_74.n0 a_27_74.t3 264.298
R5 a_27_74.n2 a_27_74.n1 218.817
R6 a_27_74.n0 a_27_74.t4 204.048
R7 a_27_74.n2 a_27_74.t0 144.663
R8 a_524_508.t0 a_524_508.t1 126.644
R9 VPWR.n23 VPWR.n22 629.155
R10 VPWR.n16 VPWR.n6 317.808
R11 VPWR.n31 VPWR.n1 313.495
R12 VPWR.n10 VPWR.t3 258.238
R13 VPWR.n9 VPWR.t2 256.252
R14 VPWR.n8 VPWR.n7 134.764
R15 VPWR.n22 VPWR.t9 110.227
R16 VPWR.n22 VPWR.t7 78.566
R17 VPWR.n7 VPWR.t8 77.0106
R18 VPWR.n7 VPWR.t4 77.0103
R19 VPWR.n1 VPWR.t5 59.1005
R20 VPWR.n1 VPWR.t6 55.271
R21 VPWR.n6 VPWR.t1 55.1136
R22 VPWR.n25 VPWR.n2 36.1417
R23 VPWR.n29 VPWR.n2 36.1417
R24 VPWR.n30 VPWR.n29 36.1417
R25 VPWR.n17 VPWR.n4 36.1417
R26 VPWR.n21 VPWR.n4 36.1417
R27 VPWR.n25 VPWR.n24 35.6194
R28 VPWR.n16 VPWR.n15 33.8829
R29 VPWR.n6 VPWR.t0 30.2812
R30 VPWR.n11 VPWR.n10 25.224
R31 VPWR.n11 VPWR.n8 25.224
R32 VPWR.n15 VPWR.n8 16.5652
R33 VPWR.n23 VPWR.n21 15.853
R34 VPWR.n17 VPWR.n16 13.5534
R35 VPWR.n32 VPWR.n31 12.5979
R36 VPWR.n12 VPWR.n11 9.3005
R37 VPWR.n15 VPWR.n14 9.3005
R38 VPWR.n16 VPWR.n5 9.3005
R39 VPWR.n18 VPWR.n17 9.3005
R40 VPWR.n19 VPWR.n4 9.3005
R41 VPWR.n21 VPWR.n20 9.3005
R42 VPWR.n24 VPWR.n3 9.3005
R43 VPWR.n26 VPWR.n25 9.3005
R44 VPWR.n27 VPWR.n2 9.3005
R45 VPWR.n29 VPWR.n28 9.3005
R46 VPWR.n30 VPWR.n0 9.3005
R47 VPWR.n10 VPWR.n9 6.88165
R48 VPWR.n13 VPWR.n8 4.62059
R49 VPWR.n24 VPWR.n23 3.57527
R50 VPWR.n31 VPWR.n30 3.01226
R51 VPWR.n12 VPWR.n9 0.610715
R52 VPWR.n13 VPWR.n12 0.184273
R53 VPWR.n14 VPWR.n13 0.184273
R54 VPWR VPWR.n32 0.163644
R55 VPWR.n32 VPWR.n0 0.144205
R56 VPWR.n14 VPWR.n5 0.122949
R57 VPWR.n18 VPWR.n5 0.122949
R58 VPWR.n19 VPWR.n18 0.122949
R59 VPWR.n20 VPWR.n19 0.122949
R60 VPWR.n20 VPWR.n3 0.122949
R61 VPWR.n26 VPWR.n3 0.122949
R62 VPWR.n27 VPWR.n26 0.122949
R63 VPWR.n28 VPWR.n27 0.122949
R64 VPWR.n28 VPWR.n0 0.122949
R65 VPB.n0 VPB 2285.62
R66 VPB.n1 VPB 1914.94
R67 VPB VPB.n2 1159.37
R68 VPB.t10 VPB.t4 564.383
R69 VPB.t9 VPB.n0 531.761
R70 VPB.t4 VPB.t3 485.216
R71 VPB.t5 VPB.t7 377.957
R72 VPB.t7 VPB 306.452
R73 VPB.t1 VPB.t0 280.914
R74 VPB.t0 VPB.t10 247.715
R75 VPB.n2 VPB.t6 232.393
R76 VPB.t3 VPB.t2 229.839
R77 VPB.n1 VPB.t9 227.044
R78 VPB.t8 VPB.t11 219.835
R79 VPB.t6 VPB.t5 214.517
R80 VPB.n2 VPB.t8 172.727
R81 VPB.t11 VPB.n1 125.621
R82 VPB.n0 VPB.t1 61.2908
R83 CLK.n3 CLK.t2 254.121
R84 CLK.n0 CLK.t1 226.809
R85 CLK.n0 CLK.t0 198.204
R86 CLK.n2 CLK.t3 196.013
R87 CLK.n4 CLK.n1 162.363
R88 CLK.n4 CLK.n3 156.382
R89 CLK.n1 CLK.n0 35.055
R90 CLK.n2 CLK.n1 25.5611
R91 CLK.n3 CLK.n2 19.7187
R92 CLK CLK.n4 2.74336
R93 VGND.n12 VGND.t3 259.137
R94 VGND.n24 VGND.n4 215.702
R95 VGND.n19 VGND.n18 211.571
R96 VGND.n33 VGND.n32 202.579
R97 VGND.n8 VGND.t1 145.184
R98 VGND.n10 VGND.n9 123.257
R99 VGND.n4 VGND.t7 120.811
R100 VGND.n32 VGND.t6 102.189
R101 VGND.n17 VGND.n6 36.1417
R102 VGND.n20 VGND.n3 36.1417
R103 VGND.n26 VGND.n25 36.1417
R104 VGND.n26 VGND.n1 36.1417
R105 VGND.n30 VGND.n1 36.1417
R106 VGND.n31 VGND.n30 36.1417
R107 VGND.n9 VGND.t0 34.0546
R108 VGND.n24 VGND.n3 32.7534
R109 VGND.n19 VGND.n17 30.8711
R110 VGND.n11 VGND.n10 28.2358
R111 VGND.n13 VGND.n11 26.7943
R112 VGND.n4 VGND.t4 22.7037
R113 VGND.n9 VGND.t2 22.7032
R114 VGND.n18 VGND.t8 22.7032
R115 VGND.n18 VGND.t9 22.7032
R116 VGND.n32 VGND.t5 22.5391
R117 VGND.n33 VGND.n31 20.7064
R118 VGND.n12 VGND.n6 17.4082
R119 VGND.n20 VGND.n19 16.5652
R120 VGND.n25 VGND.n24 14.6829
R121 VGND.n31 VGND.n0 9.3005
R122 VGND.n30 VGND.n29 9.3005
R123 VGND.n28 VGND.n1 9.3005
R124 VGND.n27 VGND.n26 9.3005
R125 VGND.n25 VGND.n2 9.3005
R126 VGND.n24 VGND.n23 9.3005
R127 VGND.n22 VGND.n3 9.3005
R128 VGND.n21 VGND.n20 9.3005
R129 VGND.n19 VGND.n5 9.3005
R130 VGND.n17 VGND.n16 9.3005
R131 VGND.n15 VGND.n6 9.3005
R132 VGND.n14 VGND.n13 9.3005
R133 VGND.n11 VGND.n7 9.3005
R134 VGND.n34 VGND.n33 7.21776
R135 VGND.n10 VGND.n8 6.70714
R136 VGND.n13 VGND.n12 1.64153
R137 VGND.n8 VGND.n7 0.645862
R138 VGND VGND.n34 0.157244
R139 VGND.n34 VGND.n0 0.150522
R140 VGND.n14 VGND.n7 0.122949
R141 VGND.n15 VGND.n14 0.122949
R142 VGND.n16 VGND.n15 0.122949
R143 VGND.n16 VGND.n5 0.122949
R144 VGND.n21 VGND.n5 0.122949
R145 VGND.n22 VGND.n21 0.122949
R146 VGND.n23 VGND.n22 0.122949
R147 VGND.n23 VGND.n2 0.122949
R148 VGND.n27 VGND.n2 0.122949
R149 VGND.n28 VGND.n27 0.122949
R150 VGND.n29 VGND.n28 0.122949
R151 VGND.n29 VGND.n0 0.122949
R152 a_1047_74.t0 a_1047_74.t1 38.9194
R153 VNB.n0 VNB 10336
R154 VNB VNB.n1 4997.95
R155 VNB.t9 VNB.t3 2852.49
R156 VNB.t7 VNB.t5 1986.35
R157 VNB.t4 VNB.n0 1760
R158 VNB.t8 VNB.t4 1613.33
R159 VNB.t12 VNB.t8 1353.85
R160 VNB.t0 VNB.t2 1154.86
R161 VNB.t5 VNB 1143.31
R162 VNB.n1 VNB.t6 1085.56
R163 VNB.t2 VNB.t1 993.177
R164 VNB.t3 VNB.t0 993.177
R165 VNB.t10 VNB.t11 993.177
R166 VNB.t11 VNB.t9 900.788
R167 VNB.t6 VNB.t7 900.788
R168 VNB.n0 VNB.t10 588.976
R169 VNB.n1 VNB.t12 372.308
R170 a_1044_368.n9 a_1044_368.n8 257.647
R171 a_1044_368.n3 a_1044_368.t4 226.809
R172 a_1044_368.n5 a_1044_368.n0 226.809
R173 a_1044_368.n7 a_1044_368.t6 226.809
R174 a_1044_368.n1 a_1044_368.t7 214.651
R175 a_1044_368.n6 a_1044_368.t9 212.081
R176 a_1044_368.n4 a_1044_368.t5 212.081
R177 a_1044_368.n2 a_1044_368.t8 212.081
R178 a_1044_368.n1 a_1044_368.t3 206.869
R179 a_1044_368.n8 a_1044_368.t0 150.623
R180 a_1044_368.n8 a_1044_368.n7 138.185
R181 a_1044_368.n4 a_1044_368.n3 80.9076
R182 a_1044_368.n2 a_1044_368.n1 71.4465
R183 a_1044_368.n6 a_1044_368.n5 71.4398
R184 a_1044_368.n9 a_1044_368.t2 32.5407
R185 a_1044_368.t1 a_1044_368.n9 26.3844
R186 a_1044_368.n7 a_1044_368.n6 8.60764
R187 a_1044_368.n3 a_1044_368.n2 5.16479
R188 a_1044_368.n5 a_1044_368.n4 2.58264
R189 GCLK GCLK.t4 295.372
R190 GCLK.n5 GCLK.n0 216.916
R191 GCLK.n3 GCLK.n1 154.645
R192 GCLK.n3 GCLK.n2 114.82
R193 GCLK.n0 GCLK.t6 26.3844
R194 GCLK.n0 GCLK.t5 26.3844
R195 GCLK.n2 GCLK.t2 22.7032
R196 GCLK.n2 GCLK.t1 22.7032
R197 GCLK.n1 GCLK.t3 22.7032
R198 GCLK.n1 GCLK.t0 22.7032
R199 GCLK.n4 GCLK 22.5396
R200 GCLK.n4 GCLK.n3 14.7144
R201 GCLK.n5 GCLK.n4 2.22659
R202 GCLK GCLK.n5 1.94833
R203 a_334_54.t5 a_334_54.t0 601.717
R204 a_334_54.t1 a_334_54.n2 463.817
R205 a_334_54.n1 a_334_54.t4 366.216
R206 a_334_54.n1 a_334_54.t2 290.442
R207 a_334_54.n0 a_334_54.t5 221.919
R208 a_334_54.n0 a_334_54.t3 199.694
R209 a_334_54.n2 a_334_54.n0 164.811
R210 a_334_54.n2 a_334_54.n1 39.2538
R211 a_84_48.n3 a_84_48.n2 730.383
R212 a_84_48.n1 a_84_48.t4 279.695
R213 a_84_48.n2 a_84_48.n0 274.027
R214 a_84_48.n1 a_84_48.t5 172.315
R215 a_84_48.n2 a_84_48.n1 152
R216 a_84_48.n3 a_84_48.t2 150.095
R217 a_84_48.t0 a_84_48.n3 112.385
R218 a_84_48.n0 a_84_48.t3 70.0005
R219 a_84_48.n0 a_84_48.t1 56.2951
R220 GATE.n0 GATE.t0 265.101
R221 GATE.n0 GATE.t1 231.629
R222 GATE GATE.n0 159.112
R223 a_286_80.t0 a_286_80.t1 45.0005
R224 a_334_338.t1 a_334_338.n1 819.091
R225 a_334_338.n0 a_334_338.t2 381.365
R226 a_334_338.n1 a_334_338.t0 314.442
R227 a_334_338.n1 a_334_338.n0 253.517
R228 a_334_338.n0 a_334_338.t3 231.361
R229 a_283_392.t0 a_283_392.t1 53.1905
R230 a_491_124.t0 a_491_124.t1 275.188
C0 VPB GATE 0.046077f
C1 VPB VGND 0.014767f
C2 VPWR GATE 0.018362f
C3 VPWR VGND 0.152132f
C4 VPB CLK 0.099346f
C5 VPB GCLK 0.014557f
C6 VPWR CLK 0.067065f
C7 GATE VGND 0.006567f
C8 VPWR GCLK 0.457838f
C9 VGND CLK 0.036932f
C10 VGND GCLK 0.306045f
C11 CLK GCLK 2.01e-19
C12 VPB VPWR 0.239121f
C13 GCLK VNB 0.057869f
C14 CLK VNB 0.232591f
C15 VGND VNB 1.03665f
C16 GATE VNB 0.115863f
C17 VPWR VNB 0.82031f
C18 VPB VNB 1.96677f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrbn_1 VNB VPB VPWR VGND Q_N Q GATE_N RESET_B D
X0 VPWR.t2 a_889_92.t3 a_1437_112.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2023 pd=1.51 as=0.231 ps=2.23 w=0.84 l=0.15
X1 VPWR.t8 RESET_B.t0 a_889_92.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2128 pd=1.5 as=0.1736 ps=1.43 w=1.12 l=0.15
X2 Q_N.t1 a_1437_112.t2 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2023 ps=1.51 w=1.12 l=0.15
X3 VGND.t6 D.t0 a_27_424.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X4 VGND.t2 a_889_92.t4 a_841_118.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1533 pd=1.57 as=0.0504 ps=0.66 w=0.42 l=0.15
X5 a_231_74.t0 GATE_N.t0 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X6 VGND RESET_B a_1133_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0888 ps=0.98 w=0.74 l=0.15
X7 a_686_74.t3 a_373_74.t2 a_611_392.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t5 a_231_74.t2 a_373_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2013 pd=1.33 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_231_74.t1 GATE_N.t1 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2562 ps=1.45 w=0.84 l=0.15
X10 a_611_392.t0 a_27_424.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.25245 ps=1.64 w=1 l=0.15
X11 a_802_508.t0 a_231_74.t3 a_686_74.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.11235 pd=0.955 as=0.1664 ps=1.385 w=0.42 l=0.15
X12 a_608_74.t1 a_27_424.t3 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2013 ps=1.33 w=0.64 l=0.15
X13 a_841_118.t0 a_373_74.t3 a_686_74.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.19175 ps=1.265 w=0.42 l=0.15
X14 VPWR.t0 a_231_74.t4 a_373_74.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.25245 pd=1.64 as=0.383 ps=2.88 w=0.84 l=0.15
X15 VPWR.t9 D.t1 a_27_424.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2562 pd=1.45 as=0.2478 ps=2.27 w=0.84 l=0.15
X16 a_1133_74# a_686_74.t4 a_889_92.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X17 a_889_92.t1 a_686_74.t5 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.239575 ps=2.025 w=1.12 l=0.15
X18 VGND.t3 a_889_92.t5 a_1437_112.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.127925 pd=1.105 as=0.1925 ps=1.8 w=0.55 l=0.15
X19 Q_N.t0 a_1437_112.t3 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.127925 ps=1.105 w=0.74 l=0.15
X20 VPWR.t3 a_889_92.t6 a_802_508.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.239575 pd=2.025 as=0.11235 ps=0.955 w=0.42 l=0.15
X21 Q.t0 a_889_92.t7 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3248 pd=2.82 as=0.2128 ps=1.5 w=1.12 l=0.15
X22 a_686_74.t1 a_231_74.t5 a_608_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.19175 pd=1.265 as=0.0768 ps=0.88 w=0.64 l=0.15
R0 a_889_92.n4 a_889_92.t4 379.413
R1 a_889_92.n0 a_889_92.t3 224.143
R2 a_889_92.n2 a_889_92.t7 218.774
R3 a_889_92.n6 a_889_92.n3 213.546
R4 a_889_92.n7 a_889_92.n6 196.673
R5 a_889_92.n5 a_889_92.t0 193.809
R6 a_889_92.n5 a_889_92.n4 176.988
R7 a_889_92.n4 a_889_92.t6 162.542
R8 a_889_92.n2 a_889_92.n1 156.249
R9 a_889_92.n0 a_889_92.t5 144.875
R10 a_889_92.n3 a_889_92.n0 84.3505
R11 a_889_92.t1 a_889_92.n7 28.1434
R12 a_889_92.n7 a_889_92.t2 26.3844
R13 a_889_92.n3 a_889_92.n2 14.7283
R14 a_889_92.n6 a_889_92.n5 9.09524
R15 a_1437_112.t1 a_1437_112.n1 420.577
R16 a_1437_112.n0 a_1437_112.t2 264.298
R17 a_1437_112.n1 a_1437_112.t0 237.19
R18 a_1437_112.n0 a_1437_112.t3 204.048
R19 a_1437_112.n1 a_1437_112.n0 176.825
R20 VPWR.n26 VPWR.n4 698.312
R21 VPWR.n19 VPWR.n18 585
R22 VPWR.n17 VPWR.n16 585
R23 VPWR.n11 VPWR.n10 323.693
R24 VPWR.n32 VPWR.n1 314.961
R25 VPWR.n18 VPWR.n17 295.5
R26 VPWR.n12 VPWR.n9 241.079
R27 VPWR.n1 VPWR.t5 107.882
R28 VPWR.n17 VPWR.t7 100.309
R29 VPWR.n18 VPWR.t3 74.5629
R30 VPWR.n4 VPWR.t0 65.6672
R31 VPWR.n9 VPWR.t2 57.0752
R32 VPWR.n30 VPWR.n2 36.1417
R33 VPWR.n31 VPWR.n30 36.1417
R34 VPWR.n20 VPWR.n5 36.1417
R35 VPWR.n24 VPWR.n5 36.1417
R36 VPWR.n25 VPWR.n24 36.1417
R37 VPWR.n15 VPWR.n8 36.1417
R38 VPWR.n4 VPWR.t4 35.5684
R39 VPWR.n1 VPWR.t9 35.1791
R40 VPWR.n10 VPWR.t8 35.1791
R41 VPWR.n10 VPWR.t1 31.6612
R42 VPWR.n9 VPWR.t6 28.4028
R43 VPWR.n26 VPWR.n2 25.977
R44 VPWR.n32 VPWR.n31 22.9652
R45 VPWR.n26 VPWR.n25 21.4593
R46 VPWR.n20 VPWR.n19 11.3956
R47 VPWR.n12 VPWR.n11 10.2312
R48 VPWR.n13 VPWR.n8 9.3005
R49 VPWR.n15 VPWR.n14 9.3005
R50 VPWR.n7 VPWR.n6 9.3005
R51 VPWR.n21 VPWR.n20 9.3005
R52 VPWR.n22 VPWR.n5 9.3005
R53 VPWR.n24 VPWR.n23 9.3005
R54 VPWR.n25 VPWR.n3 9.3005
R55 VPWR.n27 VPWR.n26 9.3005
R56 VPWR.n28 VPWR.n2 9.3005
R57 VPWR.n30 VPWR.n29 9.3005
R58 VPWR.n31 VPWR.n0 9.3005
R59 VPWR.n11 VPWR.n8 8.65932
R60 VPWR.n16 VPWR.n15 8.00733
R61 VPWR.n33 VPWR.n32 7.27223
R62 VPWR.n16 VPWR.n7 3.4329
R63 VPWR.n19 VPWR.n7 2.78933
R64 VPWR.n13 VPWR.n12 0.203538
R65 VPWR VPWR.n33 0.157962
R66 VPWR.n33 VPWR.n0 0.149814
R67 VPWR.n14 VPWR.n13 0.122949
R68 VPWR.n14 VPWR.n6 0.122949
R69 VPWR.n21 VPWR.n6 0.122949
R70 VPWR.n22 VPWR.n21 0.122949
R71 VPWR.n23 VPWR.n22 0.122949
R72 VPWR.n23 VPWR.n3 0.122949
R73 VPWR.n27 VPWR.n3 0.122949
R74 VPWR.n28 VPWR.n27 0.122949
R75 VPWR.n29 VPWR.n28 0.122949
R76 VPWR.n29 VPWR.n0 0.122949
R77 VPB.n0 VPB 3616.13
R78 VPB.n1 VPB 2398.87
R79 VPB VPB.n2 744.005
R80 VPB.n2 VPB.t2 399.873
R81 VPB.t7 VPB.t11 388.173
R82 VPB.t1 VPB.t4 332.015
R83 VPB.t2 VPB.t6 300.51
R84 VPB.t5 VPB.t8 275.807
R85 VPB.n0 VPB.t5 263.038
R86 VPB.t3 VPB.n0 260.176
R87 VPB.t0 VPB.t1 259.312
R88 VPB.t11 VPB 257.93
R89 VPB.t10 VPB.t3 253.016
R90 VPB.n1 VPB.t9 248.242
R91 VPB.t9 VPB.t10 219.599
R92 VPB.t6 VPB.t0 203.571
R93 VPB.t4 VPB.n1 196.302
R94 VPB.n2 VPB.t7 137.904
R95 RESET_B.n1 RESET_B.t0 250.909
R96 RESET_B.n1 RESET_B.n0 178.34
R97 RESET_B RESET_B.n1 159.345
R98 Q_N.n1 Q_N 589.777
R99 Q_N.n1 Q_N.n0 585
R100 Q_N.n2 Q_N.n1 585
R101 Q_N Q_N.t0 209.077
R102 Q_N.n1 Q_N.t1 26.3844
R103 Q_N Q_N.n2 12.8005
R104 Q_N Q_N.n0 11.0811
R105 Q_N Q_N.n0 3.05722
R106 Q_N.n2 Q_N 1.33781
R107 D.n0 D.t1 233.022
R108 D.n0 D.t0 179.609
R109 D D.n0 68.53
R110 a_27_424.n1 a_27_424.n0 437.741
R111 a_27_424.t1 a_27_424.n1 395.949
R112 a_27_424.n1 a_27_424.t0 303.279
R113 a_27_424.n0 a_27_424.t3 274.74
R114 a_27_424.n0 a_27_424.t2 231.629
R115 VGND.n6 VGND.t2 288.817
R116 VGND.n14 VGND.n13 185
R117 VGND.n5 VGND.n4 129.38
R118 VGND.n22 VGND.n21 119.573
R119 VGND.n13 VGND.t5 58.2861
R120 VGND.n21 VGND.t6 51.1974
R121 VGND.n13 VGND.t1 48.7505
R122 VGND.n4 VGND.t3 48.3911
R123 VGND.n7 VGND.n3 36.1417
R124 VGND.n11 VGND.n3 36.1417
R125 VGND.n12 VGND.n11 36.1417
R126 VGND.n19 VGND.n1 36.1417
R127 VGND.n20 VGND.n19 36.1417
R128 VGND.n21 VGND.t0 32.4351
R129 VGND.n4 VGND.t4 21.8154
R130 VGND.n15 VGND.n12 20.5745
R131 VGND.n14 VGND.n1 19.2555
R132 VGND.n22 VGND.n20 18.0711
R133 VGND.n7 VGND.n6 12.8005
R134 VGND.n6 VGND.n5 12.1653
R135 VGND.n8 VGND.n7 9.3005
R136 VGND.n9 VGND.n3 9.3005
R137 VGND.n11 VGND.n10 9.3005
R138 VGND.n12 VGND.n2 9.3005
R139 VGND.n16 VGND.n15 9.3005
R140 VGND.n17 VGND.n1 9.3005
R141 VGND.n19 VGND.n18 9.3005
R142 VGND.n20 VGND.n0 9.3005
R143 VGND.n23 VGND.n22 7.47871
R144 VGND.n15 VGND.n14 0.187361
R145 VGND VGND.n23 0.16068
R146 VGND.n8 VGND.n5 0.150876
R147 VGND.n23 VGND.n0 0.14713
R148 VGND.n9 VGND.n8 0.122949
R149 VGND.n10 VGND.n9 0.122949
R150 VGND.n10 VGND.n2 0.122949
R151 VGND.n16 VGND.n2 0.122949
R152 VGND.n17 VGND.n16 0.122949
R153 VGND.n18 VGND.n17 0.122949
R154 VGND.n18 VGND.n0 0.122949
R155 VNB VNB.n0 12456.3
R156 VNB.t0 VNB.t5 5007.32
R157 VNB.t8 VNB.t2 2791.14
R158 VNB.t1 VNB.t3 1889.2
R159 VNB.t4 VNB.t8 1803.88
R160 VNB.t2 VNB.t9 1413.85
R161 VNB.n0 VNB.t0 1400.56
R162 VNB.t5 VNB.t7 1276.62
R163 VNB.n0 VNB.t6 1231.02
R164 VNB.t9 VNB 1218.84
R165 VNB.t6 VNB.t1 950.693
R166 VNB.t3 VNB.t4 950.693
R167 a_841_118.t0 a_841_118.t1 68.5719
R168 GATE_N.n0 GATE_N.t1 233.054
R169 GATE_N.n0 GATE_N.t0 210.143
R170 GATE_N GATE_N.n0 69.097
R171 a_231_74.t1 a_231_74.n3 726.423
R172 a_231_74.n0 a_231_74.t3 490.748
R173 a_231_74.n0 a_231_74.t5 314.274
R174 a_231_74.n1 a_231_74.t4 270.555
R175 a_231_74.n3 a_231_74.t0 227.391
R176 a_231_74.n1 a_231_74.t2 176.03
R177 a_231_74.n2 a_231_74.n1 152
R178 a_231_74.n3 a_231_74.n2 116.014
R179 a_231_74.n2 a_231_74.n0 63.185
R180 a_373_74.t1 a_373_74.n1 920.101
R181 a_373_74.n0 a_373_74.t2 465.933
R182 a_373_74.n1 a_373_74.n0 296.493
R183 a_373_74.n0 a_373_74.t3 126.927
R184 a_373_74.n1 a_373_74.t0 118.38
R185 a_611_392.t0 a_611_392.t1 53.1905
R186 a_686_74.n3 a_686_74.n2 699.856
R187 a_686_74.n2 a_686_74.n1 274.853
R188 a_686_74.n2 a_686_74.n0 241.733
R189 a_686_74.n0 a_686_74.t5 226.809
R190 a_686_74.n0 a_686_74.t4 161.006
R191 a_686_74.n3 a_686_74.t0 110.227
R192 a_686_74.n1 a_686_74.t2 70.1791
R193 a_686_74.n1 a_686_74.t1 54.3755
R194 a_686_74.t3 a_686_74.n3 30.9107
R195 a_802_508.t0 a_802_508.t1 250.94
R196 a_608_74.t0 a_608_74.t1 45.0005
R197 Q Q.n0 595.994
R198 Q.n3 Q.n0 585
R199 Q.n2 Q.n0 585
R200 Q.n2 Q.n1 60.2513
R201 Q.n0 Q.t0 29.0228
R202 Q.n3 Q 9.78874
R203 Q.n1 Q 8.47293
R204 Q Q.n2 1.95815
R205 Q Q.n3 1.35579
R206 Q.n1 Q 0.0396059
C0 VPWR Q_N 0.130373f
C1 RESET_B Q 0.001867f
C2 VGND Q 0.117601f
C3 a_1133_74# VPWR 9.5e-19
C4 VPB D 0.064788f
C5 VGND Q_N 0.099098f
C6 VPB GATE_N 0.072896f
C7 a_1133_74# RESET_B 5.52e-19
C8 D GATE_N 0.112617f
C9 VPB VPWR 0.263324f
C10 a_1133_74# VGND 0.011028f
C11 D VPWR 0.019796f
C12 a_1133_74# Q 3.42e-19
C13 VPB RESET_B 0.032479f
C14 GATE_N VPWR 0.009263f
C15 VPB VGND 0.02429f
C16 D VGND 0.038654f
C17 VPB Q 0.018395f
C18 D Q 3.55e-21
C19 GATE_N VGND 0.020662f
C20 VPWR RESET_B 0.015249f
C21 VPB Q_N 0.013806f
C22 VPWR VGND 0.140158f
C23 VPWR Q 0.096924f
C24 RESET_B VGND 0.034455f
C25 Q_N VNB 0.111241f
C26 Q VNB 0.01974f
C27 VGND VNB 1.05182f
C28 RESET_B VNB 0.094682f
C29 VPWR VNB 0.788129f
C30 GATE_N VNB 0.122515f
C31 D VNB 0.15176f
C32 VPB VNB 2.0872f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrbp_1 VNB VPB VPWR VGND D Q_N Q GATE RESET_B
X0 a_642_392.t0 a_226_104.t2 a_564_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.405 as=0.12 ps=1.24 w=1 l=0.15
X1 a_775_124.t1 a_226_104.t3 a_642_392.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1346 ps=1.15 w=0.42 l=0.15
X2 VPWR.t3 a_226_104.t4 a_353_98.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1878 pd=1.39 as=0.2478 ps=2.27 w=0.84 l=0.15
X3 Q_N.t0 a_1342_74.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X4 VPWR.t6 D.t0 a_27_142.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.22785 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_564_392.t1 a_27_142.t2 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.1878 ps=1.39 w=1 l=0.15
X6 a_226_104.t0 GATE.t0 VGND.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2701 pd=2.21 as=0.144575 ps=1.15 w=0.74 l=0.15
X7 VGND.t5 RESET_B.t0 a_1051_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X8 a_1051_74.t0 a_642_392.t4 a_823_98.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_571_80.t0 a_27_142.t3 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.193075 ps=1.49 w=0.64 l=0.15
X10 a_642_392.t2 a_353_98.t2 a_571_80.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1346 pd=1.15 as=0.0672 ps=0.85 w=0.64 l=0.15
X11 VGND.t3 a_823_98.t2 a_1342_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.124175 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X12 VGND.t2 a_226_104.t5 a_353_98.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.193075 pd=1.49 as=0.259 ps=2.18 w=0.74 l=0.15
X13 VPWR.t4 a_823_98.t3 a_1342_74.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X14 a_753_508.t1 a_353_98.t3 a_642_392.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.10605 pd=0.925 as=0.1764 ps=1.405 w=0.42 l=0.15
X15 a_226_104.t1 GATE.t1 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3066 pd=2.41 as=0.22785 ps=1.52 w=0.84 l=0.15
X16 VGND.t1 a_823_98.t4 a_775_124.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X17 VPWR.t2 a_823_98.t5 a_753_508.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.23345 pd=1.79 as=0.10605 ps=0.925 w=0.42 l=0.15
X18 a_823_98.t1 a_642_392.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.182 pd=1.445 as=0.23345 ps=1.79 w=1.12 l=0.15
X19 VGND.t6 D.t1 a_27_142.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.144575 pd=1.15 as=0.15675 ps=1.67 w=0.55 l=0.15
R0 a_226_104.t1 a_226_104.n2 764.23
R1 a_226_104.t3 a_226_104.t2 678.014
R2 a_226_104.n0 a_226_104.t3 427.096
R3 a_226_104.n2 a_226_104.n1 277.32
R4 a_226_104.n1 a_226_104.t4 243.411
R5 a_226_104.n1 a_226_104.t5 179.947
R6 a_226_104.n0 a_226_104.t0 126.43
R7 a_226_104.n2 a_226_104.n0 26.5266
R8 a_564_392.t0 a_564_392.t1 47.2805
R9 a_642_392.n3 a_642_392.n2 653.341
R10 a_642_392.n2 a_642_392.n1 290.42
R11 a_642_392.n2 a_642_392.n0 246.938
R12 a_642_392.n1 a_642_392.t5 226.809
R13 a_642_392.n1 a_642_392.t4 198.204
R14 a_642_392.n3 a_642_392.t3 114.918
R15 a_642_392.n0 a_642_392.t1 72.8576
R16 a_642_392.n0 a_642_392.t2 60.5809
R17 a_642_392.t0 a_642_392.n3 32.8807
R18 VPB.t1 VPB.t5 1013.84
R19 VPB.t8 VPB.t3 551.614
R20 VPB.t2 VPB.t1 418.817
R21 VPB.t9 VPB.t2 334.543
R22 VPB.t7 VPB.t8 316.668
R23 VPB.t4 VPB.t9 283.469
R24 VPB.t3 VPB.t6 275.807
R25 VPB.t5 VPB.t0 257.93
R26 VPB VPB.t7 257.93
R27 VPB.t6 VPB.t4 199.195
R28 a_775_124.t0 a_775_124.t1 68.5719
R29 VNB.t8 VNB.t4 3464.57
R30 VNB.t7 VNB.t2 2621.52
R31 VNB.t1 VNB.t0 2286.61
R32 VNB.t5 VNB.t3 1524.41
R33 VNB.t2 VNB.t9 1362.73
R34 VNB.t6 VNB.t7 1293.44
R35 VNB VNB.t6 1143.31
R36 VNB.t0 VNB.t8 900.788
R37 VNB.t3 VNB.t1 900.788
R38 VNB.t9 VNB.t5 831.496
R39 a_353_98.t1 a_353_98.n1 818.976
R40 a_353_98.n0 a_353_98.t3 478.37
R41 a_353_98.n0 a_353_98.t2 314.274
R42 a_353_98.n1 a_353_98.t0 276.005
R43 a_353_98.n1 a_353_98.n0 62.7649
R44 VPWR.n24 VPWR.n1 646.029
R45 VPWR.n18 VPWR.n4 614.529
R46 VPWR.n11 VPWR.n10 585
R47 VPWR.n9 VPWR.n8 585
R48 VPWR.n7 VPWR.n6 324.065
R49 VPWR.n10 VPWR.n9 161.821
R50 VPWR.n10 VPWR.t2 70.3576
R51 VPWR.n9 VPWR.t1 58.1312
R52 VPWR.n4 VPWR.t3 56.2862
R53 VPWR.n1 VPWR.t7 55.1136
R54 VPWR.n1 VPWR.t6 55.1136
R55 VPWR.n6 VPWR.t0 43.8979
R56 VPWR.n22 VPWR.n2 36.1417
R57 VPWR.n23 VPWR.n22 36.1417
R58 VPWR.n16 VPWR.n5 36.1417
R59 VPWR.n17 VPWR.n16 36.1417
R60 VPWR.n6 VPWR.t4 35.1791
R61 VPWR.n18 VPWR.n17 32.7534
R62 VPWR.n4 VPWR.t5 30.3907
R63 VPWR.n12 VPWR.n5 27.0646
R64 VPWR.n24 VPWR.n23 16.5652
R65 VPWR.n18 VPWR.n2 14.3064
R66 VPWR.n8 VPWR.n7 9.63534
R67 VPWR.n13 VPWR.n12 9.3005
R68 VPWR.n14 VPWR.n5 9.3005
R69 VPWR.n16 VPWR.n15 9.3005
R70 VPWR.n17 VPWR.n3 9.3005
R71 VPWR.n19 VPWR.n18 9.3005
R72 VPWR.n20 VPWR.n2 9.3005
R73 VPWR.n22 VPWR.n21 9.3005
R74 VPWR.n23 VPWR.n0 9.3005
R75 VPWR.n25 VPWR.n24 7.53404
R76 VPWR.n11 VPWR.n8 5.77305
R77 VPWR.n12 VPWR.n11 0.16782
R78 VPWR VPWR.n25 0.161409
R79 VPWR.n13 VPWR.n7 0.156297
R80 VPWR.n25 VPWR.n0 0.146411
R81 VPWR.n14 VPWR.n13 0.122949
R82 VPWR.n15 VPWR.n14 0.122949
R83 VPWR.n15 VPWR.n3 0.122949
R84 VPWR.n19 VPWR.n3 0.122949
R85 VPWR.n20 VPWR.n19 0.122949
R86 VPWR.n21 VPWR.n20 0.122949
R87 VPWR.n21 VPWR.n0 0.122949
R88 a_1342_74.t1 a_1342_74.n2 440.904
R89 a_1342_74.n2 a_1342_74.t0 258.019
R90 a_1342_74.n1 a_1342_74.t2 256.933
R91 a_1342_74.n1 a_1342_74.n0 208.465
R92 a_1342_74.n2 a_1342_74.n1 176.048
R93 Q_N.n0 Q_N.t0 302.086
R94 Q_N Q_N.n0 13.3565
R95 Q_N.n0 Q_N 0.0982489
R96 D.n0 D.t0 217.934
R97 D.n0 D.t1 172.143
R98 D D.n0 153.358
R99 a_27_142.t1 a_27_142.n1 776.324
R100 a_27_142.t1 a_27_142.n2 768.644
R101 a_27_142.n1 a_27_142.n0 364.329
R102 a_27_142.n2 a_27_142.t0 284.322
R103 a_27_142.n0 a_27_142.t3 259.43
R104 a_27_142.n0 a_27_142.t2 231.629
R105 a_27_142.n2 a_27_142.n1 12.4348
R106 GATE.n0 GATE.t1 219.31
R107 GATE.n0 GATE.t0 204.048
R108 GATE GATE.n0 153.358
R109 VGND.n10 VGND.t1 257.195
R110 VGND.n17 VGND.n16 245.625
R111 VGND.n6 VGND.t3 169.094
R112 VGND.n5 VGND.t5 150.272
R113 VGND.n25 VGND.n24 125.609
R114 VGND.n24 VGND.t6 50.1666
R115 VGND.n16 VGND.t2 49.0935
R116 VGND.n9 VGND.n8 36.1417
R117 VGND.n14 VGND.n3 36.1417
R118 VGND.n15 VGND.n14 36.1417
R119 VGND.n22 VGND.n1 36.1417
R120 VGND.n23 VGND.n22 36.1417
R121 VGND.n18 VGND.n15 35.6473
R122 VGND.n10 VGND.n9 35.3887
R123 VGND.n16 VGND.t4 26.3167
R124 VGND.n24 VGND.t0 25.6983
R125 VGND.n25 VGND.n23 18.4476
R126 VGND.n17 VGND.n1 16.3142
R127 VGND.n10 VGND.n3 12.0476
R128 VGND.n6 VGND.n5 11.3522
R129 VGND.n8 VGND.n7 9.3005
R130 VGND.n9 VGND.n4 9.3005
R131 VGND.n11 VGND.n10 9.3005
R132 VGND.n12 VGND.n3 9.3005
R133 VGND.n14 VGND.n13 9.3005
R134 VGND.n15 VGND.n2 9.3005
R135 VGND.n19 VGND.n18 9.3005
R136 VGND.n20 VGND.n1 9.3005
R137 VGND.n22 VGND.n21 9.3005
R138 VGND.n23 VGND.n0 9.3005
R139 VGND.n8 VGND.n5 7.52991
R140 VGND.n26 VGND.n25 7.46433
R141 VGND.n18 VGND.n17 4.00858
R142 VGND.n7 VGND.n6 0.211603
R143 VGND VGND.n26 0.160491
R144 VGND.n26 VGND.n0 0.147317
R145 VGND.n7 VGND.n4 0.122949
R146 VGND.n11 VGND.n4 0.122949
R147 VGND.n12 VGND.n11 0.122949
R148 VGND.n13 VGND.n12 0.122949
R149 VGND.n13 VGND.n2 0.122949
R150 VGND.n19 VGND.n2 0.122949
R151 VGND.n20 VGND.n19 0.122949
R152 VGND.n21 VGND.n20 0.122949
R153 VGND.n21 VGND.n0 0.122949
R154 RESET_B.n1 RESET_B.n0 285.719
R155 RESET_B.n1 RESET_B.t0 178.34
R156 RESET_B RESET_B.n1 158.746
R157 a_1051_74.t0 a_1051_74.t1 38.9194
R158 a_823_98.n6 a_823_98.t4 376.454
R159 a_823_98.n1 a_823_98.t3 315.229
R160 a_823_98.n4 a_823_98.n0 250.909
R161 a_823_98.n3 a_823_98.n1 236.18
R162 a_823_98.t1 a_823_98.n7 229.774
R163 a_823_98.n1 a_823_98.t2 226.541
R164 a_823_98.n3 a_823_98.n2 206.969
R165 a_823_98.n5 a_823_98.n4 195.423
R166 a_823_98.n5 a_823_98.t0 194.228
R167 a_823_98.n7 a_823_98.n6 180.453
R168 a_823_98.n6 a_823_98.t5 154.508
R169 a_823_98.n4 a_823_98.n3 13.146
R170 a_823_98.n7 a_823_98.n5 7.53456
R171 a_571_80.t0 a_571_80.t1 39.3755
R172 a_753_508.t0 a_753_508.t1 236.869
C0 VPWR D 0.013018f
C1 VPB RESET_B 0.029799f
C2 VPB GATE 0.051748f
C3 VPWR RESET_B 0.016618f
C4 VPB VGND 0.0184f
C5 VPWR GATE 0.010877f
C6 VPB Q 0.015392f
C7 VPWR VGND 0.133094f
C8 D GATE 0.071943f
C9 D VGND 0.034321f
C10 VPWR Q 0.130091f
C11 VPB Q_N 0.014548f
C12 VPWR Q_N 0.112647f
C13 RESET_B VGND 0.037518f
C14 D Q 7.64e-21
C15 D Q_N 4.91e-21
C16 GATE VGND 0.022279f
C17 RESET_B Q 0.006283f
C18 GATE Q 4.34e-21
C19 GATE Q_N 1.93e-21
C20 VGND Q 0.098084f
C21 VPB VPWR 0.239602f
C22 VGND Q_N 0.088699f
C23 VPB D 0.051635f
C24 Q_N VNB 0.112664f
C25 Q VNB 0.019948f
C26 VGND VNB 1.01483f
C27 GATE VNB 0.103118f
C28 RESET_B VNB 0.105078f
C29 D VNB 0.129249f
C30 VPWR VNB 0.757122f
C31 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxbp_2 VNB VPB VPWR VGND CLK Q D Q_N
X0 VPWR.t9 a_1290_102# Q.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VGND.t6 a_1000_424.t4 a_1290_102# VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t0 CLK.t0 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 VGND a_1290_102# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t0 a_1835_368.t1 Q_N.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_1000_424.t2 a_206_368.t2 a_753_284.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.196025 pd=1.68 as=0.1935 ps=1.49 w=0.55 l=0.15
X6 VGND.t3 CLK.t1 a_27_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.20385 pd=1.355 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 a_206_368.t1 a_27_74.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3252 pd=2.59 as=0.20385 ps=1.355 w=0.74 l=0.15
X8 a_1248_128.t0 a_27_74.t3 a_1000_424.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.196025 ps=1.68 w=0.42 l=0.15
X9 Q.t1 a_1290_102# VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1988 ps=1.505 w=1.12 l=0.15
X10 a_558_445.t3 a_206_368.t3 a_451_503.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1197 pd=0.99 as=0.106225 ps=1.095 w=0.42 l=0.15
X11 a_451_503.t0 D.t0 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.35635 ps=2.6 w=0.42 l=0.15
X12 VPWR.t1 a_1835_368.t2 Q_N.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t9 a_753_284.t4 a_717_102.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.09825 pd=0.925 as=0.0504 ps=0.66 w=0.42 l=0.15
X14 Q.t0 a_1290_102# VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X15 Q_N.t1 a_1835_368.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.14385 ps=1.145 w=0.74 l=0.15
X16 a_558_445.t0 a_27_74.t4 a_451_503.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.083025 pd=0.865 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 a_717_102.t1 a_206_368.t4 a_558_445.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.083025 ps=0.865 w=0.42 l=0.15
X18 a_753_284.t0 a_558_445.t4 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1935 pd=1.49 as=0.09825 ps=0.925 w=0.55 l=0.15
X19 a_206_368.t0 a_27_74.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X20 VPWR.t5 a_753_284.t5 a_702_445.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.206525 pd=1.545 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 a_451_503.t1 D.t1 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.106225 pd=1.095 as=0.3234 ps=2.38 w=0.42 l=0.15
X22 VPWR.t6 a_1000_424.t5 a_1290_102# VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.126 ps=1.14 w=0.84 l=0.15
X23 a_702_445.t0 a_27_74.t6 a_558_445.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1197 ps=0.99 w=0.42 l=0.15
X24 a_1000_424.t1 a_27_74.t7 a_753_284.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.73 as=0.126 ps=1.14 w=0.84 l=0.15
X25 VPWR.t7 a_1290_102# a_1835_368.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.295 ps=2.59 w=1 l=0.15
X26 a_753_284.t3 a_558_445.t5 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.206525 ps=1.545 w=0.84 l=0.15
X27 VGND.t7 a_1290_102# a_1248_128.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1533 pd=1.57 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_1208_479.t0 a_206_368.t5 a_1000_424.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.24255 ps=1.73 w=0.42 l=0.15
R0 a_1000_424.n5 a_1000_424.n4 647.13
R1 a_1000_424.n0 a_1000_424.t2 330.772
R2 a_1000_424.n1 a_1000_424.t4 286.134
R3 a_1000_424.n3 a_1000_424.n2 246.892
R4 a_1000_424.n4 a_1000_424.n0 241.346
R5 a_1000_424.n4 a_1000_424.n3 217.727
R6 a_1000_424.n6 a_1000_424.n5 192.31
R7 a_1000_424.n1 a_1000_424.t5 181.821
R8 a_1000_424.n5 a_1000_424.t3 164.167
R9 a_1000_424.n7 a_1000_424.n6 52.0382
R10 a_1000_424.n0 a_1000_424.t0 40.001
R11 a_1000_424.n6 a_1000_424.t1 32.7139
R12 a_1000_424.n3 a_1000_424.n1 18.9884
R13 VPWR.n16 VPWR.t9 860.096
R14 VPWR.n2 VPWR.t3 779.655
R15 VPWR.n31 VPWR.n30 674.282
R16 VPWR.n18 VPWR.n10 606.333
R17 VPWR.n43 VPWR.n1 326.231
R18 VPWR.n12 VPWR.t7 279.082
R19 VPWR.n13 VPWR.t1 267.132
R20 VPWR.n30 VPWR.t5 131.333
R21 VPWR.n10 VPWR.t6 55.1136
R22 VPWR.n30 VPWR.t4 46.2205
R23 VPWR.n36 VPWR.n4 36.1417
R24 VPWR.n37 VPWR.n36 36.1417
R25 VPWR.n38 VPWR.n37 36.1417
R26 VPWR.n24 VPWR.n23 36.1417
R27 VPWR.n24 VPWR.n6 36.1417
R28 VPWR.n28 VPWR.n6 36.1417
R29 VPWR.n29 VPWR.n28 36.1417
R30 VPWR.n22 VPWR.n8 36.1417
R31 VPWR.n16 VPWR.n15 32.7534
R32 VPWR.n32 VPWR.n4 32.3937
R33 VPWR.n42 VPWR.n41 31.2225
R34 VPWR.n10 VPWR.t8 30.9991
R35 VPWR.n18 VPWR.n17 28.2358
R36 VPWR.n1 VPWR.t2 26.3844
R37 VPWR.n1 VPWR.t0 26.3844
R38 VPWR.n15 VPWR.n12 24.8476
R39 VPWR.n43 VPWR.n42 22.9652
R40 VPWR.n31 VPWR.n29 22.0115
R41 VPWR.n18 VPWR.n8 19.2005
R42 VPWR.n38 VPWR.n2 15.9545
R43 VPWR.n17 VPWR.n16 14.6829
R44 VPWR.n23 VPWR.n22 11.2946
R45 VPWR.n15 VPWR.n14 9.3005
R46 VPWR.n16 VPWR.n11 9.3005
R47 VPWR.n17 VPWR.n9 9.3005
R48 VPWR.n19 VPWR.n18 9.3005
R49 VPWR.n20 VPWR.n8 9.3005
R50 VPWR.n22 VPWR.n21 9.3005
R51 VPWR.n23 VPWR.n7 9.3005
R52 VPWR.n25 VPWR.n24 9.3005
R53 VPWR.n26 VPWR.n6 9.3005
R54 VPWR.n28 VPWR.n27 9.3005
R55 VPWR.n29 VPWR.n5 9.3005
R56 VPWR.n33 VPWR.n32 9.3005
R57 VPWR.n34 VPWR.n4 9.3005
R58 VPWR.n36 VPWR.n35 9.3005
R59 VPWR.n37 VPWR.n3 9.3005
R60 VPWR.n39 VPWR.n38 9.3005
R61 VPWR.n41 VPWR.n40 9.3005
R62 VPWR.n42 VPWR.n0 9.3005
R63 VPWR.n44 VPWR.n43 7.52053
R64 VPWR.n13 VPWR.n12 6.97747
R65 VPWR.n41 VPWR.n2 3.55606
R66 VPWR.n32 VPWR.n31 2.41828
R67 VPWR.n14 VPWR.n13 0.543268
R68 VPWR VPWR.n44 0.161231
R69 VPWR.n44 VPWR.n0 0.146587
R70 VPWR.n14 VPWR.n11 0.122949
R71 VPWR.n11 VPWR.n9 0.122949
R72 VPWR.n19 VPWR.n9 0.122949
R73 VPWR.n20 VPWR.n19 0.122949
R74 VPWR.n21 VPWR.n20 0.122949
R75 VPWR.n21 VPWR.n7 0.122949
R76 VPWR.n25 VPWR.n7 0.122949
R77 VPWR.n26 VPWR.n25 0.122949
R78 VPWR.n27 VPWR.n26 0.122949
R79 VPWR.n27 VPWR.n5 0.122949
R80 VPWR.n33 VPWR.n5 0.122949
R81 VPWR.n34 VPWR.n33 0.122949
R82 VPWR.n35 VPWR.n34 0.122949
R83 VPWR.n35 VPWR.n3 0.122949
R84 VPWR.n39 VPWR.n3 0.122949
R85 VPWR.n40 VPWR.n39 0.122949
R86 VPWR.n40 VPWR.n0 0.122949
R87 VPB.n0 VPB 2658.47
R88 VPB VPB.n1 2224.68
R89 VPB.t7 VPB.t10 809.543
R90 VPB.t6 VPB.t2 625.673
R91 VPB.t13 VPB.t11 515.861
R92 VPB.t11 VPB.t1 503.091
R93 VPB.n0 VPB.t7 388.173
R94 VPB.t9 VPB.t8 372.786
R95 VPB.t3 VPB.t5 367.743
R96 VPB.t10 VPB.t12 273.253
R97 VPB.t5 VPB.t6 273.253
R98 VPB.t8 VPB.t4 270.57
R99 VPB.t0 VPB 257.93
R100 VPB.t12 VPB.t13 229.839
R101 VPB.t2 VPB.t0 229.839
R102 VPB.t4 VPB.n0 168.355
R103 VPB.n1 VPB.t3 135.35
R104 VPB.n1 VPB.t9 93.1967
R105 Q Q.n0 599.011
R106 Q Q.t0 170.034
R107 Q.n0 Q.t2 26.3844
R108 Q.n0 Q.t1 26.3844
R109 VGND.n1 VGND.t5 365.2
R110 VGND.n21 VGND.t7 279.276
R111 VGND.n4 VGND.n3 204.766
R112 VGND.n41 VGND.n40 198.132
R113 VGND.n12 VGND.t0 178.81
R114 VGND.n11 VGND.t1 151.175
R115 VGND.n9 VGND.n8 117.419
R116 VGND.n3 VGND.t9 64.2862
R117 VGND.n40 VGND.t2 40.541
R118 VGND.n40 VGND.t3 39.7302
R119 VGND.n22 VGND.n6 36.1417
R120 VGND.n26 VGND.n6 36.1417
R121 VGND.n27 VGND.n26 36.1417
R122 VGND.n28 VGND.n27 36.1417
R123 VGND.n33 VGND.n32 36.1417
R124 VGND.n34 VGND.n33 36.1417
R125 VGND.n39 VGND.n38 36.1417
R126 VGND.n21 VGND.n20 34.2593
R127 VGND.n34 VGND.n1 33.8829
R128 VGND.n3 VGND.t4 32.7278
R129 VGND.n32 VGND.n4 32.377
R130 VGND.n16 VGND.n9 32.0005
R131 VGND.n15 VGND.n14 30.8711
R132 VGND.n8 VGND.t8 30.0005
R133 VGND.n14 VGND.n11 28.2358
R134 VGND.n8 VGND.t6 22.7032
R135 VGND.n16 VGND.n15 16.5652
R136 VGND.n20 VGND.n9 15.4358
R137 VGND.n28 VGND.n4 14.3064
R138 VGND.n41 VGND.n39 14.3064
R139 VGND.n38 VGND.n1 13.5534
R140 VGND.n22 VGND.n21 13.177
R141 VGND.n39 VGND.n0 9.3005
R142 VGND.n38 VGND.n37 9.3005
R143 VGND.n36 VGND.n1 9.3005
R144 VGND.n35 VGND.n34 9.3005
R145 VGND.n33 VGND.n2 9.3005
R146 VGND.n32 VGND.n31 9.3005
R147 VGND.n30 VGND.n4 9.3005
R148 VGND.n29 VGND.n28 9.3005
R149 VGND.n27 VGND.n5 9.3005
R150 VGND.n26 VGND.n25 9.3005
R151 VGND.n24 VGND.n6 9.3005
R152 VGND.n23 VGND.n22 9.3005
R153 VGND.n21 VGND.n7 9.3005
R154 VGND.n20 VGND.n19 9.3005
R155 VGND.n14 VGND.n13 9.3005
R156 VGND.n15 VGND.n10 9.3005
R157 VGND.n17 VGND.n16 9.3005
R158 VGND.n18 VGND.n9 9.3005
R159 VGND.n42 VGND.n41 7.46433
R160 VGND.n12 VGND.n11 6.79022
R161 VGND.n13 VGND.n12 0.5771
R162 VGND VGND.n42 0.160491
R163 VGND.n42 VGND.n0 0.147317
R164 VGND.n13 VGND.n10 0.122949
R165 VGND.n17 VGND.n10 0.122949
R166 VGND.n18 VGND.n17 0.122949
R167 VGND.n19 VGND.n18 0.122949
R168 VGND.n19 VGND.n7 0.122949
R169 VGND.n23 VGND.n7 0.122949
R170 VGND.n24 VGND.n23 0.122949
R171 VGND.n25 VGND.n24 0.122949
R172 VGND.n25 VGND.n5 0.122949
R173 VGND.n29 VGND.n5 0.122949
R174 VGND.n30 VGND.n29 0.122949
R175 VGND.n31 VGND.n30 0.122949
R176 VGND.n31 VGND.n2 0.122949
R177 VGND.n35 VGND.n2 0.122949
R178 VGND.n36 VGND.n35 0.122949
R179 VGND.n37 VGND.n36 0.122949
R180 VGND.n37 VGND.n0 0.122949
R181 VNB.t12 VNB.t1 4723.36
R182 VNB.t2 VNB.t7 3302.89
R183 VNB.t8 VNB.t3 2656.17
R184 VNB.t11 VNB.t10 2471.39
R185 VNB.t5 VNB.t2 1489.76
R186 VNB.t6 VNB.t8 1362.73
R187 VNB.t13 VNB.t6 1212.6
R188 VNB.t4 VNB.t9 1177.95
R189 VNB VNB.t5 1143.31
R190 VNB.t10 VNB.t12 1097.11
R191 VNB.t1 VNB.t0 993.177
R192 VNB.t7 VNB.t4 993.177
R193 VNB.t9 VNB.t13 900.788
R194 VNB.t3 VNB.t11 831.496
R195 CLK.n0 CLK.t0 285.01
R196 CLK.n0 CLK.t1 177.631
R197 CLK CLK.n0 161.168
R198 a_27_74.n1 a_27_74.t7 565.37
R199 a_27_74.n0 a_27_74.t4 293.012
R200 a_27_74.t0 a_27_74.n5 285.75
R201 a_27_74.n4 a_27_74.t5 281.017
R202 a_27_74.n3 a_27_74.n2 236.583
R203 a_27_74.n2 a_27_74.n0 218.94
R204 a_27_74.n2 a_27_74.n1 212.916
R205 a_27_74.n4 a_27_74.t2 173.638
R206 a_27_74.n3 a_27_74.t1 153.444
R207 a_27_74.n5 a_27_74.n4 152
R208 a_27_74.n0 a_27_74.t6 129.935
R209 a_27_74.n1 a_27_74.t3 76.4681
R210 a_27_74.n5 a_27_74.n3 19.1077
R211 a_1835_368.t0 a_1835_368.n3 439.978
R212 a_1835_368.n1 a_1835_368.t2 240.197
R213 a_1835_368.n3 a_1835_368.n0 240.197
R214 a_1835_368.n1 a_1835_368.t1 182.138
R215 a_1835_368.n2 a_1835_368.t3 179.947
R216 a_1835_368.n2 a_1835_368.n1 60.6157
R217 a_1835_368.n3 a_1835_368.n2 5.11262
R218 Q_N.n2 Q_N 589.385
R219 Q_N.n2 Q_N.n0 585
R220 Q_N.n3 Q_N.n2 585
R221 Q_N Q_N.n1 159.274
R222 Q_N.n2 Q_N.t0 26.3844
R223 Q_N.n1 Q_N.t2 22.7032
R224 Q_N.n1 Q_N.t1 22.7032
R225 Q_N Q_N.n3 11.7484
R226 Q_N Q_N.n0 10.1704
R227 Q_N Q_N.n0 2.80598
R228 Q_N.n3 Q_N 1.2279
R229 a_206_368.n0 a_206_368.t4 1140.73
R230 a_206_368.n0 a_206_368.t3 474.795
R231 a_206_368.n2 a_206_368.t2 418.962
R232 a_206_368.n2 a_206_368.t5 378.707
R233 a_206_368.n1 a_206_368.t1 341.94
R234 a_206_368.n3 a_206_368.n2 289.642
R235 a_206_368.t0 a_206_368.n3 216.209
R236 a_206_368.n1 a_206_368.n0 152
R237 a_206_368.n3 a_206_368.n1 23.9183
R238 a_753_284.n3 a_753_284.n2 644.038
R239 a_753_284.n2 a_753_284.n1 331.897
R240 a_753_284.n0 a_753_284.t5 310.111
R241 a_753_284.n2 a_753_284.n0 180.898
R242 a_753_284.n0 a_753_284.t4 141.946
R243 a_753_284.n1 a_753_284.t2 48.0005
R244 a_753_284.n1 a_753_284.t0 48.0005
R245 a_753_284.t1 a_753_284.n3 35.1791
R246 a_753_284.n3 a_753_284.t3 35.1791
R247 a_1248_128.t0 a_1248_128.t1 60.0005
R248 a_451_503.n1 a_451_503.n0 873.971
R249 a_451_503.n0 a_451_503.t1 220.093
R250 a_451_503.n0 a_451_503.t3 70.3576
R251 a_451_503.n1 a_451_503.t2 40.0005
R252 a_451_503.t0 a_451_503.n1 40.0005
R253 a_558_445.n2 a_558_445.n1 585
R254 a_558_445.n0 a_558_445.t4 332.699
R255 a_558_445.n3 a_558_445.n2 292.64
R256 a_558_445.n2 a_558_445.n0 270.036
R257 a_558_445.n0 a_558_445.t5 201.22
R258 a_558_445.n1 a_558_445.t3 138.369
R259 a_558_445.n1 a_558_445.t1 128.988
R260 a_558_445.n3 a_558_445.t2 69.7446
R261 a_558_445.n3 a_558_445.t0 25.6807
R262 a_558_445.n4 a_558_445.n3 16.8426
R263 D.n0 D.t0 341.587
R264 D D.t1 325.505
R265 D.n0 D 9.51845
R266 D D.n0 2.62614
R267 a_717_102.t0 a_717_102.t1 68.5719
R268 a_702_445.t0 a_702_445.t1 126.644
C0 CLK VPB 0.03313f
C1 CLK VPWR 0.016855f
C2 D VPB 0.109696f
C3 D VPWR 0.013034f
C4 VGND VPB 0.024841f
C5 D a_1290_102# 6.55e-20
C6 VGND VPWR 0.189211f
C7 Q VPB 0.002366f
C8 VGND a_1290_102# 0.304621f
C9 Q_N VPB 0.007032f
C10 Q VPWR 0.016134f
C11 Q a_1290_102# 0.220908f
C12 Q_N VPWR 0.22785f
C13 Q_N a_1290_102# 0.001958f
C14 CLK VGND 0.013211f
C15 D VGND 0.008632f
C16 VPB VPWR 0.331768f
C17 a_1290_102# VPB 0.247145f
C18 D Q_N 1.94e-21
C19 VGND Q 0.164792f
C20 a_1290_102# VPWR 0.302025f
C21 VGND Q_N 0.166564f
C22 Q_N VNB 0.030859f
C23 Q VNB 0.009808f
C24 VGND VNB 1.31949f
C25 D VNB 0.132696f
C26 CLK VNB 0.154784f
C27 VPWR VNB 1.03923f
C28 VPB VNB 2.49838f
C29 a_1290_102# VNB 0.550098f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxtp_4 VNB VPB VPWR VGND Q D CLK
X0 a_1034_424.t3 a_27_74.t2 a_696_458.t3 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2226 ps=1.37 w=0.84 l=0.15
X1 VPWR.t7 CLK.t0 a_27_74.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 a_651_503.t0 a_27_74.t3 a_544_485.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.088725 ps=0.895 w=0.42 l=0.15
X3 VPWR.t1 a_1226_296.t2 Q.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Q.t2 a_1226_296.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t3 a_1226_296.t4 Q.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_544_485.t2 a_27_74.t4 a_437_503.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.075675 pd=0.83 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 Q.t0 a_1226_296.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.203 ps=1.505 w=1.12 l=0.15
X8 a_437_503.t2 D.t0 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.088725 pd=0.895 as=0.2544 ps=2.2 w=0.42 l=0.15
X9 VGND.t7 a_1034_424.t4 a_1226_296.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 VGND.t4 CLK.t1 a_27_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.17575 pd=1.215 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 Q.t5 a_1226_296.t6 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1147 ps=1.05 w=0.74 l=0.15
X12 Q.t4 a_1226_296.t7 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.111 ps=1.04 w=0.74 l=0.15
X13 a_1034_424.t0 a_206_368.t2 a_696_458.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1076 pd=0.985 as=0.099 ps=0.985 w=0.55 l=0.15
X14 a_696_458.t0 a_544_485.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.099 pd=0.985 as=0.19715 ps=1.365 w=0.55 l=0.15
X15 a_1178_124# a_27_74.t5 a_1034_424.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.06615 pd=0.735 as=0.1076 ps=0.985 w=0.42 l=0.15
X16 VGND.t6 a_696_458.t4 a_735_102.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.19715 pd=1.365 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_1141_508.t0 a_206_368.t3 a_1034_424.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X18 a_206_368.t1 a_27_74.t6 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_544_485.t0 a_206_368.t4 a_437_503.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.088725 pd=0.895 as=0.088725 ps=0.895 w=0.42 l=0.15
X20 VPWR.t5 a_1226_296.t8 a_1141_508.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.195 as=0.09975 ps=0.895 w=0.42 l=0.15
X21 VPWR.t9 a_696_458.t5 a_651_503.t1 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.23985 pd=1.735 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 a_696_458.t1 a_544_485.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2226 pd=1.37 as=0.23985 ps=1.735 w=0.84 l=0.15
X23 VPWR.t10 a_1034_424.t5 a_1226_296.t0 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.126 ps=1.14 w=0.84 l=0.15
X24 a_206_368.t0 a_27_74.t7 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2516 pd=2.16 as=0.17575 ps=1.215 w=0.74 l=0.15
X25 a_437_503.t0 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.355025 ps=2.6 w=0.42 l=0.15
X26 a_735_102.t0 a_206_368.t5 a_544_485.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.075675 ps=0.83 w=0.42 l=0.15
R0 a_27_74.t5 a_27_74.t2 719.383
R1 a_27_74.n1 a_27_74.t5 448.339
R2 a_27_74.n2 a_27_74.n1 314.837
R3 a_27_74.n0 a_27_74.t4 313.647
R4 a_27_74.t0 a_27_74.n4 290.298
R5 a_27_74.n3 a_27_74.t6 282.012
R6 a_27_74.n1 a_27_74.n0 237.243
R7 a_27_74.n0 a_27_74.t3 208.114
R8 a_27_74.n3 a_27_74.t7 174.632
R9 a_27_74.n2 a_27_74.t1 164.523
R10 a_27_74.n4 a_27_74.n3 152
R11 a_27_74.n4 a_27_74.n2 9.46137
R12 a_696_458.n3 a_696_458.n2 667.072
R13 a_696_458.n1 a_696_458.t5 517.347
R14 a_696_458.n2 a_696_458.n0 217.018
R15 a_696_458.n2 a_696_458.n1 193.75
R16 a_696_458.n1 a_696_458.t4 155.847
R17 a_696_458.n3 a_696_458.t3 89.1195
R18 a_696_458.n0 a_696_458.t0 40.1966
R19 a_696_458.t1 a_696_458.n3 35.1791
R20 a_696_458.n0 a_696_458.t2 27.9239
R21 a_1034_424.n5 a_1034_424.n4 695.393
R22 a_1034_424.n2 a_1034_424.t5 266.707
R23 a_1034_424.n4 a_1034_424.n3 231.481
R24 a_1034_424.n3 a_1034_424.t4 223.327
R25 a_1034_424.n4 a_1034_424.n0 209.065
R26 a_1034_424.n2 a_1034_424.n1 196.013
R27 a_1034_424.n3 a_1034_424.n2 124.005
R28 a_1034_424.n5 a_1034_424.t1 112.572
R29 a_1034_424.n0 a_1034_424.t0 59.3176
R30 a_1034_424.n0 a_1034_424.t2 52.8576
R31 a_1034_424.t3 a_1034_424.n5 34.0065
R32 VPB.t10 VPB.t7 589.919
R33 VPB.t5 VPB.t14 487.769
R34 VPB.t13 VPB.t0 431.587
R35 VPB.t0 VPB.t12 347.312
R36 VPB.t9 VPB.t5 319.221
R37 VPB.t14 VPB.t4 273.253
R38 VPB.t12 VPB.t9 273.253
R39 VPB.t6 VPB.t11 273.253
R40 VPB.t7 VPB.t6 273.253
R41 VPB VPB.t8 257.93
R42 VPB.t2 VPB.t1 229.839
R43 VPB.t3 VPB.t2 229.839
R44 VPB.t4 VPB.t3 229.839
R45 VPB.t8 VPB.t10 229.839
R46 VPB.t11 VPB.t13 199.195
R47 CLK.n0 CLK.t0 259.132
R48 CLK.n0 CLK.t1 198.882
R49 CLK CLK.n0 156.934
R50 VPWR.n2 VPWR.t6 804.092
R51 VPWR.n20 VPWR.t5 683.111
R52 VPWR.n28 VPWR.n27 616.869
R53 VPWR.n13 VPWR.n11 334.173
R54 VPWR.n40 VPWR.n1 331.5
R55 VPWR.n9 VPWR.n8 326.231
R56 VPWR.n12 VPWR.t1 264.714
R57 VPWR.n27 VPWR.t0 164.47
R58 VPWR.n27 VPWR.t9 117.474
R59 VPWR.n8 VPWR.t10 55.1136
R60 VPWR.n13 VPWR.n12 40.1055
R61 VPWR.n33 VPWR.n4 36.1417
R62 VPWR.n34 VPWR.n33 36.1417
R63 VPWR.n35 VPWR.n34 36.1417
R64 VPWR.n39 VPWR.n38 36.1417
R65 VPWR.n21 VPWR.n6 36.1417
R66 VPWR.n25 VPWR.n6 36.1417
R67 VPWR.n26 VPWR.n25 36.1417
R68 VPWR.n29 VPWR.n26 36.1417
R69 VPWR.n15 VPWR.n14 36.1417
R70 VPWR.n40 VPWR.n39 35.3887
R71 VPWR.n35 VPWR.n2 31.624
R72 VPWR.n19 VPWR.n9 29.7417
R73 VPWR.n8 VPWR.t4 29.6087
R74 VPWR.n1 VPWR.t8 26.3844
R75 VPWR.n1 VPWR.t7 26.3844
R76 VPWR.n11 VPWR.t2 26.3844
R77 VPWR.n11 VPWR.t3 26.3844
R78 VPWR.n21 VPWR.n20 23.7181
R79 VPWR.n15 VPWR.n9 23.7181
R80 VPWR.n20 VPWR.n19 23.3417
R81 VPWR.n28 VPWR.n4 13.014
R82 VPWR.n14 VPWR.n10 9.3005
R83 VPWR.n16 VPWR.n15 9.3005
R84 VPWR.n17 VPWR.n9 9.3005
R85 VPWR.n19 VPWR.n18 9.3005
R86 VPWR.n20 VPWR.n7 9.3005
R87 VPWR.n22 VPWR.n21 9.3005
R88 VPWR.n23 VPWR.n6 9.3005
R89 VPWR.n25 VPWR.n24 9.3005
R90 VPWR.n26 VPWR.n5 9.3005
R91 VPWR.n30 VPWR.n29 9.3005
R92 VPWR.n31 VPWR.n4 9.3005
R93 VPWR.n33 VPWR.n32 9.3005
R94 VPWR.n34 VPWR.n3 9.3005
R95 VPWR.n36 VPWR.n35 9.3005
R96 VPWR.n38 VPWR.n37 9.3005
R97 VPWR.n39 VPWR.n0 9.3005
R98 VPWR.n41 VPWR.n40 8.45673
R99 VPWR.n29 VPWR.n28 6.99043
R100 VPWR.n38 VPWR.n2 4.51815
R101 VPWR.n12 VPWR.n10 2.0514
R102 VPWR.n14 VPWR.n13 1.50638
R103 VPWR VPWR.n41 0.163644
R104 VPWR.n41 VPWR.n0 0.144205
R105 VPWR.n16 VPWR.n10 0.122949
R106 VPWR.n17 VPWR.n16 0.122949
R107 VPWR.n18 VPWR.n17 0.122949
R108 VPWR.n18 VPWR.n7 0.122949
R109 VPWR.n22 VPWR.n7 0.122949
R110 VPWR.n23 VPWR.n22 0.122949
R111 VPWR.n24 VPWR.n23 0.122949
R112 VPWR.n24 VPWR.n5 0.122949
R113 VPWR.n30 VPWR.n5 0.122949
R114 VPWR.n31 VPWR.n30 0.122949
R115 VPWR.n32 VPWR.n31 0.122949
R116 VPWR.n32 VPWR.n3 0.122949
R117 VPWR.n36 VPWR.n3 0.122949
R118 VPWR.n37 VPWR.n36 0.122949
R119 VPWR.n37 VPWR.n0 0.122949
R120 a_544_485.n2 a_544_485.n1 600.128
R121 a_544_485.n0 a_544_485.t4 338.896
R122 a_544_485.n3 a_544_485.n2 308
R123 a_544_485.n2 a_544_485.n0 278.228
R124 a_544_485.n0 a_544_485.t5 181.821
R125 a_544_485.n1 a_544_485.t3 123.019
R126 a_544_485.n1 a_544_485.t0 70.9973
R127 a_544_485.n3 a_544_485.t2 46.4611
R128 a_544_485.n4 a_544_485.t1 25.6415
R129 a_544_485.n5 a_544_485.n4 21.6005
R130 a_544_485.n4 a_544_485.n3 16.1199
R131 a_651_503.t0 a_651_503.t1 112.572
R132 a_1226_296.t0 a_1226_296.n14 405.896
R133 a_1226_296.n3 a_1226_296.t8 291.075
R134 a_1226_296.n7 a_1226_296.t2 250.526
R135 a_1226_296.n0 a_1226_296.t3 240.197
R136 a_1226_296.n1 a_1226_296.t4 240.197
R137 a_1226_296.n10 a_1226_296.t5 240.197
R138 a_1226_296.n3 a_1226_296.n2 232.968
R139 a_1226_296.n14 a_1226_296.n3 184.257
R140 a_1226_296.n10 a_1226_296.t6 182.138
R141 a_1226_296.n7 a_1226_296.n6 179.947
R142 a_1226_296.n1 a_1226_296.n5 179.947
R143 a_1226_296.n0 a_1226_296.t7 179.947
R144 a_1226_296.n13 a_1226_296.t1 174.232
R145 a_1226_296.n8 a_1226_296.n4 165.189
R146 a_1226_296.n12 a_1226_296.n11 152
R147 a_1226_296.n9 a_1226_296.n4 152
R148 a_1226_296.n0 a_1226_296.n7 67.8456
R149 a_1226_296.n11 a_1226_296.n9 49.6611
R150 a_1226_296.n1 a_1226_296.n8 43.8187
R151 a_1226_296.n14 a_1226_296.n13 24.4711
R152 a_1226_296.n8 a_1226_296.n0 21.9096
R153 a_1226_296.n13 a_1226_296.n12 16.8732
R154 a_1226_296.n12 a_1226_296.n4 13.1884
R155 a_1226_296.n11 a_1226_296.n10 10.955
R156 a_1226_296.n9 a_1226_296.n1 5.84292
R157 Q.n5 Q.n4 585
R158 Q.n4 Q.n0 290.923
R159 Q.n3 Q.n1 250.518
R160 Q.n2 Q.t5 183.43
R161 Q.n2 Q.t4 147.944
R162 Q.n3 Q.n2 56.9923
R163 Q.n4 Q.t3 26.3844
R164 Q.n4 Q.t2 26.3844
R165 Q.n1 Q.t1 26.3844
R166 Q.n1 Q.t0 26.3844
R167 Q Q.n5 12.9944
R168 Q Q.n0 8.65194
R169 Q.n0 Q 5.59489
R170 Q Q.n3 2.52171
R171 Q.n5 Q 1.35808
R172 a_437_503.n1 a_437_503.n0 909.913
R173 a_437_503.n0 a_437_503.t2 123.659
R174 a_437_503.n0 a_437_503.t1 70.3576
R175 a_437_503.n1 a_437_503.t3 40.0005
R176 a_437_503.t0 a_437_503.n1 40.0005
R177 VNB.t7 VNB.t0 3637.8
R178 VNB.t8 VNB.t11 3360.63
R179 VNB.t4 VNB.t3 2124.93
R180 VNB.t10 VNB.t2 1836.22
R181 VNB.t5 VNB.t7 1443.57
R182 VNB.t6 VNB.t8 1351.18
R183 VNB VNB.t5 1143.31
R184 VNB.t2 VNB.t6 1097.11
R185 VNB.t9 VNB.t1 1097.11
R186 VNB.t11 VNB.t4 1062.47
R187 VNB.t0 VNB.t9 993.177
R188 VNB.t1 VNB.t10 831.496
R189 D.n0 D.t1 404.248
R190 D D.t0 317.464
R191 D.n0 D 10.3116
R192 D D.n0 2.84494
R193 VGND.n28 VGND.t0 367.163
R194 VGND.n10 VGND.t2 296.639
R195 VGND.n34 VGND.n1 221.518
R196 VGND.n21 VGND.n20 213.522
R197 VGND.n9 VGND.n8 205.559
R198 VGND.n20 VGND.t1 92.7278
R199 VGND.n1 VGND.t5 54.3248
R200 VGND.n20 VGND.t6 53.0654
R201 VGND.n35 VGND.n34 44.6887
R202 VGND.n14 VGND.n6 36.1417
R203 VGND.n18 VGND.n6 36.1417
R204 VGND.n19 VGND.n18 36.1417
R205 VGND.n22 VGND.n4 36.1417
R206 VGND.n26 VGND.n4 36.1417
R207 VGND.n27 VGND.n26 36.1417
R208 VGND.n32 VGND.n2 36.1417
R209 VGND.n33 VGND.n32 36.1417
R210 VGND.n14 VGND.n13 30.8711
R211 VGND.n8 VGND.t3 27.5681
R212 VGND.n12 VGND.n9 27.1064
R213 VGND.n28 VGND.n27 24.4711
R214 VGND.n28 VGND.n2 22.9652
R215 VGND.n8 VGND.t7 22.7032
R216 VGND.n1 VGND.t4 22.7032
R217 VGND.n13 VGND.n12 22.5887
R218 VGND.n21 VGND.n19 16.5652
R219 VGND.n33 VGND.n0 9.3005
R220 VGND.n32 VGND.n31 9.3005
R221 VGND.n30 VGND.n2 9.3005
R222 VGND.n29 VGND.n28 9.3005
R223 VGND.n27 VGND.n3 9.3005
R224 VGND.n26 VGND.n25 9.3005
R225 VGND.n24 VGND.n4 9.3005
R226 VGND.n23 VGND.n22 9.3005
R227 VGND.n19 VGND.n5 9.3005
R228 VGND.n18 VGND.n17 9.3005
R229 VGND.n16 VGND.n6 9.3005
R230 VGND.n15 VGND.n14 9.3005
R231 VGND.n13 VGND.n7 9.3005
R232 VGND.n12 VGND.n11 9.3005
R233 VGND.n10 VGND.n9 6.63016
R234 VGND.n22 VGND.n21 0.753441
R235 VGND.n34 VGND.n33 0.753441
R236 VGND.n11 VGND.n10 0.483449
R237 VGND.n11 VGND.n7 0.122949
R238 VGND.n15 VGND.n7 0.122949
R239 VGND.n16 VGND.n15 0.122949
R240 VGND.n17 VGND.n16 0.122949
R241 VGND.n17 VGND.n5 0.122949
R242 VGND.n23 VGND.n5 0.122949
R243 VGND.n24 VGND.n23 0.122949
R244 VGND.n25 VGND.n24 0.122949
R245 VGND.n25 VGND.n3 0.122949
R246 VGND.n29 VGND.n3 0.122949
R247 VGND.n30 VGND.n29 0.122949
R248 VGND.n31 VGND.n30 0.122949
R249 VGND.n31 VGND.n0 0.122949
R250 VGND.n35 VGND.n0 0.122949
R251 VGND VGND.n35 0.0617245
R252 a_206_368.n0 a_206_368.t5 1097.35
R253 a_206_368.n0 a_206_368.t4 582.323
R254 a_206_368.n2 a_206_368.t2 421.507
R255 a_206_368.n2 a_206_368.t3 364.13
R256 a_206_368.n3 a_206_368.n2 309.212
R257 a_206_368.n1 a_206_368.t0 248.32
R258 a_206_368.t1 a_206_368.n3 218.213
R259 a_206_368.n1 a_206_368.n0 152
R260 a_206_368.n3 a_206_368.n1 38.9855
R261 a_735_102.t0 a_735_102.t1 60.0005
R262 a_1141_508.t0 a_1141_508.t1 222.798
C0 a_1178_124# VPWR 7.43e-19
C1 VPB VPWR 0.258623f
C2 a_1178_124# VGND 0.004565f
C3 VPB CLK 0.0398f
C4 VPWR CLK 0.015078f
C5 VPB D 0.098058f
C6 VPWR D 0.008282f
C7 VPB VGND 0.019289f
C8 VPWR VGND 0.163639f
C9 VPB Q 0.012697f
C10 CLK VGND 0.014066f
C11 VPWR Q 0.396303f
C12 D VGND 0.008318f
C13 VGND Q 0.274629f
C14 Q VNB 0.037563f
C15 VGND VNB 1.14199f
C16 D VNB 0.147896f
C17 CLK VNB 0.163662f
C18 VPWR VNB 0.922515f
C19 VPB VNB 2.22754f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrbn_2 VNB VPB VPWR VGND D GATE_N RESET_B Q Q_N
X0 a_790_74.t1 a_363_74.t2 a_670_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.122 ps=1.09 w=0.42 l=0.15
X1 a_783_508.t1 a_230_74.t2 a_670_74.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1739 ps=1.4 w=0.42 l=0.15
X2 Q.t1 a_838_48# VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1628 ps=1.18 w=0.74 l=0.15
X3 VGND.t8 a_230_74.t3 a_363_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1917 pd=1.3 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 VPWR.t1 a_1446_368.t2 Q_N.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t4 a_838_48# a_783_508.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.745 as=0.09975 ps=0.895 w=0.42 l=0.15
X6 Q_N.t2 a_1446_368.t3 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 VGND.t3 a_838_48# Q.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1245 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_230_74.t0 GATE_N.t0 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X9 a_1446_368.t1 a_838_48# VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.1934 ps=1.475 w=1 l=0.15
X10 a_1066_74.t0 a_670_74.t4 a_838_48# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 a_670_74.t0 a_363_74.t3 a_595_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1739 pd=1.4 as=0.12 ps=1.24 w=1 l=0.15
X12 a_592_74.t0 a_27_112.t2 VGND.t10 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1917 ps=1.3 w=0.64 l=0.15
X13 VGND.t0 a_1446_368.t4 Q_N.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X14 a_230_74.t1 GATE_N.t1 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.2226 ps=1.37 w=0.84 l=0.15
X15 VPWR.t5 a_838_48# Q.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_838_48# a_670_74.t5 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.224 ps=1.745 w=1.12 l=0.15
X17 Q_N.t0 a_1446_368.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2109 ps=2.05 w=0.74 l=0.15
X18 Q a_838_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X19 a_595_392.t0 a_27_112.t3 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.25245 ps=1.64 w=1 l=0.15
X20 VPWR.t9 D.t0 a_27_112.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2226 pd=1.37 as=0.2478 ps=2.27 w=0.84 l=0.15
X21 VPWR.t8 a_230_74.t4 a_363_74.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.25245 pd=1.64 as=0.383 ps=2.88 w=0.84 l=0.15
X22 VPWR RESET_B a_838_48# VPB sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1736 ps=1.43 w=1.12 l=0.15
X23 VGND.t6 RESET_B.t0 a_1066_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1628 pd=1.18 as=0.0888 ps=0.98 w=0.74 l=0.15
X24 VGND.t9 D.t1 a_27_112.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X25 a_670_74.t3 a_230_74.t5 a_592_74.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.09 as=0.0768 ps=0.88 w=0.64 l=0.15
X26 VGND.t4 a_838_48# a_790_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 a_1446_368.t0 a_838_48# VGND.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1245 ps=1.09 w=0.64 l=0.15
R0 a_363_74.t1 a_363_74.n1 920.606
R1 a_363_74.n0 a_363_74.t3 443.44
R2 a_363_74.n1 a_363_74.n0 305.729
R3 a_363_74.n0 a_363_74.t2 231.361
R4 a_363_74.n1 a_363_74.t0 118.38
R5 a_670_74.n3 a_670_74.n2 691.846
R6 a_670_74.n2 a_670_74.n0 302.399
R7 a_670_74.n2 a_670_74.n1 239.042
R8 a_670_74.n1 a_670_74.t5 226.809
R9 a_670_74.n1 a_670_74.t4 198.204
R10 a_670_74.n3 a_670_74.t2 114.918
R11 a_670_74.n0 a_670_74.t1 64.2862
R12 a_670_74.n0 a_670_74.t3 52.0094
R13 a_670_74.t0 a_670_74.n3 30.5355
R14 a_790_74.t0 a_790_74.t1 68.5719
R15 VNB VNB.n0 5300.79
R16 VNB.t11 VNB.t9 2681.44
R17 VNB.t2 VNB.t1 2286.61
R18 VNB.t3 VNB.t7 2286.61
R19 VNB.t9 VNB.t10 1413.85
R20 VNB.t12 VNB.t6 1385.83
R21 VNB.t8 VNB.t5 1362.73
R22 VNB.n0 VNB.t13 1362.73
R23 VNB.t10 VNB 1206.65
R24 VNB.t4 VNB.t2 1154.86
R25 VNB.t1 VNB.t0 1085.56
R26 VNB.t5 VNB.t4 993.177
R27 VNB.t7 VNB.t8 900.788
R28 VNB.t6 VNB.t3 900.788
R29 VNB.t13 VNB.t12 900.788
R30 VNB.n0 VNB.t11 292.522
R31 a_230_74.t1 a_230_74.n3 756.328
R32 a_230_74.n0 a_230_74.t2 480.577
R33 a_230_74.n0 a_230_74.t5 314.274
R34 a_230_74.n1 a_230_74.t4 271.488
R35 a_230_74.n3 a_230_74.t0 218.216
R36 a_230_74.n1 a_230_74.t3 176.964
R37 a_230_74.n2 a_230_74.n1 152
R38 a_230_74.n3 a_230_74.n2 111.099
R39 a_230_74.n2 a_230_74.n0 59.9898
R40 a_783_508.t0 a_783_508.t1 222.798
R41 VPB.t7 VPB.t1 720.162
R42 VPB.t8 VPB.t9 559.274
R43 VPB.t2 VPB.t5 515.861
R44 VPB.t3 VPB.t7 395.834
R45 VPB.t11 VPB.t8 347.312
R46 VPB.t10 VPB.t3 319.221
R47 VPB.t9 VPB.t0 316.668
R48 VPB.t6 VPB.t10 280.914
R49 VPB.t1 VPB.t2 257.93
R50 VPB VPB.t11 257.93
R51 VPB.t5 VPB.t4 229.839
R52 VPB.t0 VPB.t6 199.195
R53 VGND.n20 VGND.t4 252.137
R54 VGND.n27 VGND.n26 185
R55 VGND.n9 VGND.t0 176.427
R56 VGND.n8 VGND.t1 160.286
R57 VGND.n13 VGND.n12 122.195
R58 VGND.n35 VGND.n34 120.007
R59 VGND.n6 VGND.n5 116.154
R60 VGND.n26 VGND.t8 55.4736
R61 VGND.n34 VGND.t9 51.1927
R62 VGND.n5 VGND.t2 48.6491
R63 VGND.n26 VGND.t10 45.938
R64 VGND.n12 VGND.t5 39.3755
R65 VGND.n19 VGND.n18 36.1417
R66 VGND.n24 VGND.n3 36.1417
R67 VGND.n25 VGND.n24 36.1417
R68 VGND.n32 VGND.n1 36.1417
R69 VGND.n33 VGND.n32 36.1417
R70 VGND.n14 VGND.n6 34.2593
R71 VGND.n34 VGND.t7 32.4397
R72 VGND.n13 VGND.n11 29.7417
R73 VGND.n20 VGND.n19 29.7417
R74 VGND.n11 VGND.n8 25.224
R75 VGND.n28 VGND.n25 25.1031
R76 VGND.n20 VGND.n3 23.7181
R77 VGND.n14 VGND.n13 22.9652
R78 VGND.n5 VGND.t6 22.7032
R79 VGND.n12 VGND.t3 22.6611
R80 VGND.n35 VGND.n33 18.4476
R81 VGND.n27 VGND.n1 15.2105
R82 VGND.n18 VGND.n6 13.177
R83 VGND.n11 VGND.n10 9.3005
R84 VGND.n13 VGND.n7 9.3005
R85 VGND.n15 VGND.n14 9.3005
R86 VGND.n16 VGND.n6 9.3005
R87 VGND.n18 VGND.n17 9.3005
R88 VGND.n19 VGND.n4 9.3005
R89 VGND.n21 VGND.n20 9.3005
R90 VGND.n22 VGND.n3 9.3005
R91 VGND.n24 VGND.n23 9.3005
R92 VGND.n25 VGND.n2 9.3005
R93 VGND.n29 VGND.n28 9.3005
R94 VGND.n30 VGND.n1 9.3005
R95 VGND.n32 VGND.n31 9.3005
R96 VGND.n33 VGND.n0 9.3005
R97 VGND.n36 VGND.n35 7.46433
R98 VGND.n9 VGND.n8 6.90969
R99 VGND.n28 VGND.n27 1.40196
R100 VGND.n10 VGND.n9 0.561104
R101 VGND VGND.n36 0.160491
R102 VGND.n36 VGND.n0 0.147317
R103 VGND.n10 VGND.n7 0.122949
R104 VGND.n15 VGND.n7 0.122949
R105 VGND.n16 VGND.n15 0.122949
R106 VGND.n17 VGND.n16 0.122949
R107 VGND.n17 VGND.n4 0.122949
R108 VGND.n21 VGND.n4 0.122949
R109 VGND.n22 VGND.n21 0.122949
R110 VGND.n23 VGND.n22 0.122949
R111 VGND.n23 VGND.n2 0.122949
R112 VGND.n29 VGND.n2 0.122949
R113 VGND.n30 VGND.n29 0.122949
R114 VGND.n31 VGND.n30 0.122949
R115 VGND.n31 VGND.n0 0.122949
R116 Q.n1 Q.t2 922.851
R117 Q.n1 Q.n0 185
R118 Q.n0 Q.t0 22.7032
R119 Q.n0 Q.t1 22.7032
R120 Q Q.n1 4.26717
R121 a_1446_368.n1 a_1446_368.t2 330.476
R122 a_1446_368.n0 a_1446_368.t3 264.211
R123 a_1446_368.t1 a_1446_368.n2 248.911
R124 a_1446_368.n1 a_1446_368.t4 174.898
R125 a_1446_368.n0 a_1446_368.t5 154.24
R126 a_1446_368.n2 a_1446_368.t0 146.421
R127 a_1446_368.n2 a_1446_368.n0 116.603
R128 a_1446_368.n0 a_1446_368.n1 106.478
R129 Q_N.n2 Q_N 589.572
R130 Q_N.n2 Q_N.n0 585
R131 Q_N.n3 Q_N.n2 585
R132 Q_N Q_N.n1 255.261
R133 Q_N.n2 Q_N.t3 26.3844
R134 Q_N.n2 Q_N.t2 26.3844
R135 Q_N.n1 Q_N.t1 25.9464
R136 Q_N.n1 Q_N.t0 25.9464
R137 Q_N Q_N.n3 12.2519
R138 Q_N Q_N.n0 10.6062
R139 Q_N Q_N.n0 2.92621
R140 Q_N.n3 Q_N 1.2805
R141 VPWR.n29 VPWR.n4 698.312
R142 VPWR.n35 VPWR.n1 625.283
R143 VPWR.n14 VPWR.n9 610.212
R144 VPWR.n22 VPWR.n21 585
R145 VPWR.n11 VPWR.t1 266.248
R146 VPWR.n10 VPWR.t0 259.171
R147 VPWR.n21 VPWR.t4 136.024
R148 VPWR.n21 VPWR.t6 133.179
R149 VPWR.n1 VPWR.t7 89.1195
R150 VPWR.n4 VPWR.t8 65.6672
R151 VPWR.n9 VPWR.t3 40.3855
R152 VPWR.n33 VPWR.n2 36.1417
R153 VPWR.n34 VPWR.n33 36.1417
R154 VPWR.n27 VPWR.n5 36.1417
R155 VPWR.n28 VPWR.n27 36.1417
R156 VPWR.n4 VPWR.t2 35.5684
R157 VPWR.n35 VPWR.n34 35.3887
R158 VPWR.n1 VPWR.t9 35.1791
R159 VPWR.n23 VPWR.n5 34.092
R160 VPWR.n20 VPWR.n19 30.2855
R161 VPWR.n14 VPWR.n13 30.1181
R162 VPWR.n9 VPWR.t5 27.6909
R163 VPWR.n29 VPWR.n28 27.4829
R164 VPWR.n15 VPWR.n7 25.6005
R165 VPWR.n13 VPWR.n10 25.224
R166 VPWR.n19 VPWR.n7 21.8358
R167 VPWR.n29 VPWR.n2 19.9534
R168 VPWR.n15 VPWR.n14 17.3181
R169 VPWR.n13 VPWR.n12 9.3005
R170 VPWR.n14 VPWR.n8 9.3005
R171 VPWR.n16 VPWR.n15 9.3005
R172 VPWR.n17 VPWR.n7 9.3005
R173 VPWR.n19 VPWR.n18 9.3005
R174 VPWR.n20 VPWR.n6 9.3005
R175 VPWR.n24 VPWR.n23 9.3005
R176 VPWR.n25 VPWR.n5 9.3005
R177 VPWR.n27 VPWR.n26 9.3005
R178 VPWR.n28 VPWR.n3 9.3005
R179 VPWR.n30 VPWR.n29 9.3005
R180 VPWR.n31 VPWR.n2 9.3005
R181 VPWR.n33 VPWR.n32 9.3005
R182 VPWR.n34 VPWR.n0 9.3005
R183 VPWR.n36 VPWR.n35 8.45673
R184 VPWR.n11 VPWR.n10 6.95806
R185 VPWR.n23 VPWR.n22 4.51815
R186 VPWR.n22 VPWR.n20 3.51423
R187 VPWR.n12 VPWR.n11 0.546775
R188 VPWR VPWR.n36 0.163644
R189 VPWR.n36 VPWR.n0 0.144205
R190 VPWR.n12 VPWR.n8 0.122949
R191 VPWR.n16 VPWR.n8 0.122949
R192 VPWR.n17 VPWR.n16 0.122949
R193 VPWR.n18 VPWR.n17 0.122949
R194 VPWR.n18 VPWR.n6 0.122949
R195 VPWR.n24 VPWR.n6 0.122949
R196 VPWR.n25 VPWR.n24 0.122949
R197 VPWR.n26 VPWR.n25 0.122949
R198 VPWR.n26 VPWR.n3 0.122949
R199 VPWR.n30 VPWR.n3 0.122949
R200 VPWR.n31 VPWR.n30 0.122949
R201 VPWR.n32 VPWR.n31 0.122949
R202 VPWR.n32 VPWR.n0 0.122949
R203 GATE_N.n0 GATE_N.t1 235.516
R204 GATE_N.n0 GATE_N.t0 212.588
R205 GATE_N GATE_N.n0 68.7712
R206 a_1066_74.t0 a_1066_74.t1 38.9194
R207 a_595_392.t0 a_595_392.t1 47.2805
R208 a_27_112.n1 a_27_112.n0 411.488
R209 a_27_112.t1 a_27_112.n1 391.995
R210 a_27_112.n1 a_27_112.t0 304.394
R211 a_27_112.n0 a_27_112.t2 274.74
R212 a_27_112.n0 a_27_112.t3 231.629
R213 a_592_74.t0 a_592_74.t1 45.0005
R214 D.n0 D.t0 234.22
R215 D.n0 D.t1 180.798
R216 D D.n0 68.4106
R217 RESET_B.n1 RESET_B.n0 285.719
R218 RESET_B.n1 RESET_B.t0 178.34
R219 RESET_B RESET_B.n1 158.227
C0 a_838_48# Q_N 5.16e-19
C1 VPWR Q 0.016789f
C2 RESET_B VGND 0.056102f
C3 VPWR Q_N 0.223435f
C4 RESET_B Q 0.033419f
C5 VGND Q 0.0675f
C6 VPB D 0.062839f
C7 VGND Q_N 0.063967f
C8 a_838_48# VPB 0.243544f
C9 VPB GATE_N 0.070318f
C10 a_838_48# D 2.75e-20
C11 VPB VPWR 0.278575f
C12 D GATE_N 0.12289f
C13 a_838_48# GATE_N 4.64e-19
C14 VPB RESET_B 0.03063f
C15 D VPWR 0.015701f
C16 a_838_48# VPWR 0.333316f
C17 GATE_N VPWR 0.009111f
C18 VPB VGND 0.020771f
C19 a_838_48# RESET_B 0.139236f
C20 VPB Q 0.003926f
C21 D VGND 0.036328f
C22 a_838_48# VGND 0.224843f
C23 VPB Q_N 0.007069f
C24 GATE_N VGND 0.021641f
C25 VPWR RESET_B 0.019078f
C26 a_838_48# Q 0.160408f
C27 VPWR VGND 0.163088f
C28 Q_N VNB 0.036197f
C29 Q VNB 0.010076f
C30 VGND VNB 1.13751f
C31 RESET_B VNB 0.107678f
C32 VPWR VNB 0.870523f
C33 GATE_N VNB 0.119399f
C34 D VNB 0.150131f
C35 VPB VNB 2.13048f
C36 a_838_48# VNB 0.486029f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrbp_2 VNB VPB VPWR VGND GATE D RESET_B Q_N Q
X0 a_569_80.t1 a_27_112.t2 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.188225 ps=1.415 w=0.64 l=0.15
X1 VPWR.t0 D.t0 a_27_112.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.22785 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 VGND.t2 a_230_74.t2 a_363_82.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.188225 pd=1.415 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 VPWR.t4 a_1449_368.t2 Q_N.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Q_N.t2 a_1449_368.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2159 ps=1.52 w=1.12 l=0.15
X5 VGND.t3 a_821_98.t3 Q.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VPWR.t8 RESET_B.t0 a_821_98.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2128 pd=1.5 as=0.196 ps=1.47 w=1.12 l=0.15
X7 a_230_74.t0 GATE.t0 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X8 VPWR.t6 a_230_74.t3 a_363_82.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2028 pd=1.42 as=0.2478 ps=2.27 w=0.84 l=0.15
X9 VGND.t4 a_821_98.t4 a_1449_368.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1469 pd=1.16 as=0.1824 ps=1.85 w=0.64 l=0.15
X10 a_641_80.t3 a_230_74.t4 a_566_392.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1664 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND RESET_B a_1049_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0888 ps=0.98 w=0.74 l=0.15
X12 VGND.t0 a_1449_368.t4 Q_N.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_821_98.t2 a_641_80.t4 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.22085 ps=1.73 w=1.12 l=0.15
X14 a_566_392.t1 a_27_112.t3 VPWR.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.2028 ps=1.42 w=1 l=0.15
X15 a_757_508.t0 a_363_82.t2 a_641_80.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.10605 pd=0.925 as=0.1664 ps=1.385 w=0.42 l=0.15
X16 VGND.t5 a_821_98.t5 a_773_124.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X17 VPWR.t7 a_821_98.t6 a_757_508.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.22085 pd=1.73 as=0.10605 ps=0.925 w=0.42 l=0.15
X18 VPWR.t1 a_821_98.t7 a_1449_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2159 pd=1.52 as=0.295 ps=2.59 w=1 l=0.15
X19 a_641_80.t0 a_363_82.t3 a_569_80.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1346 pd=1.15 as=0.0672 ps=0.85 w=0.64 l=0.15
X20 a_773_124.t0 a_230_74.t5 a_641_80.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1346 ps=1.15 w=0.42 l=0.15
X21 Q_N.t0 a_1449_368.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1469 ps=1.16 w=0.74 l=0.15
X22 a_230_74.t1 GATE.t1 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.2898 pd=2.37 as=0.22785 ps=1.52 w=0.84 l=0.15
X23 VGND.t7 D.t1 a_27_112.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X24 VPWR.t2 a_821_98.t8 Q.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X25 a_1049_74# a_641_80.t5 a_821_98.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X26 Q.t1 a_821_98.t9 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2128 ps=1.5 w=1.12 l=0.15
R0 a_27_112.t0 a_27_112.n1 776.111
R1 a_27_112.t0 a_27_112.n2 761.966
R2 a_27_112.n1 a_27_112.n0 338
R3 a_27_112.n2 a_27_112.t1 293.642
R4 a_27_112.n0 a_27_112.t2 263.092
R5 a_27_112.n0 a_27_112.t3 229.619
R6 a_27_112.n2 a_27_112.n1 11.7338
R7 VGND.n19 VGND.t5 257.195
R8 VGND.n12 VGND.t3 242.715
R9 VGND.n26 VGND.n25 218.752
R10 VGND.n9 VGND.t0 178.799
R11 VGND.n8 VGND.n7 119.629
R12 VGND.n34 VGND.n33 119.475
R13 VGND.n33 VGND.t7 51.1943
R14 VGND.n25 VGND.t2 45.7097
R15 VGND.n7 VGND.t4 39.3755
R16 VGND.n13 VGND.n5 36.1417
R17 VGND.n18 VGND.n17 36.1417
R18 VGND.n19 VGND.n18 36.1417
R19 VGND.n23 VGND.n3 36.1417
R20 VGND.n24 VGND.n23 36.1417
R21 VGND.n27 VGND.n24 36.1417
R22 VGND.n31 VGND.n1 36.1417
R23 VGND.n32 VGND.n31 36.1417
R24 VGND.n7 VGND.t1 35.7861
R25 VGND.n12 VGND.n11 34.6358
R26 VGND.n33 VGND.t8 32.4381
R27 VGND.n25 VGND.t6 26.0934
R28 VGND.n11 VGND.n8 22.9652
R29 VGND.n34 VGND.n32 18.4476
R30 VGND.n26 VGND.n1 15.1848
R31 VGND.n13 VGND.n12 12.8005
R32 VGND.n17 VGND.n5 11.2946
R33 VGND.n19 VGND.n3 11.2946
R34 VGND.n11 VGND.n10 9.3005
R35 VGND.n12 VGND.n6 9.3005
R36 VGND.n14 VGND.n13 9.3005
R37 VGND.n15 VGND.n5 9.3005
R38 VGND.n17 VGND.n16 9.3005
R39 VGND.n18 VGND.n4 9.3005
R40 VGND.n20 VGND.n19 9.3005
R41 VGND.n21 VGND.n3 9.3005
R42 VGND.n23 VGND.n22 9.3005
R43 VGND.n24 VGND.n2 9.3005
R44 VGND.n28 VGND.n27 9.3005
R45 VGND.n29 VGND.n1 9.3005
R46 VGND.n31 VGND.n30 9.3005
R47 VGND.n32 VGND.n0 9.3005
R48 VGND.n35 VGND.n34 7.46433
R49 VGND.n9 VGND.n8 6.74444
R50 VGND.n27 VGND.n26 4.39646
R51 VGND.n10 VGND.n9 0.585372
R52 VGND VGND.n35 0.160491
R53 VGND.n35 VGND.n0 0.147317
R54 VGND.n10 VGND.n6 0.122949
R55 VGND.n14 VGND.n6 0.122949
R56 VGND.n15 VGND.n14 0.122949
R57 VGND.n16 VGND.n15 0.122949
R58 VGND.n16 VGND.n4 0.122949
R59 VGND.n20 VGND.n4 0.122949
R60 VGND.n21 VGND.n20 0.122949
R61 VGND.n22 VGND.n21 0.122949
R62 VGND.n22 VGND.n2 0.122949
R63 VGND.n28 VGND.n2 0.122949
R64 VGND.n29 VGND.n28 0.122949
R65 VGND.n30 VGND.n29 0.122949
R66 VGND.n30 VGND.n0 0.122949
R67 a_569_80.t0 a_569_80.t1 39.3755
R68 VNB.t9 VNB.t5 3141.21
R69 VNB.t11 VNB.t3 2540.68
R70 VNB.t5 VNB.t6 2529.13
R71 VNB.t7 VNB.t9 2286.61
R72 VNB.t2 VNB.t4 1524.41
R73 VNB.t3 VNB.t8 1374.28
R74 VNB.t10 VNB.t11 1339.63
R75 VNB.t6 VNB.t1 1316.54
R76 VNB VNB.t10 1143.31
R77 VNB.t1 VNB.t0 993.177
R78 VNB.t4 VNB.t7 900.788
R79 VNB.t8 VNB.t2 831.496
R80 D.n0 D.t1 221.012
R81 D.n0 D.t0 210.569
R82 D D.n0 153.745
R83 VPWR.n36 VPWR.n1 647.192
R84 VPWR.n30 VPWR.n4 604.112
R85 VPWR.n23 VPWR.n22 585
R86 VPWR.n15 VPWR.t2 343.724
R87 VPWR.n12 VPWR.t4 265.976
R88 VPWR.n11 VPWR.n10 227.118
R89 VPWR.n8 VPWR.n7 221.766
R90 VPWR.n22 VPWR.t7 143.06
R91 VPWR.n22 VPWR.t10 119.108
R92 VPWR.n4 VPWR.t6 58.6315
R93 VPWR.n1 VPWR.t11 55.1136
R94 VPWR.n1 VPWR.t0 55.1136
R95 VPWR.n10 VPWR.t1 39.4005
R96 VPWR.n10 VPWR.t5 37.4007
R97 VPWR.n34 VPWR.n2 36.1417
R98 VPWR.n35 VPWR.n34 36.1417
R99 VPWR.n28 VPWR.n5 36.1417
R100 VPWR.n29 VPWR.n28 36.1417
R101 VPWR.n7 VPWR.t8 35.1791
R102 VPWR.n21 VPWR.n20 34.6776
R103 VPWR.n4 VPWR.t9 33.6733
R104 VPWR.n15 VPWR.n14 33.5064
R105 VPWR.n30 VPWR.n29 32.0005
R106 VPWR.n7 VPWR.t3 31.6612
R107 VPWR.n16 VPWR.n8 31.2476
R108 VPWR.n24 VPWR.n5 28.2358
R109 VPWR.n14 VPWR.n11 21.4593
R110 VPWR.n36 VPWR.n35 16.5652
R111 VPWR.n20 VPWR.n8 16.1887
R112 VPWR.n16 VPWR.n15 13.9299
R113 VPWR.n30 VPWR.n2 12.8005
R114 VPWR.n14 VPWR.n13 9.3005
R115 VPWR.n15 VPWR.n9 9.3005
R116 VPWR.n17 VPWR.n16 9.3005
R117 VPWR.n18 VPWR.n8 9.3005
R118 VPWR.n20 VPWR.n19 9.3005
R119 VPWR.n21 VPWR.n6 9.3005
R120 VPWR.n25 VPWR.n24 9.3005
R121 VPWR.n26 VPWR.n5 9.3005
R122 VPWR.n28 VPWR.n27 9.3005
R123 VPWR.n29 VPWR.n3 9.3005
R124 VPWR.n31 VPWR.n30 9.3005
R125 VPWR.n32 VPWR.n2 9.3005
R126 VPWR.n34 VPWR.n33 9.3005
R127 VPWR.n35 VPWR.n0 9.3005
R128 VPWR.n37 VPWR.n36 7.53404
R129 VPWR.n12 VPWR.n11 6.8344
R130 VPWR.n23 VPWR.n21 4.93645
R131 VPWR.n24 VPWR.n23 3.09592
R132 VPWR.n13 VPWR.n12 0.569119
R133 VPWR VPWR.n37 0.161409
R134 VPWR.n37 VPWR.n0 0.146411
R135 VPWR.n13 VPWR.n9 0.122949
R136 VPWR.n17 VPWR.n9 0.122949
R137 VPWR.n18 VPWR.n17 0.122949
R138 VPWR.n19 VPWR.n18 0.122949
R139 VPWR.n19 VPWR.n6 0.122949
R140 VPWR.n25 VPWR.n6 0.122949
R141 VPWR.n26 VPWR.n25 0.122949
R142 VPWR.n27 VPWR.n26 0.122949
R143 VPWR.n27 VPWR.n3 0.122949
R144 VPWR.n31 VPWR.n3 0.122949
R145 VPWR.n32 VPWR.n31 0.122949
R146 VPWR.n33 VPWR.n32 0.122949
R147 VPWR.n33 VPWR.n0 0.122949
R148 VPB.t13 VPB.t6 541.399
R149 VPB.t2 VPB.t1 515.861
R150 VPB.t8 VPB.t12 388.173
R151 VPB.t11 VPB.t8 334.543
R152 VPB.t0 VPB.t13 316.668
R153 VPB.t6 VPB.t10 291.13
R154 VPB.t1 VPB.t5 280.914
R155 VPB.t7 VPB.t11 273.253
R156 VPB.t9 VPB.t3 270.7
R157 VPB VPB.t0 257.93
R158 VPB.t12 VPB.t9 255.376
R159 VPB.t5 VPB.t4 229.839
R160 VPB.t3 VPB.t2 229.839
R161 VPB.t10 VPB.t7 214.517
R162 a_230_74.t1 a_230_74.n2 775.958
R163 a_230_74.t5 a_230_74.t4 661.947
R164 a_230_74.n0 a_230_74.t5 425.043
R165 a_230_74.n1 a_230_74.t3 284.916
R166 a_230_74.n2 a_230_74.n1 250.007
R167 a_230_74.n1 a_230_74.t2 194.751
R168 a_230_74.n0 a_230_74.t0 133.702
R169 a_230_74.n2 a_230_74.n0 35.4488
R170 a_363_82.t1 a_363_82.n1 828.385
R171 a_363_82.n0 a_363_82.t2 476.577
R172 a_363_82.n0 a_363_82.t3 314.274
R173 a_363_82.n1 a_363_82.t0 296.377
R174 a_363_82.n1 a_363_82.n0 61.0989
R175 a_1449_368.t0 a_1449_368.n3 247.167
R176 a_1449_368.n0 a_1449_368.t2 240.197
R177 a_1449_368.n2 a_1449_368.t3 240.197
R178 a_1449_368.n3 a_1449_368.n2 190.792
R179 a_1449_368.n0 a_1449_368.t4 181.407
R180 a_1449_368.n1 a_1449_368.t5 179.947
R181 a_1449_368.n3 a_1449_368.t1 146.071
R182 a_1449_368.n1 a_1449_368.n0 61.346
R183 a_1449_368.n2 a_1449_368.n1 4.38232
R184 Q_N Q_N.n0 204.428
R185 Q_N Q_N.n1 159.339
R186 Q_N.n0 Q_N.t3 26.3844
R187 Q_N.n0 Q_N.t2 26.3844
R188 Q_N.n1 Q_N.t1 22.7032
R189 Q_N.n1 Q_N.t0 22.7032
R190 a_821_98.n7 a_821_98.t5 373.579
R191 a_821_98.n1 a_821_98.t8 240.197
R192 a_821_98.n4 a_821_98.t9 240.197
R193 a_821_98.n0 a_821_98.t7 220.917
R194 a_821_98.n9 a_821_98.n8 199.038
R195 a_821_98.n6 a_821_98.t1 194.022
R196 a_821_98.n4 a_821_98.n3 187.981
R197 a_821_98.n8 a_821_98.n7 180.145
R198 a_821_98.n2 a_821_98.t3 179.947
R199 a_821_98.n0 a_821_98.t4 165.341
R200 a_821_98.n7 a_821_98.t6 154.508
R201 a_821_98.n1 a_821_98.n0 147.522
R202 a_821_98.n6 a_821_98.n5 116.805
R203 a_821_98.n9 a_821_98.t2 35.1791
R204 a_821_98.t0 a_821_98.n9 26.3844
R205 a_821_98.n5 a_821_98.n4 25.6895
R206 a_821_98.n5 a_821_98.n2 22.3626
R207 a_821_98.n2 a_821_98.n1 10.955
R208 a_821_98.n8 a_821_98.n6 7.93372
R209 Q Q.n0 285.245
R210 Q Q.t0 184.716
R211 Q.n0 Q.t2 26.3844
R212 Q.n0 Q.t1 26.3844
R213 RESET_B.n1 RESET_B.t0 285.719
R214 RESET_B.n1 RESET_B.n0 178.34
R215 RESET_B RESET_B.n1 158.4
R216 GATE.n0 GATE.t1 272.866
R217 GATE.n0 GATE.t0 178.34
R218 GATE GATE.n0 159.226
R219 a_566_392.t0 a_566_392.t1 53.1905
R220 a_641_80.n3 a_641_80.n2 386
R221 a_641_80.n2 a_641_80.n1 284.182
R222 a_641_80.n2 a_641_80.n0 251.636
R223 a_641_80.n1 a_641_80.t4 226.809
R224 a_641_80.n1 a_641_80.t5 203.762
R225 a_641_80.n3 a_641_80.t1 123.823
R226 a_641_80.n0 a_641_80.t2 72.8576
R227 a_641_80.n0 a_641_80.t0 60.5809
R228 a_641_80.t3 a_641_80.n3 17.9641
R229 a_757_508.t0 a_757_508.t1 236.869
R230 a_773_124.t0 a_773_124.t1 68.5719
C0 a_1049_74# RESET_B 9.21e-19
C1 VGND Q 0.168631f
C2 VPB VPWR 0.287186f
C3 VGND Q_N 0.168325f
C4 VPB RESET_B 0.030658f
C5 VPWR RESET_B 0.019514f
C6 VPB D 0.049924f
C7 a_1049_74# VGND 0.009369f
C8 a_1049_74# Q 3.96e-19
C9 VPWR D 0.012906f
C10 VPB GATE 0.047181f
C11 VPB VGND 0.021656f
C12 VPWR GATE 0.010471f
C13 VPWR VGND 0.16235f
C14 VPB Q 0.009483f
C15 VPWR Q 0.191634f
C16 VPB Q_N 0.007005f
C17 D GATE 0.056963f
C18 RESET_B VGND 0.036718f
C19 RESET_B Q 0.003154f
C20 VPWR Q_N 0.234553f
C21 D VGND 0.027167f
C22 GATE VGND 0.021211f
C23 a_1049_74# VPWR 8.71e-19
C24 Q_N VNB 0.03086f
C25 Q VNB 0.020048f
C26 VGND VNB 1.14353f
C27 GATE VNB 0.11975f
C28 D VNB 0.142924f
C29 RESET_B VNB 0.105935f
C30 VPWR VNB 0.876328f
C31 VPB VNB 2.1204f
.ends

* NGSPICE file created from sky130_fd_sc_hs__dlrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtn_1 VNB VPB VPWR VGND D GATE_N RESET_B Q
X0 VGND.t0 RESET_B.t0 a_1139_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.163525 pd=1.185 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 Q.t0 a_897_406.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2382 ps=1.555 w=1.12 l=0.15
X2 a_681_74.t1 a_27_136.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.398075 ps=1.925 w=0.64 l=0.15
X3 a_654_392.t3 a_357_392.t2 a_570_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.20145 pd=1.545 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t5 a_897_406.t3 a_854_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1239 pd=1.43 as=0.05775 ps=0.695 w=0.42 l=0.15
X5 a_570_392.t0 a_27_136.t3 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.24665 ps=1.6 w=1 l=0.15
X6 VPWR.t1 a_897_406.t4 a_793_508.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2234 pd=1.885 as=0.11235 ps=0.955 w=0.42 l=0.15
X7 a_897_406.t1 a_654_392.t4 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.235 pd=1.47 as=0.2234 ps=1.885 w=1 l=0.15
X8 VGND.t4 a_232_98.t2 a_357_392.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.398075 pd=1.925 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 VPWR.t7 a_232_98.t3 a_357_392.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.24665 pd=1.6 as=0.2478 ps=2.27 w=0.84 l=0.15
X10 VPWR.t2 RESET_B.t1 a_897_406.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.235 ps=1.47 w=1 l=0.15
X11 VGND.t3 D.t0 a_27_136.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.200625 pd=1.49 as=0.15675 ps=1.67 w=0.55 l=0.15
X12 a_232_98.t1 GATE_N.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.198125 ps=1.315 w=0.84 l=0.15
X13 a_793_508.t1 a_232_98.t4 a_654_392.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.11235 pd=0.955 as=0.20145 ps=1.545 w=0.42 l=0.15
X14 a_232_98.t0 GATE_N.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.200625 ps=1.49 w=0.74 l=0.15
X15 a_854_74.t1 a_357_392.t3 a_654_392.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.05775 pd=0.695 as=0.09575 ps=0.965 w=0.42 l=0.15
X16 VPWR.t6 D.t1 a_27_136.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.198125 pd=1.315 as=0.2478 ps=2.27 w=0.84 l=0.15
X17 a_654_392.t0 a_232_98.t5 a_681_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.09575 pd=0.965 as=0.0768 ps=0.88 w=0.64 l=0.15
R0 RESET_B.n0 RESET_B.t1 266.44
R1 RESET_B.n0 RESET_B.t0 178.34
R2 RESET_B RESET_B.n0 158.4
R3 VGND.n1 VGND.n0 275.382
R4 VGND.n7 VGND.t5 245.817
R5 VGND.n16 VGND.n15 185
R6 VGND.n14 VGND.n3 185
R7 VGND.n6 VGND.t0 156.952
R8 VGND.n15 VGND.n14 74.4583
R9 VGND.n0 VGND.t3 55.6369
R10 VGND.n8 VGND.n5 36.1417
R11 VGND.n12 VGND.n5 36.1417
R12 VGND.n21 VGND.n20 36.1417
R13 VGND.n22 VGND.n21 36.1417
R14 VGND.n15 VGND.t2 35.0269
R15 VGND.n13 VGND.n12 32.1868
R16 VGND.n14 VGND.t4 31.3528
R17 VGND.n0 VGND.t1 30.0005
R18 VGND.n22 VGND.n1 22.7142
R19 VGND.n20 VGND.n3 18.9495
R20 VGND.n17 VGND.n16 10.2146
R21 VGND.n7 VGND.n6 9.82037
R22 VGND.n24 VGND.n1 9.36437
R23 VGND.n23 VGND.n22 9.3005
R24 VGND.n21 VGND.n2 9.3005
R25 VGND.n20 VGND.n19 9.3005
R26 VGND.n18 VGND.n17 9.3005
R27 VGND.n13 VGND.n4 9.3005
R28 VGND.n12 VGND.n11 9.3005
R29 VGND.n10 VGND.n5 9.3005
R30 VGND.n9 VGND.n8 9.3005
R31 VGND.n8 VGND.n7 8.28285
R32 VGND.n17 VGND.n3 3.10353
R33 VGND.n16 VGND.n13 2.19848
R34 VGND.n9 VGND.n6 0.237019
R35 VGND VGND.n24 0.161675
R36 VGND.n24 VGND.n23 0.146149
R37 VGND.n10 VGND.n9 0.122949
R38 VGND.n11 VGND.n10 0.122949
R39 VGND.n11 VGND.n4 0.122949
R40 VGND.n18 VGND.n4 0.122949
R41 VGND.n19 VGND.n18 0.122949
R42 VGND.n19 VGND.n2 0.122949
R43 VGND.n23 VGND.n2 0.122949
R44 VNB.t7 VNB.t1 3210.5
R45 VNB.t2 VNB.t5 2633.07
R46 VNB.t5 VNB.t3 2552.23
R47 VNB.t4 VNB.t2 1362.73
R48 VNB VNB.t4 1143.31
R49 VNB.t0 VNB.t6 1097.11
R50 VNB.t6 VNB.t7 981.628
R51 VNB.t3 VNB.t0 900.788
R52 a_897_406.n2 a_897_406.t3 482
R53 a_897_406.n1 a_897_406.t2 258.233
R54 a_897_406.n3 a_897_406.n1 211.562
R55 a_897_406.n1 a_897_406.n0 209.764
R56 a_897_406.n4 a_897_406.n3 196.912
R57 a_897_406.n3 a_897_406.n2 185.423
R58 a_897_406.n2 a_897_406.t4 143.798
R59 a_897_406.t0 a_897_406.n4 46.2955
R60 a_897_406.n4 a_897_406.t1 46.2955
R61 VPWR.n20 VPWR.n19 675.105
R62 VPWR.n12 VPWR.n11 585
R63 VPWR.n10 VPWR.n9 585
R64 VPWR.n27 VPWR.n1 323.387
R65 VPWR.n11 VPWR.n10 305.351
R66 VPWR.n8 VPWR.n7 227.428
R67 VPWR.n11 VPWR.t1 74.11
R68 VPWR.n19 VPWR.t7 65.6672
R69 VPWR.n10 VPWR.t3 65.3869
R70 VPWR.n1 VPWR.t4 55.1136
R71 VPWR.n1 VPWR.t6 55.1136
R72 VPWR.n7 VPWR.t2 46.2955
R73 VPWR.n25 VPWR.n2 36.1417
R74 VPWR.n26 VPWR.n25 36.1417
R75 VPWR.n13 VPWR.n4 36.1417
R76 VPWR.n17 VPWR.n4 36.1417
R77 VPWR.n18 VPWR.n17 36.1417
R78 VPWR.n21 VPWR.n18 36.1417
R79 VPWR.n19 VPWR.t5 35.5684
R80 VPWR.n7 VPWR.t0 35.2408
R81 VPWR.n9 VPWR.n8 16.4473
R82 VPWR.n27 VPWR.n26 16.1887
R83 VPWR.n20 VPWR.n2 10.5417
R84 VPWR.n6 VPWR.n5 9.3005
R85 VPWR.n14 VPWR.n13 9.3005
R86 VPWR.n15 VPWR.n4 9.3005
R87 VPWR.n17 VPWR.n16 9.3005
R88 VPWR.n18 VPWR.n3 9.3005
R89 VPWR.n22 VPWR.n21 9.3005
R90 VPWR.n23 VPWR.n2 9.3005
R91 VPWR.n25 VPWR.n24 9.3005
R92 VPWR.n26 VPWR.n0 9.3005
R93 VPWR.n13 VPWR.n12 8.034
R94 VPWR.n28 VPWR.n27 7.54736
R95 VPWR.n12 VPWR.n6 3.47169
R96 VPWR.n9 VPWR.n6 3.25474
R97 VPWR.n21 VPWR.n20 0.753441
R98 VPWR.n8 VPWR.n5 0.491584
R99 VPWR VPWR.n28 0.161584
R100 VPWR.n28 VPWR.n0 0.146238
R101 VPWR.n14 VPWR.n5 0.122949
R102 VPWR.n15 VPWR.n14 0.122949
R103 VPWR.n16 VPWR.n15 0.122949
R104 VPWR.n16 VPWR.n3 0.122949
R105 VPWR.n22 VPWR.n3 0.122949
R106 VPWR.n23 VPWR.n22 0.122949
R107 VPWR.n24 VPWR.n23 0.122949
R108 VPWR.n24 VPWR.n0 0.122949
R109 Q.n1 Q 589.444
R110 Q.n1 Q.n0 585
R111 Q.n2 Q.n1 585
R112 Q.n1 Q.t0 26.3844
R113 Q Q.n2 11.9116
R114 Q Q.n0 10.3116
R115 Q Q.n0 2.84494
R116 Q.n2 Q 1.24494
R117 VPB.t5 VPB.t9 523.521
R118 VPB.t0 VPB.t4 467.339
R119 VPB.t2 VPB.t7 354.974
R120 VPB.t7 VPB.t0 349.866
R121 VPB.t4 VPB.t3 316.668
R122 VPB.t9 VPB.t6 316.668
R123 VPB.t8 VPB.t5 316.668
R124 VPB.t3 VPB.t1 298.791
R125 VPB VPB.t8 260.485
R126 VPB.t6 VPB.t2 214.517
R127 a_27_136.t1 a_27_136.n1 458.661
R128 a_27_136.n1 a_27_136.n0 349.45
R129 a_27_136.n0 a_27_136.t2 332.58
R130 a_27_136.n0 a_27_136.t3 287.861
R131 a_27_136.n1 a_27_136.t0 215.546
R132 a_681_74.t0 a_681_74.t1 45.0005
R133 a_357_392.t1 a_357_392.n1 747.706
R134 a_357_392.n0 a_357_392.t3 411.678
R135 a_357_392.n0 a_357_392.t2 390.322
R136 a_357_392.n1 a_357_392.t0 335.464
R137 a_357_392.n1 a_357_392.n0 76.8461
R138 a_570_392.t0 a_570_392.t1 53.1905
R139 a_654_392.t3 a_654_392.n3 864.467
R140 a_654_392.n3 a_654_392.n0 288.447
R141 a_654_392.n2 a_654_392.n1 277.37
R142 a_654_392.n2 a_654_392.t4 276.322
R143 a_654_392.t3 a_654_392.t1 215.351
R144 a_654_392.n3 a_654_392.n2 152
R145 a_654_392.n0 a_654_392.t0 40.5809
R146 a_654_392.n0 a_654_392.t2 40.0005
R147 a_854_74.t0 a_854_74.t1 78.5719
R148 a_793_508.t0 a_793_508.t1 250.94
R149 a_232_98.t1 a_232_98.n1 770.229
R150 a_232_98.t1 a_232_98.n4 768.644
R151 a_232_98.n0 a_232_98.t5 450.065
R152 a_232_98.n1 a_232_98.n0 336.562
R153 a_232_98.n3 a_232_98.t0 287.55
R154 a_232_98.n2 a_232_98.t3 216.632
R155 a_232_98.n3 a_232_98.n2 212.615
R156 a_232_98.n2 a_232_98.t2 192.102
R157 a_232_98.n0 a_232_98.t4 137.57
R158 a_232_98.n4 a_232_98.n3 30.7175
R159 a_232_98.n4 a_232_98.n1 12.9325
R160 D.n0 D.t1 212.907
R161 D.n0 D.t0 182.113
R162 D D.n0 153.358
R163 GATE_N.n0 GATE_N.t0 213.954
R164 GATE_N.n0 GATE_N.t1 213.688
R165 GATE_N GATE_N.n0 154.133
C0 VPB VGND 0.01559f
C1 GATE_N Q 7.82e-21
C2 RESET_B VGND 0.031218f
C3 VPB Q 0.01375f
C4 RESET_B Q 0.005796f
C5 VGND Q 0.089148f
C6 VPWR D 0.039213f
C7 VPWR GATE_N 0.020271f
C8 VPB VPWR 0.222834f
C9 D GATE_N 0.068911f
C10 VPWR RESET_B 0.017757f
C11 VPB D 0.050977f
C12 VPWR VGND 0.119084f
C13 VPB GATE_N 0.051581f
C14 VPWR Q 0.119302f
C15 D VGND 0.008329f
C16 VPB RESET_B 0.03558f
C17 GATE_N VGND 0.007185f
C18 D Q 1.05e-20
C19 Q VNB 0.114741f
C20 VGND VNB 0.875657f
C21 RESET_B VNB 0.111822f
C22 GATE_N VNB 0.105192f
C23 D VNB 0.131408f
C24 VPWR VNB 0.678966f
C25 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2111o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111o_4 VNB VPB VPWR VGND X D1 C1 B1 A2 A1
X0 VGND.t4 a_137_260.t9 X.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_137_260.t8 B1.t0 VGND.t10 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0928 ps=0.93 w=0.64 l=0.15
X2 VGND.t7 B1.t1 a_137_260.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 VPWR.t3 a_137_260.t10 X.t7 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_549_392.t1 C1.t0 a_814_392.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X5 X.t6 a_137_260.t11 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_814_392.t2 C1.t1 a_549_392.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X7 VPWR.t1 a_137_260.t12 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t4 a_137_260.t13 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X9 a_549_392.t3 D1.t0 a_137_260.t7 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X10 VGND.t5 C1.t2 a_137_260.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.0896 ps=0.92 w=0.64 l=0.15
X11 VGND.t0 A2.t0 a_1210_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X12 VGND.t3 a_137_260.t14 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_1013_392.t4 A2.t1 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X14 VPWR.t6 A2.t2 a_1013_392.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X15 a_1013_392.t5 A1.t0 VPWR.t7 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X16 a_137_260.t0 A1.t1 a_1210_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X17 a_137_260.t6 D1.t1 a_549_392.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X18 VPWR.t4 A1.t2 a_1013_392.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X19 VGND.t9 D1.t2 a_137_260.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.0896 ps=0.92 w=0.64 l=0.15
X20 a_1013_392.t1 B1.t2 a_814_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X21 a_814_392.t0 B1.t3 a_1013_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X22 a_137_260.t2 C1.t3 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0928 ps=0.93 w=0.64 l=0.15
X23 X.t1 a_137_260.t15 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 X.t0 a_137_260.t16 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X25 a_137_260.t4 D1.t3 VGND.t8 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1165 ps=1.065 w=0.64 l=0.15
R0 a_137_260.n1 a_137_260.t0 344.507
R1 a_137_260.n21 a_137_260.n20 339.134
R2 a_137_260.n8 a_137_260.t13 278.173
R3 a_137_260.n16 a_137_260.t10 240.197
R4 a_137_260.n7 a_137_260.t11 240.197
R5 a_137_260.n9 a_137_260.t12 240.197
R6 a_137_260.n18 a_137_260.t14 193.093
R7 a_137_260.n14 a_137_260.t9 179.947
R8 a_137_260.n10 a_137_260.t16 179.947
R9 a_137_260.n17 a_137_260.t15 179.947
R10 a_137_260.n12 a_137_260.n8 165.189
R11 a_137_260.n12 a_137_260.n11 152
R12 a_137_260.n14 a_137_260.n13 152
R13 a_137_260.n15 a_137_260.n6 152
R14 a_137_260.n19 a_137_260.n18 152
R15 a_137_260.n1 a_137_260.n0 117.099
R16 a_137_260.n3 a_137_260.n2 102.793
R17 a_137_260.n5 a_137_260.n4 101.909
R18 a_137_260.n3 a_137_260.n1 67.0123
R19 a_137_260.n5 a_137_260.n3 59.1064
R20 a_137_260.n18 a_137_260.n17 49.6611
R21 a_137_260.n15 a_137_260.n14 49.6611
R22 a_137_260.n11 a_137_260.n7 43.8187
R23 a_137_260.n21 a_137_260.t7 29.5505
R24 a_137_260.t6 a_137_260.n21 29.5505
R25 a_137_260.n9 a_137_260.n8 27.752
R26 a_137_260.n4 a_137_260.t5 26.2505
R27 a_137_260.n4 a_137_260.t4 26.2505
R28 a_137_260.n2 a_137_260.t1 26.2505
R29 a_137_260.n2 a_137_260.t2 26.2505
R30 a_137_260.n0 a_137_260.t3 26.2505
R31 a_137_260.n0 a_137_260.t8 26.2505
R32 a_137_260.n20 a_137_260.n19 25.0187
R33 a_137_260.n20 a_137_260.n5 19.3795
R34 a_137_260.n19 a_137_260.n6 16.6793
R35 a_137_260.n13 a_137_260.n6 13.1884
R36 a_137_260.n13 a_137_260.n12 13.1884
R37 a_137_260.n11 a_137_260.n10 13.146
R38 a_137_260.n16 a_137_260.n15 10.2247
R39 a_137_260.n10 a_137_260.n9 8.76414
R40 a_137_260.n14 a_137_260.n7 5.84292
R41 a_137_260.n17 a_137_260.n16 2.92171
R42 X.n2 X.n0 250.518
R43 X.n2 X.n1 207.6
R44 X.n5 X.n3 141.925
R45 X.n5 X.n4 102.019
R46 X X.n5 61.6234
R47 X.n0 X.t7 26.3844
R48 X.n0 X.t6 26.3844
R49 X.n1 X.t5 26.3844
R50 X.n1 X.t4 26.3844
R51 X.n3 X.t2 22.7032
R52 X.n3 X.t1 22.7032
R53 X.n4 X.t3 22.7032
R54 X.n4 X.t0 22.7032
R55 X X.n2 21.3661
R56 VGND.n7 VGND.t0 240.243
R57 VGND.n23 VGND.t1 231.946
R58 VGND.n21 VGND.n1 225.66
R59 VGND.n15 VGND.n14 205.707
R60 VGND.n8 VGND.t7 154.23
R61 VGND.n3 VGND.n2 123.141
R62 VGND.n6 VGND.n5 114.404
R63 VGND.n20 VGND.n3 35.0123
R64 VGND.n2 VGND.t8 34.688
R65 VGND.n23 VGND.n22 33.5064
R66 VGND.n16 VGND.n15 30.8711
R67 VGND.n5 VGND.t10 27.188
R68 VGND.n5 VGND.t5 27.188
R69 VGND.n14 VGND.t6 27.188
R70 VGND.n14 VGND.t9 27.188
R71 VGND.n13 VGND.n6 24.0946
R72 VGND.n1 VGND.t2 22.7032
R73 VGND.n1 VGND.t4 22.7032
R74 VGND.n2 VGND.t3 22.6611
R75 VGND.n9 VGND.n6 22.5887
R76 VGND.n22 VGND.n21 18.824
R77 VGND.n16 VGND.n3 18.4476
R78 VGND.n9 VGND.n8 17.3181
R79 VGND.n21 VGND.n20 17.3181
R80 VGND.n15 VGND.n13 15.8123
R81 VGND.n22 VGND.n0 9.3005
R82 VGND.n20 VGND.n19 9.3005
R83 VGND.n18 VGND.n3 9.3005
R84 VGND.n10 VGND.n9 9.3005
R85 VGND.n11 VGND.n6 9.3005
R86 VGND.n13 VGND.n12 9.3005
R87 VGND.n15 VGND.n4 9.3005
R88 VGND.n17 VGND.n16 9.3005
R89 VGND.n8 VGND.n7 7.43028
R90 VGND.n24 VGND.n23 6.47485
R91 VGND VGND.n24 0.264179
R92 VGND.n24 VGND.n0 0.166455
R93 VGND.n10 VGND.n7 0.16238
R94 VGND.n11 VGND.n10 0.122949
R95 VGND.n12 VGND.n11 0.122949
R96 VGND.n12 VGND.n4 0.122949
R97 VGND.n17 VGND.n4 0.122949
R98 VGND.n18 VGND.n17 0.122949
R99 VGND.n19 VGND.n18 0.122949
R100 VGND.n19 VGND.n0 0.122949
R101 VNB VNB.t2 2967.98
R102 VNB.t8 VNB.t1 2702.36
R103 VNB.t1 VNB.t0 1986.35
R104 VNB.t4 VNB.t9 1097.11
R105 VNB.t6 VNB.t11 1016.27
R106 VNB.t10 VNB.t7 1016.27
R107 VNB.t11 VNB.t8 993.177
R108 VNB.t7 VNB.t6 993.177
R109 VNB.t9 VNB.t10 993.177
R110 VNB.t3 VNB.t4 993.177
R111 VNB.t5 VNB.t3 993.177
R112 VNB.t2 VNB.t5 993.177
R113 B1.n1 B1.t0 266.707
R114 B1.n0 B1.t2 215.44
R115 B1.n0 B1.t3 212.883
R116 B1.n3 B1.n2 152
R117 B1.n1 B1.t1 128.534
R118 B1.n2 B1.n1 69.8905
R119 B1 B1.n3 13.3823
R120 B1.n2 B1.n0 13.2555
R121 B1.n3 B1 5.23686
R122 A2.n2 A2.t2 268.873
R123 A2.n1 A2.t1 263.762
R124 A2.n1 A2.n0 185.351
R125 A2.n2 A2.t0 183.161
R126 A2.n4 A2.n3 152
R127 A2.n3 A2.n1 37.246
R128 A2.n3 A2.n2 23.3702
R129 A2.n4 A2 10.462
R130 A2 A2.n4 1.35435
R131 a_1210_74.t1 a_1210_74.t0 332.997
R132 VPWR.n31 VPWR.t0 351.637
R133 VPWR.n2 VPWR.n1 334.173
R134 VPWR.n9 VPWR.n8 329.149
R135 VPWR.n11 VPWR.n10 316.447
R136 VPWR.n24 VPWR.t3 259.171
R137 VPWR.n26 VPWR.n25 36.1417
R138 VPWR.n30 VPWR.n29 36.1417
R139 VPWR.n13 VPWR.n12 36.1417
R140 VPWR.n13 VPWR.n6 36.1417
R141 VPWR.n17 VPWR.n6 36.1417
R142 VPWR.n18 VPWR.n17 36.1417
R143 VPWR.n19 VPWR.n18 36.1417
R144 VPWR.n19 VPWR.n4 36.1417
R145 VPWR.n23 VPWR.n4 36.1417
R146 VPWR.n10 VPWR.t7 29.5505
R147 VPWR.n10 VPWR.t4 29.5505
R148 VPWR.n8 VPWR.t5 29.5505
R149 VPWR.n8 VPWR.t6 29.5505
R150 VPWR.n12 VPWR.n11 28.2358
R151 VPWR.n1 VPWR.t2 26.3844
R152 VPWR.n1 VPWR.t1 26.3844
R153 VPWR.n32 VPWR.n31 20.2181
R154 VPWR.n29 VPWR.n2 18.824
R155 VPWR.n26 VPWR.n2 17.3181
R156 VPWR.n24 VPWR.n23 9.41227
R157 VPWR.n12 VPWR.n7 9.3005
R158 VPWR.n14 VPWR.n13 9.3005
R159 VPWR.n15 VPWR.n6 9.3005
R160 VPWR.n17 VPWR.n16 9.3005
R161 VPWR.n18 VPWR.n5 9.3005
R162 VPWR.n20 VPWR.n19 9.3005
R163 VPWR.n21 VPWR.n4 9.3005
R164 VPWR.n23 VPWR.n22 9.3005
R165 VPWR.n25 VPWR.n3 9.3005
R166 VPWR.n27 VPWR.n26 9.3005
R167 VPWR.n29 VPWR.n28 9.3005
R168 VPWR.n30 VPWR.n0 9.3005
R169 VPWR.n25 VPWR.n24 7.90638
R170 VPWR.n31 VPWR.n30 6.4005
R171 VPWR.n11 VPWR.n9 6.39895
R172 VPWR.n9 VPWR.n7 0.609313
R173 VPWR.n14 VPWR.n7 0.122949
R174 VPWR.n15 VPWR.n14 0.122949
R175 VPWR.n16 VPWR.n15 0.122949
R176 VPWR.n16 VPWR.n5 0.122949
R177 VPWR.n20 VPWR.n5 0.122949
R178 VPWR.n21 VPWR.n20 0.122949
R179 VPWR.n22 VPWR.n21 0.122949
R180 VPWR.n22 VPWR.n3 0.122949
R181 VPWR.n27 VPWR.n3 0.122949
R182 VPWR.n28 VPWR.n27 0.122949
R183 VPWR.n28 VPWR.n0 0.122949
R184 VPWR.n32 VPWR.n0 0.122949
R185 VPWR VPWR.n32 0.0617245
R186 VPB.t7 VPB.t0 495.43
R187 VPB.t5 VPB.t8 495.43
R188 VPB VPB.t2 395.834
R189 VPB.t9 VPB.t10 229.839
R190 VPB.t13 VPB.t9 229.839
R191 VPB.t6 VPB.t13 229.839
R192 VPB.t1 VPB.t6 229.839
R193 VPB.t0 VPB.t1 229.839
R194 VPB.t11 VPB.t7 229.839
R195 VPB.t12 VPB.t11 229.839
R196 VPB.t8 VPB.t12 229.839
R197 VPB.t4 VPB.t5 229.839
R198 VPB.t3 VPB.t4 229.839
R199 VPB.t2 VPB.t3 229.839
R200 C1.n1 C1.t3 259.502
R201 C1.n3 C1.t2 238.543
R202 C1.n4 C1.t0 212.883
R203 C1.n1 C1.t1 212.883
R204 C1.n5 C1.n4 154.191
R205 C1.n2 C1.n0 152
R206 C1.n3 C1.n2 36.5157
R207 C1.n2 C1.n1 18.2581
R208 C1.n5 C1.n0 13.1884
R209 C1.n4 C1.n3 10.955
R210 C1.n0 C1 4.84898
R211 C1 C1.n5 0.582318
R212 a_814_392.n1 a_814_392.n0 695.787
R213 a_814_392.n0 a_814_392.t3 29.5505
R214 a_814_392.n0 a_814_392.t2 29.5505
R215 a_814_392.n1 a_814_392.t1 29.5505
R216 a_814_392.t0 a_814_392.n1 29.5505
R217 a_549_392.t1 a_549_392.n1 375.207
R218 a_549_392.n1 a_549_392.t2 375.205
R219 a_549_392.n1 a_549_392.n0 209.173
R220 a_549_392.n0 a_549_392.t0 29.5505
R221 a_549_392.n0 a_549_392.t3 29.5505
R222 D1.n0 D1.t0 273.255
R223 D1.n1 D1.t1 263.762
R224 D1.n1 D1.t3 190.957
R225 D1.n0 D1.t2 183.161
R226 D1 D1.n2 158.012
R227 D1.n2 D1.n1 54.7732
R228 D1.n2 D1.n0 1.46111
R229 a_1013_392.n2 a_1013_392.t0 425.094
R230 a_1013_392.n1 a_1013_392.t4 290.378
R231 a_1013_392.n1 a_1013_392.n0 208.897
R232 a_1013_392.n3 a_1013_392.n2 183.911
R233 a_1013_392.n2 a_1013_392.n1 92.7514
R234 a_1013_392.n0 a_1013_392.t3 29.5505
R235 a_1013_392.n0 a_1013_392.t5 29.5505
R236 a_1013_392.n3 a_1013_392.t2 29.5505
R237 a_1013_392.t1 a_1013_392.n3 29.5505
R238 A1.n1 A1.n0 254.827
R239 A1.n2 A1.t1 244.214
R240 A1.n2 A1.t2 223.839
R241 A1.n1 A1.t0 212.883
R242 A1.n4 A1.n3 152
R243 A1.n3 A1.n1 46.0096
R244 A1.n4 A1 16.4853
R245 A1.n3 A1.n2 8.76414
R246 A1 A1.n4 2.13383
C0 VPB A1 0.074914f
C1 D1 B1 4.65e-19
C2 X VGND 0.32034f
C3 D1 A1 1.05e-19
C4 VPB A2 0.080357f
C5 C1 B1 0.067148f
C6 VPB VPWR 0.228371f
C7 D1 A2 0.00121f
C8 B1 A1 0.082424f
C9 C1 A2 9.18e-20
C10 VPB X 0.02517f
C11 D1 VPWR 0.012748f
C12 C1 VPWR 0.013417f
C13 B1 A2 6.32e-19
C14 VPB VGND 0.01658f
C15 D1 X 0.001825f
C16 A1 A2 0.106035f
C17 B1 VPWR 0.013247f
C18 D1 VGND 0.026702f
C19 C1 VGND 0.037648f
C20 A1 VPWR 0.040862f
C21 B1 VGND 0.043562f
C22 A2 VPWR 0.036154f
C23 VPB D1 0.081848f
C24 A1 VGND 0.013483f
C25 VPB C1 0.091205f
C26 A2 VGND 0.034691f
C27 VPWR X 0.427109f
C28 D1 C1 0.101108f
C29 VPB B1 0.093128f
C30 VPWR VGND 0.129828f
C31 VGND VNB 0.991903f
C32 X VNB 0.093808f
C33 VPWR VNB 0.788037f
C34 A2 VNB 0.265334f
C35 A1 VNB 0.209566f
C36 B1 VNB 0.272832f
C37 C1 VNB 0.225331f
C38 D1 VNB 0.212602f
C39 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2111oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111oi_1 VNB VPB VPWR VGND D1 C1 B1 A2 A1 Y
X0 a_342_368.t1 A2.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.2184 ps=1.51 w=1.12 l=0.15
X1 a_461_74.t1 A1.t0 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VGND.t3 C1.t0 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.185 pd=1.24 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t0 D1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 Y.t2 B1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.185 ps=1.24 w=0.74 l=0.15
X5 VGND.t1 A2.t1 a_461_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X6 a_234_368.t0 C1.t1 a_156_368.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1344 ps=1.36 w=1.12 l=0.15
X7 a_342_368.t0 B1.t1 a_234_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.2184 ps=1.51 w=1.12 l=0.15
X8 a_156_368.t0 D1.t1 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.36 as=0.308 ps=2.79 w=1.12 l=0.15
X9 VPWR.t1 A1.t1 a_342_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.2184 ps=1.51 w=1.12 l=0.15
R0 A2.n0 A2.t0 285.719
R1 A2.n0 A2.t1 178.34
R2 A2 A2.n0 160.476
R3 VPWR VPWR.n0 320.175
R4 VPWR.n0 VPWR.t0 38.6969
R5 VPWR.n0 VPWR.t1 29.9023
R6 a_342_368.n0 a_342_368.t1 485.421
R7 a_342_368.n0 a_342_368.t2 38.6969
R8 a_342_368.t0 a_342_368.n0 29.9023
R9 VPB VPB.t4 360.082
R10 VPB.t3 VPB.t2 275.807
R11 VPB.t1 VPB.t3 275.807
R12 VPB.t0 VPB.t1 275.807
R13 VPB.t4 VPB.t0 199.195
R14 A1.n0 A1.t1 250.909
R15 A1.n0 A1.t0 220.113
R16 A1 A1.n0 157.209
R17 Y.n4 Y.t3 221.385
R18 Y.n2 Y.n0 158.181
R19 Y.n3 Y.n2 106.165
R20 Y.n2 Y.n1 104.579
R21 Y.n0 Y.t4 22.7032
R22 Y.n0 Y.t2 22.7032
R23 Y.n1 Y.t1 22.7032
R24 Y.n1 Y.t0 22.7032
R25 Y.n4 Y.n3 3.35584
R26 Y Y.n4 1.92671
R27 Y.n3 Y 0.683995
R28 a_461_74.t0 a_461_74.t1 51.8924
R29 VNB VNB.t0 1662.99
R30 VNB.t2 VNB.t3 1501.31
R31 VNB.t4 VNB.t1 1085.56
R32 VNB.t3 VNB.t4 993.177
R33 VNB.t0 VNB.t2 993.177
R34 C1.n0 C1.t1 250.909
R35 C1.n0 C1.t0 220.113
R36 C1 C1.n0 154.522
R37 VGND.n7 VGND.t0 233.886
R38 VGND.n2 VGND.n1 206.073
R39 VGND.n3 VGND.t1 163.734
R40 VGND.n1 VGND.t2 40.541
R41 VGND.n1 VGND.t3 40.541
R42 VGND.n6 VGND.n5 36.1417
R43 VGND.n8 VGND.n7 16.8299
R44 VGND.n6 VGND.n0 9.3005
R45 VGND.n5 VGND.n4 9.3005
R46 VGND.n3 VGND.n2 7.52945
R47 VGND.n5 VGND.n2 5.27109
R48 VGND.n7 VGND.n6 3.76521
R49 VGND.n4 VGND.n3 0.269269
R50 VGND.n4 VGND.n0 0.122949
R51 VGND.n8 VGND.n0 0.122949
R52 VGND VGND.n8 0.0617245
R53 D1.n0 D1.t1 250.909
R54 D1.n0 D1.t0 220.113
R55 D1 D1.n0 154.25
R56 B1.n0 B1.t1 250.909
R57 B1.n0 B1.t0 220.113
R58 B1 B1.n0 155.423
R59 a_156_368.t0 a_156_368.t1 42.2148
R60 a_234_368.t0 a_234_368.t1 68.5987
C0 VPB VPWR 0.090017f
C1 C1 A2 1.82e-19
C2 B1 A1 0.094641f
C3 D1 Y 0.133922f
C4 B1 A2 4.66e-19
C5 D1 VPWR 0.003988f
C6 VPB VGND 0.008648f
C7 C1 Y 0.090787f
C8 A1 A2 0.073708f
C9 B1 Y 0.051493f
C10 D1 VGND 0.014698f
C11 C1 VPWR 0.004785f
C12 C1 VGND 0.013036f
C13 A1 Y 0.02161f
C14 B1 VPWR 0.010557f
C15 B1 VGND 0.015663f
C16 A2 Y 0.00532f
C17 A1 VPWR 0.017069f
C18 VPB D1 0.035917f
C19 A2 VPWR 0.017897f
C20 A1 VGND 0.016746f
C21 VPB C1 0.031725f
C22 Y VPWR 0.133272f
C23 A2 VGND 0.054266f
C24 D1 C1 0.10227f
C25 VPB B1 0.034193f
C26 Y VGND 0.311402f
C27 VPB A1 0.035485f
C28 VPWR VGND 0.054652f
C29 VPB A2 0.038364f
C30 C1 B1 0.080858f
C31 VPB Y 0.030098f
C32 D1 A2 1.14e-19
C33 VGND VNB 0.498057f
C34 VPWR VNB 0.351926f
C35 Y VNB 0.117654f
C36 A2 VNB 0.159694f
C37 A1 VNB 0.108544f
C38 B1 VNB 0.103701f
C39 C1 VNB 0.103701f
C40 D1 VNB 0.132239f
C41 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2111oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111oi_2 VNB VPB VPWR VGND D1 B1 Y C1 A2 A1
X0 Y.t1 A1.t0 a_722_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X1 a_69_368.t2 C1.t0 a_334_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VPWR.t1 A2.t0 a_533_368.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t2 B1.t0 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X4 a_533_368.t3 A1.t1 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_533_368.t0 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t2 A1.t2 a_533_368.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_722_74.t0 A2.t2 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1073 ps=1.03 w=0.74 l=0.15
X8 a_334_368.t1 C1.t1 a_69_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_69_368.t0 D1.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_533_368.t5 B1.t1 a_334_368.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_334_368.t0 B1.t2 a_533_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X12 Y.t4 D1.t1 a_69_368.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X13 a_722_74.t1 A1.t3 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VGND.t0 A2.t3 a_722_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VGND.t2 C1.t2 Y.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X16 Y.t5 D1.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.2109 ps=2.05 w=0.74 l=0.15
R0 A1.n1 A1.t2 231.921
R1 A1.n0 A1.t1 226.809
R2 A1.n0 A1.t3 198.204
R3 A1.n1 A1.t0 196.013
R4 A1.n3 A1.n2 152
R5 A1.n2 A1.n0 34.3247
R6 A1.n2 A1.n1 26.2914
R7 A1 A1.n3 10.2703
R8 A1.n3 A1 4.0191
R9 a_722_74.n1 a_722_74.t2 343.711
R10 a_722_74.t0 a_722_74.n1 230.924
R11 a_722_74.n1 a_722_74.n0 86.1054
R12 a_722_74.n0 a_722_74.t3 22.7032
R13 a_722_74.n0 a_722_74.t1 22.7032
R14 Y Y.n0 355.39
R15 Y.n2 Y.n1 286.401
R16 Y.n2 Y.t2 145.892
R17 Y.n4 Y.n3 101.71
R18 Y Y.n4 67.0123
R19 Y.n4 Y.n2 58.0315
R20 Y.n3 Y.t5 34.0546
R21 Y.n3 Y.t6 29.1897
R22 Y.n0 Y.t3 26.3844
R23 Y.n0 Y.t4 26.3844
R24 Y.n1 Y.t0 22.7032
R25 Y.n1 Y.t1 22.7032
R26 VNB.t3 VNB.t2 4226.77
R27 VNB VNB.t4 2402.1
R28 VNB.t6 VNB.t3 1247.24
R29 VNB.t4 VNB.t6 1247.24
R30 VNB.t5 VNB.t0 1016.27
R31 VNB.t1 VNB.t5 993.177
R32 VNB.t2 VNB.t1 993.177
R33 C1.n0 C1.t0 273.401
R34 C1.n0 C1.t1 225.713
R35 C1.n1 C1.t2 220.113
R36 C1.n2 C1.n1 152
R37 C1.n1 C1.n0 19.7187
R38 C1.n2 C1 12.0563
R39 C1 C1.n2 2.23306
R40 a_334_368.n1 a_334_368.n0 681.883
R41 a_334_368.n0 a_334_368.t2 26.3844
R42 a_334_368.n0 a_334_368.t1 26.3844
R43 a_334_368.n1 a_334_368.t3 26.3844
R44 a_334_368.t0 a_334_368.n1 26.3844
R45 a_69_368.t2 a_69_368.n1 393.747
R46 a_69_368.n1 a_69_368.t3 393.745
R47 a_69_368.n1 a_69_368.n0 215.829
R48 a_69_368.n0 a_69_368.t1 26.3844
R49 a_69_368.n0 a_69_368.t0 26.3844
R50 VPB.t6 VPB.t4 495.43
R51 VPB VPB.t8 354.974
R52 VPB.t7 VPB.t0 229.839
R53 VPB.t2 VPB.t7 229.839
R54 VPB.t1 VPB.t2 229.839
R55 VPB.t9 VPB.t1 229.839
R56 VPB.t4 VPB.t9 229.839
R57 VPB.t5 VPB.t6 229.839
R58 VPB.t3 VPB.t5 229.839
R59 VPB.t8 VPB.t3 229.839
R60 A2.n0 A2.t1 228.47
R61 A2.n1 A2.t0 226.809
R62 A2.n1 A2.t3 196.744
R63 A2.n0 A2.t2 196.013
R64 A2 A2.n2 154.522
R65 A2.n2 A2.n0 34.3247
R66 A2.n2 A2.n1 29.2126
R67 a_533_368.n1 a_533_368.t4 398.909
R68 a_533_368.t0 a_533_368.n3 287.007
R69 a_533_368.n3 a_533_368.n2 206.078
R70 a_533_368.n1 a_533_368.n0 188.462
R71 a_533_368.n3 a_533_368.n1 57.9149
R72 a_533_368.n0 a_533_368.t2 26.3844
R73 a_533_368.n0 a_533_368.t5 26.3844
R74 a_533_368.n2 a_533_368.t1 26.3844
R75 a_533_368.n2 a_533_368.t3 26.3844
R76 VPWR.n2 VPWR.n1 340.33
R77 VPWR.n2 VPWR.n0 322.077
R78 VPWR.n1 VPWR.t3 26.3844
R79 VPWR.n1 VPWR.t2 26.3844
R80 VPWR.n0 VPWR.t0 26.3844
R81 VPWR.n0 VPWR.t1 26.3844
R82 VPWR VPWR.n2 1.46047
R83 B1.n0 B1.t0 413.553
R84 B1.n1 B1.t1 271.524
R85 B1.n0 B1.t2 261.62
R86 B1.n2 B1.n1 152
R87 B1.n1 B1.n0 49.521
R88 B1 B1.n2 12.2816
R89 B1.n2 B1 4.32482
R90 VGND.n6 VGND.t3 233.886
R91 VGND.n2 VGND.n1 217.041
R92 VGND.n4 VGND.n3 210.412
R93 VGND.n3 VGND.t4 34.8654
R94 VGND.n5 VGND.n4 34.6358
R95 VGND.n3 VGND.t2 28.3789
R96 VGND.n1 VGND.t1 23.514
R97 VGND.n1 VGND.t0 23.514
R98 VGND.n6 VGND.n5 15.8123
R99 VGND.n5 VGND.n0 9.3005
R100 VGND.n7 VGND.n6 7.56047
R101 VGND.n4 VGND.n2 6.2859
R102 VGND.n2 VGND.n0 0.171074
R103 VGND VGND.n7 0.161757
R104 VGND.n7 VGND.n0 0.146068
R105 D1.n0 D1.t1 277.2
R106 D1.n1 D1.t0 229
R107 D1.n0 D1.t2 196.013
R108 D1 D1.n1 152.447
R109 D1.n1 D1.n0 13.146
C0 C1 VGND 0.02233f
C1 A1 Y 0.043271f
C2 B1 VPWR 0.013215f
C3 B1 VGND 0.021101f
C4 A2 Y 9.53e-21
C5 A1 VPWR 0.031648f
C6 VPB D1 0.068546f
C7 A1 VGND 0.014741f
C8 A2 VPWR 0.041167f
C9 VPB C1 0.06923f
C10 A2 VGND 0.035374f
C11 Y VPWR 0.019059f
C12 VPB B1 0.083446f
C13 D1 C1 0.089907f
C14 Y VGND 0.344107f
C15 VPB A1 0.061602f
C16 D1 B1 1.08e-19
C17 VPWR VGND 0.089263f
C18 VPB A2 0.064123f
C19 C1 B1 0.067756f
C20 C1 A1 0.004699f
C21 VPB Y 0.01668f
C22 VPB VPWR 0.135324f
C23 D1 Y 0.176016f
C24 B1 A1 0.065837f
C25 VPB VGND 0.009942f
C26 D1 VPWR 0.011189f
C27 B1 A2 4.72e-19
C28 C1 Y 0.113433f
C29 B1 Y 0.088542f
C30 A1 A2 0.097245f
C31 C1 VPWR 0.012865f
C32 D1 VGND 0.022012f
C33 VGND VNB 0.735087f
C34 VPWR VNB 0.550971f
C35 Y VNB 0.135372f
C36 A2 VNB 0.232883f
C37 A1 VNB 0.196864f
C38 B1 VNB 0.275418f
C39 C1 VNB 0.162552f
C40 D1 VNB 0.190278f
C41 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2111oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111oi_4 VNB VPB VPWR VGND Y D1 C1 B1 A2 A1
X0 a_29_368.t7 C1.t0 a_474_368.t7 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t8 C1.t1 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 Y.t9 B1.t0 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.4366 ps=1.92 w=0.74 l=0.15
X3 a_474_368.t6 C1.t2 a_29_368.t6 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_474_368.t0 B1.t1 a_853_368.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 a_29_368.t5 C1.t3 a_474_368.t5 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_853_368.t5 B1.t2 a_474_368.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t4 D1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X8 a_474_368.t4 C1.t4 a_29_368.t4 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_29_368.t0 D1.t1 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_1228_74.t3 A2.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 Y.t1 D1.t2 a_29_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_29_368.t2 D1.t3 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_1228_74.t2 A2.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_853_368.t9 A2.t2 VPWR.t7 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_1228_74.t1 A1.t0 Y.t10 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VPWR.t6 A2.t3 a_853_368.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_853_368.t11 A2.t4 VPWR.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_1228_74.t0 A1.t1 Y.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 VPWR.t4 A2.t5 a_853_368.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_853_368.t0 A1.t2 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 VPWR.t3 A1.t3 a_853_368.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_853_368.t1 A1.t4 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 Y.t3 D1.t4 a_29_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X24 VGND.t4 C1.t5 Y.t7 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.4366 pd=1.92 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 VPWR.t2 A1.t5 a_853_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 a_853_368.t4 B1.t3 a_474_368.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 VGND.t2 B1.t4 Y.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 a_474_368.t3 B1.t5 a_853_368.t3 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 VGND.t7 D1.t5 Y.t11 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 C1.n1 C1.t0 246.583
R1 C1.n5 C1.t4 228.877
R2 C1.n4 C1.t3 226.809
R3 C1.n2 C1.t2 218.774
R4 C1.n5 C1.t1 195.495
R5 C1.n7 C1.t5 186.374
R6 C1.n1 C1.n0 162.121
R7 C1.n6 C1 156.614
R8 C1.n3 C1.n0 152
R9 C1.n9 C1.n8 152
R10 C1.n4 C1.n3 44.8533
R11 C1.n7 C1.n6 38.8283
R12 C1.n2 C1.n1 27.8082
R13 C1.n3 C1.n2 14.4708
R14 C1.n6 C1.n5 12.0505
R15 C1 C1.n9 8.7819
R16 C1.n8 C1.n7 6.69494
R17 C1.n9 C1 5.50748
R18 C1 C1.n0 1.34003
R19 C1.n8 C1.n4 0.669944
R20 a_474_368.n2 a_474_368.n0 348.139
R21 a_474_368.n4 a_474_368.n3 345.543
R22 a_474_368.n5 a_474_368.n4 302.625
R23 a_474_368.n2 a_474_368.n1 302.483
R24 a_474_368.n4 a_474_368.n2 83.577
R25 a_474_368.n3 a_474_368.t2 26.3844
R26 a_474_368.n3 a_474_368.t3 26.3844
R27 a_474_368.n0 a_474_368.t5 26.3844
R28 a_474_368.n0 a_474_368.t4 26.3844
R29 a_474_368.n1 a_474_368.t7 26.3844
R30 a_474_368.n1 a_474_368.t6 26.3844
R31 a_474_368.n5 a_474_368.t1 26.3844
R32 a_474_368.t0 a_474_368.n5 26.3844
R33 a_29_368.n2 a_29_368.t3 472.947
R34 a_29_368.n4 a_29_368.t7 442.921
R35 a_29_368.n2 a_29_368.n1 309.978
R36 a_29_368.n5 a_29_368.n4 299.76
R37 a_29_368.n3 a_29_368.n0 188.462
R38 a_29_368.n3 a_29_368.n2 76.3752
R39 a_29_368.n4 a_29_368.n3 61.9285
R40 a_29_368.n0 a_29_368.t4 26.3844
R41 a_29_368.n0 a_29_368.t0 26.3844
R42 a_29_368.n1 a_29_368.t1 26.3844
R43 a_29_368.n1 a_29_368.t2 26.3844
R44 a_29_368.t6 a_29_368.n5 26.3844
R45 a_29_368.n5 a_29_368.t5 26.3844
R46 VPB.t19 VPB.t8 505.646
R47 VPB VPB.t3 252.823
R48 VPB.t14 VPB.t13 229.839
R49 VPB.t15 VPB.t14 229.839
R50 VPB.t7 VPB.t15 229.839
R51 VPB.t4 VPB.t7 229.839
R52 VPB.t12 VPB.t4 229.839
R53 VPB.t5 VPB.t12 229.839
R54 VPB.t6 VPB.t5 229.839
R55 VPB.t10 VPB.t6 229.839
R56 VPB.t11 VPB.t10 229.839
R57 VPB.t9 VPB.t11 229.839
R58 VPB.t8 VPB.t9 229.839
R59 VPB.t18 VPB.t19 229.839
R60 VPB.t17 VPB.t18 229.839
R61 VPB.t16 VPB.t17 229.839
R62 VPB.t0 VPB.t16 229.839
R63 VPB.t1 VPB.t0 229.839
R64 VPB.t2 VPB.t1 229.839
R65 VPB.t3 VPB.t2 229.839
R66 VGND.n37 VGND.t0 292.372
R67 VGND.n10 VGND.t1 239.349
R68 VGND.n9 VGND.t3 233.886
R69 VGND.n5 VGND.t2 232.528
R70 VGND.n35 VGND.n2 206.333
R71 VGND.n30 VGND.n29 185
R72 VGND.n28 VGND.n4 185
R73 VGND.n27 VGND.n26 185
R74 VGND.n28 VGND.n27 72.9735
R75 VGND.n29 VGND.n28 72.9735
R76 VGND.n13 VGND.n12 36.1417
R77 VGND.n14 VGND.n13 36.1417
R78 VGND.n14 VGND.n7 36.1417
R79 VGND.n18 VGND.n7 36.1417
R80 VGND.n19 VGND.n18 36.1417
R81 VGND.n20 VGND.n19 36.1417
R82 VGND.n35 VGND.n1 32.377
R83 VGND.n24 VGND.n5 31.624
R84 VGND.n12 VGND.n9 26.3534
R85 VGND.n37 VGND.n36 24.8476
R86 VGND.n27 VGND.t6 22.7032
R87 VGND.n29 VGND.t4 22.7032
R88 VGND.n2 VGND.t5 22.7032
R89 VGND.n2 VGND.t7 22.7032
R90 VGND.n20 VGND.n5 15.8123
R91 VGND.n36 VGND.n35 15.0593
R92 VGND.n26 VGND.n24 14.868
R93 VGND.n30 VGND.n1 14.1151
R94 VGND.n36 VGND.n0 9.3005
R95 VGND.n35 VGND.n34 9.3005
R96 VGND.n33 VGND.n1 9.3005
R97 VGND.n32 VGND.n31 9.3005
R98 VGND.n25 VGND.n3 9.3005
R99 VGND.n12 VGND.n11 9.3005
R100 VGND.n13 VGND.n8 9.3005
R101 VGND.n15 VGND.n14 9.3005
R102 VGND.n16 VGND.n7 9.3005
R103 VGND.n18 VGND.n17 9.3005
R104 VGND.n19 VGND.n6 9.3005
R105 VGND.n21 VGND.n20 9.3005
R106 VGND.n22 VGND.n5 9.3005
R107 VGND.n24 VGND.n23 9.3005
R108 VGND.n38 VGND.n37 7.09071
R109 VGND.n10 VGND.n9 6.46493
R110 VGND.n25 VGND.n4 3.39077
R111 VGND.n31 VGND.n4 3.25239
R112 VGND.n31 VGND.n30 2.97564
R113 VGND.n26 VGND.n25 2.83726
R114 VGND.n11 VGND.n10 0.645984
R115 VGND VGND.n38 0.273695
R116 VGND.n38 VGND.n0 0.157083
R117 VGND.n11 VGND.n8 0.122949
R118 VGND.n15 VGND.n8 0.122949
R119 VGND.n16 VGND.n15 0.122949
R120 VGND.n17 VGND.n16 0.122949
R121 VGND.n17 VGND.n6 0.122949
R122 VGND.n21 VGND.n6 0.122949
R123 VGND.n22 VGND.n21 0.122949
R124 VGND.n23 VGND.n22 0.122949
R125 VGND.n23 VGND.n3 0.122949
R126 VGND.n32 VGND.n3 0.122949
R127 VGND.n33 VGND.n32 0.122949
R128 VGND.n34 VGND.n33 0.122949
R129 VGND.n34 VGND.n0 0.122949
R130 Y.n2 Y.n0 351.935
R131 Y.n4 Y.t10 317.572
R132 Y.n2 Y.n1 305.048
R133 Y.n4 Y.t5 275
R134 Y.n6 Y.n4 144.391
R135 Y.n8 Y.n6 116.316
R136 Y Y.n9 110.731
R137 Y.n6 Y.n5 103.555
R138 Y.n9 Y.n3 98.5686
R139 Y.n8 Y.n7 96.9594
R140 Y.n9 Y.n8 59.4273
R141 Y Y.n2 27.5811
R142 Y.n0 Y.t0 26.3844
R143 Y.n0 Y.t1 26.3844
R144 Y.n1 Y.t2 26.3844
R145 Y.n1 Y.t3 26.3844
R146 Y.n3 Y.t11 22.7032
R147 Y.n3 Y.t4 22.7032
R148 Y.n7 Y.t7 22.7032
R149 Y.n7 Y.t8 22.7032
R150 Y.n5 Y.t6 22.7032
R151 Y.n5 Y.t9 22.7032
R152 VNB.t3 VNB.t2 5728.08
R153 VNB VNB.t0 3233.6
R154 VNB.t5 VNB.t7 3071.92
R155 VNB.t4 VNB.t1 1986.35
R156 VNB.t8 VNB.t4 1986.35
R157 VNB.t2 VNB.t8 1986.35
R158 VNB.t7 VNB.t3 993.177
R159 VNB.t6 VNB.t5 993.177
R160 VNB.t9 VNB.t6 993.177
R161 VNB.t0 VNB.t9 993.177
R162 B1.n4 B1.t0 267.613
R163 B1.n0 B1.t3 261.921
R164 B1.n1 B1.t5 226.809
R165 B1.n7 B1.t2 226.809
R166 B1.n2 B1.t1 226.809
R167 B1.n3 B1.t4 196.013
R168 B1 B1.n4 153.042
R169 B1.n9 B1.n8 152
R170 B1.n6 B1.n5 152
R171 B1 B1.n0 70.0185
R172 B1.n8 B1.n1 56.2338
R173 B1.n7 B1.n6 44.549
R174 B1.n3 B1.n2 27.0217
R175 B1.n1 B1.n0 22.5061
R176 B1.n6 B1.n2 21.1793
R177 B1.n8 B1.n7 9.49444
R178 B1.n5 B1 9.07957
R179 B1 B1.n9 8.48422
R180 B1.n9 B1 5.80515
R181 B1.n5 B1 5.2098
R182 B1.n4 B1.n3 1.46111
R183 a_853_368.t6 a_853_368.n9 436.579
R184 a_853_368.n9 a_853_368.n8 299.76
R185 a_853_368.n4 a_853_368.t9 280.983
R186 a_853_368.n7 a_853_368.n0 208.065
R187 a_853_368.n6 a_853_368.n1 208.065
R188 a_853_368.n5 a_853_368.n2 208.065
R189 a_853_368.n4 a_853_368.n3 203.27
R190 a_853_368.n6 a_853_368.n5 67.7652
R191 a_853_368.n7 a_853_368.n6 67.7652
R192 a_853_368.n9 a_853_368.n7 59.1064
R193 a_853_368.n5 a_853_368.n4 55.3417
R194 a_853_368.n0 a_853_368.t2 26.3844
R195 a_853_368.n0 a_853_368.t4 26.3844
R196 a_853_368.n1 a_853_368.t8 26.3844
R197 a_853_368.n1 a_853_368.t1 26.3844
R198 a_853_368.n2 a_853_368.t7 26.3844
R199 a_853_368.n2 a_853_368.t0 26.3844
R200 a_853_368.n3 a_853_368.t10 26.3844
R201 a_853_368.n3 a_853_368.t11 26.3844
R202 a_853_368.n8 a_853_368.t3 26.3844
R203 a_853_368.n8 a_853_368.t5 26.3844
R204 D1.n8 D1.t4 294.483
R205 D1.n1 D1.t1 264.183
R206 D1.n5 D1.t2 261.62
R207 D1.n7 D1.t3 261.62
R208 D1 D1.n2 157.017
R209 D1.n4 D1.t0 154.24
R210 D1.n1 D1.t5 154.24
R211 D1.n4 D1.n3 152
R212 D1.n6 D1.n0 152
R213 D1.n9 D1.n8 152
R214 D1.n4 D1.n2 49.6611
R215 D1.n6 D1.n5 48.9308
R216 D1.n8 D1.n7 32.8641
R217 D1.n7 D1.n6 16.7975
R218 D1.n2 D1.n1 13.146
R219 D1.n9 D1.n0 11.7627
R220 D1.n3 D1 9.85996
R221 D1.n3 D1 6.74645
R222 D1 D1.n9 2.94104
R223 D1 D1.n0 1.9032
R224 D1.n5 D1.n4 0.730803
R225 A2.n0 A2.t2 237.762
R226 A2.n3 A2.t3 226.809
R227 A2.n5 A2.t4 226.809
R228 A2.n8 A2.t5 226.809
R229 A2.n8 A2.n7 198.204
R230 A2.n6 A2.t1 196.013
R231 A2.n4 A2.n2 196.013
R232 A2.n0 A2.t0 196.013
R233 A2 A2.n1 155.423
R234 A2.n14 A2.n13 152
R235 A2.n12 A2.n11 152
R236 A2.n10 A2.n9 152
R237 A2.n13 A2.n12 49.6611
R238 A2.n9 A2.n6 40.8975
R239 A2.n3 A2.n1 37.246
R240 A2.n9 A2.n8 19.7187
R241 A2.n1 A2.n0 17.5278
R242 A2.n11 A2.n10 10.1214
R243 A2.n4 A2.n3 8.03383
R244 A2.n14 A2 7.5912
R245 A2 A2.n14 6.69817
R246 A2.n6 A2.n5 5.11262
R247 A2.n13 A2.n4 4.38232
R248 A2.n12 A2.n5 3.65202
R249 A2.n11 A2 2.53073
R250 A2.n10 A2 1.63771
R251 a_1228_74.n0 a_1228_74.t0 338.563
R252 a_1228_74.n1 a_1228_74.t3 210.411
R253 a_1228_74.t2 a_1228_74.n1 152.094
R254 a_1228_74.n0 a_1228_74.t1 134.165
R255 a_1228_74.n1 a_1228_74.n0 81.2437
R256 VPWR.n7 VPWR.n6 329.325
R257 VPWR.n5 VPWR.n4 323.406
R258 VPWR.n10 VPWR.n3 316.683
R259 VPWR.n12 VPWR.n1 316.682
R260 VPWR.n11 VPWR.n10 32.7534
R261 VPWR.n9 VPWR.n5 28.2358
R262 VPWR.n1 VPWR.t1 26.3844
R263 VPWR.n1 VPWR.t2 26.3844
R264 VPWR.n3 VPWR.t0 26.3844
R265 VPWR.n3 VPWR.t3 26.3844
R266 VPWR.n4 VPWR.t5 26.3844
R267 VPWR.n4 VPWR.t4 26.3844
R268 VPWR.n6 VPWR.t7 26.3844
R269 VPWR.n6 VPWR.t6 26.3844
R270 VPWR.n10 VPWR.n9 14.6829
R271 VPWR.n12 VPWR.n11 10.1652
R272 VPWR.n9 VPWR.n8 9.3005
R273 VPWR.n10 VPWR.n2 9.3005
R274 VPWR.n11 VPWR.n0 9.3005
R275 VPWR.n13 VPWR.n12 8.77986
R276 VPWR.n7 VPWR.n5 6.89176
R277 VPWR VPWR.n13 1.6348
R278 VPWR.n8 VPWR.n7 0.477517
R279 VPWR.n13 VPWR.n0 0.149471
R280 VPWR.n8 VPWR.n2 0.122949
R281 VPWR.n2 VPWR.n0 0.122949
R282 A1.n6 A1.t5 236.303
R283 A1.n1 A1.t2 226.809
R284 A1.n10 A1.t3 226.809
R285 A1.n4 A1.t4 226.809
R286 A1.n1 A1.t0 196.744
R287 A1.n6 A1.n5 196.013
R288 A1.n3 A1.t1 196.013
R289 A1.n11 A1.n2 196.013
R290 A1 A1.n7 157.507
R291 A1.n14 A1.n13 152
R292 A1.n12 A1.n0 152
R293 A1.n9 A1.n8 152
R294 A1.n13 A1.n12 49.6611
R295 A1.n10 A1.n9 44.549
R296 A1.n7 A1.n4 28.4823
R297 A1.n7 A1.n6 27.752
R298 A1.n9 A1.n3 14.6066
R299 A1.n13 A1.n1 10.955
R300 A1.n14 A1.n0 10.1214
R301 A1.n8 A1 9.67492
R302 A1.n4 A1.n3 6.57323
R303 A1.n8 A1 4.61445
R304 A1 A1.n14 3.72143
R305 A1.n11 A1.n10 3.65202
R306 A1.n12 A1.n11 1.46111
R307 A1 A1.n0 0.447012
C0 B1 A1 0.061978f
C1 D1 Y 0.353978f
C2 VPB VPWR 0.218939f
C3 VPB VGND 0.01084f
C4 C1 Y 0.150939f
C5 D1 VPWR 0.022826f
C6 B1 Y 0.193066f
C7 D1 VGND 0.040716f
C8 A1 A2 0.09536f
C9 C1 VPWR 0.026803f
C10 A1 Y 0.141012f
C11 C1 VGND 0.041927f
C12 B1 VPWR 0.025656f
C13 B1 VGND 0.042372f
C14 A1 VPWR 0.076774f
C15 A2 Y 8.18e-21
C16 VPB D1 0.126921f
C17 A2 VPWR 0.073871f
C18 A1 VGND 0.027212f
C19 VPB C1 0.138813f
C20 A2 VGND 0.072648f
C21 Y VPWR 0.026137f
C22 VPB B1 0.167401f
C23 D1 C1 0.071476f
C24 Y VGND 0.617667f
C25 VPB A1 0.133327f
C26 D1 B1 1.6e-19
C27 VPWR VGND 0.157514f
C28 C1 B1 0.049553f
C29 VPB A2 0.136946f
C30 D1 A1 6.61e-20
C31 D1 A2 3.72e-20
C32 VPB Y 0.0169f
C33 VGND VNB 1.19877f
C34 VPWR VNB 0.911146f
C35 Y VNB 0.165241f
C36 A2 VNB 0.4349f
C37 A1 VNB 0.40232f
C38 B1 VNB 0.395117f
C39 C1 VNB 0.330976f
C40 D1 VNB 0.376209f
C41 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2_1 VNB VPB VPWR VGND A B X
X0 VGND.t0 B.t0 a_143_136.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X1 X.t0 a_56_136.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X2 VPWR.t0 B.t1 a_56_136.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X3 a_143_136.t1 A.t0 a_56_136.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X4 a_56_136.t1 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X5 X.t1 a_56_136.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
R0 B.n0 B.t1 280.899
R1 B B.n0 163.831
R2 B.n0 B.t0 162.274
R3 a_143_136.n0 a_143_136.t1 58.1616
R4 a_143_136.n0 a_143_136.t0 21.7331
R5 a_143_136.n1 a_143_136.n0 19.2005
R6 VGND VGND.n0 223.911
R7 VGND.n0 VGND.t0 41.2505
R8 VGND.n0 VGND.t1 30.2643
R9 VNB VNB.t2 1478.22
R10 VNB.t0 VNB.t1 1339.63
R11 VNB.t2 VNB.t0 1316.54
R12 a_56_136.n2 a_56_136.n1 310.726
R13 a_56_136.n1 a_56_136.t2 266.307
R14 a_56_136.n0 a_56_136.t4 250.909
R15 a_56_136.n1 a_56_136.n0 206.288
R16 a_56_136.n0 a_56_136.t3 178.34
R17 a_56_136.n2 a_56_136.t1 46.9053
R18 a_56_136.t0 a_56_136.n2 35.1791
R19 X X.n0 589.052
R20 X.n2 X.n0 585
R21 X.n1 X.n0 585
R22 X X.t0 194.166
R23 X.n0 X.t1 26.3844
R24 X X.n1 9.88404
R25 X X.n2 8.91189
R26 X.n2 X 3.07898
R27 X.n1 X 2.10683
R28 VPWR.n1 VPWR.t1 408.699
R29 VPWR.n1 VPWR.n0 322.483
R30 VPWR.n0 VPWR.t0 55.1136
R31 VPWR.n0 VPWR.t2 30.9991
R32 VPWR VPWR.n1 0.41117
R33 VPB VPB.t1 380.512
R34 VPB.t0 VPB.t2 273.253
R35 VPB.t1 VPB.t0 255.376
R36 A.t0 A.t1 446.654
R37 A.n0 A.t0 226.732
R38 A.n0 A 9.35543
R39 A A.n0 5.14939
C0 VPB A 0.060048f
C1 B VPB 0.05551f
C2 VPWR VPB 0.082423f
C3 B A 0.060516f
C4 VPWR A 0.020238f
C5 X VPB 0.019336f
C6 B VPWR 0.016027f
C7 VGND VPB 0.007978f
C8 X A 3.75e-19
C9 B X 0.007749f
C10 VGND A 0.114134f
C11 B VGND 0.025943f
C12 VPWR X 0.108372f
C13 VPWR VGND 0.039835f
C14 X VGND 0.088401f
C15 VGND VNB 0.344552f
C16 X VNB 0.113887f
C17 VPWR VNB 0.294908f
C18 B VNB 0.110132f
C19 A VNB 0.244567f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2_2 VNB VPB VPWR VGND A B X
X0 X.t2 a_31_74.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1332 ps=1.1 w=0.74 l=0.15
X1 a_118_74.t1 A.t0 a_31_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 VPWR.t3 a_31_74.t4 X.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X.t3 a_31_74.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1934 ps=1.475 w=1.12 l=0.15
X4 VGND.t0 B.t0 a_118_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X5 VPWR.t0 B.t1 a_31_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1934 pd=1.475 as=0.15 ps=1.3 w=1 l=0.15
X6 VGND.t1 a_31_74.t6 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 a_31_74.t2 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.29 ps=2.58 w=1 l=0.15
R0 a_31_74.n4 a_31_74.n3 277.866
R1 a_31_74.n0 a_31_74.t4 270.384
R2 a_31_74.n1 a_31_74.t5 261.62
R3 a_31_74.n3 a_31_74.t1 224.952
R4 a_31_74.n1 a_31_74.t3 160.083
R5 a_31_74.n0 a_31_74.t6 154.24
R6 a_31_74.n3 a_31_74.n2 152
R7 a_31_74.n2 a_31_74.n0 49.6611
R8 a_31_74.t0 a_31_74.n4 29.5505
R9 a_31_74.n4 a_31_74.t2 29.5505
R10 a_31_74.n2 a_31_74.n1 7.30353
R11 VGND.n1 VGND.t1 291.466
R12 VGND.n1 VGND.n0 212.487
R13 VGND.n0 VGND.t2 35.6762
R14 VGND.n0 VGND.t0 22.7032
R15 VGND VGND.n1 0.625231
R16 X.n2 X 591.4
R17 X.n2 X.n0 585
R18 X.n3 X.n2 585
R19 X X.n1 285.452
R20 X.n2 X.t0 26.3844
R21 X.n2 X.t3 26.3844
R22 X.n1 X.t1 22.7032
R23 X.n1 X.t2 22.7032
R24 X X.n3 17.1525
R25 X X.n0 14.8485
R26 X X.n0 4.0965
R27 X.n3 X 1.7925
R28 VNB VNB.t3 1189.5
R29 VNB.t0 VNB.t2 1177.95
R30 VNB.t2 VNB.t1 993.177
R31 VNB.t3 VNB.t0 900.788
R32 A.n0 A.t1 269.449
R33 A.n0 A.t0 196.345
R34 A A.n0 155.067
R35 a_118_74.t0 a_118_74.t1 38.9194
R36 VPWR.n1 VPWR.t3 432.55
R37 VPWR.n3 VPWR.n2 315.928
R38 VPWR.n5 VPWR.t1 251.91
R39 VPWR.n2 VPWR.t0 39.4005
R40 VPWR.n2 VPWR.t2 28.5357
R41 VPWR.n4 VPWR.n3 25.6005
R42 VPWR.n5 VPWR.n4 21.0829
R43 VPWR.n4 VPWR.n0 9.3005
R44 VPWR.n6 VPWR.n5 9.3005
R45 VPWR.n3 VPWR.n1 6.57989
R46 VPWR.n1 VPWR.n0 0.608915
R47 VPWR.n6 VPWR.n0 0.122949
R48 VPWR VPWR.n6 0.0617245
R49 VPB.t0 VPB.t2 257.93
R50 VPB VPB.t1 255.376
R51 VPB.t2 VPB.t3 229.839
R52 VPB.t1 VPB.t0 229.839
R53 B.n0 B.t1 277.151
R54 B.n0 B.t0 204.048
R55 B B.n0 160.8
C0 X VGND 0.115705f
C1 VPB A 0.051525f
C2 VPB B 0.0428f
C3 VPB VPWR 0.086824f
C4 A B 0.119367f
C5 A VPWR 0.055467f
C6 VPB X 0.006802f
C7 VPB VGND 0.006415f
C8 A X 2.51e-19
C9 B VPWR 0.019833f
C10 A VGND 0.01424f
C11 B X 0.001552f
C12 VPWR X 0.161582f
C13 B VGND 0.018046f
C14 VPWR VGND 0.048577f
C15 VGND VNB 0.348341f
C16 X VNB 0.056229f
C17 VPWR VNB 0.335572f
C18 B VNB 0.104639f
C19 A VNB 0.16975f
C20 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2_4 VNB VPB VPWR VGND X A B
X0 X.t3 a_83_269.t6 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_83_269.t1 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1365 pd=1.165 as=0.199925 ps=1.505 w=0.84 l=0.15
X2 a_83_269.t5 A.t0 a_504_119.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.0976 ps=0.945 w=0.64 l=0.15
X3 VPWR.t6 a_83_269.t7 X.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.199925 pd=1.505 as=0.1792 ps=1.44 w=1.12 l=0.15
X4 VGND.t5 a_83_269.t8 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.1591 ps=1.17 w=0.74 l=0.15
X5 X.t6 a_83_269.t9 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 X.t1 a_83_269.t10 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VPWR.t4 a_83_269.t11 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t2 B.t1 a_83_269.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
X9 a_83_269.t4 A.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1365 ps=1.165 w=0.84 l=0.15
X10 VGND.t3 a_83_269.t12 X.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t0 A.t2 a_83_269.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1365 pd=1.165 as=0.1365 ps=1.165 w=0.84 l=0.15
X12 VGND.t1 B.t2 a_504_119.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.096 ps=0.94 w=0.64 l=0.15
X13 a_504_119.t0 A.t3 a_83_269.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.096 pd=0.94 as=0.104 ps=0.965 w=0.64 l=0.15
X14 X.t4 a_83_269.t13 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1591 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_504_119.t2 B.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0976 pd=0.945 as=0.12945 ps=1.1 w=0.64 l=0.15
R0 a_83_269.n13 a_83_269.n11 307.771
R1 a_83_269.n15 a_83_269.n14 303.752
R2 a_83_269.n1 a_83_269.t7 228.148
R3 a_83_269.n7 a_83_269.t10 228.148
R4 a_83_269.n4 a_83_269.t11 228.148
R5 a_83_269.n2 a_83_269.t6 228.148
R6 a_83_269.n13 a_83_269.n12 169.456
R7 a_83_269.n5 a_83_269.n0 165.189
R8 a_83_269.n1 a_83_269.t8 163.005
R9 a_83_269.n2 a_83_269.t9 155.702
R10 a_83_269.n3 a_83_269.t12 154.24
R11 a_83_269.n6 a_83_269.t13 154.24
R12 a_83_269.n8 a_83_269.n0 152
R13 a_83_269.n10 a_83_269.n9 152
R14 a_83_269.n14 a_83_269.n10 63.008
R15 a_83_269.n3 a_83_269.n2 61.346
R16 a_83_269.n14 a_83_269.n13 59.1064
R17 a_83_269.n9 a_83_269.n8 49.6611
R18 a_83_269.t0 a_83_269.n15 41.0422
R19 a_83_269.n11 a_83_269.t2 35.1791
R20 a_83_269.n11 a_83_269.t4 35.1791
R21 a_83_269.n15 a_83_269.t1 35.1791
R22 a_83_269.n12 a_83_269.t5 34.688
R23 a_83_269.n5 a_83_269.n4 31.4035
R24 a_83_269.n6 a_83_269.n5 27.0217
R25 a_83_269.n12 a_83_269.t3 26.2505
R26 a_83_269.n8 a_83_269.n7 15.3369
R27 a_83_269.n10 a_83_269.n0 13.1884
R28 a_83_269.n7 a_83_269.n6 7.30353
R29 a_83_269.n4 a_83_269.n3 4.38232
R30 a_83_269.n9 a_83_269.n1 3.65202
R31 VPWR.n5 VPWR.t2 419.036
R32 VPWR.n13 VPWR.n2 324.702
R33 VPWR.n7 VPWR.n6 318.065
R34 VPWR.n4 VPWR.n3 315.928
R35 VPWR.n15 VPWR.t7 259.171
R36 VPWR.n3 VPWR.t1 55.1136
R37 VPWR.n6 VPWR.t0 41.0422
R38 VPWR.n6 VPWR.t3 35.1791
R39 VPWR.n13 VPWR.n12 31.2476
R40 VPWR.n3 VPWR.t6 29.339
R41 VPWR.n8 VPWR.n4 28.2358
R42 VPWR.n15 VPWR.n14 26.7299
R43 VPWR.n2 VPWR.t5 26.3844
R44 VPWR.n2 VPWR.t4 26.3844
R45 VPWR.n8 VPWR.n7 24.8476
R46 VPWR.n14 VPWR.n13 22.2123
R47 VPWR.n12 VPWR.n4 19.2005
R48 VPWR.n9 VPWR.n8 9.3005
R49 VPWR.n10 VPWR.n4 9.3005
R50 VPWR.n12 VPWR.n11 9.3005
R51 VPWR.n13 VPWR.n1 9.3005
R52 VPWR.n14 VPWR.n0 9.3005
R53 VPWR.n16 VPWR.n15 9.3005
R54 VPWR.n7 VPWR.n5 6.5258
R55 VPWR.n9 VPWR.n5 0.686454
R56 VPWR.n10 VPWR.n9 0.122949
R57 VPWR.n11 VPWR.n10 0.122949
R58 VPWR.n11 VPWR.n1 0.122949
R59 VPWR.n1 VPWR.n0 0.122949
R60 VPWR.n16 VPWR.n0 0.122949
R61 VPWR VPWR.n16 0.0617245
R62 X.n2 X.n0 257.577
R63 X.n2 X.n1 208.775
R64 X.n5 X.n3 152.303
R65 X.n5 X.n4 97.9238
R66 X.n3 X.t7 35.6762
R67 X.n3 X.t4 34.0546
R68 X.n0 X.t2 29.9023
R69 X.n0 X.t1 26.3844
R70 X.n1 X.t0 26.3844
R71 X.n1 X.t3 26.3844
R72 X X.n5 24.8766
R73 X.n4 X.t5 22.7032
R74 X.n4 X.t6 22.7032
R75 X X.n2 15.4488
R76 VPB.t6 VPB.t1 273.253
R77 VPB VPB.t7 257.93
R78 VPB.t0 VPB.t3 242.608
R79 VPB.t1 VPB.t0 242.608
R80 VPB.t5 VPB.t6 240.054
R81 VPB.t3 VPB.t2 229.839
R82 VPB.t4 VPB.t5 229.839
R83 VPB.t7 VPB.t4 229.839
R84 B.t3 B.t2 867.601
R85 B.t2 B.t1 462.721
R86 B.n0 B.t0 262.154
R87 B.n0 B.t3 162.274
R88 B B.n0 155.972
R89 A.n1 A.t2 175.344
R90 A.n0 A.t1 173.788
R91 A.n0 A.t3 173.469
R92 A.n1 A.t0 171.913
R93 A A.n2 154.133
R94 A.n2 A.n0 27.9876
R95 A.n2 A.n1 19.6951
R96 a_504_119.n1 a_504_119.n0 377.872
R97 a_504_119.t1 a_504_119.n1 30.938
R98 a_504_119.n0 a_504_119.t3 30.0005
R99 a_504_119.n0 a_504_119.t0 26.2505
R100 a_504_119.n1 a_504_119.t2 26.2505
R101 VNB.t4 VNB.t7 1339.63
R102 VNB.t7 VNB.t2 1177.95
R103 VNB VNB.t6 1143.31
R104 VNB.t1 VNB.t0 1097.11
R105 VNB.t2 VNB.t1 1050.92
R106 VNB.t0 VNB.t3 1039.37
R107 VNB.t5 VNB.t4 993.177
R108 VNB.t6 VNB.t5 993.177
R109 VGND.n8 VGND.n2 210.988
R110 VGND.n10 VGND.t4 178.171
R111 VGND.n5 VGND.t1 168.736
R112 VGND.n4 VGND.n3 123.285
R113 VGND.n3 VGND.t0 41.2505
R114 VGND.n8 VGND.n1 28.2358
R115 VGND.n10 VGND.n9 26.7299
R116 VGND.n4 VGND.n1 22.9652
R117 VGND.n2 VGND.t2 22.7032
R118 VGND.n2 VGND.t3 22.7032
R119 VGND.n3 VGND.t5 21.3263
R120 VGND.n9 VGND.n8 19.2005
R121 VGND.n11 VGND.n10 9.3005
R122 VGND.n6 VGND.n1 9.3005
R123 VGND.n8 VGND.n7 9.3005
R124 VGND.n9 VGND.n0 9.3005
R125 VGND.n5 VGND.n4 7.17186
R126 VGND.n6 VGND.n5 0.171952
R127 VGND.n7 VGND.n6 0.122949
R128 VGND.n7 VGND.n0 0.122949
R129 VGND.n11 VGND.n0 0.122949
R130 VGND VGND.n11 0.0617245
C0 A VGND 0.009894f
C1 VPB VPWR 0.145815f
C2 VPB X 0.010553f
C3 VPWR X 0.370488f
C4 VPB B 0.098707f
C5 VPB A 0.08246f
C6 VPWR B 0.040592f
C7 X B 0.002512f
C8 VPB VGND 0.011479f
C9 VPWR A 0.039125f
C10 VPWR VGND 0.095958f
C11 X A 1.2e-19
C12 B A 0.184741f
C13 X VGND 0.265557f
C14 B VGND 0.097732f
C15 VGND VNB 0.621534f
C16 A VNB 0.158972f
C17 B VNB 0.411672f
C18 X VNB 0.036453f
C19 VPWR VNB 0.500911f
C20 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2b_4 VNB VPB VPWR VGND A_N B X
X0 a_233_74.t2 a_27_392.t2 a_218_424.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.096 pd=0.94 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 a_233_74.t3 B.t0 VGND.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.112 ps=0.99 w=0.64 l=0.15
X2 VGND.t5 a_218_424.t6 X.t7 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1073 ps=1.03 w=0.74 l=0.15
X3 VPWR.t7 a_27_392.t3 a_218_424.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1554 pd=1.21 as=0.126 ps=1.14 w=0.84 l=0.15
X4 a_218_424.t2 a_27_392.t4 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1778 ps=1.37 w=0.84 l=0.15
X5 VGND.t4 a_218_424.t7 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VPWR.t5 a_218_424.t8 X.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X7 X.t2 a_218_424.t9 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t3 a_218_424.t10 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VGND.t0 A_N.t0 a_27_392.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X10 X.t0 a_218_424.t11 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1925 ps=1.49 w=1.12 l=0.15
X11 X.t5 a_218_424.t12 VGND.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1197 ps=1.075 w=0.74 l=0.15
X12 VPWR.t1 B.t1 a_218_424.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1925 pd=1.49 as=0.126 ps=1.14 w=0.84 l=0.15
X13 X.t4 a_218_424.t13 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11655 ps=1.055 w=0.74 l=0.15
X14 a_218_424.t1 B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1554 ps=1.21 w=0.84 l=0.15
X15 VGND.t1 B.t3 a_233_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.075 as=0.096 ps=0.94 w=0.64 l=0.15
X16 VPWR.t8 A_N.t1 a_27_392.t1 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1778 pd=1.37 as=0.285 ps=2.57 w=1 l=0.15
X17 a_218_424.t4 a_27_392.t5 a_233_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
R0 a_27_392.n0 a_27_392.t4 303.661
R1 a_27_392.t1 a_27_392.n3 295.322
R2 a_27_392.n3 a_27_392.n2 231.362
R3 a_27_392.n2 a_27_392.n0 207.261
R4 a_27_392.n1 a_27_392.t2 194.407
R5 a_27_392.n0 a_27_392.t3 159.06
R6 a_27_392.n1 a_27_392.t5 149.129
R7 a_27_392.n3 a_27_392.t0 140.62
R8 a_27_392.n2 a_27_392.n1 13.146
R9 a_218_424.n13 a_218_424.n3 354.461
R10 a_218_424.n5 a_218_424.t8 319.192
R11 a_218_424.n14 a_218_424.n13 306.272
R12 a_218_424.n12 a_218_424.n4 292.671
R13 a_218_424.n7 a_218_424.t9 264.647
R14 a_218_424.n9 a_218_424.t11 237.095
R15 a_218_424.n1 a_218_424.t10 234.841
R16 a_218_424.n9 a_218_424.t12 187.079
R17 a_218_424.n2 a_218_424.t6 186.374
R18 a_218_424.n6 a_218_424.t13 165.588
R19 a_218_424.n8 a_218_424.n0 165.189
R20 a_218_424.n11 a_218_424.n10 152
R21 a_218_424.n2 a_218_424.n0 152
R22 a_218_424.n5 a_218_424.t7 142.994
R23 a_218_424.n6 a_218_424.n5 110.861
R24 a_218_424.n7 a_218_424.n6 68.2656
R25 a_218_424.n13 a_218_424.n12 58.3534
R26 a_218_424.n10 a_218_424.n2 49.6611
R27 a_218_424.n1 a_218_424.n8 46.7399
R28 a_218_424.n3 a_218_424.t3 35.1791
R29 a_218_424.n3 a_218_424.t2 35.1791
R30 a_218_424.t0 a_218_424.n14 35.1791
R31 a_218_424.n14 a_218_424.t1 35.1791
R32 a_218_424.n4 a_218_424.t5 26.2505
R33 a_218_424.n4 a_218_424.t4 26.2505
R34 a_218_424.n11 a_218_424.n0 13.1884
R35 a_218_424.n10 a_218_424.n9 12.4399
R36 a_218_424.n8 a_218_424.n7 8.27067
R37 a_218_424.n12 a_218_424.n11 7.95202
R38 a_218_424.n2 a_218_424.n1 2.92171
R39 a_233_74.n1 a_233_74.n0 418.276
R40 a_233_74.n0 a_233_74.t1 33.7505
R41 a_233_74.n0 a_233_74.t3 31.8755
R42 a_233_74.n1 a_233_74.t0 30.0005
R43 a_233_74.t2 a_233_74.n1 26.2505
R44 VNB VNB.t0 1362.73
R45 VNB.t8 VNB.t6 1154.86
R46 VNB.t0 VNB.t8 1154.86
R47 VNB.t5 VNB.t2 1120.21
R48 VNB.t4 VNB.t1 1074.02
R49 VNB.t7 VNB.t5 1039.37
R50 VNB.t2 VNB.t4 1016.27
R51 VNB.t1 VNB.t3 993.177
R52 VNB.t6 VNB.t7 993.177
R53 B B.t0 455.644
R54 B.n0 B.t2 285.988
R55 B.n1 B.t3 194.407
R56 B.n0 B.t1 176.733
R57 B.n2 B.n1 152
R58 B.n1 B.n0 134.96
R59 B B.n2 4.62272
R60 B.n2 B 4.14865
R61 VGND.n3 VGND.t4 239.328
R62 VGND.n5 VGND.n4 218.024
R63 VGND.n8 VGND.n7 204.394
R64 VGND.n15 VGND.n14 114.885
R65 VGND.n14 VGND.t0 39.3755
R66 VGND.n12 VGND.n1 36.1417
R67 VGND.n13 VGND.n12 36.1417
R68 VGND.n7 VGND.t1 35.6255
R69 VGND.n8 VGND.n1 30.8711
R70 VGND.n4 VGND.t3 28.3789
R71 VGND.n14 VGND.t2 26.2505
R72 VGND.n6 VGND.n5 24.4711
R73 VGND.n7 VGND.t6 23.5986
R74 VGND.n4 VGND.t5 22.7032
R75 VGND.n8 VGND.n6 16.5652
R76 VGND.n15 VGND.n13 12.0476
R77 VGND.n6 VGND.n2 9.3005
R78 VGND.n9 VGND.n8 9.3005
R79 VGND.n10 VGND.n1 9.3005
R80 VGND.n12 VGND.n11 9.3005
R81 VGND.n13 VGND.n0 9.3005
R82 VGND.n16 VGND.n15 7.68156
R83 VGND.n5 VGND.n3 6.90487
R84 VGND.n3 VGND.n2 0.616746
R85 VGND VGND.n16 0.163351
R86 VGND.n16 VGND.n0 0.144494
R87 VGND.n9 VGND.n2 0.122949
R88 VGND.n10 VGND.n9 0.122949
R89 VGND.n11 VGND.n10 0.122949
R90 VGND.n11 VGND.n0 0.122949
R91 X.n2 X.n1 279.149
R92 X.n2 X.n0 211.383
R93 X.n5 X.n3 156.356
R94 X.n5 X.n4 103.043
R95 X X.n2 60.0394
R96 X X.n5 29.5289
R97 X.n1 X.t1 26.3844
R98 X.n1 X.t0 26.3844
R99 X.n0 X.t3 26.3844
R100 X.n0 X.t2 26.3844
R101 X.n3 X.t5 24.3248
R102 X.n3 X.t7 22.7032
R103 X.n4 X.t6 22.7032
R104 X.n4 X.t4 22.7032
R105 VPWR.n14 VPWR.n3 323.281
R106 VPWR.n16 VPWR.n1 317.714
R107 VPWR.n8 VPWR.n7 317.152
R108 VPWR.n5 VPWR.n4 315.832
R109 VPWR.n6 VPWR.t5 256.714
R110 VPWR.n1 VPWR.t6 51.5957
R111 VPWR.n3 VPWR.t0 51.5957
R112 VPWR.n4 VPWR.t1 51.5957
R113 VPWR.n3 VPWR.t7 35.1791
R114 VPWR.n1 VPWR.t8 31.2164
R115 VPWR.n4 VPWR.t2 30.9991
R116 VPWR.n15 VPWR.n14 30.4946
R117 VPWR.n13 VPWR.n5 30.4946
R118 VPWR.n7 VPWR.t4 26.3844
R119 VPWR.n7 VPWR.t3 26.3844
R120 VPWR.n9 VPWR.n8 25.977
R121 VPWR.n16 VPWR.n15 23.7181
R122 VPWR.n14 VPWR.n13 22.9652
R123 VPWR.n9 VPWR.n5 16.9417
R124 VPWR.n10 VPWR.n9 9.3005
R125 VPWR.n11 VPWR.n5 9.3005
R126 VPWR.n13 VPWR.n12 9.3005
R127 VPWR.n14 VPWR.n2 9.3005
R128 VPWR.n15 VPWR.n0 9.3005
R129 VPWR.n17 VPWR.n16 7.23624
R130 VPWR.n8 VPWR.n6 6.46335
R131 VPWR.n10 VPWR.n6 0.686829
R132 VPWR VPWR.n17 0.157488
R133 VPWR.n17 VPWR.n0 0.150282
R134 VPWR.n11 VPWR.n10 0.122949
R135 VPWR.n12 VPWR.n11 0.122949
R136 VPWR.n12 VPWR.n2 0.122949
R137 VPWR.n2 VPWR.n0 0.122949
R138 VPB.t1 VPB.t2 265.591
R139 VPB.t7 VPB.t0 265.591
R140 VPB.t8 VPB.t6 265.591
R141 VPB VPB.t8 252.823
R142 VPB.t4 VPB.t5 229.839
R143 VPB.t3 VPB.t4 229.839
R144 VPB.t2 VPB.t3 229.839
R145 VPB.t0 VPB.t1 229.839
R146 VPB.t6 VPB.t7 229.839
R147 A_N.n0 A_N.t0 267.604
R148 A_N.n0 A_N.t1 236.275
R149 A_N A_N.n0 154.133
C0 VPB B 0.118332f
C1 VPB VPWR 0.140781f
C2 A_N B 0.071552f
C3 A_N VPWR 0.040758f
C4 VPB X 0.011177f
C5 VPB VGND 0.008056f
C6 B VPWR 0.040395f
C7 B X 0.003355f
C8 A_N VGND 0.015647f
C9 B VGND 0.034044f
C10 VPWR X 0.387746f
C11 VPWR VGND 0.080539f
C12 X VGND 0.25939f
C13 VPB A_N 0.0507f
C14 VGND VNB 0.608242f
C15 X VNB 0.070166f
C16 VPWR VNB 0.499432f
C17 B VNB 0.255529f
C18 A_N VNB 0.146471f
C19 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3b_1 VNB VPB VPWR VGND X A_N C B
X0 X.t1 a_266_94.t4 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.19855 ps=1.305 w=0.74 l=0.15
X1 a_431_94.t0 B.t0 a_353_94.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
X2 VPWR.t3 a_114_74.t2 a_266_94.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1659 pd=1.235 as=0.2478 ps=2.27 w=0.84 l=0.15
X3 X.t0 a_266_94.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.231 ps=1.555 w=1.12 l=0.15
X4 a_114_74.t0 A_N.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.19525 pd=1.81 as=0.15675 ps=1.67 w=0.55 l=0.15
X5 a_266_94.t0 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1281 pd=1.145 as=0.1659 ps=1.235 w=0.84 l=0.15
X6 VGND.t2 C.t0 a_431_94.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.19855 pd=1.305 as=0.1248 ps=1.03 w=0.64 l=0.15
X7 VPWR.t1 C.t1 a_266_94.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.1281 ps=1.145 w=0.84 l=0.15
X8 a_353_94.t0 a_114_74.t3 a_266_94.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X9 a_114_74.t1 A_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2856 pd=2.36 as=0.252 ps=2.28 w=0.84 l=0.15
R0 a_266_94.n2 a_266_94.t1 388.627
R1 a_266_94.n3 a_266_94.n2 351.048
R2 a_266_94.n1 a_266_94.n0 275.921
R3 a_266_94.n0 a_266_94.t5 264.298
R4 a_266_94.n0 a_266_94.t4 204.048
R5 a_266_94.n1 a_266_94.t2 139.244
R6 a_266_94.t0 a_266_94.n3 36.3517
R7 a_266_94.n3 a_266_94.t3 35.1791
R8 a_266_94.n2 a_266_94.n1 33.9271
R9 VGND.n1 VGND.t0 247.54
R10 VGND.n1 VGND.n0 98.2965
R11 VGND.n0 VGND.t2 49.1757
R12 VGND.n0 VGND.t1 41.4991
R13 VGND VGND.n1 0.099922
R14 X.n1 X 588.903
R15 X.n1 X.n0 585
R16 X.n2 X.n1 585
R17 X X.t1 205.376
R18 X.n1 X.t0 26.3844
R19 X X.n2 10.459
R20 X X.n0 9.05416
R21 X X.n0 2.49806
R22 X.n2 X 1.09318
R23 VNB.t0 VNB.t2 2760.1
R24 VNB.t4 VNB.t3 1651.44
R25 VNB.t1 VNB.t4 1247.24
R26 VNB VNB.t0 1143.31
R27 VNB.t2 VNB.t1 900.788
R28 B.n0 B.t1 205.922
R29 B.n0 B.t0 204.048
R30 B B.n0 155.119
R31 a_353_94.t0 a_353_94.t1 45.0005
R32 a_431_94.t0 a_431_94.t1 73.1255
R33 a_114_74.t1 a_114_74.n1 426
R34 a_114_74.n0 a_114_74.t2 297.527
R35 a_114_74.n1 a_114_74.t0 260.091
R36 a_114_74.n1 a_114_74.n0 235.916
R37 a_114_74.n0 a_114_74.t3 150.25
R38 VPWR.n4 VPWR.n3 618.939
R39 VPWR.n10 VPWR.t0 408.029
R40 VPWR.n5 VPWR.n2 332.841
R41 VPWR.n2 VPWR.t1 55.1136
R42 VPWR.n3 VPWR.t3 46.9053
R43 VPWR.n3 VPWR.t2 45.7326
R44 VPWR.n2 VPWR.t4 38.522
R45 VPWR.n8 VPWR.n1 36.1417
R46 VPWR.n9 VPWR.n8 36.1417
R47 VPWR.n10 VPWR.n9 20.7064
R48 VPWR.n4 VPWR.n1 9.78874
R49 VPWR.n6 VPWR.n1 9.3005
R50 VPWR.n8 VPWR.n7 9.3005
R51 VPWR.n9 VPWR.n0 9.3005
R52 VPWR.n11 VPWR.n10 9.3005
R53 VPWR.n5 VPWR.n4 8.73405
R54 VPWR.n6 VPWR.n5 0.539371
R55 VPWR.n7 VPWR.n6 0.122949
R56 VPWR.n7 VPWR.n0 0.122949
R57 VPWR.n11 VPWR.n0 0.122949
R58 VPWR VPWR.n11 0.0617245
R59 VPB.t0 VPB.t3 607.797
R60 VPB.t1 VPB.t4 298.791
R61 VPB.t3 VPB.t2 278.361
R62 VPB VPB.t0 260.485
R63 VPB.t2 VPB.t1 232.393
R64 A_N.n0 A_N.t1 265.247
R65 A_N.n1 A_N.t0 173.52
R66 A_N A_N.n0 153.007
R67 A_N.n2 A_N.n1 152
R68 A_N.n1 A_N.n0 49.6611
R69 A_N A_N.n2 8.77353
R70 A_N.n2 A_N 1.87016
R71 C.n0 C.t1 205.922
R72 C.n0 C.t0 204.048
R73 C C.n0 157.088
C0 VPWR B 0.013278f
C1 VPB X 0.017871f
C2 VPWR C 0.022148f
C3 VPB VGND 0.012223f
C4 A_N X 1.45e-19
C5 A_N VGND 0.05189f
C6 B C 0.086536f
C7 VPWR X 0.133261f
C8 B X 5.06e-19
C9 VPWR VGND 0.065276f
C10 C X 0.006442f
C11 B VGND 0.009914f
C12 C VGND 0.015655f
C13 X VGND 0.087896f
C14 VPB A_N 0.073781f
C15 VPB VPWR 0.147981f
C16 A_N VPWR 0.045207f
C17 VPB B 0.034166f
C18 VPB C 0.038707f
C19 VGND VNB 0.53103f
C20 X VNB 0.112796f
C21 C VNB 0.109088f
C22 B VNB 0.099723f
C23 VPWR VNB 0.425258f
C24 A_N VNB 0.201149f
C25 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3_4 VNB VPB VPWR VGND X A B C
X0 VPWR.t7 C.t0 a_83_260.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.273 pd=1.49 as=0.126 ps=1.14 w=0.84 l=0.15
X1 X.t7 a_83_260.t8 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t2 a_83_260.t9 X.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_83_260.t3 C.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.2051 ps=1.52 w=0.84 l=0.15
X4 X.t5 a_83_260.t10 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X5 X.t3 a_83_260.t11 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 a_686_74.t1 A.t0 a_83_260.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2144 pd=1.95 as=0.1184 ps=1.01 w=0.64 l=0.15
X7 a_489_74.t1 C.t2 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1245 ps=1.09 w=0.64 l=0.15
X8 X.t2 a_83_260.t12 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 a_83_260.t2 B.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.18 as=0.273 ps=1.49 w=0.84 l=0.15
X10 VGND.t1 a_83_260.t13 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1245 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_489_74.t3 B.t1 a_686_74.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1824 ps=1.85 w=0.64 l=0.15
X12 VPWR.t0 a_83_260.t14 X.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t0 a_83_260.t15 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_83_260.t0 A.t1 a_686_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.01 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 VPWR.t4 B.t2 a_83_260.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.2 as=0.1428 ps=1.18 w=0.84 l=0.15
X16 a_83_260.t7 A.t2 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1512 ps=1.2 w=0.84 l=0.15
X17 VPWR.t8 A.t3 a_83_260.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2898 pd=2.37 as=0.126 ps=1.14 w=0.84 l=0.15
X18 VGND.t4 C.t3 a_489_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X19 a_686_74.t2 B.t3 a_489_74.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1024 ps=0.96 w=0.64 l=0.15
R0 C.n1 C.t2 274.442
R1 C.n3 C.t3 244.214
R2 C.n4 C.t0 230.022
R3 C.n1 C.t1 230.022
R4 C.n5 C.n4 162.956
R5 C.n2 C.n0 152
R6 C.n2 C.n1 27.0217
R7 C.n4 C.n3 22.6399
R8 C.n3 C.n2 16.0672
R9 C.n5 C.n0 13.1884
R10 C.n0 C 5.23686
R11 C C.n5 0.194439
R12 a_83_260.n14 a_83_260.n12 312.18
R13 a_83_260.n11 a_83_260.n10 306.661
R14 a_83_260.n14 a_83_260.n13 306.659
R15 a_83_260.n16 a_83_260.n15 306.659
R16 a_83_260.n0 a_83_260.t9 251.151
R17 a_83_260.n2 a_83_260.t8 240.928
R18 a_83_260.n7 a_83_260.t10 240.197
R19 a_83_260.n4 a_83_260.t14 240.197
R20 a_83_260.n2 a_83_260.t11 179.947
R21 a_83_260.n3 a_83_260.t15 179.947
R22 a_83_260.n6 a_83_260.t12 179.947
R23 a_83_260.n0 a_83_260.t13 179.947
R24 a_83_260.n5 a_83_260.n1 165.189
R25 a_83_260.n8 a_83_260.n1 152
R26 a_83_260.n9 a_83_260.n0 152
R27 a_83_260.n15 a_83_260.n11 69.2711
R28 a_83_260.n11 a_83_260.n9 65.8144
R29 a_83_260.n3 a_83_260.n2 62.8066
R30 a_83_260.n15 a_83_260.n14 50.4476
R31 a_83_260.n0 a_83_260.n8 49.6611
R32 a_83_260.t1 a_83_260.n16 44.56
R33 a_83_260.n12 a_83_260.t0 39.3755
R34 a_83_260.n5 a_83_260.n4 35.7853
R35 a_83_260.n13 a_83_260.t6 35.1791
R36 a_83_260.n13 a_83_260.t7 35.1791
R37 a_83_260.n10 a_83_260.t4 35.1791
R38 a_83_260.n10 a_83_260.t3 35.1791
R39 a_83_260.n16 a_83_260.t2 35.1791
R40 a_83_260.n6 a_83_260.n5 35.055
R41 a_83_260.n12 a_83_260.t5 30.0005
R42 a_83_260.n9 a_83_260.n1 13.1884
R43 a_83_260.n7 a_83_260.n6 9.49444
R44 a_83_260.n8 a_83_260.n7 5.11262
R45 a_83_260.n4 a_83_260.n3 2.19141
R46 VPWR.n9 VPWR.t8 369.536
R47 VPWR.n18 VPWR.n2 317.341
R48 VPWR.n4 VPWR.n3 315.928
R49 VPWR.n8 VPWR.n7 315.928
R50 VPWR.n20 VPWR.t3 259.171
R51 VPWR.n12 VPWR.n6 142.032
R52 VPWR.n6 VPWR.t7 71.4398
R53 VPWR.n6 VPWR.t5 71.4395
R54 VPWR.n3 VPWR.t6 46.9053
R55 VPWR.n7 VPWR.t9 46.9053
R56 VPWR.n3 VPWR.t2 43.0102
R57 VPWR.n7 VPWR.t4 37.5243
R58 VPWR.n2 VPWR.t1 35.1791
R59 VPWR.n2 VPWR.t0 35.1791
R60 VPWR.n12 VPWR.n11 32.7534
R61 VPWR.n13 VPWR.n12 32.0005
R62 VPWR.n17 VPWR.n4 28.9887
R63 VPWR.n20 VPWR.n19 26.7299
R64 VPWR.n19 VPWR.n18 25.977
R65 VPWR.n18 VPWR.n17 21.4593
R66 VPWR.n13 VPWR.n4 18.4476
R67 VPWR.n11 VPWR.n8 17.6946
R68 VPWR.n11 VPWR.n10 9.3005
R69 VPWR.n14 VPWR.n13 9.3005
R70 VPWR.n15 VPWR.n4 9.3005
R71 VPWR.n17 VPWR.n16 9.3005
R72 VPWR.n18 VPWR.n1 9.3005
R73 VPWR.n19 VPWR.n0 9.3005
R74 VPWR.n21 VPWR.n20 9.3005
R75 VPWR.n9 VPWR.n8 6.96039
R76 VPWR.n12 VPWR.n5 4.62059
R77 VPWR.n10 VPWR.n9 0.594857
R78 VPWR.n10 VPWR.n5 0.184273
R79 VPWR.n14 VPWR.n5 0.184273
R80 VPWR.n15 VPWR.n14 0.122949
R81 VPWR.n16 VPWR.n15 0.122949
R82 VPWR.n16 VPWR.n1 0.122949
R83 VPWR.n1 VPWR.n0 0.122949
R84 VPWR.n21 VPWR.n0 0.122949
R85 VPWR VPWR.n21 0.0617245
R86 VPB.t7 VPB.t5 408.603
R87 VPB.t2 VPB.t6 280.914
R88 VPB.t0 VPB.t1 280.914
R89 VPB.t4 VPB.t9 260.485
R90 VPB VPB.t3 257.93
R91 VPB.t5 VPB.t4 250.269
R92 VPB.t9 VPB.t8 229.839
R93 VPB.t6 VPB.t7 229.839
R94 VPB.t1 VPB.t2 229.839
R95 VPB.t3 VPB.t0 229.839
R96 X.n3 X 589.777
R97 X.n3 X.n2 585
R98 X.n4 X.n3 585
R99 X.n5 X.n1 258.046
R100 X.n8 X.n7 185
R101 X.n9 X.n8 185
R102 X.n6 X.n0 147.196
R103 X.n3 X.t4 26.3844
R104 X.n3 X.t7 26.3844
R105 X.n1 X.t6 26.3844
R106 X.n1 X.t5 26.3844
R107 X.n8 X.t0 22.7032
R108 X.n8 X.t3 22.7032
R109 X.n0 X.t1 22.7032
R110 X.n0 X.t2 22.7032
R111 X X.n5 13.4883
R112 X.n4 X 12.8005
R113 X.n9 X 12.6066
R114 X.n2 X 11.0811
R115 X.n6 X 7.02111
R116 X.n7 X 4.84898
R117 X.n7 X.n6 3.10353
R118 X.n2 X 3.05722
R119 X.n5 X 2.48408
R120 X X.n9 1.74595
R121 X X.n4 1.33781
R122 VGND.n5 VGND.t4 241.863
R123 VGND.n8 VGND.n2 217
R124 VGND.n10 VGND.t3 171.77
R125 VGND.n4 VGND.n3 115.751
R126 VGND.n3 VGND.t5 39.3755
R127 VGND.n2 VGND.t2 34.0546
R128 VGND.n8 VGND.n1 27.1064
R129 VGND.n9 VGND.n8 26.3534
R130 VGND.n10 VGND.n9 25.6005
R131 VGND.n2 VGND.t0 22.7032
R132 VGND.n3 VGND.t1 22.6611
R133 VGND.n4 VGND.n1 18.0711
R134 VGND.n11 VGND.n10 9.3005
R135 VGND.n6 VGND.n1 9.3005
R136 VGND.n8 VGND.n7 9.3005
R137 VGND.n9 VGND.n0 9.3005
R138 VGND.n5 VGND.n4 6.92854
R139 VGND.n6 VGND.n5 0.592857
R140 VGND.n7 VGND.n6 0.122949
R141 VGND.n7 VGND.n0 0.122949
R142 VGND.n11 VGND.n0 0.122949
R143 VGND VGND.n11 0.0617245
R144 VNB.t5 VNB.t9 2286.61
R145 VNB.t4 VNB.t7 1201.05
R146 VNB VNB.t3 1177.95
R147 VNB.t1 VNB.t6 1154.86
R148 VNB.t0 VNB.t2 1154.86
R149 VNB.t9 VNB.t8 1085.56
R150 VNB.t8 VNB.t4 993.177
R151 VNB.t6 VNB.t5 993.177
R152 VNB.t2 VNB.t1 993.177
R153 VNB.t3 VNB.t0 993.177
R154 A.n2 A.t1 257.36
R155 A.n0 A.t0 257.36
R156 A.n1 A.t3 200.894
R157 A.n1 A.t2 199.076
R158 A A.n2 158.788
R159 A A.n0 158.4
R160 A.n2 A.n1 28.4823
R161 A.n1 A.n0 21.1793
R162 a_686_74.n1 a_686_74.t3 266.192
R163 a_686_74.t1 a_686_74.n1 188.543
R164 a_686_74.n1 a_686_74.n0 102.562
R165 a_686_74.n0 a_686_74.t0 26.2505
R166 a_686_74.n0 a_686_74.t2 26.2505
R167 a_489_74.n1 a_489_74.n0 405.964
R168 a_489_74.n0 a_489_74.t2 33.7505
R169 a_489_74.n0 a_489_74.t3 26.2505
R170 a_489_74.n1 a_489_74.t0 26.2505
R171 a_489_74.t1 a_489_74.n1 26.2505
R172 B.n2 B.t0 268.606
R173 B.n0 B.t2 263.493
R174 B.n0 B.t3 206.238
R175 B.n2 B.t1 204.048
R176 B B.n1 156.923
R177 B.n4 B.n3 152
R178 B.n3 B.n1 49.6611
R179 B.n1 B.n0 10.955
R180 B.n4 B 8.86204
R181 B.n3 B.n2 5.84292
R182 B B.n4 4.64226
C0 C VPWR 0.039232f
C1 VPB X 0.01234f
C2 B A 0.094545f
C3 C X 0.003669f
C4 B VPWR 0.038986f
C5 VPB VGND 0.010675f
C6 A VPWR 0.037385f
C7 C VGND 0.037728f
C8 B X 7.41e-20
C9 B VGND 0.013635f
C10 A X 2.79e-20
C11 VPWR X 0.409606f
C12 A VGND 0.012406f
C13 VPWR VGND 0.106737f
C14 X VGND 0.29919f
C15 VPB C 0.121851f
C16 VPB B 0.107163f
C17 VPB A 0.099409f
C18 C B 0.057723f
C19 VPB VPWR 0.169045f
C20 VGND VNB 0.721217f
C21 X VNB 0.039185f
C22 VPWR VNB 0.605124f
C23 A VNB 0.250205f
C24 B VNB 0.223975f
C25 C VNB 0.242613f
C26 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3_2 VNB VPB VPWR VGND C X A B
X0 a_247_136.t1 B.t0 a_133_136.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1344 ps=1.06 w=0.64 l=0.15
X1 VGND.t2 a_41_384.t4 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.3552 pd=2.44 as=0.1184 ps=1.06 w=0.74 l=0.15
X2 VPWR.t0 A.t0 a_41_384.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.26 as=0.2478 ps=2.27 w=0.84 l=0.15
X3 VPWR.t4 C.t0 a_41_384.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2845 pd=1.69 as=0.126 ps=1.14 w=0.84 l=0.15
X4 a_41_384.t1 B.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1764 ps=1.26 w=0.84 l=0.15
X5 VGND.t0 C.t1 a_247_136.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.170225 pd=1.34 as=0.0768 ps=0.88 w=0.64 l=0.15
X6 VPWR.t2 a_41_384.t5 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.4088 pd=2.97 as=0.168 ps=1.42 w=1.12 l=0.15
X7 X.t0 a_41_384.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2845 ps=1.69 w=1.12 l=0.15
X8 a_133_136.t1 A.t1 a_41_384.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.1824 ps=1.85 w=0.64 l=0.15
X9 X.t2 a_41_384.t7 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.170225 ps=1.34 w=0.74 l=0.15
R0 B.n0 B.t1 205.922
R1 B.n0 B.t0 162.274
R2 B B.n0 152.469
R3 a_133_136.t0 a_133_136.t1 78.7505
R4 a_247_136.t0 a_247_136.t1 45.0005
R5 VNB VNB.t4 1362.73
R6 VNB.t0 VNB.t2 1339.63
R7 VNB.t4 VNB.t3 1316.54
R8 VNB.t2 VNB.t1 1085.56
R9 VNB.t3 VNB.t0 900.788
R10 a_41_384.t0 a_41_384.n5 390.748
R11 a_41_384.n4 a_41_384.n3 300.373
R12 a_41_384.n0 a_41_384.t5 253.587
R13 a_41_384.n5 a_41_384.t2 247.905
R14 a_41_384.n1 a_41_384.t6 229.487
R15 a_41_384.n4 a_41_384.n2 223.165
R16 a_41_384.n2 a_41_384.t7 193.093
R17 a_41_384.n0 a_41_384.t4 179.947
R18 a_41_384.n5 a_41_384.n4 51.9534
R19 a_41_384.n1 a_41_384.n0 41.6278
R20 a_41_384.n3 a_41_384.t3 35.1791
R21 a_41_384.n3 a_41_384.t1 35.1791
R22 a_41_384.n2 a_41_384.n1 13.8763
R23 X.n2 X.n0 264.964
R24 X.n2 X.n1 94.1587
R25 X.n1 X.t3 29.1897
R26 X.n0 X.t1 26.3844
R27 X.n0 X.t0 26.3844
R28 X.n1 X.t2 22.7032
R29 X X.n2 1.87043
R30 VGND.n1 VGND.t2 162.044
R31 VGND.n1 VGND.n0 125.224
R32 VGND.n0 VGND.t0 50.1733
R33 VGND.n0 VGND.t1 32.9025
R34 VGND VGND.n1 0.665547
R35 A.t1 A.t0 406.488
R36 A.n0 A.t1 223.054
R37 A.n0 A 9.80404
R38 A A.n0 4.70078
R39 VPWR.n8 VPWR.n1 618.939
R40 VPWR.n3 VPWR.n2 322.298
R41 VPWR.n4 VPWR.t2 269.017
R42 VPWR.n2 VPWR.t4 89.6504
R43 VPWR.n1 VPWR.t3 51.5957
R44 VPWR.n1 VPWR.t0 46.9053
R45 VPWR.n7 VPWR.n6 36.1417
R46 VPWR.n2 VPWR.t1 35.3598
R47 VPWR.n6 VPWR.n3 14.6829
R48 VPWR.n8 VPWR.n7 13.9299
R49 VPWR.n6 VPWR.n5 9.3005
R50 VPWR.n7 VPWR.n0 9.3005
R51 VPWR.n9 VPWR.n8 7.6232
R52 VPWR.n4 VPWR.n3 7.08285
R53 VPWR.n5 VPWR.n4 0.583515
R54 VPWR VPWR.n9 0.162583
R55 VPWR.n9 VPWR.n0 0.145253
R56 VPWR.n5 VPWR.n0 0.122949
R57 VPB.t4 VPB.t1 367.743
R58 VPB VPB.t0 293.683
R59 VPB.t0 VPB.t3 291.13
R60 VPB.t1 VPB.t2 229.839
R61 VPB.t3 VPB.t4 229.839
R62 C.n0 C.t0 205.213
R63 C.n0 C.t1 161.565
R64 C C.n0 154.012
C0 A X 1.53e-19
C1 VPWR VGND 0.071407f
C2 B C 0.085872f
C3 A VGND 0.171937f
C4 B X 0.002968f
C5 B VGND 0.009103f
C6 C X 0.001873f
C7 C VGND 0.029116f
C8 X VGND 0.176522f
C9 VPB VPWR 0.12489f
C10 VPB A 0.041045f
C11 VPB B 0.039891f
C12 VPWR A 0.015096f
C13 VPWR B 0.013594f
C14 VPB C 0.04553f
C15 A B 0.07209f
C16 VPB X 0.006168f
C17 VPWR C 0.012269f
C18 VPB VGND 0.011495f
C19 A C 0.001187f
C20 VPWR X 0.197401f
C21 VGND VNB 0.480628f
C22 X VNB 0.029878f
C23 C VNB 0.095896f
C24 B VNB 0.092096f
C25 A VNB 0.241796f
C26 VPWR VNB 0.394908f
C27 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3_1 VNB VPB VPWR VGND A B C X
X0 VPWR.t0 A.t0 a_27_398.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 VPWR.t3 C.t0 a_27_398.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.363225 pd=1.84 as=0.126 ps=1.14 w=0.84 l=0.15
X2 a_27_398.t2 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X3 VGND.t0 C.t1 a_233_136.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.111 ps=1.045 w=0.64 l=0.15
X4 a_233_136.t1 B.t1 a_121_136.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.045 as=0.1312 ps=1.05 w=0.64 l=0.15
X5 X.t1 a_27_398.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X6 a_121_136.t0 A.t1 a_27_398.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1312 pd=1.05 as=0.1824 ps=1.85 w=0.64 l=0.15
X7 X.t0 a_27_398.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.363225 ps=1.84 w=1.12 l=0.15
R0 A.t1 A.t0 423.118
R1 A A.t1 249.47
R2 a_27_398.t0 a_27_398.n3 393.147
R3 a_27_398.n2 a_27_398.n1 303.039
R4 a_27_398.n3 a_27_398.t1 248.774
R5 a_27_398.n0 a_27_398.t5 246.942
R6 a_27_398.n2 a_27_398.n0 235.577
R7 a_27_398.n0 a_27_398.t4 174.375
R8 a_27_398.n3 a_27_398.n2 47.8123
R9 a_27_398.n1 a_27_398.t3 35.1791
R10 a_27_398.n1 a_27_398.t2 35.1791
R11 VPWR.n6 VPWR.n5 624.508
R12 VPWR.n3 VPWR.n1 587.927
R13 VPWR.n4 VPWR.n0 585
R14 VPWR.n3 VPWR.n2 297.137
R15 VPWR.n2 VPWR.n0 70.3025
R16 VPWR.n5 VPWR.t1 46.9053
R17 VPWR.n5 VPWR.t0 46.9053
R18 VPWR.n1 VPWR.t3 36.3517
R19 VPWR.n2 VPWR.t2 21.8518
R20 VPWR.n6 VPWR.n4 14.3287
R21 VPWR.n1 VPWR.n0 12.8993
R22 VPWR.n4 VPWR.n3 2.92683
R23 VPWR VPWR.n6 0.401709
R24 VPB.t3 VPB.t2 444.356
R25 VPB.t0 VPB.t1 280.914
R26 VPB VPB.t0 257.93
R27 VPB.t1 VPB.t3 229.839
R28 C.n0 C.t0 215.093
R29 C.n0 C.t1 190.19
R30 C C.n0 154.133
R31 B.n0 B.t0 224.667
R32 B.n0 B.t1 162.274
R33 B B.n0 152.41
R34 a_233_136.n0 a_233_136.t1 37.8045
R35 a_233_136.n0 a_233_136.t0 21.7331
R36 a_233_136.n1 a_233_136.n0 19.2005
R37 VGND VGND.n0 127.731
R38 VGND.n0 VGND.t0 41.2505
R39 VGND.n0 VGND.t1 30.2643
R40 VNB.t0 VNB.t2 1339.63
R41 VNB.t1 VNB.t3 1293.44
R42 VNB VNB.t1 1224.15
R43 VNB.t3 VNB.t0 1097.11
R44 a_121_136.t0 a_121_136.t1 76.8755
R45 X X.n0 590.615
R46 X.n2 X.n0 585
R47 X.n1 X.n0 585
R48 X X.t1 203.68
R49 X.n0 X.t0 26.3844
R50 X X.n1 13.6987
R51 X X.n2 12.3514
R52 X.n2 X 4.26717
R53 X.n1 X 2.9198
C0 VPB C 0.054761f
C1 A B 0.07502f
C2 A C 0.004285f
C3 VPB VPWR 0.091247f
C4 VPB X 0.012715f
C5 A VPWR 0.015835f
C6 B C 0.082699f
C7 VPB VGND 0.008493f
C8 B VPWR 0.01686f
C9 B X 0.003414f
C10 A VGND 0.168609f
C11 C VPWR 0.019564f
C12 C X 0.00155f
C13 B VGND 0.009385f
C14 C VGND 0.0291f
C15 VPWR X 0.09515f
C16 VPWR VGND 0.048262f
C17 X VGND 0.094092f
C18 VPB A 0.044791f
C19 VPB B 0.044093f
C20 VGND VNB 0.392833f
C21 X VNB 0.110557f
C22 VPWR VNB 0.305242f
C23 C VNB 0.111723f
C24 B VNB 0.097478f
C25 A VNB 0.2408f
C26 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4_1 VNB VPB VPWR VGND A B C D X
X0 a_257_74.t1 B.t0 a_179_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.0768 ps=0.88 w=0.64 l=0.15
X1 a_96_74.t1 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2898 ps=2.37 w=0.84 l=0.15
X2 VGND.t1 D.t0 a_335_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1277 pd=1.1 as=0.1344 ps=1.06 w=0.64 l=0.15
X3 VPWR.t3 D.t1 a_96_74.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2198 pd=1.555 as=0.147 ps=1.19 w=0.84 l=0.15
X4 VPWR.t4 B.t1 a_96_74.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.4 as=0.147 ps=1.19 w=0.84 l=0.15
X5 X.t1 a_96_74.t5 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2198 ps=1.555 w=1.12 l=0.15
X6 a_335_74.t0 C.t0 a_257_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
X7 X.t0 a_96_74.t6 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1277 ps=1.1 w=0.74 l=0.15
X8 a_179_74.t0 A.t1 a_96_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1696 ps=1.81 w=0.64 l=0.15
X9 a_96_74.t2 C.t1 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2352 ps=1.4 w=0.84 l=0.15
R0 B.n0 B.t0 274.971
R1 B.n0 B.t1 246.05
R2 B B.n0 154.327
R3 a_179_74.t0 a_179_74.t1 45.0005
R4 a_257_74.t0 a_257_74.t1 45.0005
R5 VNB VNB.t3 1893.96
R6 VNB.t0 VNB.t2 1316.54
R7 VNB.t2 VNB.t1 1177.95
R8 VNB.t4 VNB.t0 900.788
R9 VNB.t3 VNB.t4 900.788
R10 A.n0 A.t0 251.444
R11 A.n1 A.t1 165.482
R12 A A.n0 153.477
R13 A.n2 A.n1 152
R14 A.n1 A.n0 49.6611
R15 A A.n2 9.68255
R16 A.n2 A 2.46204
R17 VPWR.n6 VPWR.t1 363.021
R18 VPWR.n2 VPWR.n1 321.678
R19 VPWR.n4 VPWR.n3 305.721
R20 VPWR.n3 VPWR.t2 65.6672
R21 VPWR.n3 VPWR.t4 65.6672
R22 VPWR.n1 VPWR.t3 55.1136
R23 VPWR.n1 VPWR.t0 42.7253
R24 VPWR.n5 VPWR.n4 29.7417
R25 VPWR.n6 VPWR.n5 20.7064
R26 VPWR.n5 VPWR.n0 9.3005
R27 VPWR.n7 VPWR.n6 9.3005
R28 VPWR.n4 VPWR.n2 3.93908
R29 VPWR.n2 VPWR.n0 0.402172
R30 VPWR.n7 VPWR.n0 0.122949
R31 VPWR VPWR.n7 0.0617245
R32 a_96_74.n4 a_96_74.n3 306.132
R33 a_96_74.n2 a_96_74.n0 306.132
R34 a_96_74.n1 a_96_74.t5 258.582
R35 a_96_74.n3 a_96_74.t0 252.165
R36 a_96_74.n2 a_96_74.n1 215.593
R37 a_96_74.n1 a_96_74.t6 210.114
R38 a_96_74.n3 a_96_74.n2 70.024
R39 a_96_74.n0 a_96_74.t2 46.9053
R40 a_96_74.n4 a_96_74.t4 46.9053
R41 a_96_74.n0 a_96_74.t3 35.1791
R42 a_96_74.t1 a_96_74.n4 35.1791
R43 VPB.t3 VPB.t1 362.635
R44 VPB.t2 VPB.t4 298.791
R45 VPB VPB.t0 283.469
R46 VPB.t1 VPB.t2 255.376
R47 VPB.t0 VPB.t3 255.376
R48 D.n0 D.t1 280.899
R49 D.n0 D.t0 236.18
R50 D D.n0 156.614
R51 a_335_74.t0 a_335_74.t1 78.7505
R52 VGND VGND.n0 122.925
R53 VGND.n0 VGND.t0 37.6611
R54 VGND.n0 VGND.t1 26.2505
R55 X.n0 X.t1 290.902
R56 X.t0 X.n0 279.738
R57 X.n1 X.t0 279.738
R58 X.n1 X 7.63353
R59 X.n0 X 2.93628
R60 X X.n1 1.05738
R61 C.n0 C.t1 251.444
R62 C.n1 C.t0 162.274
R63 C C.n0 153.745
R64 C.n2 C.n1 152
R65 C.n1 C.n0 49.6611
R66 C C.n2 11.4429
R67 C.n2 C 2.90959
C0 VPB A 0.061237f
C1 VPWR VGND 0.055104f
C2 VPB B 0.055609f
C3 X VGND 0.114748f
C4 VPB C 0.05463f
C5 A B 0.144096f
C6 VPB D 0.057473f
C7 B C 0.176247f
C8 VPB VPWR 0.098563f
C9 A VPWR 0.018982f
C10 VPB X 0.014028f
C11 B D 4.01e-20
C12 B VPWR 0.02169f
C13 C D 0.117129f
C14 VPB VGND 0.008852f
C15 A VGND 0.012387f
C16 C VPWR 0.019733f
C17 D VPWR 0.016952f
C18 C X 0.005998f
C19 B VGND 0.033555f
C20 C VGND 0.064837f
C21 D X 0.003097f
C22 VPWR X 0.100254f
C23 D VGND 0.030937f
C24 VGND VNB 0.436836f
C25 X VNB 0.121725f
C26 VPWR VNB 0.365279f
C27 D VNB 0.116599f
C28 C VNB 0.117081f
C29 B VNB 0.111803f
C30 A VNB 0.170773f
C31 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3b_4 VNB VPB VPWR VGND X B C A_N
X0 a_239_98.t2 a_27_74.t2 a_298_368.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 VGND.t5 a_298_368.t8 X.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_498_98.t3 C.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 X.t2 a_298_368.t9 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.12945 ps=1.1 w=0.74 l=0.15
X4 a_498_98.t0 B.t0 a_239_98.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 VGND.t1 A_N.t0 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1888 pd=1.87 as=0.1824 ps=1.85 w=0.64 l=0.15
X6 VPWR.t7 B.t1 a_298_368.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.23 pd=1.46 as=0.15 ps=1.3 w=1 l=0.15
X7 a_298_368.t7 B.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X8 a_298_368.t0 a_27_74.t3 a_239_98.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X9 X.t1 a_298_368.t10 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.111 ps=1.04 w=0.74 l=0.15
X10 VPWR.t5 a_298_368.t11 X.t6 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X11 X.t5 a_298_368.t12 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2382 ps=1.555 w=1.12 l=0.15
X12 VPWR.t0 A_N.t1 a_27_74.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.295 ps=2.59 w=1 l=0.15
X13 VPWR.t9 C.t1 a_298_368.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.15 ps=1.3 w=1 l=0.15
X14 a_298_368.t6 C.t2 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.23 ps=1.46 w=1 l=0.15
X15 VGND.t2 a_298_368.t13 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1295 ps=1.09 w=0.74 l=0.15
X16 VGND.t6 C.t3 a_498_98.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.12945 pd=1.1 as=0.0896 ps=0.92 w=0.64 l=0.15
X17 VPWR.t2 a_27_74.t4 a_298_368.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X18 a_298_368.t2 a_27_74.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X19 X.t4 a_298_368.t14 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X20 a_239_98.t3 B.t3 a_498_98.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.112 ps=0.99 w=0.64 l=0.15
R0 a_27_74.t1 a_27_74.n3 240.571
R1 a_27_74.n0 a_27_74.t4 215.561
R2 a_27_74.n2 a_27_74.t5 215.561
R3 a_27_74.n3 a_27_74.t0 213.233
R4 a_27_74.n3 a_27_74.n2 198.956
R5 a_27_74.n0 a_27_74.t2 188.161
R6 a_27_74.n1 a_27_74.t3 163.881
R7 a_27_74.n1 a_27_74.n0 45.2793
R8 a_27_74.n2 a_27_74.n1 20.449
R9 a_298_368.n11 a_298_368.t12 289.041
R10 a_298_368.n17 a_298_368.n0 261.849
R11 a_298_368.n4 a_298_368.t8 245.929
R12 a_298_368.n4 a_298_368.n3 209.403
R13 a_298_368.n7 a_298_368.t14 209.403
R14 a_298_368.n10 a_298_368.t11 209.403
R15 a_298_368.n16 a_298_368.n15 202.178
R16 a_298_368.n14 a_298_368.n1 201.501
R17 a_298_368.n18 a_298_368.n17 201.069
R18 a_298_368.n11 a_298_368.t9 179.947
R19 a_298_368.n8 a_298_368.t13 179.947
R20 a_298_368.n5 a_298_368.t10 179.947
R21 a_298_368.n6 a_298_368.n2 165.189
R22 a_298_368.n13 a_298_368.n12 152
R23 a_298_368.n9 a_298_368.n2 152
R24 a_298_368.n14 a_298_368.n13 104.251
R25 a_298_368.n16 a_298_368.n14 54.9652
R26 a_298_368.n17 a_298_368.n16 46.4944
R27 a_298_368.n10 a_298_368.n9 32.4949
R28 a_298_368.n1 a_298_368.t5 29.5505
R29 a_298_368.n1 a_298_368.t6 29.5505
R30 a_298_368.n15 a_298_368.t4 29.5505
R31 a_298_368.n15 a_298_368.t7 29.5505
R32 a_298_368.n18 a_298_368.t3 29.5505
R33 a_298_368.t2 a_298_368.n18 29.5505
R34 a_298_368.n0 a_298_368.t1 26.2505
R35 a_298_368.n0 a_298_368.t0 26.2505
R36 a_298_368.n6 a_298_368.n5 21.1218
R37 a_298_368.n5 a_298_368.n4 17.8724
R38 a_298_368.n8 a_298_368.n7 17.8724
R39 a_298_368.n13 a_298_368.n2 13.1884
R40 a_298_368.n7 a_298_368.n6 9.74881
R41 a_298_368.n9 a_298_368.n8 9.20724
R42 a_298_368.n12 a_298_368.n11 8.1241
R43 a_298_368.n12 a_298_368.n10 4.33308
R44 a_239_98.n0 a_239_98.t3 297.853
R45 a_239_98.n0 a_239_98.t1 193.889
R46 a_239_98.n1 a_239_98.n0 97.3258
R47 a_239_98.n1 a_239_98.t0 26.2505
R48 a_239_98.t2 a_239_98.n1 26.2505
R49 VNB.t1 VNB.t3 2448.29
R50 VNB.t10 VNB.t0 2286.61
R51 VNB.t9 VNB.t7 1177.95
R52 VNB.t7 VNB.t5 1154.86
R53 VNB.t2 VNB.t10 1154.86
R54 VNB VNB.t1 1143.31
R55 VNB.t5 VNB.t6 1039.37
R56 VNB.t6 VNB.t8 993.177
R57 VNB.t0 VNB.t9 993.177
R58 VNB.t4 VNB.t2 993.177
R59 VNB.t3 VNB.t4 993.177
R60 X.n4 X.n3 258.046
R61 X.n4 X.t4 233.983
R62 X.n2 X.n0 155.478
R63 X.n2 X.n1 105.553
R64 X.n5 X.n2 56.492
R65 X X.n5 42.9509
R66 X.n0 X.t2 34.0546
R67 X.n3 X.t6 26.3844
R68 X.n3 X.t5 26.3844
R69 X.n1 X.t3 22.7032
R70 X.n1 X.t1 22.7032
R71 X.n0 X.t0 22.7032
R72 X.n5 X.n4 9.03579
R73 VGND.n14 VGND.t0 237.433
R74 VGND.n7 VGND.n6 209.243
R75 VGND.n5 VGND.t5 170.638
R76 VGND.n22 VGND.t1 156.772
R77 VGND.n10 VGND.n9 116.819
R78 VGND.n9 VGND.t6 41.0701
R79 VGND.n16 VGND.n15 36.1417
R80 VGND.n16 VGND.n1 36.1417
R81 VGND.n20 VGND.n1 36.1417
R82 VGND.n21 VGND.n20 36.1417
R83 VGND.n15 VGND.n14 30.4946
R84 VGND.n10 VGND.n3 28.9887
R85 VGND.n8 VGND.n7 26.7299
R86 VGND.n6 VGND.t3 25.9464
R87 VGND.n22 VGND.n21 24.4711
R88 VGND.n6 VGND.t2 22.7032
R89 VGND.n9 VGND.t4 21.1849
R90 VGND.n10 VGND.n8 18.4476
R91 VGND.n14 VGND.n3 16.9417
R92 VGND.n21 VGND.n0 9.3005
R93 VGND.n20 VGND.n19 9.3005
R94 VGND.n18 VGND.n1 9.3005
R95 VGND.n17 VGND.n16 9.3005
R96 VGND.n15 VGND.n2 9.3005
R97 VGND.n14 VGND.n13 9.3005
R98 VGND.n12 VGND.n3 9.3005
R99 VGND.n11 VGND.n10 9.3005
R100 VGND.n8 VGND.n4 9.3005
R101 VGND.n23 VGND.n22 7.43488
R102 VGND.n7 VGND.n5 6.39244
R103 VGND.n5 VGND.n4 0.709244
R104 VGND VGND.n23 0.160103
R105 VGND.n23 VGND.n0 0.1477
R106 VGND.n11 VGND.n4 0.122949
R107 VGND.n12 VGND.n11 0.122949
R108 VGND.n13 VGND.n12 0.122949
R109 VGND.n13 VGND.n2 0.122949
R110 VGND.n17 VGND.n2 0.122949
R111 VGND.n18 VGND.n17 0.122949
R112 VGND.n19 VGND.n18 0.122949
R113 VGND.n19 VGND.n0 0.122949
R114 C.n0 C.t3 245.314
R115 C.n0 C.t1 207.529
R116 C.n2 C.t2 207.529
R117 C C.n2 170.834
R118 C.n1 C.t0 133.353
R119 C.n2 C.n1 43.6342
R120 C.n1 C.n0 2.02997
R121 a_498_98.n1 a_498_98.n0 383.808
R122 a_498_98.n0 a_498_98.t0 39.3755
R123 a_498_98.n0 a_498_98.t1 26.2505
R124 a_498_98.t2 a_498_98.n1 26.2505
R125 a_498_98.n1 a_498_98.t3 26.2505
R126 B.n0 B.t1 207.529
R127 B.n1 B.t2 207.529
R128 B.n0 B.t3 181.797
R129 B.n1 B.t0 173.52
R130 B.n3 B.n2 152
R131 B.n2 B.n0 54.7732
R132 B.n3 B 12.354
R133 B.n2 B.n1 10.955
R134 B B.n3 1.93538
R135 A_N.n0 A_N.t1 279.341
R136 A_N.n0 A_N.t0 183.014
R137 A_N A_N.n0 157.237
R138 VPWR.n7 VPWR.n6 323.93
R139 VPWR.n1 VPWR.n0 322.322
R140 VPWR.n15 VPWR.n3 319.616
R141 VPWR.n5 VPWR.n4 319.616
R142 VPWR.n9 VPWR.n8 223.696
R143 VPWR.n4 VPWR.t8 51.2205
R144 VPWR.n8 VPWR.t9 46.2955
R145 VPWR.n0 VPWR.t1 39.4005
R146 VPWR.n0 VPWR.t0 39.4005
R147 VPWR.n3 VPWR.t6 39.4005
R148 VPWR.n3 VPWR.t2 39.4005
R149 VPWR.n4 VPWR.t7 39.4005
R150 VPWR.n10 VPWR.n9 35.3887
R151 VPWR.n8 VPWR.t4 35.2408
R152 VPWR.n6 VPWR.t3 35.1791
R153 VPWR.n6 VPWR.t5 35.1791
R154 VPWR.n16 VPWR.n1 28.2358
R155 VPWR.n14 VPWR.n5 25.224
R156 VPWR.n15 VPWR.n14 25.224
R157 VPWR.n16 VPWR.n15 22.2123
R158 VPWR.n10 VPWR.n5 22.2123
R159 VPWR.n11 VPWR.n10 9.3005
R160 VPWR.n12 VPWR.n5 9.3005
R161 VPWR.n14 VPWR.n13 9.3005
R162 VPWR.n15 VPWR.n2 9.3005
R163 VPWR.n17 VPWR.n16 9.3005
R164 VPWR.n18 VPWR.n1 6.88467
R165 VPWR.n9 VPWR.n7 5.96665
R166 VPWR.n11 VPWR.n7 0.485762
R167 VPWR VPWR.n18 0.270511
R168 VPWR.n18 VPWR.n17 0.160218
R169 VPWR.n12 VPWR.n11 0.122949
R170 VPWR.n13 VPWR.n12 0.122949
R171 VPWR.n13 VPWR.n2 0.122949
R172 VPWR.n17 VPWR.n2 0.122949
R173 VPB VPB.t0 441.801
R174 VPB.t7 VPB.t8 311.56
R175 VPB.t9 VPB.t4 298.791
R176 VPB.t5 VPB.t3 280.914
R177 VPB.t2 VPB.t6 280.914
R178 VPB.t0 VPB.t1 280.914
R179 VPB.t4 VPB.t5 229.839
R180 VPB.t8 VPB.t9 229.839
R181 VPB.t6 VPB.t7 229.839
R182 VPB.t1 VPB.t2 229.839
C0 X A_N 3.94e-20
C1 X B 7.08e-20
C2 VGND VPB 0.013536f
C3 X C 0.001514f
C4 VGND A_N 0.044106f
C5 X VPWR 0.46756f
C6 VGND B 0.014478f
C7 VPB A_N 0.043959f
C8 VGND C 0.038575f
C9 VPB B 0.066959f
C10 VGND VPWR 0.112987f
C11 VPB C 0.086707f
C12 VPB VPWR 0.219147f
C13 A_N C 1.96e-19
C14 A_N VPWR 0.018446f
C15 B C 0.080178f
C16 B VPWR 0.033297f
C17 X VGND 0.31573f
C18 C VPWR 0.03868f
C19 X VPB 0.021155f
C20 VGND VNB 0.852692f
C21 X VNB 0.055363f
C22 VPWR VNB 0.655188f
C23 C VNB 0.258255f
C24 B VNB 0.197056f
C25 A_N VNB 0.177115f
C26 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3b_2 VNB VPB VPWR VGND A_N C B X
X0 X.t1 a_284_368.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1 VGND.t1 a_284_368.t5 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t3 a_27_88.t2 a_284_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.295 ps=2.59 w=1 l=0.15
X3 VGND.t3 A_N.t0 a_27_88.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.16225 pd=1.69 as=0.15675 ps=1.67 w=0.55 l=0.15
X4 VPWR.t5 C.t0 a_284_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2127 pd=1.51 as=0.15 ps=1.3 w=1 l=0.15
X5 a_284_368.t1 B.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.21 ps=1.42 w=1 l=0.15
X6 X.t3 a_284_368.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.2127 ps=1.51 w=1.12 l=0.15
X7 a_376_74.t0 a_27_88.t3 a_284_368.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VPWR.t0 A_N.t1 a_27_88.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2562 pd=2.29 as=0.2478 ps=2.27 w=0.84 l=0.15
X9 VGND.t2 C.t1 a_454_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X10 a_454_74.t1 B.t1 a_376_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X11 VPWR.t1 a_284_368.t7 X.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
R0 a_284_368.n4 a_284_368.n3 346.307
R1 a_284_368.n3 a_284_368.t7 240.197
R2 a_284_368.n1 a_284_368.t6 240.197
R3 a_284_368.n0 a_284_368.t3 230.7
R4 a_284_368.n5 a_284_368.n4 194.815
R5 a_284_368.n1 a_284_368.t4 182.138
R6 a_284_368.n0 a_284_368.t0 181.769
R7 a_284_368.n2 a_284_368.t5 179.947
R8 a_284_368.n2 a_284_368.n1 60.6157
R9 a_284_368.n4 a_284_368.n0 58.053
R10 a_284_368.n5 a_284_368.t2 29.5505
R11 a_284_368.t1 a_284_368.n5 29.5505
R12 a_284_368.n3 a_284_368.n2 7.30353
R13 VGND.n11 VGND.t3 239.595
R14 VGND.n2 VGND.t1 178.633
R15 VGND.n4 VGND.n3 116.644
R16 VGND.n3 VGND.t0 45.4059
R17 VGND.n5 VGND.n1 36.1417
R18 VGND.n9 VGND.n1 36.1417
R19 VGND.n10 VGND.n9 36.1417
R20 VGND.n11 VGND.n10 24.4711
R21 VGND.n3 VGND.t2 22.7032
R22 VGND.n5 VGND.n4 13.177
R23 VGND.n10 VGND.n0 9.3005
R24 VGND.n9 VGND.n8 9.3005
R25 VGND.n7 VGND.n1 9.3005
R26 VGND.n6 VGND.n5 9.3005
R27 VGND.n12 VGND.n11 7.19894
R28 VGND.n4 VGND.n2 7.18692
R29 VGND.n6 VGND.n2 0.537296
R30 VGND VGND.n12 0.156997
R31 VGND.n12 VGND.n0 0.150766
R32 VGND.n7 VGND.n6 0.122949
R33 VGND.n8 VGND.n7 0.122949
R34 VGND.n8 VGND.n0 0.122949
R35 X X.n0 601.997
R36 X.n2 X.n1 185
R37 X.n3 X.n2 185
R38 X.n0 X.t2 28.1434
R39 X.n0 X.t3 27.2639
R40 X.n2 X.t0 22.7032
R41 X.n2 X.t1 22.7032
R42 X.n3 X 12.6066
R43 X.n1 X 9.75788
R44 X.n1 X 4.84898
R45 X X.n3 1.74595
R46 VNB.t3 VNB.t4 3025.72
R47 VNB.t2 VNB.t1 1316.54
R48 VNB.t5 VNB.t2 1316.54
R49 VNB VNB.t3 1143.31
R50 VNB.t1 VNB.t0 993.177
R51 VNB.t4 VNB.t5 900.788
R52 a_27_88.t0 a_27_88.n1 469.452
R53 a_27_88.n1 a_27_88.t1 288.829
R54 a_27_88.n0 a_27_88.t2 226.273
R55 a_27_88.n1 a_27_88.n0 157.877
R56 a_27_88.n0 a_27_88.t3 144.696
R57 VPWR.n3 VPWR.t1 825.821
R58 VPWR.n12 VPWR.t0 649.472
R59 VPWR.n5 VPWR.n4 608.856
R60 VPWR.n2 VPWR.n1 319.616
R61 VPWR.n4 VPWR.t5 47.2805
R62 VPWR.n1 VPWR.t4 43.3405
R63 VPWR.n1 VPWR.t3 39.4005
R64 VPWR.n11 VPWR.n10 36.1417
R65 VPWR.n6 VPWR.n2 30.8711
R66 VPWR.n4 VPWR.t2 26.8503
R67 VPWR.n6 VPWR.n5 24.0946
R68 VPWR.n12 VPWR.n11 22.5887
R69 VPWR.n10 VPWR.n2 16.5652
R70 VPWR.n7 VPWR.n6 9.3005
R71 VPWR.n8 VPWR.n2 9.3005
R72 VPWR.n10 VPWR.n9 9.3005
R73 VPWR.n11 VPWR.n0 9.3005
R74 VPWR.n13 VPWR.n12 7.28976
R75 VPWR.n5 VPWR.n3 6.58468
R76 VPWR.n7 VPWR.n3 0.670526
R77 VPWR VPWR.n13 0.158192
R78 VPWR.n13 VPWR.n0 0.149586
R79 VPWR.n8 VPWR.n7 0.122949
R80 VPWR.n9 VPWR.n8 0.122949
R81 VPWR.n9 VPWR.n0 0.122949
R82 VPB.t0 VPB.t3 656.317
R83 VPB.t3 VPB.t4 291.13
R84 VPB.t5 VPB.t2 275.807
R85 VPB VPB.t0 257.93
R86 VPB.t2 VPB.t1 237.5
R87 VPB.t4 VPB.t5 229.839
R88 A_N.n0 A_N.t1 235.811
R89 A_N.n0 A_N.t0 218.167
R90 A_N A_N.n0 68.3727
R91 C.n0 C.t0 231.629
R92 C.n0 C.t1 220.113
R93 C C.n0 157.358
R94 B.n0 B.t0 266.44
R95 B.n0 B.t1 178.34
R96 B.n1 B.n0 152
R97 B B.n1 6.16346
R98 B.n1 B 5.53136
R99 a_376_74.t0 a_376_74.t1 38.9194
R100 a_454_74.t0 a_454_74.t1 68.1086
C0 C VGND 0.051637f
C1 X VGND 0.156708f
C2 VPB A_N 0.075204f
C3 VPB VPWR 0.150356f
C4 A_N VPWR 0.018523f
C5 VPB B 0.033064f
C6 VPB C 0.036846f
C7 A_N B 1.35e-19
C8 VPB X 0.00345f
C9 VPWR B 0.017864f
C10 VPB VGND 0.012547f
C11 A_N X 1.26e-19
C12 VPWR C 0.017707f
C13 A_N VGND 0.015577f
C14 B C 0.090714f
C15 VPWR X 0.019181f
C16 VPWR VGND 0.073612f
C17 B X 0.005424f
C18 B VGND 0.075761f
C19 C X 0.03679f
C20 VGND VNB 0.5999f
C21 X VNB 0.01388f
C22 C VNB 0.10895f
C23 B VNB 0.111276f
C24 VPWR VNB 0.442844f
C25 A_N VNB 0.198284f
C26 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2b_2 VNB VPB VPWR VGND X B A_N
X0 VPWR.t4 A_N.t0 a_27_74.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.25205 pd=1.6 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 a_198_48.t2 a_27_74.t2 a_505_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2 VGND.t3 A_N.t1 a_27_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.13925 pd=1.16 as=0.15675 ps=1.67 w=0.55 l=0.15
X3 VGND.t0 a_198_48.t3 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.29785 pd=1.545 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VPWR.t3 a_27_74.t3 a_198_48.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X5 a_198_48.t0 B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.367275 ps=1.8 w=1 l=0.15
X6 VPWR.t1 a_198_48.t4 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.367275 pd=1.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7 X.t0 a_198_48.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.25205 ps=1.6 w=1.12 l=0.15
X8 X.t2 a_198_48.t6 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.13925 ps=1.16 w=0.74 l=0.15
X9 a_505_74.t1 B.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.29785 ps=1.545 w=0.74 l=0.15
R0 A_N.n0 A_N.t1 247.749
R1 A_N.n0 A_N.t0 203.03
R2 A_N A_N.n0 158.847
R3 a_27_74.n1 a_27_74.n0 374.312
R4 a_27_74.t1 a_27_74.n1 340.56
R5 a_27_74.n1 a_27_74.t0 318.082
R6 a_27_74.n0 a_27_74.t3 258.406
R7 a_27_74.n0 a_27_74.t2 204.048
R8 VPWR.n4 VPWR.t3 851.471
R9 VPWR.n8 VPWR.n1 679.76
R10 VPWR.n3 VPWR.n2 585
R11 VPWR.n2 VPWR.t0 75.8455
R12 VPWR.n1 VPWR.t4 65.6672
R13 VPWR.n2 VPWR.t1 41.9945
R14 VPWR.n1 VPWR.t2 34.0942
R15 VPWR.n7 VPWR.n6 33.5164
R16 VPWR.n8 VPWR.n7 16.5652
R17 VPWR.n4 VPWR.n3 10.6337
R18 VPWR.n6 VPWR.n5 9.3005
R19 VPWR.n7 VPWR.n0 9.3005
R20 VPWR.n9 VPWR.n8 7.53404
R21 VPWR.n6 VPWR.n3 4.49322
R22 VPWR.n5 VPWR.n4 0.58916
R23 VPWR VPWR.n9 0.161409
R24 VPWR.n9 VPWR.n0 0.146411
R25 VPWR.n5 VPWR.n0 0.122949
R26 VPB.t1 VPB.t0 423.925
R27 VPB.t4 VPB.t2 316.668
R28 VPB VPB.t4 257.93
R29 VPB.t0 VPB.t3 229.839
R30 VPB.t2 VPB.t1 229.839
R31 a_505_74.t0 a_505_74.t1 38.9194
R32 a_198_48.n4 a_198_48.n3 647.665
R33 a_198_48.n3 a_198_48.t2 255.589
R34 a_198_48.n2 a_198_48.t4 240.197
R35 a_198_48.n0 a_198_48.t5 240.197
R36 a_198_48.n0 a_198_48.t6 190.712
R37 a_198_48.n1 a_198_48.t3 179.947
R38 a_198_48.n3 a_198_48.n2 158.573
R39 a_198_48.n1 a_198_48.n0 54.0429
R40 a_198_48.n4 a_198_48.t1 29.5505
R41 a_198_48.t0 a_198_48.n4 29.5505
R42 a_198_48.n2 a_198_48.n1 11.6853
R43 VNB.t1 VNB.t3 2205.77
R44 VNB.t4 VNB.t0 1316.54
R45 VNB VNB.t4 1143.31
R46 VNB.t0 VNB.t1 993.177
R47 VNB.t3 VNB.t2 900.788
R48 VGND.n9 VGND.n8 209.631
R49 VGND.n4 VGND.n3 186.024
R50 VGND.n2 VGND.n1 185
R51 VGND.n3 VGND.n2 73.7843
R52 VGND.n8 VGND.t3 45.8187
R53 VGND.n8 VGND.t1 39.2753
R54 VGND.n2 VGND.t0 34.0546
R55 VGND.n7 VGND.n6 32.4622
R56 VGND.n3 VGND.t2 22.7032
R57 VGND.n9 VGND.n7 19.2005
R58 VGND.n6 VGND.n5 9.3005
R59 VGND.n7 VGND.n0 9.3005
R60 VGND.n10 VGND.n9 7.43488
R61 VGND.n4 VGND.n1 7.43002
R62 VGND.n5 VGND.n4 6.91664
R63 VGND.n6 VGND.n1 1.86911
R64 VGND VGND.n10 0.160103
R65 VGND.n10 VGND.n0 0.1477
R66 VGND.n5 VGND.n0 0.122949
R67 X.n2 X.n1 590.818
R68 X.n2 X.n0 155.022
R69 X.n1 X.t1 26.3844
R70 X.n1 X.t0 26.3844
R71 X.n0 X.t3 22.7032
R72 X.n0 X.t2 22.7032
R73 X X.n2 3.29747
R74 B.n0 B.t0 279.829
R75 B.n0 B.t1 178.34
R76 B B.n0 161.859
C0 VPB VPWR 0.108773f
C1 VPB A_N 0.045021f
C2 VPWR A_N 0.008482f
C3 VPB X 0.002925f
C4 VPWR X 0.015498f
C5 VPB B 0.039778f
C6 A_N X 0.001264f
C7 VPWR B 0.015082f
C8 VPB VGND 0.008271f
C9 VPWR VGND 0.058649f
C10 A_N VGND 0.015497f
C11 X B 6.29e-19
C12 X VGND 0.106619f
C13 B VGND 0.017476f
C14 VGND VNB 0.43222f
C15 B VNB 0.119342f
C16 X VNB 0.00647f
C17 A_N VNB 0.18386f
C18 VPWR VNB 0.363803f
C19 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and2b_1 VNB VPB VPWR VGND B A_N X
X0 VPWR.t3 B.t0 a_266_98.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.555 as=0.126 ps=1.14 w=0.84 l=0.15
X1 a_266_98.t0 a_27_74.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X2 VPWR.t0 A_N.t0 a_27_74.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.8526 ps=3.71 w=0.84 l=0.15
X3 VGND.t2 A_N.t1 a_27_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.19525 pd=1.81 as=0.15675 ps=1.67 w=0.55 l=0.15
X4 VGND.t1 B.t1 a_353_98.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2157 pd=1.375 as=0.0768 ps=0.88 w=0.64 l=0.15
X5 X.t1 a_266_98.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2157 ps=1.375 w=0.74 l=0.15
X6 X.t0 a_266_98.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.231 ps=1.555 w=1.12 l=0.15
X7 a_353_98.t1 a_27_74.t3 a_266_98.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
R0 B.n0 B.t0 203.316
R1 B.n0 B.t1 195.016
R2 B B.n0 156.019
R3 a_266_98.n2 a_266_98.n1 362.289
R4 a_266_98.n0 a_266_98.t4 257.245
R5 a_266_98.n1 a_266_98.n0 236.518
R6 a_266_98.n0 a_266_98.t3 202.35
R7 a_266_98.n1 a_266_98.t1 147.048
R8 a_266_98.n2 a_266_98.t2 35.1791
R9 a_266_98.t0 a_266_98.n2 35.1791
R10 VPWR.n2 VPWR.n1 368.43
R11 VPWR.n2 VPWR.n0 235.833
R12 VPWR.n0 VPWR.t3 56.9954
R13 VPWR.n0 VPWR.t1 36.6056
R14 VPWR.n1 VPWR.t2 35.1791
R15 VPWR.n1 VPWR.t0 35.1791
R16 VPWR VPWR.n2 0.69755
R17 VPB VPB.t0 625.673
R18 VPB.t3 VPB.t1 298.791
R19 VPB.t2 VPB.t3 229.839
R20 VPB.t0 VPB.t2 229.839
R21 a_27_74.n1 a_27_74.n0 319.094
R22 a_27_74.t0 a_27_74.n1 289.599
R23 a_27_74.n0 a_27_74.t2 287.594
R24 a_27_74.n1 a_27_74.t1 264.361
R25 a_27_74.n0 a_27_74.t3 148.618
R26 A_N.n0 A_N.t0 388.94
R27 A_N.n0 A_N.t1 249.263
R28 A_N A_N.n0 153.958
R29 VGND.n1 VGND.t2 259.659
R30 VGND.n1 VGND.n0 95.9164
R31 VGND.n0 VGND.t1 54.4579
R32 VGND.n0 VGND.t0 50.8684
R33 VGND VGND.n1 0.228996
R34 VNB.t3 VNB.t2 2760.1
R35 VNB.t1 VNB.t0 1813.12
R36 VNB VNB.t3 1143.31
R37 VNB.t2 VNB.t1 900.788
R38 a_353_98.t0 a_353_98.t1 45.0005
R39 X.n1 X 588.299
R40 X.n1 X.n0 585
R41 X.n2 X.n1 585
R42 X X.t1 204.071
R43 X.n1 X.t0 26.3844
R44 X X.n2 8.84174
R45 X X.n0 7.65411
R46 X X.n0 2.11184
R47 X.n2 X 0.924211
C0 X VGND 0.076373f
C1 X VPB 0.021944f
C2 VGND VPB 0.009145f
C3 X VPWR 0.140859f
C4 X A_N 4.83e-20
C5 VGND VPWR 0.056817f
C6 VPB VPWR 0.121946f
C7 X B 0.005784f
C8 VGND A_N 0.018743f
C9 VPB A_N 0.085833f
C10 VGND B 0.015253f
C11 VPWR A_N 0.015898f
C12 VPB B 0.040465f
C13 VPWR B 0.028993f
C14 VGND VNB 0.456563f
C15 X VNB 0.109473f
C16 B VNB 0.109839f
C17 A_N VNB 0.225851f
C18 VPWR VNB 0.367254f
C19 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__buf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__buf_2 VNB VPB VPWR VGND A X
X0 a_21_260.t0 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.64 as=0.2102 ps=1.505 w=1 l=0.15
X1 VGND.t1 a_21_260.t2 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR.t0 a_21_260.t3 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X.t0 a_21_260.t4 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.756 ps=3.59 w=1.12 l=0.15
X4 a_21_260.t1 A.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.15535 ps=1.17 w=0.64 l=0.15
X5 X.t2 a_21_260.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
R0 A.n0 A.t0 228.737
R1 A.n0 A.t1 201.155
R2 A A.n0 154.53
R3 VPWR.n1 VPWR.n0 612.011
R4 VPWR.n1 VPWR.t1 215.78
R5 VPWR.n0 VPWR.t2 46.2955
R6 VPWR.n0 VPWR.t0 27.0196
R7 VPWR VPWR.n1 0.347023
R8 a_21_260.t0 a_21_260.n2 256.697
R9 a_21_260.n2 a_21_260.t1 252.517
R10 a_21_260.n2 a_21_260.n0 250.502
R11 a_21_260.n1 a_21_260.t3 242.162
R12 a_21_260.n0 a_21_260.t4 240.197
R13 a_21_260.n1 a_21_260.t2 180.631
R14 a_21_260.n0 a_21_260.t5 179.947
R15 a_21_260.n0 a_21_260.n1 63.582
R16 VPB VPB.t0 452.017
R17 VPB.t1 VPB.t2 273.253
R18 VPB.t0 VPB.t1 229.839
R19 X X.n0 586.212
R20 X X.n1 106.046
R21 X.n0 X.t1 26.3844
R22 X.n0 X.t0 26.3844
R23 X.n1 X.t3 22.7032
R24 X.n1 X.t2 22.7032
R25 VGND.n1 VGND.n0 216.882
R26 VGND.n1 VGND.t0 177.453
R27 VGND.n0 VGND.t2 41.2505
R28 VGND.n0 VGND.t1 30.6984
R29 VGND VGND.n1 0.481408
R30 VNB VNB.t0 2067.19
R31 VNB.t1 VNB.t2 1339.63
R32 VNB.t0 VNB.t1 993.177
C0 VPB VPWR 0.080872f
C1 VPB X 0.002197f
C2 VPWR X 0.015598f
C3 VPB A 0.043503f
C4 VPB VGND 0.005736f
C5 VPWR A 0.012333f
C6 VPWR VGND 0.042955f
C7 X A 9.2e-19
C8 X VGND 0.145698f
C9 A VGND 0.014195f
C10 VGND VNB 0.379666f
C11 A VNB 0.163061f
C12 X VNB 0.011471f
C13 VPWR VNB 0.308452f
C14 VPB VNB 0.620496f
.ends

* NGSPICE file created from sky130_fd_sc_hs__buf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__buf_1 VNB VPB VPWR VGND A X
X0 VGND.t1 A.t0 a_27_164.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.24915 ps=2.37 w=0.55 l=0.15
X1 X.t1 a_27_164.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X2 X.t0 a_27_164.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2051 ps=1.52 w=1.12 l=0.15
X3 VPWR.t1 A.t1 a_27_164.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2051 pd=1.52 as=0.2478 ps=2.27 w=0.84 l=0.15
R0 A.n0 A.t1 234.841
R1 A.n0 A.t0 197.62
R2 A.n1 A.n0 100.508
R3 A.n1 A 14.6021
R4 A A.n1 3.80117
R5 a_27_164.t0 a_27_164.n1 459.712
R6 a_27_164.n0 a_27_164.t3 263.589
R7 a_27_164.n0 a_27_164.t2 203.339
R8 a_27_164.n1 a_27_164.t1 196.582
R9 a_27_164.n1 a_27_164.n0 152
R10 VGND VGND.n0 124.972
R11 VGND.n0 VGND.t1 51.1752
R12 VGND.n0 VGND.t0 32.4566
R13 VNB VNB.t1 1951.71
R14 VNB.t1 VNB.t0 1339.63
R15 X.n1 X 589.444
R16 X.n1 X.n0 585
R17 X.n2 X.n1 585
R18 X X.t1 206.337
R19 X.n1 X.t0 26.3844
R20 X X.n2 11.9116
R21 X X.n0 10.3116
R22 X X.n0 2.84494
R23 X.n2 X 1.24494
R24 VPWR VPWR.n0 322.007
R25 VPWR.n0 VPWR.t1 46.9053
R26 VPWR.n0 VPWR.t0 42.7253
R27 VPB VPB.t1 439.248
R28 VPB.t1 VPB.t0 280.914
C0 VPB A 0.097814f
C1 VPB VPWR 0.063751f
C2 A VPWR 0.024849f
C3 VPB X 0.013871f
C4 A X 0.002797f
C5 VPB VGND 0.00763f
C6 VPWR X 0.09996f
C7 A VGND 0.014584f
C8 VPWR VGND 0.031858f
C9 X VGND 0.090589f
C10 VGND VNB 0.301636f
C11 X VNB 0.111672f
C12 VPWR VNB 0.227682f
C13 A VNB 0.191502f
C14 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4bb_4 VNB VPB VPWR VGND B_N A_N D C X
X0 VPWR.t11 B_N.t0 a_27_74.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.295 ps=2.59 w=1 l=0.15
X1 VPWR.t13 a_200_74.t2 a_472_388.t7 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.235 ps=1.47 w=1 l=0.15
X2 VPWR.t0 a_472_388.t10 X.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_685_140.t1 a_27_74.t2 a_412_140.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 VPWR.t4 C.t0 a_472_388.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.61 pd=2.22 as=0.15 ps=1.3 w=1 l=0.15
X5 X.t2 a_472_388.t11 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_200_74.t1 A_N.t0 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2 ps=1.4 w=1 l=0.15
X7 a_472_388.t6 a_200_74.t3 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.235 pd=1.47 as=0.32 ps=2.64 w=1 l=0.15
X8 VPWR.t2 a_472_388.t12 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_472_388.t1 C.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X10 X.t0 a_472_388.t13 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2102 ps=1.505 w=1.12 l=0.15
X11 a_882_137# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X12 VPWR.t6 D.t0 a_472_388.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2102 pd=1.505 as=0.18625 ps=1.455 w=1 l=0.15
X13 VGND.t4 B_N.t1 a_27_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X14 X.t5 a_472_388.t14 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1245 ps=1.09 w=0.74 l=0.15
X15 a_412_140.t0 a_27_74.t3 a_685_140.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 a_685_140.t2 C.t2 a_882_137# VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2272 ps=1.99 w=0.64 l=0.15
X17 X.t4 a_472_388.t15 VGND.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1406 ps=1.12 w=0.74 l=0.15
X18 a_472_388.t9 a_200_74.t4 a_412_140.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2272 ps=1.99 w=0.64 l=0.15
X19 a_472_388.t5 a_27_74.t4 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR.t8 a_27_74.t5 a_472_388.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.165 ps=1.33 w=1 l=0.15
X21 a_200_74.t0 A_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1915 pd=1.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X22 a_472_388.t3 D.t1 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.18625 pd=1.455 as=0.61 ps=2.22 w=1 l=0.15
X23 a_412_140.t2 a_200_74.t5 a_472_388.t8 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X24 a_882_137# C.t3 a_685_140.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X25 VGND.t1 D.t2 a_882_137# VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1245 pd=1.09 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 B_N.n0 B_N.t1 268.313
R1 B_N.n0 B_N.t0 239.54
R2 B_N.n1 B_N.n0 152
R3 B_N.n1 B_N 9.69747
R4 B_N B_N.n1 8.92171
R5 a_27_74.t2 a_27_74.t4 430.079
R6 a_27_74.t3 a_27_74.t5 422.152
R7 a_27_74.t0 a_27_74.n1 371.697
R8 a_27_74.n1 a_27_74.n0 257.995
R9 a_27_74.n1 a_27_74.t1 242.804
R10 a_27_74.n0 a_27_74.t3 220.113
R11 a_27_74.n0 a_27_74.t2 152.925
R12 VPWR.n2 VPWR.t10 798.005
R13 VPWR.n13 VPWR.t0 349.373
R14 VPWR.n17 VPWR.n12 315.928
R15 VPWR.n40 VPWR.n1 315.926
R16 VPWR.n15 VPWR.n14 315.812
R17 VPWR.n26 VPWR.n25 292.5
R18 VPWR.n24 VPWR.n23 292.5
R19 VPWR.n22 VPWR.n9 292.5
R20 VPWR.n33 VPWR.n4 223.115
R21 VPWR.n6 VPWR.n5 223.115
R22 VPWR.n24 VPWR.n9 85.6955
R23 VPWR.n25 VPWR.n24 85.6955
R24 VPWR.n12 VPWR.t6 46.2955
R25 VPWR.n25 VPWR.t4 39.4005
R26 VPWR.n1 VPWR.t12 39.4005
R27 VPWR.n1 VPWR.t11 39.4005
R28 VPWR.n5 VPWR.t5 39.4005
R29 VPWR.n5 VPWR.t8 39.4005
R30 VPWR.n39 VPWR.n38 36.1417
R31 VPWR.n4 VPWR.t9 33.4905
R32 VPWR.n28 VPWR.n27 31.348
R33 VPWR.n34 VPWR.n2 31.2476
R34 VPWR.n17 VPWR.n10 29.7417
R35 VPWR.n9 VPWR.t7 29.5505
R36 VPWR.n4 VPWR.t13 29.5505
R37 VPWR.n32 VPWR.n6 27.4829
R38 VPWR.n12 VPWR.t3 26.8503
R39 VPWR.n14 VPWR.t1 26.3844
R40 VPWR.n14 VPWR.t2 26.3844
R41 VPWR.n22 VPWR.n10 25.5955
R42 VPWR.n16 VPWR.n15 25.224
R43 VPWR.n34 VPWR.n33 24.4711
R44 VPWR.n33 VPWR.n32 22.9652
R45 VPWR.n28 VPWR.n6 19.9534
R46 VPWR.n40 VPWR.n39 19.2005
R47 VPWR.n17 VPWR.n16 17.6946
R48 VPWR.n38 VPWR.n2 15.8123
R49 VPWR.n16 VPWR.n11 9.3005
R50 VPWR.n18 VPWR.n17 9.3005
R51 VPWR.n19 VPWR.n10 9.3005
R52 VPWR.n22 VPWR.n21 9.3005
R53 VPWR.n20 VPWR.n8 9.3005
R54 VPWR.n27 VPWR.n7 9.3005
R55 VPWR.n29 VPWR.n28 9.3005
R56 VPWR.n30 VPWR.n6 9.3005
R57 VPWR.n32 VPWR.n31 9.3005
R58 VPWR.n33 VPWR.n3 9.3005
R59 VPWR.n35 VPWR.n34 9.3005
R60 VPWR.n36 VPWR.n2 9.3005
R61 VPWR.n38 VPWR.n37 9.3005
R62 VPWR.n39 VPWR.n0 9.3005
R63 VPWR.n41 VPWR.n40 7.43488
R64 VPWR.n15 VPWR.n13 6.50549
R65 VPWR.n23 VPWR.n22 4.94983
R66 VPWR.n26 VPWR.n8 4.43783
R67 VPWR.n27 VPWR.n26 1.0245
R68 VPWR.n13 VPWR.n11 0.686474
R69 VPWR.n23 VPWR.n8 0.5125
R70 VPWR VPWR.n41 0.160103
R71 VPWR.n41 VPWR.n0 0.1477
R72 VPWR.n18 VPWR.n11 0.122949
R73 VPWR.n19 VPWR.n18 0.122949
R74 VPWR.n21 VPWR.n19 0.122949
R75 VPWR.n21 VPWR.n20 0.122949
R76 VPWR.n20 VPWR.n7 0.122949
R77 VPWR.n29 VPWR.n7 0.122949
R78 VPWR.n30 VPWR.n29 0.122949
R79 VPWR.n31 VPWR.n30 0.122949
R80 VPWR.n31 VPWR.n3 0.122949
R81 VPWR.n35 VPWR.n3 0.122949
R82 VPWR.n36 VPWR.n35 0.122949
R83 VPWR.n37 VPWR.n36 0.122949
R84 VPWR.n37 VPWR.n0 0.122949
R85 VPB.n0 VPB 3049.19
R86 VPB VPB.n1 928.409
R87 VPB.t4 VPB.n0 601.847
R88 VPB.n1 VPB.t12 339.651
R89 VPB.t10 VPB.t13 334.659
R90 VPB.n1 VPB.t10 304.973
R91 VPB.t8 VPB.t5 296.875
R92 VPB.t12 VPB.t11 280.914
R93 VPB.t6 VPB.t3 273.253
R94 VPB.t9 VPB.t8 259.091
R95 VPB.t7 VPB.t6 257.93
R96 VPB.t11 VPB 257.93
R97 VPB.t13 VPB.t9 253.694
R98 VPB.t5 VPB.t4 242.899
R99 VPB.t1 VPB.t0 229.839
R100 VPB.t2 VPB.t1 229.839
R101 VPB.t3 VPB.t2 229.839
R102 VPB.n0 VPB.t7 130.243
R103 a_200_74.t5 a_200_74.t0 1042.52
R104 a_200_74.t1 a_200_74.n2 572.039
R105 a_200_74.n0 a_200_74.t2 207.529
R106 a_200_74.n2 a_200_74.t3 207.529
R107 a_200_74.n0 a_200_74.t5 130.542
R108 a_200_74.n1 a_200_74.t4 128.534
R109 a_200_74.n1 a_200_74.n0 55.5644
R110 a_200_74.n2 a_200_74.n1 27.4477
R111 a_472_388.n18 a_472_388.n17 299.649
R112 a_472_388.n8 a_472_388.t10 236.654
R113 a_472_388.n9 a_472_388.t11 234.841
R114 a_472_388.n1 a_472_388.t12 234.841
R115 a_472_388.n14 a_472_388.t13 234.841
R116 a_472_388.n4 a_472_388.n2 218.196
R117 a_472_388.n22 a_472_388.n21 218.196
R118 a_472_388.n4 a_472_388.n3 208.758
R119 a_472_388.n20 a_472_388.n19 204.427
R120 a_472_388.n14 a_472_388.t14 200.195
R121 a_472_388.n8 a_472_388.n7 187.834
R122 a_472_388.n13 a_472_388.n5 186.374
R123 a_472_388.n6 a_472_388.t15 186.374
R124 a_472_388.n11 a_472_388.n10 165.189
R125 a_472_388.n16 a_472_388.n15 152
R126 a_472_388.n1 a_472_388.n0 152
R127 a_472_388.n12 a_472_388.n11 152
R128 a_472_388.n20 a_472_388.n18 115.954
R129 a_472_388.n18 a_472_388.n16 68.0276
R130 a_472_388.n21 a_472_388.n20 64.2173
R131 a_472_388.n21 a_472_388.n4 53.0829
R132 a_472_388.n1 a_472_388.n12 49.6611
R133 a_472_388.n2 a_472_388.t7 46.2955
R134 a_472_388.n2 a_472_388.t6 46.2955
R135 a_472_388.n17 a_472_388.t3 41.2931
R136 a_472_388.t5 a_472_388.n22 35.4605
R137 a_472_388.n15 a_472_388.n13 35.055
R138 a_472_388.n10 a_472_388.n9 34.3247
R139 a_472_388.n17 a_472_388.t2 31.2572
R140 a_472_388.n10 a_472_388.n8 30.6732
R141 a_472_388.n19 a_472_388.t0 29.5505
R142 a_472_388.n19 a_472_388.t1 29.5505
R143 a_472_388.n22 a_472_388.t4 29.5505
R144 a_472_388.n3 a_472_388.t8 26.2505
R145 a_472_388.n3 a_472_388.t9 26.2505
R146 a_472_388.n15 a_472_388.n14 16.7975
R147 a_472_388.n13 a_472_388.n1 14.6066
R148 a_472_388.n11 a_472_388.n0 13.1884
R149 a_472_388.n16 a_472_388.n0 13.1884
R150 a_472_388.n12 a_472_388.n6 13.146
R151 a_472_388.n9 a_472_388.n6 2.19141
R152 X.n2 X.n1 585
R153 X.n3 X.t4 263.75
R154 X.n2 X.n0 241.315
R155 X.n3 X.t5 204.832
R156 X.n0 X.t1 26.3844
R157 X.n0 X.t0 26.3844
R158 X.n1 X.t3 26.3844
R159 X.n1 X.t2 26.3844
R160 X X.n2 15.7096
R161 X X.n3 13.1373
R162 a_412_140.n0 a_412_140.t0 328.262
R163 a_412_140.n0 a_412_140.t3 314.454
R164 a_412_140.n1 a_412_140.n0 185
R165 a_412_140.n1 a_412_140.t1 26.2505
R166 a_412_140.t2 a_412_140.n1 26.2505
R167 a_685_140.n1 a_685_140.n0 474.342
R168 a_685_140.n0 a_685_140.t3 26.2505
R169 a_685_140.n0 a_685_140.t2 26.2505
R170 a_685_140.n1 a_685_140.t0 26.2505
R171 a_685_140.t1 a_685_140.n1 26.2505
R172 VNB.n0 VNB 13789
R173 VNB VNB.n1 3774.56
R174 VNB.t2 VNB.t6 2326.18
R175 VNB.t9 VNB.t8 2217.32
R176 VNB.n1 VNB.t0 1836.22
R177 VNB.n1 VNB.t5 1689.78
R178 VNB.n0 VNB.t1 1662.99
R179 VNB.t7 VNB.n0 1536.16
R180 VNB.t1 VNB.t9 1154.86
R181 VNB.t10 VNB 1143.31
R182 VNB.t0 VNB.t10 993.177
R183 VNB.t6 VNB.t7 943.641
R184 VNB.t3 VNB.t2 943.641
R185 VNB.t4 VNB.t3 943.641
R186 VNB.t5 VNB.t4 943.641
R187 C.n2 C.t1 271.065
R188 C.n3 C.t0 207.529
R189 C.n1 C.n0 181.213
R190 C C.n4 163.831
R191 C.n2 C.t2 142.994
R192 C.n1 C.t3 142.994
R193 C.n4 C.n3 40.1672
R194 C.n4 C.n1 20.449
R195 C.n0 C 17.2611
R196 C.n3 C.n2 2.19141
R197 C C.n0 1.35808
R198 A_N.n0 A_N.t1 260.611
R199 A_N.n0 A_N.t0 229.281
R200 A_N A_N.n0 154.133
R201 D.n1 D.t1 239.418
R202 D.n3 D.t0 210.45
R203 D.n1 D.n0 179.947
R204 D.n2 D.t2 179.947
R205 D D.n3 161.377
R206 D.n2 D.n1 62.8066
R207 D.n3 D.n2 2.92171
R208 VGND.n6 VGND.t2 243.202
R209 VGND.n8 VGND.n7 119.629
R210 VGND.n28 VGND.n27 114.885
R211 VGND.n14 VGND.n13 36.1417
R212 VGND.n15 VGND.n14 36.1417
R213 VGND.n15 VGND.n3 36.1417
R214 VGND.n19 VGND.n3 36.1417
R215 VGND.n20 VGND.n19 36.1417
R216 VGND.n21 VGND.n20 36.1417
R217 VGND.n21 VGND.n1 36.1417
R218 VGND.n25 VGND.n1 36.1417
R219 VGND.n26 VGND.n25 36.1417
R220 VGND.n7 VGND.t3 35.7861
R221 VGND.n13 VGND.n5 27.1064
R222 VGND.n9 VGND.n5 26.3534
R223 VGND.n7 VGND.t1 26.2505
R224 VGND.n27 VGND.t0 26.2505
R225 VGND.n27 VGND.t4 26.2505
R226 VGND.n28 VGND.n26 24.4711
R227 VGND.n9 VGND.n8 19.577
R228 VGND.n26 VGND.n0 9.3005
R229 VGND.n25 VGND.n24 9.3005
R230 VGND.n23 VGND.n1 9.3005
R231 VGND.n22 VGND.n21 9.3005
R232 VGND.n20 VGND.n2 9.3005
R233 VGND.n19 VGND.n18 9.3005
R234 VGND.n17 VGND.n3 9.3005
R235 VGND.n16 VGND.n15 9.3005
R236 VGND.n14 VGND.n4 9.3005
R237 VGND.n13 VGND.n12 9.3005
R238 VGND.n11 VGND.n5 9.3005
R239 VGND.n10 VGND.n9 9.3005
R240 VGND.n29 VGND.n28 7.19894
R241 VGND.n8 VGND.n6 6.96194
R242 VGND.n10 VGND.n6 0.513528
R243 VGND VGND.n29 0.156997
R244 VGND.n29 VGND.n0 0.150766
R245 VGND.n11 VGND.n10 0.122949
R246 VGND.n12 VGND.n11 0.122949
R247 VGND.n12 VGND.n4 0.122949
R248 VGND.n16 VGND.n4 0.122949
R249 VGND.n17 VGND.n16 0.122949
R250 VGND.n18 VGND.n17 0.122949
R251 VGND.n18 VGND.n2 0.122949
R252 VGND.n22 VGND.n2 0.122949
R253 VGND.n23 VGND.n22 0.122949
R254 VGND.n24 VGND.n23 0.122949
R255 VGND.n24 VGND.n0 0.122949
C0 VPB D 0.091083f
C1 a_882_137# VGND 0.183499f
C2 A_N VPWR 0.019732f
C3 VPB X 0.013752f
C4 A_N C 6.37e-20
C5 VPWR C 0.048037f
C6 VPB VGND 0.014943f
C7 A_N D 6.63e-19
C8 B_N VGND 0.018798f
C9 A_N X 3.52e-20
C10 VPWR D 0.038903f
C11 a_882_137# VPB 3.96e-19
C12 VPWR X 0.238965f
C13 A_N VGND 0.018587f
C14 C D 0.046659f
C15 VPWR VGND 0.149266f
C16 C X 9.61e-20
C17 a_882_137# A_N 1.83e-19
C18 C VGND 0.016723f
C19 D X 0.001869f
C20 VPB B_N 0.049238f
C21 a_882_137# VPWR 0.003441f
C22 D VGND 0.046712f
C23 a_882_137# C 0.115907f
C24 VPB A_N 0.057801f
C25 X VGND 0.259552f
C26 a_882_137# D 0.045293f
C27 VPB VPWR 0.261254f
C28 B_N A_N 0.096618f
C29 a_882_137# X 0.002003f
C30 B_N VPWR 0.018579f
C31 VPB C 0.104361f
C32 VGND VNB 1.08958f
C33 X VNB 0.078924f
C34 D VNB 0.223121f
C35 C VNB 0.265739f
C36 VPWR VNB 0.830956f
C37 A_N VNB 0.136509f
C38 B_N VNB 0.160472f
C39 VPB VNB 2.0694f
C40 a_882_137# VNB 0.030059f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4bb_2 VNB VPB VPWR VGND X B_N A_N D C
X0 VPWR.t5 D.t0 a_225_82.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3284 pd=1.745 as=0.15 ps=1.3 w=1 l=0.15
X1 a_390_82.t0 a_354_252.t2 a_312_82.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0888 ps=0.98 w=0.74 l=0.15
X2 a_225_82.t3 C.t0 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.255 ps=1.51 w=1 l=0.15
X3 X.t3 a_225_82.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2553 ps=1.43 w=0.74 l=0.15
X4 VPWR.t7 A_N.t0 a_27_74.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.42 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 VGND.t4 A_N.t1 a_27_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X6 a_225_82.t1 a_27_74.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.285 pd=1.57 as=0.2 ps=1.42 w=1 l=0.15
X7 a_354_252.t1 B_N.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2604 pd=2.3 as=0.203 ps=1.505 w=0.84 l=0.15
X8 VPWR.t1 a_225_82.t6 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_498_82.t0 C.t1 a_390_82.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.1443 ps=1.13 w=0.74 l=0.15
X10 X.t0 a_225_82.t7 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3284 ps=1.745 w=1.12 l=0.15
X11 a_354_252.t0 B_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.189025 ps=1.41 w=0.55 l=0.15
X12 a_312_82.t1 a_27_74.t3 a_225_82.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X13 VGND.t3 D.t1 a_498_82.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=1.43 as=0.1332 ps=1.1 w=0.74 l=0.15
X14 VPWR.t0 a_354_252.t3 a_225_82.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.255 pd=1.51 as=0.285 ps=1.57 w=1 l=0.15
X15 VGND.t2 a_225_82.t8 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.189025 pd=1.41 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 D.n0 D.t0 240.554
R1 D.n0 D.t1 225.291
R2 D D.n0 153.957
R3 a_225_82.n3 a_225_82.n0 238.093
R4 a_225_82.n1 a_225_82.t6 233.868
R5 a_225_82.n0 a_225_82.t7 229.487
R6 a_225_82.n4 a_225_82.t4 208.648
R7 a_225_82.n3 a_225_82.n2 205.487
R8 a_225_82.n5 a_225_82.n4 205.202
R9 a_225_82.n0 a_225_82.t5 179.947
R10 a_225_82.n1 a_225_82.t8 179.947
R11 a_225_82.n5 a_225_82.t1 68.9505
R12 a_225_82.n4 a_225_82.n3 64.0005
R13 a_225_82.n0 a_225_82.n1 62.8066
R14 a_225_82.t0 a_225_82.n5 43.3405
R15 a_225_82.n2 a_225_82.t2 29.5505
R16 a_225_82.n2 a_225_82.t3 29.5505
R17 VPWR.n7 VPWR.n6 353.276
R18 VPWR.n16 VPWR.n1 319.238
R19 VPWR.n3 VPWR.n2 316.353
R20 VPWR.n8 VPWR.n5 315.812
R21 VPWR.n5 VPWR.t2 63.9957
R22 VPWR.n1 VPWR.t7 63.3219
R23 VPWR.n5 VPWR.t5 57.1305
R24 VPWR.n6 VPWR.t4 55.6717
R25 VPWR.n2 VPWR.t0 52.2055
R26 VPWR.n2 VPWR.t6 48.2655
R27 VPWR.n15 VPWR.n14 36.1417
R28 VPWR.n10 VPWR.n9 36.1417
R29 VPWR.n1 VPWR.t3 30.4598
R30 VPWR.n6 VPWR.t1 29.3881
R31 VPWR.n14 VPWR.n3 28.9887
R32 VPWR.n10 VPWR.n3 18.4476
R33 VPWR.n8 VPWR.n7 12.5764
R34 VPWR.n17 VPWR.n16 12.2214
R35 VPWR.n9 VPWR.n4 9.3005
R36 VPWR.n11 VPWR.n10 9.3005
R37 VPWR.n12 VPWR.n3 9.3005
R38 VPWR.n14 VPWR.n13 9.3005
R39 VPWR.n15 VPWR.n0 9.3005
R40 VPWR.n16 VPWR.n15 6.77697
R41 VPWR.n9 VPWR.n8 6.02403
R42 VPWR.n7 VPWR.n4 0.474878
R43 VPWR VPWR.n17 0.163644
R44 VPWR.n17 VPWR.n0 0.144205
R45 VPWR.n11 VPWR.n4 0.122949
R46 VPWR.n12 VPWR.n11 0.122949
R47 VPWR.n13 VPWR.n12 0.122949
R48 VPWR.n13 VPWR.n0 0.122949
R49 VPB.t5 VPB.t1 395.834
R50 VPB.t3 VPB.t0 367.743
R51 VPB.t0 VPB.t6 337.098
R52 VPB VPB.t7 306.452
R53 VPB.t7 VPB.t3 291.13
R54 VPB.t2 VPB.t4 273.253
R55 VPB.t1 VPB.t2 229.839
R56 VPB.t6 VPB.t5 229.839
R57 a_354_252.t1 a_354_252.n1 494.014
R58 a_354_252.n1 a_354_252.n0 360.954
R59 a_354_252.n0 a_354_252.t3 287.861
R60 a_354_252.n1 a_354_252.t0 249.446
R61 a_354_252.n0 a_354_252.t2 178.34
R62 a_312_82.t0 a_312_82.t1 38.9194
R63 a_390_82.t0 a_390_82.t1 63.2437
R64 VNB.t6 VNB.t7 2286.61
R65 VNB.t5 VNB.t2 1940.16
R66 VNB.t1 VNB.t0 1362.73
R67 VNB.t3 VNB.t4 1247.24
R68 VNB.t4 VNB.t5 1177.95
R69 VNB VNB.t6 1143.31
R70 VNB.t2 VNB.t1 993.177
R71 VNB.t7 VNB.t3 900.788
R72 C.n0 C.t0 245.018
R73 C.n0 C.t1 229.754
R74 C C.n0 154.845
R75 VGND.n3 VGND.n2 252.788
R76 VGND.n12 VGND.t4 240.565
R77 VGND.n5 VGND.n4 210.794
R78 VGND.n4 VGND.t1 89.1897
R79 VGND.n2 VGND.t0 56.7278
R80 VGND.n6 VGND.n1 36.1417
R81 VGND.n10 VGND.n1 36.1417
R82 VGND.n11 VGND.n10 36.1417
R83 VGND.n2 VGND.t2 29.1897
R84 VGND.n6 VGND.n5 25.224
R85 VGND.n12 VGND.n11 24.4711
R86 VGND.n4 VGND.t3 22.7032
R87 VGND.n7 VGND.n6 9.3005
R88 VGND.n8 VGND.n1 9.3005
R89 VGND.n10 VGND.n9 9.3005
R90 VGND.n11 VGND.n0 9.3005
R91 VGND.n13 VGND.n12 7.19894
R92 VGND.n5 VGND.n3 6.97701
R93 VGND.n7 VGND.n3 0.246479
R94 VGND VGND.n13 0.156997
R95 VGND.n13 VGND.n0 0.150766
R96 VGND.n8 VGND.n7 0.122949
R97 VGND.n9 VGND.n8 0.122949
R98 VGND.n9 VGND.n0 0.122949
R99 X.n2 X 589.444
R100 X.n2 X.n0 585
R101 X.n3 X.n2 585
R102 X X.n1 244.917
R103 X.n2 X.t1 26.3844
R104 X.n2 X.t0 26.3844
R105 X.n1 X.t2 22.7032
R106 X.n1 X.t3 22.7032
R107 X X.n3 11.2005
R108 X X.n0 9.95606
R109 X X.n0 3.2005
R110 X.n3 X 1.95606
R111 A_N.n0 A_N.t1 276.748
R112 A_N.n0 A_N.t0 207.809
R113 A_N A_N.n0 160.922
R114 a_27_74.t0 a_27_74.n1 439.56
R115 a_27_74.n1 a_27_74.t1 289.007
R116 a_27_74.n0 a_27_74.t2 266.44
R117 a_27_74.n0 a_27_74.t3 265.392
R118 a_27_74.n1 a_27_74.n0 152
R119 B_N.n0 B_N.t0 222.32
R120 B_N B_N.n0 160.339
R121 B_N.n0 B_N.t1 140.112
R122 a_498_82.t0 a_498_82.t1 58.3789
C0 A_N B_N 2e-20
C1 VPWR X 0.162213f
C2 D VGND 0.017483f
C3 A_N VGND 0.019449f
C4 VPWR B_N 0.014526f
C5 VPWR VGND 0.088533f
C6 X B_N 0.001236f
C7 VPB C 0.04368f
C8 X VGND 0.008758f
C9 VPB D 0.049968f
C10 B_N VGND 0.007255f
C11 C D 0.094082f
C12 VPB A_N 0.061811f
C13 VPB VPWR 0.159173f
C14 VPB X 0.004527f
C15 C VPWR 0.017099f
C16 D VPWR 0.017101f
C17 VPB B_N 0.046192f
C18 C X 1.56e-19
C19 VPB VGND 0.011803f
C20 D X 0.001042f
C21 A_N VPWR 0.01566f
C22 A_N X 9.65e-20
C23 C VGND 0.012605f
C24 VGND VNB 0.670229f
C25 B_N VNB 0.171022f
C26 X VNB 0.00634f
C27 VPWR VNB 0.524175f
C28 A_N VNB 0.189991f
C29 D VNB 0.11295f
C30 C VNB 0.101649f
C31 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4bb_1 VNB VPB VPWR VGND D B_N X C A_N
X0 a_179_48.t1 C.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X1 VPWR.t2 A_N.t0 a_27_74.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 a_503_48.t0 B_N.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1764 ps=1.26 w=0.84 l=0.15
X3 a_647_74.t1 C.t1 a_533_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1152 pd=1 as=0.1344 ps=1.06 w=0.64 l=0.15
X4 VGND.t2 A_N.t1 a_27_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.113125 pd=1.065 as=0.15675 ps=1.67 w=0.55 l=0.15
X5 a_533_74.t1 a_503_48.t2 a_455_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
X6 X.t1 a_179_48.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.113125 ps=1.065 w=0.74 l=0.15
X7 VPWR.t4 a_503_48.t3 a_179_48.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.147 ps=1.19 w=0.84 l=0.15
X8 X.t0 a_179_48.t6 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.4816 pd=3.1 as=0.203 ps=1.505 w=1.12 l=0.15
X9 VGND.t0 D.t0 a_647_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.151825 pd=1.125 as=0.1152 ps=1 w=0.64 l=0.15
X10 a_179_48.t3 a_27_74.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.2478 ps=2.27 w=0.84 l=0.15
X11 a_455_74.t0 a_27_74.t3 a_179_48.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X12 a_503_48.t1 B_N.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.151825 ps=1.125 w=0.55 l=0.15
X13 VPWR.t1 D.t1 a_179_48.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.26 as=0.126 ps=1.14 w=0.84 l=0.15
R0 C.n0 C.t0 253.881
R1 C.n0 C.t1 206.525
R2 C C.n0 68.5511
R3 VPWR.n2 VPWR.t6 766.605
R4 VPWR.n14 VPWR.n1 673.114
R5 VPWR.n5 VPWR.n4 322.065
R6 VPWR.n7 VPWR.n6 315.341
R7 VPWR.n1 VPWR.t2 55.1136
R8 VPWR.n4 VPWR.t1 51.5957
R9 VPWR.n6 VPWR.t3 46.9053
R10 VPWR.n6 VPWR.t4 46.9053
R11 VPWR.n4 VPWR.t5 46.9053
R12 VPWR.n13 VPWR.n12 36.1417
R13 VPWR.n9 VPWR.n8 36.1417
R14 VPWR.n1 VPWR.t0 29.6087
R15 VPWR.n14 VPWR.n13 16.5652
R16 VPWR.n8 VPWR.n7 11.6711
R17 VPWR.n8 VPWR.n3 9.3005
R18 VPWR.n10 VPWR.n9 9.3005
R19 VPWR.n12 VPWR.n11 9.3005
R20 VPWR.n13 VPWR.n0 9.3005
R21 VPWR.n12 VPWR.n2 8.65932
R22 VPWR.n15 VPWR.n14 7.53404
R23 VPWR.n7 VPWR.n5 7.22544
R24 VPWR.n9 VPWR.n2 2.63579
R25 VPWR.n5 VPWR.n3 0.531941
R26 VPWR VPWR.n15 0.161409
R27 VPWR.n15 VPWR.n0 0.146411
R28 VPWR.n10 VPWR.n3 0.122949
R29 VPWR.n11 VPWR.n10 0.122949
R30 VPWR.n11 VPWR.n0 0.122949
R31 a_179_48.n4 a_179_48.n3 366.428
R32 a_179_48.n3 a_179_48.n0 300.26
R33 a_179_48.n2 a_179_48.n1 250.069
R34 a_179_48.n1 a_179_48.t6 240.197
R35 a_179_48.n1 a_179_48.t5 192.792
R36 a_179_48.n2 a_179_48.t4 133.108
R37 a_179_48.n3 a_179_48.n2 89.2673
R38 a_179_48.n0 a_179_48.t3 46.9053
R39 a_179_48.n0 a_179_48.t2 35.1791
R40 a_179_48.t0 a_179_48.n4 35.1791
R41 a_179_48.n4 a_179_48.t1 35.1791
R42 VPB.t0 VPB.t6 584.812
R43 VPB.t1 VPB.t5 291.13
R44 VPB.t4 VPB.t3 280.914
R45 VPB.t2 VPB.t0 273.253
R46 VPB VPB.t2 257.93
R47 VPB.t6 VPB.t4 255.376
R48 VPB.t3 VPB.t1 229.839
R49 A_N.n0 A_N.t1 226.704
R50 A_N.n0 A_N.t0 211.441
R51 A_N A_N.n0 155.067
R52 a_27_74.t0 a_27_74.n1 327.072
R53 a_27_74.n1 a_27_74.t1 325.928
R54 a_27_74.n0 a_27_74.t3 223.178
R55 a_27_74.n0 a_27_74.t2 210.727
R56 a_27_74.n1 a_27_74.n0 183.476
R57 B_N.n0 B_N.t0 285.193
R58 B_N.n0 B_N.t1 196.56
R59 B_N B_N.n0 156.99
R60 a_503_48.t0 a_503_48.n1 480.575
R61 a_503_48.n0 a_503_48.t3 273.94
R62 a_503_48.n1 a_503_48.t1 238.43
R63 a_503_48.n0 a_503_48.t2 182.75
R64 a_503_48.n1 a_503_48.n0 181.833
R65 a_533_74.t0 a_533_74.t1 78.7505
R66 a_647_74.t0 a_647_74.t1 67.5005
R67 VNB.t2 VNB.t1 2840.95
R68 VNB.t0 VNB.t4 1466.67
R69 VNB.t6 VNB.t5 1316.54
R70 VNB.t5 VNB.t0 1177.95
R71 VNB VNB.t3 1143.31
R72 VNB.t3 VNB.t2 1097.11
R73 VNB.t1 VNB.t6 900.788
R74 VGND.n2 VGND.n1 215.097
R75 VGND.n2 VGND.n0 208.353
R76 VGND.n0 VGND.t3 61.7473
R77 VGND.n1 VGND.t1 33.8208
R78 VGND.n1 VGND.t2 30.546
R79 VGND.n0 VGND.t0 26.2181
R80 VGND VGND.n2 0.189802
R81 a_455_74.t0 a_455_74.t1 45.0005
R82 X X.t0 783.467
R83 X X.t1 224.583
R84 D.n0 D.t1 253.899
R85 D.n0 D.t0 206.477
R86 D D.n0 68.1655
C0 B_N VPWR 0.019316f
C1 VGND VPWR 0.077619f
C2 X A_N 0.002022f
C3 VGND A_N 0.017316f
C4 VPWR A_N 0.008859f
C5 VPB C 0.051209f
C6 VPB D 0.052185f
C7 X VPB 0.006246f
C8 C D 0.144841f
C9 VPB B_N 0.068034f
C10 VGND VPB 0.012367f
C11 VPB VPWR 0.149529f
C12 VGND C 0.010118f
C13 C VPWR 0.01726f
C14 D B_N 0.065761f
C15 VPB A_N 0.049117f
C16 X B_N 1.51e-20
C17 VGND D 0.015253f
C18 X VGND 0.066115f
C19 D VPWR 0.026946f
C20 VGND B_N 0.013217f
C21 X VPWR 0.021092f
C22 VGND VNB 0.60703f
C23 X VNB 0.01241f
C24 A_N VNB 0.192876f
C25 VPWR VNB 0.478689f
C26 B_N VNB 0.19314f
C27 D VNB 0.116874f
C28 C VNB 0.111229f
C29 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4b_4 VNB VPB VPWR VGND A_N D C B X
X0 VGND.t6 D.t0 a_751_125.t3 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.174875 pd=1.315 as=0.104 ps=0.965 w=0.64 l=0.15
X1 VPWR.t1 A_N.t0 a_27_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2354 pd=1.55 as=0.295 ps=2.59 w=1 l=0.15
X2 a_199_294.t1 B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.16 ps=1.32 w=1 l=0.15
X3 VPWR.t3 a_199_294.t8 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X4 X.t7 a_199_294.t9 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1421 ps=1.145 w=0.74 l=0.15
X5 X.t2 a_199_294.t10 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2296 pd=1.53 as=0.1848 ps=1.45 w=1.12 l=0.15
X6 VPWR.t5 a_199_294.t11 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2159 pd=1.52 as=0.2296 ps=1.53 w=1.12 l=0.15
X7 a_751_125.t1 C.t0 a_664_125.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.178725 ps=1.85 w=0.64 l=0.15
X8 a_664_125.t2 C.t1 a_751_125.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 VGND.t1 a_199_294.t12 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1813 pd=1.23 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VGND.t2 a_199_294.t13 X.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t2 C.t2 a_199_294.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.43 ps=1.86 w=1 l=0.15
X12 X.t0 a_199_294.t14 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2354 ps=1.55 w=1.12 l=0.15
X13 a_1136_125.t1 B.t1 a_664_125.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X14 a_199_294.t2 a_27_368.t2 a_1136_125.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 a_199_294.t6 D.t1 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.43 pd=1.86 as=0.1925 ps=1.385 w=1 l=0.15
X16 VPWR.t8 D.t2 a_199_294.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1925 pd=1.385 as=0.15 ps=1.3 w=1 l=0.15
X17 a_199_294.t7 C.t3 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2159 ps=1.52 w=1 l=0.15
X18 X.t4 a_199_294.t15 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1813 ps=1.23 w=0.74 l=0.15
X19 a_199_294.t4 a_27_368.t3 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X20 a_1136_125.t2 a_27_368.t4 a_199_294.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.16 pd=1.14 as=0.0896 ps=0.92 w=0.64 l=0.15
X21 a_751_125.t2 D.t3 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.174875 ps=1.315 w=0.64 l=0.15
X22 a_664_125.t0 B.t2 a_1136_125.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1792 pd=1.84 as=0.16 ps=1.14 w=0.64 l=0.15
X23 VGND.t4 A_N.t1 a_27_368.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1421 pd=1.145 as=0.1824 ps=1.85 w=0.64 l=0.15
R0 D.n0 D.t2 346.8
R1 D.n0 D.t1 209.776
R2 D.n5 D.n4 152
R3 D.n3 D.n2 152
R4 D.n4 D.t3 147.621
R5 D.n1 D.t0 128.534
R6 D.n4 D.n3 36.0181
R7 D D.n5 14.352
R8 D.n2 D 9.69747
R9 D.n3 D.n1 9.53457
R10 D.n2 D 8.92171
R11 D.n5 D 4.26717
R12 D.n1 D.n0 2.47952
R13 a_751_125.n1 a_751_125.n0 435.272
R14 a_751_125.n0 a_751_125.t3 30.938
R15 a_751_125.n0 a_751_125.t1 30.0005
R16 a_751_125.t0 a_751_125.n1 26.2505
R17 a_751_125.n1 a_751_125.t2 26.2505
R18 VGND.n4 VGND.n3 248.887
R19 VGND.n10 VGND.n2 210.018
R20 VGND.n5 VGND.t2 154.727
R21 VGND.n13 VGND.n12 118.763
R22 VGND.n12 VGND.t0 46.0986
R23 VGND.n3 VGND.t5 41.2505
R24 VGND.n3 VGND.t6 41.2505
R25 VGND.n2 VGND.t3 40.541
R26 VGND.n2 VGND.t1 38.9194
R27 VGND.n6 VGND.n1 36.1417
R28 VGND.n11 VGND.n10 35.3887
R29 VGND.n12 VGND.t4 26.2505
R30 VGND.n13 VGND.n11 21.4593
R31 VGND.n5 VGND.n4 13.6052
R32 VGND.n10 VGND.n1 12.0476
R33 VGND.n11 VGND.n0 9.3005
R34 VGND.n10 VGND.n9 9.3005
R35 VGND.n8 VGND.n1 9.3005
R36 VGND.n7 VGND.n6 9.3005
R37 VGND.n14 VGND.n13 7.34058
R38 VGND.n6 VGND.n5 5.27109
R39 VGND.n7 VGND.n4 0.217259
R40 VGND VGND.n14 0.158861
R41 VGND.n14 VGND.n0 0.148926
R42 VGND.n8 VGND.n7 0.122949
R43 VGND.n9 VGND.n8 0.122949
R44 VGND.n9 VGND.n0 0.122949
R45 VNB.t4 VNB.t6 2517.59
R46 VNB.t9 VNB.t0 1501.31
R47 VNB.t3 VNB.t5 1478.22
R48 VNB.t12 VNB.t11 1362.73
R49 VNB.t8 VNB.t2 1281.89
R50 VNB VNB.t8 1235.7
R51 VNB.t6 VNB.t12 1097.11
R52 VNB.t10 VNB.t9 993.177
R53 VNB.t7 VNB.t10 993.177
R54 VNB.t1 VNB.t7 993.177
R55 VNB.t11 VNB.t1 993.177
R56 VNB.t5 VNB.t4 993.177
R57 VNB.t2 VNB.t3 993.177
R58 A_N.n0 A_N.t0 265.731
R59 A_N.n0 A_N.t1 161.565
R60 A_N A_N.n0 157.464
R61 a_27_368.n4 a_27_368.n3 850.918
R62 a_27_368.n4 a_27_368.t1 298.175
R63 a_27_368.t0 a_27_368.n4 221.603
R64 a_27_368.n0 a_27_368.t3 211.179
R65 a_27_368.n2 a_27_368.n1 187.585
R66 a_27_368.n2 a_27_368.t2 170.153
R67 a_27_368.n0 a_27_368.t4 168.701
R68 a_27_368.n3 a_27_368.n2 54.0495
R69 a_27_368.n3 a_27_368.n0 7.30353
R70 VPWR.n9 VPWR.t7 844.048
R71 VPWR.n17 VPWR.n7 604.976
R72 VPWR.n5 VPWR.n4 604.107
R73 VPWR.n11 VPWR.n10 603.835
R74 VPWR.n24 VPWR.n3 603.312
R75 VPWR.n26 VPWR.n1 602.58
R76 VPWR.n1 VPWR.t1 50.2355
R77 VPWR.n4 VPWR.t10 48.2655
R78 VPWR.n7 VPWR.t8 46.2955
R79 VPWR.n19 VPWR.n18 36.1417
R80 VPWR.n12 VPWR.n8 36.1417
R81 VPWR.n16 VPWR.n8 36.1417
R82 VPWR.n23 VPWR.n5 35.7652
R83 VPWR.n10 VPWR.t0 31.5205
R84 VPWR.n10 VPWR.t2 31.5205
R85 VPWR.n1 VPWR.t6 30.5869
R86 VPWR.n25 VPWR.n24 29.7417
R87 VPWR.n7 VPWR.t9 29.5505
R88 VPWR.n3 VPWR.t4 29.0228
R89 VPWR.n3 VPWR.t3 29.0228
R90 VPWR.n4 VPWR.t5 28.6759
R91 VPWR.n24 VPWR.n23 15.4358
R92 VPWR.n26 VPWR.n25 13.177
R93 VPWR.n19 VPWR.n5 10.5417
R94 VPWR.n12 VPWR.n11 10.5417
R95 VPWR.n13 VPWR.n12 9.3005
R96 VPWR.n14 VPWR.n8 9.3005
R97 VPWR.n16 VPWR.n15 9.3005
R98 VPWR.n18 VPWR.n6 9.3005
R99 VPWR.n20 VPWR.n19 9.3005
R100 VPWR.n21 VPWR.n5 9.3005
R101 VPWR.n23 VPWR.n22 9.3005
R102 VPWR.n24 VPWR.n2 9.3005
R103 VPWR.n25 VPWR.n0 9.3005
R104 VPWR.n18 VPWR.n17 9.03579
R105 VPWR.n27 VPWR.n26 7.53404
R106 VPWR.n11 VPWR.n9 6.89633
R107 VPWR.n17 VPWR.n16 2.25932
R108 VPWR.n13 VPWR.n9 0.834264
R109 VPWR VPWR.n27 0.161409
R110 VPWR.n27 VPWR.n0 0.146411
R111 VPWR.n14 VPWR.n13 0.122949
R112 VPWR.n15 VPWR.n14 0.122949
R113 VPWR.n15 VPWR.n6 0.122949
R114 VPWR.n20 VPWR.n6 0.122949
R115 VPWR.n21 VPWR.n20 0.122949
R116 VPWR.n22 VPWR.n21 0.122949
R117 VPWR.n22 VPWR.n2 0.122949
R118 VPWR.n2 VPWR.n0 0.122949
R119 VPB.t9 VPB.t2 515.861
R120 VPB.t0 VPB.t7 459.678
R121 VPB.t1 VPB.t6 296.238
R122 VPB.t4 VPB.t5 286.022
R123 VPB.t5 VPB.t10 280.914
R124 VPB.t8 VPB.t9 273.253
R125 VPB VPB.t1 257.93
R126 VPB.t3 VPB.t4 245.161
R127 VPB.t2 VPB.t0 240.054
R128 VPB.t10 VPB.t8 229.839
R129 VPB.t6 VPB.t3 229.839
R130 B.t2 B.t1 928.654
R131 B.t1 B.t0 460.579
R132 B.n1 B.n0 230.919
R133 B.n1 B.t2 192.091
R134 B B.n1 157.43
R135 a_199_294.n1 a_199_294.t4 834.814
R136 a_199_294.t1 a_199_294.n17 808.268
R137 a_199_294.n12 a_199_294.n11 585
R138 a_199_294.n14 a_199_294.n13 585
R139 a_199_294.n16 a_199_294.n15 585
R140 a_199_294.n2 a_199_294.t14 305.635
R141 a_199_294.n1 a_199_294.n0 245.55
R142 a_199_294.n6 a_199_294.t11 234.841
R143 a_199_294.n7 a_199_294.t10 234.841
R144 a_199_294.n4 a_199_294.t8 234.841
R145 a_199_294.n2 a_199_294.t9 208.968
R146 a_199_294.n6 a_199_294.t13 188.565
R147 a_199_294.n3 a_199_294.t12 186.374
R148 a_199_294.n8 a_199_294.t15 186.374
R149 a_199_294.n10 a_199_294.n9 152
R150 a_199_294.n15 a_199_294.n14 110.32
R151 a_199_294.n3 a_199_294.n2 97.715
R152 a_199_294.n10 a_199_294.n5 81.6328
R153 a_199_294.n12 a_199_294.n10 68.0998
R154 a_199_294.n13 a_199_294.n12 49.8067
R155 a_199_294.n17 a_199_294.n16 46.1994
R156 a_199_294.n5 a_199_294.n4 39.1596
R157 a_199_294.n9 a_199_294.n6 35.7853
R158 a_199_294.n15 a_199_294.t0 29.5505
R159 a_199_294.n14 a_199_294.t6 29.5505
R160 a_199_294.n11 a_199_294.t5 29.5505
R161 a_199_294.n11 a_199_294.t7 29.5505
R162 a_199_294.n16 a_199_294.n13 28.6725
R163 a_199_294.n0 a_199_294.t3 26.2505
R164 a_199_294.n0 a_199_294.t2 26.2505
R165 a_199_294.n9 a_199_294.n8 24.8308
R166 a_199_294.n7 a_199_294.n5 24.2289
R167 a_199_294.n8 a_199_294.n7 21.1793
R168 a_199_294.n17 a_199_294.n1 8.22907
R169 a_199_294.n4 a_199_294.n3 2.19141
R170 X.n3 X.n1 614.76
R171 X.n3 X.n2 585
R172 X.n7 X.n6 185
R173 X.n8 X.n7 185
R174 X.n5 X.n0 156.264
R175 X.n1 X.t1 45.7326
R176 X.n2 X.t3 26.3844
R177 X.n2 X.t0 26.3844
R178 X.n1 X.t2 26.3844
R179 X.n7 X.t6 22.7032
R180 X.n7 X.t7 22.7032
R181 X.n0 X.t5 22.7032
R182 X.n0 X.t4 22.7032
R183 X X.n4 13.357
R184 X.n8 X 10.8057
R185 X.n5 X 6.1656
R186 X.n6 X 4.15634
R187 X.n4 X.n3 3.5205
R188 X.n6 X.n5 3.32518
R189 X.n4 X 2.7205
R190 X X.n8 1.4966
R191 C.n0 C.t1 702.114
R192 C.n1 C.n0 539.841
R193 C.t1 C.t2 468.639
R194 C.n1 C.t3 263.762
R195 C.n0 C.t0 221.72
R196 C C.n1 154.522
R197 a_664_125.n0 a_664_125.t0 444.705
R198 a_664_125.n0 a_664_125.t3 380.454
R199 a_664_125.n1 a_664_125.n0 86.3508
R200 a_664_125.n1 a_664_125.t1 26.2505
R201 a_664_125.t2 a_664_125.n1 26.2505
R202 a_1136_125.n1 a_1136_125.n0 435.545
R203 a_1136_125.n0 a_1136_125.t0 46.8755
R204 a_1136_125.n0 a_1136_125.t2 46.8755
R205 a_1136_125.n1 a_1136_125.t3 26.2505
R206 a_1136_125.t1 a_1136_125.n1 26.2505
C0 B VGND 0.042289f
C1 VPWR X 0.043503f
C2 VPB A_N 0.039443f
C3 VPWR VGND 0.126951f
C4 VPB C 0.083017f
C5 X VGND 0.326669f
C6 A_N C 6.44e-19
C7 VPB D 0.124813f
C8 VPB B 0.080929f
C9 C D 0.144731f
C10 VPB VPWR 0.210991f
C11 C B 0.075327f
C12 A_N VPWR 0.014428f
C13 VPB X 0.008024f
C14 D B 0.002217f
C15 A_N X 0.027744f
C16 C VPWR 0.024239f
C17 VPB VGND 0.013857f
C18 A_N VGND 0.044423f
C19 C X 0.004822f
C20 D VPWR 0.026886f
C21 C VGND 0.118816f
C22 B VPWR 0.028723f
C23 D X 1.07e-20
C24 B X 2.81e-21
C25 D VGND 0.016559f
C26 VGND VNB 0.88959f
C27 X VNB 0.019812f
C28 VPWR VNB 0.723381f
C29 B VNB 0.409109f
C30 D VNB 0.206063f
C31 C VNB 0.558288f
C32 A_N VNB 0.143307f
C33 VPB VNB 1.79899f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4b_2 VNB VPB VPWR VGND X A_N D C B
X0 VPWR.t4 A_N.t0 a_27_112.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2086 pd=1.515 as=0.2478 ps=2.27 w=0.84 l=0.15
X1 a_186_48.t4 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.2578 ps=1.59 w=1 l=0.15
X2 VPWR.t2 a_27_112.t2 a_186_48.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.43335 pd=2.99 as=0.17 ps=1.34 w=1 l=0.15
X3 a_537_74.t1 C.t0 a_459_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0888 ps=0.98 w=0.74 l=0.15
X4 a_645_74.t1 B.t0 a_537_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X5 a_186_48.t2 a_27_112.t3 a_645_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1443 ps=1.13 w=0.74 l=0.15
X6 VGND.t1 a_186_48.t5 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.23495 pd=1.375 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 X.t3 a_186_48.t6 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.126075 ps=1.1 w=0.74 l=0.15
X8 a_459_74.t0 D.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.23495 ps=1.375 w=0.74 l=0.15
X9 a_186_48.t3 B.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.17 pd=1.34 as=0.24805 ps=1.56 w=1 l=0.15
X10 VPWR.t0 C.t1 a_186_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.24805 pd=1.56 as=0.1625 ps=1.325 w=1 l=0.15
X11 VPWR.t6 a_186_48.t7 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2578 pd=1.59 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VGND.t2 A_N.t1 a_27_112.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X13 X.t0 a_186_48.t8 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2086 ps=1.515 w=1.12 l=0.15
R0 A_N.n0 A_N.t0 212.131
R1 A_N.n0 A_N.t1 166.341
R2 A_N A_N.n0 155.601
R3 a_27_112.n1 a_27_112.n0 446.637
R4 a_27_112.t0 a_27_112.n1 326.464
R5 a_27_112.n1 a_27_112.t1 311.671
R6 a_27_112.n0 a_27_112.t2 231.629
R7 a_27_112.n0 a_27_112.t3 220.113
R8 VPWR.n7 VPWR.t2 836.747
R9 VPWR.n13 VPWR.n1 686.101
R10 VPWR.n11 VPWR.n3 605.365
R11 VPWR.n6 VPWR.n5 605.365
R12 VPWR.n1 VPWR.t4 56.2862
R13 VPWR.n3 VPWR.t1 46.2955
R14 VPWR.n5 VPWR.t5 46.2955
R15 VPWR.n5 VPWR.t0 46.2955
R16 VPWR.n3 VPWR.t6 41.0193
R17 VPWR.n10 VPWR.n4 36.1417
R18 VPWR.n12 VPWR.n11 33.5064
R19 VPWR.n1 VPWR.t3 30.268
R20 VPWR.n13 VPWR.n12 16.5652
R21 VPWR.n11 VPWR.n10 13.9299
R22 VPWR.n7 VPWR.n6 10.9855
R23 VPWR.n8 VPWR.n4 9.3005
R24 VPWR.n10 VPWR.n9 9.3005
R25 VPWR.n11 VPWR.n2 9.3005
R26 VPWR.n12 VPWR.n0 9.3005
R27 VPWR.n14 VPWR.n13 7.53404
R28 VPWR.n6 VPWR.n4 7.52991
R29 VPWR.n8 VPWR.n7 0.558158
R30 VPWR VPWR.n14 0.161409
R31 VPWR.n14 VPWR.n0 0.146411
R32 VPWR.n9 VPWR.n8 0.122949
R33 VPWR.n9 VPWR.n2 0.122949
R34 VPWR.n2 VPWR.n0 0.122949
R35 VPB.t0 VPB.t5 316.668
R36 VPB.t6 VPB.t1 316.668
R37 VPB.t4 VPB.t3 278.361
R38 VPB VPB.t4 257.93
R39 VPB.t5 VPB.t2 250.269
R40 VPB.t1 VPB.t0 242.608
R41 VPB.t3 VPB.t6 229.839
R42 D.n0 D.t0 231.629
R43 D.n0 D.t1 220.113
R44 D D.n0 154.522
R45 a_186_48.n5 a_186_48.n0 641.577
R46 a_186_48.n6 a_186_48.n5 585
R47 a_186_48.n4 a_186_48.t2 319.466
R48 a_186_48.n3 a_186_48.t7 240.197
R49 a_186_48.n1 a_186_48.t8 240.197
R50 a_186_48.n1 a_186_48.t6 187.412
R51 a_186_48.n2 a_186_48.t5 179.947
R52 a_186_48.n4 a_186_48.n3 160.764
R53 a_186_48.n5 a_186_48.n4 63.3723
R54 a_186_48.n2 a_186_48.n1 56.2338
R55 a_186_48.n0 a_186_48.t1 33.4905
R56 a_186_48.n0 a_186_48.t3 33.4905
R57 a_186_48.t0 a_186_48.n6 32.5055
R58 a_186_48.n6 a_186_48.t4 31.5205
R59 a_186_48.n3 a_186_48.n2 9.49444
R60 C.n0 C.t1 231.629
R61 C.n0 C.t0 220.113
R62 C C.n0 155.423
R63 a_459_74.t0 a_459_74.t1 38.9194
R64 a_537_74.t0 a_537_74.t1 63.2437
R65 VNB.t3 VNB.t5 1813.12
R66 VNB.t1 VNB.t0 1247.24
R67 VNB.t6 VNB.t1 1247.24
R68 VNB.t4 VNB.t2 1177.95
R69 VNB VNB.t4 1143.31
R70 VNB.t2 VNB.t3 993.177
R71 VNB.t5 VNB.t6 900.788
R72 B.n0 B.t1 231.629
R73 B.n0 B.t0 220.113
R74 B B.n0 158.102
R75 a_645_74.t0 a_645_74.t1 63.2437
R76 X X.n0 586.995
R77 X X.n1 159.344
R78 X.n0 X.t1 26.3844
R79 X.n0 X.t0 26.3844
R80 X.n1 X.t2 22.7032
R81 X.n1 X.t3 22.7032
R82 VGND.n2 VGND.n0 223.137
R83 VGND.n2 VGND.n1 96.9483
R84 VGND.n0 VGND.t2 47.6797
R85 VGND.n1 VGND.t3 47.612
R86 VGND.n1 VGND.t1 47.612
R87 VGND.n0 VGND.t0 21.551
R88 VGND VGND.n2 0.380058
C0 VGND B 0.008325f
C1 X C 2.51e-19
C2 D C 0.096059f
C3 X B 1.32e-19
C4 C B 0.083778f
C5 VPB VPWR 0.141701f
C6 VGND VPB 0.009469f
C7 VPB A_N 0.048104f
C8 VGND VPWR 0.074609f
C9 VPWR A_N 0.007625f
C10 VPB X 0.002988f
C11 VGND A_N 0.012087f
C12 VPWR X 0.0141f
C13 VPB D 0.037313f
C14 VGND X 0.114983f
C15 A_N X 0.001169f
C16 VPWR D 0.010428f
C17 VPB C 0.034694f
C18 VGND D 0.015655f
C19 VPWR C 0.010801f
C20 VPB B 0.035349f
C21 VGND C 0.009916f
C22 VPWR B 0.011438f
C23 X D 4.58e-19
C24 VGND VNB 0.549173f
C25 B VNB 0.105294f
C26 C VNB 0.10133f
C27 D VNB 0.105286f
C28 X VNB 0.006422f
C29 A_N VNB 0.173026f
C30 VPWR VNB 0.446775f
C31 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4b_1 VNB VPB VPWR VGND X A_N D C B
X0 VGND.t2 D.t0 a_526_139.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1709 ps=1.275 w=0.64 l=0.15
X1 X.t1 a_226_424.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X2 VPWR.t3 D.t1 a_226_424.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2513 pd=1.63 as=0.147 ps=1.19 w=0.84 l=0.15
X3 a_526_139.t1 C.t0 a_448_139.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1709 pd=1.275 as=0.0768 ps=0.88 w=0.64 l=0.15
X4 VGND.t0 A_N.t0 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.15675 ps=1.67 w=0.55 l=0.15
X5 a_353_124.t1 a_27_74.t2 a_226_424.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.11055 pd=1.04 as=0.1824 ps=1.85 w=0.64 l=0.15
X6 a_226_424.t2 C.t1 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.3864 ps=1.76 w=0.84 l=0.15
X7 VPWR.t4 A_N.t1 a_27_74.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X8 a_448_139.t0 B.t0 a_353_124.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.11055 ps=1.04 w=0.64 l=0.15
X9 VPWR.t1 B.t1 a_226_424.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=1.76 as=0.1596 ps=1.22 w=0.84 l=0.15
X10 a_226_424.t0 a_27_74.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1596 pd=1.22 as=0.168 ps=1.24 w=0.84 l=0.15
X11 X.t0 a_226_424.t6 VPWR.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2513 ps=1.63 w=1.12 l=0.15
R0 D.n0 D.t1 226.984
R1 D.n0 D.t0 226.18
R2 D D.n0 157.237
R3 a_526_139.n0 a_526_139.t1 85.7871
R4 a_526_139.n1 a_526_139.n0 24.0005
R5 a_526_139.n0 a_526_139.t0 21.9339
R6 VGND.n1 VGND.t0 243.446
R7 VGND.n1 VGND.n0 225.452
R8 VGND.n0 VGND.t2 41.2505
R9 VGND.n0 VGND.t1 30.2643
R10 VGND VGND.n1 0.191614
R11 VNB.t1 VNB.t4 2760.1
R12 VNB.t5 VNB.t3 1593.7
R13 VNB.t3 VNB.t2 1339.63
R14 VNB VNB.t1 1143.31
R15 VNB.t4 VNB.t0 1097.11
R16 VNB.t0 VNB.t5 900.788
R17 a_226_424.n4 a_226_424.n3 658.567
R18 a_226_424.n3 a_226_424.n0 299.289
R19 a_226_424.n1 a_226_424.t6 249.861
R20 a_226_424.n2 a_226_424.n1 233.718
R21 a_226_424.n2 a_226_424.t4 217.939
R22 a_226_424.n1 a_226_424.t5 177.292
R23 a_226_424.n3 a_226_424.n2 63.624
R24 a_226_424.n4 a_226_424.t1 50.4231
R25 a_226_424.n0 a_226_424.t2 46.9053
R26 a_226_424.t0 a_226_424.n4 38.6969
R27 a_226_424.n0 a_226_424.t3 35.1791
R28 X X.n0 589.508
R29 X.n2 X.n0 585
R30 X.n1 X.n0 585
R31 X X.t1 193.761
R32 X.n0 X.t0 26.3844
R33 X X.n1 10.9977
R34 X X.n2 9.91599
R35 X.n2 X 3.42585
R36 X.n1 X 2.34416
R37 VPWR.n5 VPWR.n2 585
R38 VPWR.n7 VPWR.n6 585
R39 VPWR.n4 VPWR.n3 323.243
R40 VPWR.n13 VPWR.n1 315.339
R41 VPWR.n6 VPWR.n5 145.405
R42 VPWR.n3 VPWR.t3 63.3219
R43 VPWR.n3 VPWR.t5 52.1063
R44 VPWR.n1 VPWR.t0 46.9053
R45 VPWR.n1 VPWR.t4 46.9053
R46 VPWR.n6 VPWR.t2 35.1791
R47 VPWR.n5 VPWR.t1 35.1791
R48 VPWR.n12 VPWR.n11 34.0155
R49 VPWR.n13 VPWR.n12 19.2005
R50 VPWR.n7 VPWR.n4 13.0286
R51 VPWR.n9 VPWR.n8 9.3005
R52 VPWR.n11 VPWR.n10 9.3005
R53 VPWR.n12 VPWR.n0 9.3005
R54 VPWR.n14 VPWR.n13 7.43488
R55 VPWR.n8 VPWR.n2 5.09141
R56 VPWR.n8 VPWR.n7 3.92777
R57 VPWR.n11 VPWR.n2 1.89141
R58 VPWR.n9 VPWR.n4 0.528998
R59 VPWR VPWR.n14 0.160103
R60 VPWR.n14 VPWR.n0 0.1477
R61 VPWR.n10 VPWR.n9 0.122949
R62 VPWR.n10 VPWR.n0 0.122949
R63 VPB VPB.t0 110.16
R64 VPB.t0 VPB.t1 28.2984
R65 C.t0 C.t1 443.142
R66 C C.t0 317.05
R67 a_448_139.t0 a_448_139.t1 45.0005
R68 A_N.n0 A_N.t1 253.928
R69 A_N.n0 A_N.t0 220.865
R70 A_N A_N.n0 67.5934
R71 a_27_74.n0 a_27_74.t2 637.847
R72 a_27_74.t1 a_27_74.n1 442.344
R73 a_27_74.n1 a_27_74.t0 306.911
R74 a_27_74.n0 a_27_74.t3 227.344
R75 a_27_74.n1 a_27_74.n0 152
R76 a_353_124.t0 a_353_124.t1 59.2478
R77 B.n0 B.t0 210.766
R78 B.n1 B.t1 203
R79 B.n0 B 152
R80 B.n2 B.n1 152
R81 B.n1 B.n0 50.3914
R82 B.n2 B 10.7712
R83 B B.n2 4.21513
C0 A_N VPWR 0.017932f
C1 VPB VGND 0.008766f
C2 B VPWR 0.023628f
C3 VPB X 0.016264f
C4 C D 0.053836f
C5 A_N VGND 0.016584f
C6 B VGND 0.006502f
C7 C VPWR 0.013876f
C8 C VGND 0.119137f
C9 B X 1.35e-19
C10 D VPWR 0.022345f
C11 D VGND 0.013467f
C12 C X 3.39e-19
C13 VPWR VGND 0.071231f
C14 D X 0.0088f
C15 VPB A_N 0.061355f
C16 VPWR X 0.107784f
C17 VPB B 0.061238f
C18 VGND X 0.078884f
C19 VPB C 0.031265f
C20 VPB D 0.049481f
C21 A_N C 0.0011f
C22 VPB VPWR 0.119974f
C23 B C 0.057031f
C24 X VNB 0.105386f
C25 VGND VNB 0.569019f
C26 VPWR VNB 0.425583f
C27 D VNB 0.115939f
C28 C VNB 0.171745f
C29 B VNB 0.146921f
C30 A_N VNB 0.201381f
C31 VPB VNB 0.98688f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4_4 VNB VPB VPWR VGND D C B A X
X0 a_116_392.t9 B.t0 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X1 a_116_392.t2 A.t0 a_119_119.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 VGND.t4 D.t0 a_463_119.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.170525 pd=1.285 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 VPWR.t10 B.t1 a_116_392.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.1575 ps=1.315 w=1 l=0.15
X4 a_116_392.t3 D.t1 VPWR.t6 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.3675 ps=1.735 w=1 l=0.15
X5 a_119_119.t3 B.t2 a_32_119.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X6 a_32_119.t1 C.t0 a_463_119.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1705 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X7 VGND.t2 a_116_392.t10 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1147 ps=1.05 w=0.74 l=0.15
X8 a_119_119.t0 A.t1 a_116_392.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 VPWR.t0 a_116_392.t11 X.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X10 X.t2 a_116_392.t12 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t2 a_116_392.t13 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X12 a_32_119.t2 B.t3 a_119_119.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X13 a_116_392.t0 A.t2 VPWR.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.315 as=0.15 ps=1.3 w=1 l=0.15
X14 X.t0 a_116_392.t14 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2209 ps=1.53 w=1.12 l=0.15
X15 VPWR.t5 A.t3 a_116_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X16 VPWR.t7 D.t2 a_116_392.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3675 pd=1.735 as=0.15 ps=1.3 w=1 l=0.15
X17 X.t5 a_116_392.t15 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.2405 ps=2.13 w=0.74 l=0.15
X18 a_116_392.t5 C.t1 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X19 a_463_119.t0 C.t2 a_32_119.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X20 VPWR.t9 C.t3 a_116_392.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2209 pd=1.53 as=0.175 ps=1.35 w=1 l=0.15
X21 X.t4 a_116_392.t16 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X22 a_463_119.t1 D.t3 VGND.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.170525 ps=1.285 w=0.64 l=0.15
R0 B.t2 B.t3 838.681
R1 B.t3 B.t1 475.43
R2 B.n0 B.t0 234.091
R3 B.n0 B.t2 193.121
R4 B B.n0 160.922
R5 VPWR.n11 VPWR.n10 325.255
R6 VPWR.n8 VPWR.n7 315.928
R7 VPWR.n23 VPWR.n2 314.962
R8 VPWR.n9 VPWR.t0 265.527
R9 VPWR.n25 VPWR.t11 256.836
R10 VPWR.n4 VPWR.n3 222.464
R11 VPWR.n17 VPWR.n6 138.477
R12 VPWR.n6 VPWR.t7 67.5347
R13 VPWR.n6 VPWR.t6 66.5494
R14 VPWR.n3 VPWR.t8 39.4005
R15 VPWR.n7 VPWR.t9 39.4005
R16 VPWR.n7 VPWR.t3 39.3707
R17 VPWR.n17 VPWR.n16 32.7534
R18 VPWR.n12 VPWR.n8 29.7417
R19 VPWR.n2 VPWR.t4 29.5505
R20 VPWR.n2 VPWR.t5 29.5505
R21 VPWR.n3 VPWR.t10 29.5505
R22 VPWR.n18 VPWR.n4 28.6123
R23 VPWR.n12 VPWR.n11 27.4829
R24 VPWR.n10 VPWR.t1 26.3844
R25 VPWR.n10 VPWR.t2 26.3844
R26 VPWR.n23 VPWR.n22 25.224
R27 VPWR.n25 VPWR.n24 24.4711
R28 VPWR.n24 VPWR.n23 22.2123
R29 VPWR.n18 VPWR.n17 21.8358
R30 VPWR.n22 VPWR.n4 18.824
R31 VPWR.n16 VPWR.n8 17.6946
R32 VPWR.n13 VPWR.n12 9.3005
R33 VPWR.n14 VPWR.n8 9.3005
R34 VPWR.n16 VPWR.n15 9.3005
R35 VPWR.n19 VPWR.n18 9.3005
R36 VPWR.n20 VPWR.n4 9.3005
R37 VPWR.n22 VPWR.n21 9.3005
R38 VPWR.n23 VPWR.n1 9.3005
R39 VPWR.n24 VPWR.n0 9.3005
R40 VPWR.n26 VPWR.n25 9.3005
R41 VPWR.n11 VPWR.n9 6.75308
R42 VPWR.n17 VPWR.n5 4.62059
R43 VPWR.n13 VPWR.n9 0.636608
R44 VPWR.n15 VPWR.n5 0.184273
R45 VPWR.n19 VPWR.n5 0.184273
R46 VPWR.n14 VPWR.n13 0.122949
R47 VPWR.n15 VPWR.n14 0.122949
R48 VPWR.n20 VPWR.n19 0.122949
R49 VPWR.n21 VPWR.n20 0.122949
R50 VPWR.n21 VPWR.n1 0.122949
R51 VPWR.n1 VPWR.n0 0.122949
R52 VPWR.n26 VPWR.n0 0.122949
R53 VPWR VPWR.n26 0.0617245
R54 a_116_392.n19 a_116_392.n18 588.311
R55 a_116_392.n18 a_116_392.n1 255.762
R56 a_116_392.n5 a_116_392.t11 243.849
R57 a_116_392.n0 a_116_392.t12 240.197
R58 a_116_392.n7 a_116_392.t13 240.197
R59 a_116_392.n10 a_116_392.t14 240.197
R60 a_116_392.n17 a_116_392.n16 205.004
R61 a_116_392.n13 a_116_392.n2 204.712
R62 a_116_392.n15 a_116_392.n14 204.427
R63 a_116_392.n10 a_116_392.t15 182.138
R64 a_116_392.n8 a_116_392.t10 179.947
R65 a_116_392.n0 a_116_392.t16 179.947
R66 a_116_392.n5 a_116_392.n4 179.947
R67 a_116_392.n6 a_116_392.n3 165.189
R68 a_116_392.n12 a_116_392.n11 152
R69 a_116_392.n9 a_116_392.n3 152
R70 a_116_392.n17 a_116_392.n15 87.0108
R71 a_116_392.n15 a_116_392.n13 79.4358
R72 a_116_392.n13 a_116_392.n12 69.1684
R73 a_116_392.n0 a_116_392.n5 62.0763
R74 a_116_392.n11 a_116_392.n9 49.6611
R75 a_116_392.n2 a_116_392.t3 39.4005
R76 a_116_392.n7 a_116_392.n6 37.246
R77 a_116_392.n18 a_116_392.n17 37.0764
R78 a_116_392.n16 a_116_392.t0 32.5055
R79 a_116_392.n16 a_116_392.t8 29.5505
R80 a_116_392.n14 a_116_392.t4 29.5505
R81 a_116_392.n14 a_116_392.t5 29.5505
R82 a_116_392.n2 a_116_392.t7 29.5505
R83 a_116_392.n19 a_116_392.t1 29.5505
R84 a_116_392.t9 a_116_392.n19 29.5505
R85 a_116_392.n6 a_116_392.n0 28.4823
R86 a_116_392.n1 a_116_392.t6 26.2505
R87 a_116_392.n1 a_116_392.t2 26.2505
R88 a_116_392.n12 a_116_392.n3 13.1884
R89 a_116_392.n11 a_116_392.n10 10.955
R90 a_116_392.n8 a_116_392.n7 8.03383
R91 a_116_392.n9 a_116_392.n8 4.38232
R92 VPB.t3 VPB.t2 452.017
R93 VPB.t9 VPB.t4 286.022
R94 VPB VPB.t11 257.93
R95 VPB.t4 VPB.t5 255.376
R96 VPB.t2 VPB.t9 255.376
R97 VPB.t10 VPB.t8 255.376
R98 VPB.t0 VPB.t10 237.5
R99 VPB.t6 VPB.t7 229.839
R100 VPB.t5 VPB.t6 229.839
R101 VPB.t8 VPB.t3 229.839
R102 VPB.t1 VPB.t0 229.839
R103 VPB.t11 VPB.t1 229.839
R104 A.n0 A.t2 216.536
R105 A.n1 A.t3 214.537
R106 A.n1 A.t0 173.375
R107 A.n0 A.t1 171.913
R108 A A.n2 156.268
R109 A.n2 A.n1 38.7066
R110 A.n2 A.n0 22.6399
R111 a_119_119.n1 a_119_119.n0 431.156
R112 a_119_119.n0 a_119_119.t2 26.2505
R113 a_119_119.n0 a_119_119.t0 26.2505
R114 a_119_119.t1 a_119_119.n1 26.2505
R115 a_119_119.n1 a_119_119.t3 26.2505
R116 VNB.t8 VNB.t3 2448.29
R117 VNB.t1 VNB.t0 1362.73
R118 VNB VNB.t10 1201.05
R119 VNB.t4 VNB.t2 1154.86
R120 VNB.t3 VNB.t4 1062.47
R121 VNB.t0 VNB.t8 993.177
R122 VNB.t5 VNB.t1 993.177
R123 VNB.t9 VNB.t5 993.177
R124 VNB.t6 VNB.t9 993.177
R125 VNB.t7 VNB.t6 993.177
R126 VNB.t10 VNB.t7 993.177
R127 D.n0 D.t1 325.531
R128 D.n1 D.t2 207.529
R129 D.n1 D.t0 166.597
R130 D D.n2 154.327
R131 D.n0 D.t3 138.173
R132 D.n2 D.n1 29.1324
R133 D.n2 D.n0 17.4796
R134 a_463_119.n1 a_463_119.n0 442.875
R135 a_463_119.n0 a_463_119.t3 26.2505
R136 a_463_119.n0 a_463_119.t1 26.2505
R137 a_463_119.n1 a_463_119.t2 26.2505
R138 a_463_119.t0 a_463_119.n1 26.2505
R139 VGND.n8 VGND.n7 230.579
R140 VGND.n3 VGND.n2 214.662
R141 VGND.n1 VGND.t1 158.242
R142 VGND.n7 VGND.t3 41.2505
R143 VGND.n7 VGND.t4 41.2505
R144 VGND.n6 VGND.n5 36.1417
R145 VGND.n8 VGND.n6 35.3887
R146 VGND.n2 VGND.t0 34.0546
R147 VGND.n2 VGND.t2 22.7032
R148 VGND.n5 VGND.n1 18.824
R149 VGND.n6 VGND.n0 9.3005
R150 VGND.n5 VGND.n4 9.3005
R151 VGND.n3 VGND.n1 6.90401
R152 VGND.n9 VGND.n8 6.28599
R153 VGND VGND.n9 0.751719
R154 VGND.n4 VGND.n3 0.587719
R155 VGND.n9 VGND.n0 0.170982
R156 VGND.n4 VGND.n0 0.122949
R157 a_32_119.n0 a_32_119.t1 365.24
R158 a_32_119.n0 a_32_119.t3 305.688
R159 a_32_119.n1 a_32_119.n0 86.3508
R160 a_32_119.n1 a_32_119.t0 26.2505
R161 a_32_119.t2 a_32_119.n1 26.2505
R162 C.n0 C.t2 678.014
R163 C.n1 C.n0 538.234
R164 C.t2 C.t1 465.058
R165 C.n1 C.t3 265.101
R166 C.n0 C.t0 212.081
R167 C C.n1 158.032
R168 X.n2 X.n0 256.541
R169 X.n2 X.n1 211.54
R170 X.n4 X.n3 153.22
R171 X.n4 X.t4 148.052
R172 X X.n2 55.7175
R173 X.n0 X.t0 35.1791
R174 X X.n4 29.889
R175 X.n3 X.t5 27.5681
R176 X.n1 X.t3 26.3844
R177 X.n1 X.t2 26.3844
R178 X.n0 X.t1 26.3844
R179 X.n3 X.t6 22.7032
C0 VPB C 0.08297f
C1 B A 0.138112f
C2 VPB D 0.112826f
C3 B C 0.07531f
C4 B D 2.38e-19
C5 VPB VPWR 0.197105f
C6 A C 6.22e-19
C7 A D 0.002393f
C8 B VPWR 0.078001f
C9 VPB X 0.013172f
C10 C D 0.149799f
C11 A VPWR 0.040124f
C12 VPB VGND 0.010483f
C13 C VPWR 0.041713f
C14 B VGND 0.041033f
C15 D VPWR 0.043915f
C16 C X 0.005062f
C17 A VGND 0.006942f
C18 C VGND 0.112895f
C19 D VGND 0.015765f
C20 VPWR X 0.412555f
C21 VPB B 0.083289f
C22 VPWR VGND 0.112554f
C23 VPB A 0.070724f
C24 X VGND 0.309709f
C25 VGND VNB 0.79707f
C26 X VNB 0.068591f
C27 VPWR VNB 0.689866f
C28 D VNB 0.196151f
C29 C VNB 0.553537f
C30 A VNB 0.157805f
C31 B VNB 0.403264f
C32 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__and4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4_2 VNB VPB VPWR VGND D C B A X
X0 a_221_74.t1 B.t0 a_143_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 VGND.t1 a_56_74.t5 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2738 pd=2.22 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_56_74.t3 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.385 ps=2.77 w=1 l=0.15
X3 VPWR.t2 a_56_74.t6 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.4536 pd=3.05 as=0.168 ps=1.42 w=1.12 l=0.15
X4 X.t2 a_56_74.t7 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2509 ps=1.59 w=1.12 l=0.15
X5 VPWR.t5 D.t0 a_56_74.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2509 pd=1.59 as=0.15 ps=1.3 w=1 l=0.15
X6 a_56_74.t0 C.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.255 ps=1.51 w=1 l=0.15
X7 a_143_74.t0 A.t1 a_56_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VGND.t2 D.t1 a_335_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 a_335_74.t0 C.t1 a_221_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X10 VPWR.t4 B.t1 a_56_74.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.255 pd=1.51 as=0.15 ps=1.3 w=1 l=0.15
X11 X.t0 a_56_74.t8 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
R0 B.n0 B.t1 298.572
R1 B.n0 B.t0 178.34
R2 B B.n0 158.222
R3 a_143_74.t0 a_143_74.t1 38.9194
R4 a_221_74.t0 a_221_74.t1 68.1086
R5 VNB VNB.t1 1478.22
R6 VNB.t5 VNB.t4 1316.54
R7 VNB.t0 VNB.t5 1316.54
R8 VNB.t2 VNB.t0 1316.54
R9 VNB.t4 VNB.t3 993.177
R10 VNB.t1 VNB.t2 900.788
R11 a_56_74.n5 a_56_74.n4 341.365
R12 a_56_74.n2 a_56_74.t7 248.231
R13 a_56_74.n4 a_56_74.t6 240.197
R14 a_56_74.n1 a_56_74.n0 212.072
R15 a_56_74.n1 a_56_74.t1 202.851
R16 a_56_74.n6 a_56_74.n5 194.877
R17 a_56_74.n2 a_56_74.t8 185.571
R18 a_56_74.n3 a_56_74.t5 177.897
R19 a_56_74.n5 a_56_74.n1 77.9755
R20 a_56_74.n3 a_56_74.n2 62.3209
R21 a_56_74.n0 a_56_74.t2 29.5505
R22 a_56_74.n0 a_56_74.t3 29.5505
R23 a_56_74.n6 a_56_74.t4 29.5505
R24 a_56_74.t0 a_56_74.n6 29.5505
R25 a_56_74.n4 a_56_74.n3 7.91068
R26 X X.n0 586.12
R27 X.n2 X.n1 185
R28 X.n0 X.t3 26.3844
R29 X.n0 X.t2 26.3844
R30 X.n1 X.t1 22.7032
R31 X.n1 X.t0 22.7032
R32 X X.n2 9.6005
R33 X.n2 X 2.2405
R34 VGND.n1 VGND.t1 150.351
R35 VGND.n1 VGND.n0 121.74
R36 VGND.n0 VGND.t0 38.1086
R37 VGND.n0 VGND.t2 30.0005
R38 VGND VGND.n1 0.978455
R39 A.n0 A.t0 253.05
R40 A A.n0 201.343
R41 A.n0 A.t1 187.412
R42 VPWR.n5 VPWR.t2 803.058
R43 VPWR.n6 VPWR.n4 605.753
R44 VPWR.n2 VPWR.n1 318.368
R45 VPWR.n13 VPWR.t0 269.639
R46 VPWR.n1 VPWR.t4 51.2205
R47 VPWR.n1 VPWR.t3 49.2505
R48 VPWR.n4 VPWR.t5 46.2955
R49 VPWR.n4 VPWR.t1 44.2957
R50 VPWR.n12 VPWR.n11 36.1417
R51 VPWR.n8 VPWR.n7 36.1417
R52 VPWR.n13 VPWR.n12 20.7064
R53 VPWR.n7 VPWR.n6 10.5417
R54 VPWR.n8 VPWR.n2 10.1652
R55 VPWR.n7 VPWR.n3 9.3005
R56 VPWR.n9 VPWR.n8 9.3005
R57 VPWR.n11 VPWR.n10 9.3005
R58 VPWR.n12 VPWR.n0 9.3005
R59 VPWR.n14 VPWR.n13 9.3005
R60 VPWR.n6 VPWR.n5 7.97372
R61 VPWR.n11 VPWR.n2 1.12991
R62 VPWR.n5 VPWR.n3 0.558158
R63 VPWR.n9 VPWR.n3 0.122949
R64 VPWR.n10 VPWR.n9 0.122949
R65 VPWR.n10 VPWR.n0 0.122949
R66 VPWR.n14 VPWR.n0 0.122949
R67 VPWR VPWR.n14 0.0617245
R68 VPB.t4 VPB.t3 337.098
R69 VPB.t5 VPB.t1 316.668
R70 VPB VPB.t0 303.899
R71 VPB.t1 VPB.t2 229.839
R72 VPB.t3 VPB.t5 229.839
R73 VPB.t0 VPB.t4 229.839
R74 D.n0 D.t0 313.738
R75 D.n0 D.t1 178.34
R76 D D.n0 158.4
R77 C.n0 C.t0 298.572
R78 C.n0 C.t1 178.34
R79 C C.n0 158.788
R80 a_335_74.t0 a_335_74.t1 68.1086
C0 A B 0.071095f
C1 VPB C 0.039584f
C2 VPB D 0.042244f
C3 VPB VPWR 0.118636f
C4 B C 0.13038f
C5 A VPWR 0.049047f
C6 VPB X 0.004598f
C7 C D 0.094802f
C8 B VPWR 0.020646f
C9 VPB VGND 0.007241f
C10 A VGND 0.011706f
C11 C VPWR 0.01632f
C12 B X 1.54e-19
C13 C X 0.00433f
C14 B VGND 0.037237f
C15 D VPWR 0.012977f
C16 D X 0.020344f
C17 C VGND 0.061851f
C18 D VGND 0.036256f
C19 VPWR X 0.01864f
C20 VPB A 0.057533f
C21 VPWR VGND 0.067078f
C22 VPB B 0.039326f
C23 X VGND 0.081655f
C24 VGND VNB 0.530772f
C25 X VNB 0.017256f
C26 VPWR VNB 0.43526f
C27 D VNB 0.111424f
C28 C VNB 0.11085f
C29 B VNB 0.10867f
C30 A VNB 0.182778f
C31 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__buf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__buf_4 VNB VPB VPWR VGND A X
X0 a_86_260.t2 A.t0 VPWR.t5 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.203 ps=1.505 w=0.84 l=0.15
X1 VPWR.t0 a_86_260.t3 X.t7 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_86_260.t0 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2664 ps=1.46 w=0.74 l=0.15
X3 X.t6 a_86_260.t4 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t2 a_86_260.t5 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VGND.t4 a_86_260.t6 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2664 pd=1.46 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 X.t3 a_86_260.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X7 X.t2 a_86_260.t8 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8 X.t4 a_86_260.t9 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X9 VGND.t1 a_86_260.t10 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VPWR.t4 A.t2 a_86_260.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.126 ps=1.14 w=0.84 l=0.15
R0 A.n0 A.t0 227.612
R1 A.n1 A.t1 217.508
R2 A.n0 A.t2 191.591
R3 A A.n1 157.507
R4 A.n1 A.n0 11.7248
R5 VPWR.n5 VPWR.t4 806.17
R6 VPWR.n8 VPWR.n2 318.089
R7 VPWR.n10 VPWR.t3 250.081
R8 VPWR.n4 VPWR.n3 233.377
R9 VPWR.n3 VPWR.t5 55.4847
R10 VPWR.n3 VPWR.t0 29.5747
R11 VPWR.n2 VPWR.t1 26.3844
R12 VPWR.n2 VPWR.t2 26.3844
R13 VPWR.n8 VPWR.n7 24.0946
R14 VPWR.n9 VPWR.n8 23.3417
R15 VPWR.n10 VPWR.n9 19.577
R16 VPWR.n7 VPWR.n4 18.824
R17 VPWR.n7 VPWR.n6 9.3005
R18 VPWR.n8 VPWR.n1 9.3005
R19 VPWR.n9 VPWR.n0 9.3005
R20 VPWR.n11 VPWR.n10 9.3005
R21 VPWR.n5 VPWR.n4 6.90183
R22 VPWR.n6 VPWR.n5 0.606651
R23 VPWR.n6 VPWR.n1 0.122949
R24 VPWR.n1 VPWR.n0 0.122949
R25 VPWR.n11 VPWR.n0 0.122949
R26 VPWR VPWR.n11 0.0617245
R27 a_86_260.n11 a_86_260.n10 677.174
R28 a_86_260.n1 a_86_260.t9 302.858
R29 a_86_260.n7 a_86_260.t3 240.197
R30 a_86_260.n5 a_86_260.t4 240.197
R31 a_86_260.n2 a_86_260.t5 240.197
R32 a_86_260.n8 a_86_260.t6 193.093
R33 a_86_260.n6 a_86_260.t8 179.947
R34 a_86_260.n1 a_86_260.t7 179.947
R35 a_86_260.n3 a_86_260.t10 179.947
R36 a_86_260.n4 a_86_260.n0 165.189
R37 a_86_260.n6 a_86_260.n0 152
R38 a_86_260.n9 a_86_260.n8 152
R39 a_86_260.n10 a_86_260.t0 147.204
R40 a_86_260.n2 a_86_260.n1 114.365
R41 a_86_260.n10 a_86_260.n9 78.0782
R42 a_86_260.n7 a_86_260.n6 44.549
R43 a_86_260.n11 a_86_260.t1 35.1791
R44 a_86_260.t2 a_86_260.n11 35.1791
R45 a_86_260.n4 a_86_260.n3 33.5944
R46 a_86_260.n5 a_86_260.n4 28.4823
R47 a_86_260.n6 a_86_260.n5 21.1793
R48 a_86_260.n9 a_86_260.n0 13.1884
R49 a_86_260.n8 a_86_260.n7 5.11262
R50 a_86_260.n3 a_86_260.n2 3.65202
R51 VPB.t5 VPB.t1 273.253
R52 VPB VPB.t2 265.591
R53 VPB.t1 VPB.t0 229.839
R54 VPB.t4 VPB.t5 229.839
R55 VPB.t3 VPB.t4 229.839
R56 VPB.t2 VPB.t3 229.839
R57 X.n2 X.n0 273.656
R58 X.n2 X.n1 218.403
R59 X.n5 X.n3 150.219
R60 X.n5 X.n4 99.7716
R61 X X.n2 45.8738
R62 X.n1 X.t5 26.3844
R63 X.n1 X.t4 26.3844
R64 X.n0 X.t7 26.3844
R65 X.n0 X.t6 26.3844
R66 X.n4 X.t1 22.7032
R67 X.n4 X.t3 22.7032
R68 X.n3 X.t0 22.7032
R69 X.n3 X.t2 22.7032
R70 X X.n5 7.87613
R71 VGND.n6 VGND.t3 245.43
R72 VGND.n4 VGND.n3 207.109
R73 VGND.n2 VGND.n1 190.769
R74 VGND.n1 VGND.t0 58.3789
R75 VGND.n1 VGND.t4 58.3789
R76 VGND.n3 VGND.t2 34.0546
R77 VGND.n3 VGND.t1 34.0546
R78 VGND.n5 VGND.n4 29.7417
R79 VGND.n6 VGND.n5 20.7064
R80 VGND.n7 VGND.n6 9.3005
R81 VGND.n5 VGND.n0 9.3005
R82 VGND.n4 VGND.n2 6.55244
R83 VGND.n2 VGND.n0 0.375476
R84 VGND.n7 VGND.n0 0.122949
R85 VGND VGND.n7 0.0617245
R86 VNB.t4 VNB.t0 2009.45
R87 VNB.t1 VNB.t2 1316.54
R88 VNB VNB.t3 1304.99
R89 VNB.t2 VNB.t4 993.177
R90 VNB.t3 VNB.t1 993.177
C0 VGND VPB 0.008477f
C1 VGND VPWR 0.070266f
C2 VGND X 0.284968f
C3 VPB VPWR 0.125485f
C4 VGND A 0.018043f
C5 VPB X 0.010946f
C6 VPB A 0.071758f
C7 VPWR X 0.398463f
C8 VPWR A 0.034577f
C9 X A 0.003282f
C10 VGND VNB 0.461471f
C11 A VNB 0.184833f
C12 X VNB 0.048717f
C13 VPWR VNB 0.411367f
C14 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__buf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__buf_8 VNB VPB VPWR VGND X A
X0 VGND.t7 a_27_74.t6 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VPWR.t7 a_27_74.t7 X.t15 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t10 A.t0 a_27_74.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 X.t14 a_27_74.t8 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 VPWR.t8 A.t1 a_27_74.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 X.t6 a_27_74.t9 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6 VGND.t8 A.t2 a_27_74.t1 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 VGND.t5 a_27_74.t10 X.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.10545 ps=1.025 w=0.74 l=0.15
X8 VPWR.t5 a_27_74.t11 X.t13 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X9 a_27_74.t2 A.t3 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X10 VGND.t4 a_27_74.t12 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t4 a_27_74.t13 X.t12 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X12 X.t11 a_27_74.t14 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VPWR.t2 a_27_74.t15 X.t10 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.168 ps=1.42 w=1.12 l=0.15
X14 X.t3 a_27_74.t16 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X15 X.t2 a_27_74.t17 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 VPWR.t9 A.t4 a_27_74.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 X.t9 a_27_74.t18 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X18 a_27_74.t4 A.t5 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 X.t1 a_27_74.t19 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 X.t8 a_27_74.t20 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
X21 VGND.t0 a_27_74.t21 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_27_74.t0 a_27_74.n32 274.788
R1 a_27_74.n6 a_27_74.t13 242.388
R2 a_27_74.n8 a_27_74.t20 240.197
R3 a_27_74.n10 a_27_74.t15 240.197
R4 a_27_74.n12 a_27_74.t18 240.197
R5 a_27_74.n17 a_27_74.t7 240.197
R6 a_27_74.n20 a_27_74.t8 240.197
R7 a_27_74.n25 a_27_74.t11 240.197
R8 a_27_74.n27 a_27_74.t14 240.197
R9 a_27_74.n1 a_27_74.t1 213.799
R10 a_27_74.n32 a_27_74.n31 205.487
R11 a_27_74.n27 a_27_74.t19 184.328
R12 a_27_74.n26 a_27_74.t6 179.947
R13 a_27_74.n3 a_27_74.t16 179.947
R14 a_27_74.n19 a_27_74.t12 179.947
R15 a_27_74.n5 a_27_74.t9 179.947
R16 a_27_74.n11 a_27_74.t21 179.947
R17 a_27_74.n7 a_27_74.t17 179.947
R18 a_27_74.n6 a_27_74.t10 179.947
R19 a_27_74.n29 a_27_74.n28 152
R20 a_27_74.n26 a_27_74.n2 152
R21 a_27_74.n24 a_27_74.n23 152
R22 a_27_74.n22 a_27_74.n21 152
R23 a_27_74.n18 a_27_74.n4 152
R24 a_27_74.n16 a_27_74.n15 152
R25 a_27_74.n14 a_27_74.n13 152
R26 a_27_74.n1 a_27_74.n0 103.65
R27 a_27_74.n14 a_27_74.n9 81.6328
R28 a_27_74.n7 a_27_74.n6 63.5369
R29 a_27_74.n28 a_27_74.n26 49.6611
R30 a_27_74.n32 a_27_74.n30 49.3181
R31 a_27_74.n30 a_27_74.n1 46.6829
R32 a_27_74.n17 a_27_74.n16 45.2793
R33 a_27_74.n9 a_27_74.n8 37.699
R34 a_27_74.n21 a_27_74.n19 36.5157
R35 a_27_74.n25 a_27_74.n24 35.055
R36 a_27_74.n13 a_27_74.n11 33.5944
R37 a_27_74.n10 a_27_74.n9 26.4198
R38 a_27_74.n31 a_27_74.t3 26.3844
R39 a_27_74.n31 a_27_74.t4 26.3844
R40 a_27_74.n24 a_27_74.n3 23.3702
R41 a_27_74.n0 a_27_74.t5 22.7032
R42 a_27_74.n0 a_27_74.t2 22.7032
R43 a_27_74.n13 a_27_74.n12 21.9096
R44 a_27_74.n16 a_27_74.n5 20.449
R45 a_27_74.n20 a_27_74.n3 14.6066
R46 a_27_74.n26 a_27_74.n25 14.6066
R47 a_27_74.n15 a_27_74.n14 13.1884
R48 a_27_74.n15 a_27_74.n4 13.1884
R49 a_27_74.n22 a_27_74.n4 13.1884
R50 a_27_74.n23 a_27_74.n22 13.1884
R51 a_27_74.n23 a_27_74.n2 13.1884
R52 a_27_74.n29 a_27_74.n2 13.1884
R53 a_27_74.n19 a_27_74.n18 13.146
R54 a_27_74.n21 a_27_74.n20 11.6853
R55 a_27_74.n11 a_27_74.n10 10.2247
R56 a_27_74.n30 a_27_74.n29 9.11565
R57 a_27_74.n28 a_27_74.n27 8.76414
R58 a_27_74.n12 a_27_74.n5 7.30353
R59 a_27_74.n18 a_27_74.n17 4.38232
R60 a_27_74.n8 a_27_74.n7 2.19141
R61 X.n15 X.n14 585
R62 X.n14 X.n0 290.945
R63 X.n3 X.n1 254.282
R64 X.n3 X.n2 207.6
R65 X.n5 X.n4 207.6
R66 X.n8 X.n6 157.781
R67 X.n8 X.n7 99.7716
R68 X.n10 X.n9 99.7716
R69 X.n12 X.n11 99.6658
R70 X.n13 X.n12 56.9431
R71 X.n10 X.n8 50.4476
R72 X.n12 X.n10 50.4476
R73 X.n5 X.n3 46.6829
R74 X.n13 X.n5 46.6829
R75 X.n1 X.t11 35.1791
R76 X.n14 X.t8 29.0228
R77 X.n14 X.t12 26.3844
R78 X.n1 X.t13 26.3844
R79 X.n2 X.t15 26.3844
R80 X.n2 X.t14 26.3844
R81 X.n4 X.t10 26.3844
R82 X.n4 X.t9 26.3844
R83 X.n11 X.t5 23.514
R84 X.n11 X.t2 22.7032
R85 X.n6 X.t7 22.7032
R86 X.n6 X.t1 22.7032
R87 X.n7 X.t4 22.7032
R88 X.n7 X.t3 22.7032
R89 X.n9 X.t0 22.7032
R90 X.n9 X.t6 22.7032
R91 X X.n15 12.8005
R92 X X.n0 8.52393
R93 X.n0 X 5.51184
R94 X X.n13 2.48408
R95 X.n15 X 1.33781
R96 VGND.n18 VGND.n2 211.183
R97 VGND.n21 VGND.n20 211.183
R98 VGND.n7 VGND.n6 209.243
R99 VGND.n11 VGND.n5 209.243
R100 VGND.n14 VGND.n13 209.243
R101 VGND.n8 VGND.t5 161.438
R102 VGND.n14 VGND.n12 36.1417
R103 VGND.n6 VGND.t2 34.0546
R104 VGND.n6 VGND.t0 34.0546
R105 VGND.n5 VGND.t6 34.0546
R106 VGND.n5 VGND.t4 34.0546
R107 VGND.n13 VGND.t3 34.0546
R108 VGND.n11 VGND.n4 33.1299
R109 VGND.n20 VGND.t9 30.0005
R110 VGND.n18 VGND.n1 28.6123
R111 VGND.n21 VGND.n19 24.4711
R112 VGND.n13 VGND.t7 22.7032
R113 VGND.n2 VGND.t1 22.7032
R114 VGND.n2 VGND.t10 22.7032
R115 VGND.n20 VGND.t8 22.7032
R116 VGND.n19 VGND.n18 18.824
R117 VGND.n7 VGND.n4 17.3181
R118 VGND.n12 VGND.n11 14.3064
R119 VGND.n14 VGND.n1 11.2946
R120 VGND.n19 VGND.n0 9.3005
R121 VGND.n18 VGND.n17 9.3005
R122 VGND.n16 VGND.n1 9.3005
R123 VGND.n15 VGND.n14 9.3005
R124 VGND.n12 VGND.n3 9.3005
R125 VGND.n11 VGND.n10 9.3005
R126 VGND.n9 VGND.n4 9.3005
R127 VGND.n22 VGND.n21 7.19894
R128 VGND.n8 VGND.n7 6.97928
R129 VGND.n9 VGND.n8 0.591052
R130 VGND VGND.n22 0.156997
R131 VGND.n22 VGND.n0 0.150766
R132 VGND.n10 VGND.n9 0.122949
R133 VGND.n10 VGND.n3 0.122949
R134 VGND.n15 VGND.n3 0.122949
R135 VGND.n16 VGND.n15 0.122949
R136 VGND.n17 VGND.n16 0.122949
R137 VGND.n17 VGND.n0 0.122949
R138 VNB.t0 VNB.t2 1316.54
R139 VNB.t4 VNB.t6 1316.54
R140 VNB.t7 VNB.t3 1154.86
R141 VNB VNB.t8 1143.31
R142 VNB.t8 VNB.t9 1097.11
R143 VNB.t2 VNB.t5 1004.72
R144 VNB.t6 VNB.t0 993.177
R145 VNB.t3 VNB.t4 993.177
R146 VNB.t1 VNB.t7 993.177
R147 VNB.t10 VNB.t1 993.177
R148 VNB.t9 VNB.t10 993.177
R149 VPWR.n21 VPWR.n1 331.5
R150 VPWR.n5 VPWR.n4 325.255
R151 VPWR.n13 VPWR.n7 325.255
R152 VPWR.n9 VPWR.n8 325.255
R153 VPWR.n19 VPWR.n3 323.406
R154 VPWR.n10 VPWR.t4 266.057
R155 VPWR.n4 VPWR.t6 35.1791
R156 VPWR.n7 VPWR.t1 35.1791
R157 VPWR.n21 VPWR.n20 35.0123
R158 VPWR.n8 VPWR.t0 32.5407
R159 VPWR.n13 VPWR.n12 28.6123
R160 VPWR.n14 VPWR.n5 27.8593
R161 VPWR.n19 VPWR.n18 27.1064
R162 VPWR.n1 VPWR.t10 26.3844
R163 VPWR.n1 VPWR.t8 26.3844
R164 VPWR.n3 VPWR.t3 26.3844
R165 VPWR.n3 VPWR.t9 26.3844
R166 VPWR.n4 VPWR.t5 26.3844
R167 VPWR.n7 VPWR.t7 26.3844
R168 VPWR.n8 VPWR.t2 26.3844
R169 VPWR.n20 VPWR.n19 26.3534
R170 VPWR.n18 VPWR.n5 25.6005
R171 VPWR.n14 VPWR.n13 24.8476
R172 VPWR.n12 VPWR.n9 24.0946
R173 VPWR.n12 VPWR.n11 9.3005
R174 VPWR.n13 VPWR.n6 9.3005
R175 VPWR.n15 VPWR.n14 9.3005
R176 VPWR.n16 VPWR.n5 9.3005
R177 VPWR.n18 VPWR.n17 9.3005
R178 VPWR.n19 VPWR.n2 9.3005
R179 VPWR.n20 VPWR.n0 9.3005
R180 VPWR.n22 VPWR.n21 8.8332
R181 VPWR.n10 VPWR.n9 6.97636
R182 VPWR.n11 VPWR.n10 0.569174
R183 VPWR VPWR.n22 0.163644
R184 VPWR.n22 VPWR.n0 0.144205
R185 VPWR.n11 VPWR.n6 0.122949
R186 VPWR.n15 VPWR.n6 0.122949
R187 VPWR.n16 VPWR.n15 0.122949
R188 VPWR.n17 VPWR.n16 0.122949
R189 VPWR.n17 VPWR.n2 0.122949
R190 VPWR.n2 VPWR.n0 0.122949
R191 VPB VPB.t8 260.485
R192 VPB.t7 VPB.t1 255.376
R193 VPB.t5 VPB.t6 255.376
R194 VPB.t3 VPB.t5 255.376
R195 VPB.t2 VPB.t0 247.715
R196 VPB.t0 VPB.t4 237.5
R197 VPB.t1 VPB.t2 229.839
R198 VPB.t6 VPB.t7 229.839
R199 VPB.t9 VPB.t3 229.839
R200 VPB.t10 VPB.t9 229.839
R201 VPB.t8 VPB.t10 229.839
R202 A.n0 A.t4 228.268
R203 A.n3 A.t5 226.809
R204 A.n4 A.t1 226.809
R205 A.n4 A.t2 198.204
R206 A.n2 A.t3 196.013
R207 A.n0 A.t0 196.013
R208 A A.n1 156.465
R209 A.n8 A.n7 152
R210 A.n6 A.n5 152
R211 A.n7 A.n6 49.6611
R212 A.n2 A.n1 43.0884
R213 A.n1 A.n0 19.7187
R214 A.n5 A 12.8005
R215 A.n6 A.n4 10.955
R216 A.n8 A 8.63306
R217 A A.n8 5.65631
R218 A.n7 A.n3 5.11262
R219 A.n5 A 1.48887
R220 A.n3 A.n2 1.46111
C0 VPB A 0.101906f
C1 VPB VPWR 0.167621f
C2 VPB X 0.02402f
C3 A VPWR 0.047631f
C4 A X 8.64e-19
C5 VPB VGND 0.010497f
C6 A VGND 0.055075f
C7 VPWR X 0.815992f
C8 VPWR VGND 0.109066f
C9 X VGND 0.601117f
C10 VGND VNB 0.721381f
C11 X VNB 0.052843f
C12 VPWR VNB 0.585362f
C13 A VNB 0.341587f
C14 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__bufbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__bufbuf_8 VNB VPB VPWR VGND A X
X0 a_334_368.t2 a_221_368.t2 VGND.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VPWR.t11 A.t0 a_27_112.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1946 pd=1.495 as=0.2478 ps=2.27 w=0.84 l=0.15
X2 VGND.t5 a_334_368.t6 X.t15 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 X.t14 a_334_368.t7 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_221_368.t1 a_27_112.t2 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1946 ps=1.495 w=1.12 l=0.15
X5 VPWR.t1 a_334_368.t8 X.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_221_368.t0 a_27_112.t3 VGND.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.151975 ps=1.17 w=0.74 l=0.15
X7 X.t6 a_334_368.t9 VPWR.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t7 a_334_368.t10 X.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X9 VGND.t3 a_221_368.t3 a_334_368.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 VPWR.t6 a_334_368.t11 X.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X11 X.t3 a_334_368.t12 VPWR.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 X.t13 a_334_368.t13 VGND.t7 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 VPWR.t4 a_334_368.t14 X.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VGND.t8 a_334_368.t15 X.t12 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.25955 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 X.t1 a_334_368.t16 VPWR.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1708 ps=1.425 w=1.12 l=0.15
X16 X.t11 a_334_368.t17 VGND.t9 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X17 X.t0 a_334_368.t18 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X18 VGND.t10 a_334_368.t19 X.t10 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 VGND.t2 a_221_368.t4 a_334_368.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 X.t9 a_334_368.t20 VGND.t11 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X21 VPWR.t10 a_221_368.t5 a_334_368.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X22 VGND.t0 A.t1 a_27_112.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.151975 pd=1.17 as=0.15675 ps=1.67 w=0.55 l=0.15
X23 a_334_368.t4 a_221_368.t6 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 VGND.t12 a_334_368.t21 X.t8 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1258 ps=1.08 w=0.74 l=0.15
X25 VPWR.t8 a_221_368.t7 a_334_368.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 a_221_368.t1 a_221_368.n6 248.513
R1 a_221_368.n2 a_221_368.t5 242.388
R2 a_221_368.n0 a_221_368.t6 240.197
R3 a_221_368.n1 a_221_368.t7 240.197
R4 a_221_368.n3 a_221_368.t3 179.947
R5 a_221_368.n0 a_221_368.t2 179.947
R6 a_221_368.n2 a_221_368.t4 179.947
R7 a_221_368.n5 a_221_368.n4 170.654
R8 a_221_368.n6 a_221_368.t0 162.561
R9 a_221_368.n5 a_221_368.n1 85.0177
R10 a_221_368.n0 a_221_368.n2 62.8066
R11 a_221_368.n4 a_221_368.n3 44.549
R12 a_221_368.n6 a_221_368.n5 18.6929
R13 a_221_368.n4 a_221_368.n0 18.2581
R14 a_221_368.n3 a_221_368.n1 3.65202
R15 VGND.n28 VGND.n27 211.183
R16 VGND.n8 VGND.n7 206.139
R17 VGND.n13 VGND.n12 206.139
R18 VGND.n5 VGND.n4 206.139
R19 VGND.n20 VGND.n19 206.139
R20 VGND.n2 VGND.n1 206.139
R21 VGND.n9 VGND.t8 156.154
R22 VGND.n27 VGND.t0 48.0005
R23 VGND.n26 VGND.n25 36.1417
R24 VGND.n27 VGND.t1 35.7351
R25 VGND.n7 VGND.t11 34.0546
R26 VGND.n4 VGND.t10 34.0546
R27 VGND.n19 VGND.t9 34.0546
R28 VGND.n25 VGND.n2 32.7534
R29 VGND.n18 VGND.n5 28.2358
R30 VGND.n13 VGND.n11 26.7299
R31 VGND.n21 VGND.n20 25.224
R32 VGND.n7 VGND.t12 22.7032
R33 VGND.n12 VGND.t6 22.7032
R34 VGND.n12 VGND.t5 22.7032
R35 VGND.n4 VGND.t7 22.7032
R36 VGND.n19 VGND.t2 22.7032
R37 VGND.n1 VGND.t4 22.7032
R38 VGND.n1 VGND.t3 22.7032
R39 VGND.n20 VGND.n18 22.2123
R40 VGND.n14 VGND.n13 20.7064
R41 VGND.n14 VGND.n5 19.2005
R42 VGND.n28 VGND.n26 18.4476
R43 VGND.n11 VGND.n8 17.6946
R44 VGND.n21 VGND.n2 14.6829
R45 VGND.n26 VGND.n0 9.3005
R46 VGND.n25 VGND.n24 9.3005
R47 VGND.n23 VGND.n2 9.3005
R48 VGND.n22 VGND.n21 9.3005
R49 VGND.n20 VGND.n3 9.3005
R50 VGND.n18 VGND.n17 9.3005
R51 VGND.n16 VGND.n5 9.3005
R52 VGND.n15 VGND.n14 9.3005
R53 VGND.n13 VGND.n6 9.3005
R54 VGND.n11 VGND.n10 9.3005
R55 VGND.n29 VGND.n28 7.46433
R56 VGND.n9 VGND.n8 6.96039
R57 VGND.n10 VGND.n9 0.594857
R58 VGND VGND.n29 0.160491
R59 VGND.n29 VGND.n0 0.147317
R60 VGND.n10 VGND.n6 0.122949
R61 VGND.n15 VGND.n6 0.122949
R62 VGND.n16 VGND.n15 0.122949
R63 VGND.n17 VGND.n16 0.122949
R64 VGND.n17 VGND.n3 0.122949
R65 VGND.n22 VGND.n3 0.122949
R66 VGND.n23 VGND.n22 0.122949
R67 VGND.n24 VGND.n23 0.122949
R68 VGND.n24 VGND.n0 0.122949
R69 a_334_368.n28 a_334_368.t3 276.125
R70 a_334_368.n4 a_334_368.t11 241.657
R71 a_334_368.n6 a_334_368.t12 240.197
R72 a_334_368.n8 a_334_368.t14 240.197
R73 a_334_368.n3 a_334_368.t16 240.197
R74 a_334_368.n15 a_334_368.t8 240.197
R75 a_334_368.n17 a_334_368.t9 240.197
R76 a_334_368.n22 a_334_368.t10 240.197
R77 a_334_368.n24 a_334_368.t18 240.197
R78 a_334_368.n28 a_334_368.n27 206.823
R79 a_334_368.n30 a_334_368.t1 186.852
R80 a_334_368.n31 a_334_368.n30 186.125
R81 a_334_368.n24 a_334_368.t17 182.138
R82 a_334_368.n13 a_334_368.t7 179.947
R83 a_334_368.n23 a_334_368.t19 179.947
R84 a_334_368.n1 a_334_368.t13 179.947
R85 a_334_368.n16 a_334_368.t6 179.947
R86 a_334_368.n9 a_334_368.t21 179.947
R87 a_334_368.n5 a_334_368.t20 179.947
R88 a_334_368.n4 a_334_368.t15 179.947
R89 a_334_368.n11 a_334_368.n7 165.189
R90 a_334_368.n26 a_334_368.n25 152
R91 a_334_368.n23 a_334_368.n0 152
R92 a_334_368.n21 a_334_368.n20 152
R93 a_334_368.n19 a_334_368.n18 152
R94 a_334_368.n14 a_334_368.n2 152
R95 a_334_368.n13 a_334_368.n12 152
R96 a_334_368.n11 a_334_368.n10 152
R97 a_334_368.n5 a_334_368.n4 62.8066
R98 a_334_368.n14 a_334_368.n13 49.6611
R99 a_334_368.n25 a_334_368.n23 49.6611
R100 a_334_368.n7 a_334_368.n6 43.8187
R101 a_334_368.n10 a_334_368.n3 37.9763
R102 a_334_368.n22 a_334_368.n21 37.246
R103 a_334_368.n18 a_334_368.n16 36.5157
R104 a_334_368.n27 a_334_368.t5 26.3844
R105 a_334_368.n27 a_334_368.t4 26.3844
R106 a_334_368.n21 a_334_368.n1 23.3702
R107 a_334_368.n31 a_334_368.t0 22.7032
R108 a_334_368.t2 a_334_368.n31 22.7032
R109 a_334_368.n8 a_334_368.n7 21.9096
R110 a_334_368.n10 a_334_368.n9 21.9096
R111 a_334_368.n18 a_334_368.n17 21.1793
R112 a_334_368.n29 a_334_368.n28 19.5202
R113 a_334_368.n29 a_334_368.n26 15.1278
R114 a_334_368.n12 a_334_368.n11 13.1884
R115 a_334_368.n12 a_334_368.n2 13.1884
R116 a_334_368.n19 a_334_368.n2 13.1884
R117 a_334_368.n20 a_334_368.n19 13.1884
R118 a_334_368.n20 a_334_368.n0 13.1884
R119 a_334_368.n26 a_334_368.n0 13.1884
R120 a_334_368.n30 a_334_368.n29 12.9412
R121 a_334_368.n23 a_334_368.n22 12.4157
R122 a_334_368.n13 a_334_368.n3 11.6853
R123 a_334_368.n25 a_334_368.n24 10.955
R124 a_334_368.n16 a_334_368.n15 8.03383
R125 a_334_368.n9 a_334_368.n8 5.84292
R126 a_334_368.n15 a_334_368.n14 5.11262
R127 a_334_368.n17 a_334_368.n1 5.11262
R128 a_334_368.n6 a_334_368.n5 1.46111
R129 VNB.t9 VNB.t11 2286.61
R130 VNB.t8 VNB.t9 1339.63
R131 VNB.t0 VNB.t1 1154.86
R132 VNB.t2 VNB.t5 1154.86
R133 VNB.t10 VNB.t3 1154.86
R134 VNB VNB.t8 1143.31
R135 VNB.t6 VNB.t0 1131.76
R136 VNB.t1 VNB.t4 993.177
R137 VNB.t7 VNB.t6 993.177
R138 VNB.t5 VNB.t7 993.177
R139 VNB.t3 VNB.t2 993.177
R140 VNB.t12 VNB.t10 993.177
R141 VNB.t11 VNB.t12 993.177
R142 A.n0 A.t0 207.99
R143 A.n0 A.t1 189.588
R144 A A.n0 159.442
R145 a_27_112.t1 a_27_112.n1 429.495
R146 a_27_112.n1 a_27_112.t0 269.447
R147 a_27_112.n0 a_27_112.t2 263.589
R148 a_27_112.n0 a_27_112.t3 203.339
R149 a_27_112.n1 a_27_112.n0 152
R150 VPWR.n28 VPWR.n1 613.665
R151 VPWR.n3 VPWR.n2 327.825
R152 VPWR.n7 VPWR.n6 324.615
R153 VPWR.n11 VPWR.n10 324.279
R154 VPWR.n15 VPWR.n9 322.288
R155 VPWR.n12 VPWR.t6 258.418
R156 VPWR.n21 VPWR.n5 223.696
R157 VPWR.n1 VPWR.t12 46.2432
R158 VPWR.n1 VPWR.t11 37.5243
R159 VPWR.n27 VPWR.n26 36.1417
R160 VPWR.n26 VPWR.n3 35.3887
R161 VPWR.n5 VPWR.t10 35.1791
R162 VPWR.n20 VPWR.n7 32.7534
R163 VPWR.n22 VPWR.n21 30.8711
R164 VPWR.n16 VPWR.n15 27.8593
R165 VPWR.n9 VPWR.t3 27.2639
R166 VPWR.n2 VPWR.t9 26.3844
R167 VPWR.n2 VPWR.t8 26.3844
R168 VPWR.n5 VPWR.t2 26.3844
R169 VPWR.n6 VPWR.t0 26.3844
R170 VPWR.n6 VPWR.t7 26.3844
R171 VPWR.n9 VPWR.t1 26.3844
R172 VPWR.n10 VPWR.t5 26.3844
R173 VPWR.n10 VPWR.t4 26.3844
R174 VPWR.n14 VPWR.n11 23.7181
R175 VPWR.n15 VPWR.n14 23.7181
R176 VPWR.n28 VPWR.n27 21.0829
R177 VPWR.n16 VPWR.n7 20.3299
R178 VPWR.n22 VPWR.n3 19.577
R179 VPWR.n21 VPWR.n20 16.5652
R180 VPWR.n14 VPWR.n13 9.3005
R181 VPWR.n15 VPWR.n8 9.3005
R182 VPWR.n17 VPWR.n16 9.3005
R183 VPWR.n18 VPWR.n7 9.3005
R184 VPWR.n20 VPWR.n19 9.3005
R185 VPWR.n21 VPWR.n4 9.3005
R186 VPWR.n23 VPWR.n22 9.3005
R187 VPWR.n24 VPWR.n3 9.3005
R188 VPWR.n26 VPWR.n25 9.3005
R189 VPWR.n27 VPWR.n0 9.3005
R190 VPWR.n29 VPWR.n28 7.27223
R191 VPWR.n12 VPWR.n11 6.85856
R192 VPWR.n13 VPWR.n12 0.630035
R193 VPWR VPWR.n29 0.157962
R194 VPWR.n29 VPWR.n0 0.149814
R195 VPWR.n13 VPWR.n8 0.122949
R196 VPWR.n17 VPWR.n8 0.122949
R197 VPWR.n18 VPWR.n17 0.122949
R198 VPWR.n19 VPWR.n18 0.122949
R199 VPWR.n19 VPWR.n4 0.122949
R200 VPWR.n23 VPWR.n4 0.122949
R201 VPWR.n24 VPWR.n23 0.122949
R202 VPWR.n25 VPWR.n24 0.122949
R203 VPWR.n25 VPWR.n0 0.122949
R204 VPB.t12 VPB.t8 515.861
R205 VPB.t11 VPB.t12 268.146
R206 VPB VPB.t11 257.93
R207 VPB.t0 VPB.t5 255.376
R208 VPB.t10 VPB.t0 255.376
R209 VPB.t7 VPB.t1 232.393
R210 VPB.t3 VPB.t4 229.839
R211 VPB.t2 VPB.t3 229.839
R212 VPB.t1 VPB.t2 229.839
R213 VPB.t6 VPB.t7 229.839
R214 VPB.t5 VPB.t6 229.839
R215 VPB.t9 VPB.t10 229.839
R216 VPB.t8 VPB.t9 229.839
R217 X.n2 X.n0 260.695
R218 X.n2 X.n1 211.54
R219 X.n4 X.n3 210.34
R220 X.n6 X.n5 209.938
R221 X.n11 X.n10 185
R222 X.n9 X.n8 185
R223 X.n9 X.n7 137.388
R224 X.n13 X.n12 98.2201
R225 X.n4 X.n2 48.1887
R226 X.n11 X.n9 45.5685
R227 X.n6 X.n4 45.177
R228 X.n13 X.n11 40.7045
R229 X.n0 X.t0 35.1791
R230 X.n10 X.t8 27.5681
R231 X.n10 X.t14 27.5681
R232 X.n0 X.t5 26.3844
R233 X.n1 X.t7 26.3844
R234 X.n1 X.t6 26.3844
R235 X.n3 X.t2 26.3844
R236 X.n3 X.t1 26.3844
R237 X.n5 X.t4 26.3844
R238 X.n5 X.t3 26.3844
R239 X.n12 X.t12 22.7032
R240 X.n12 X.t9 22.7032
R241 X.n8 X.t15 22.7032
R242 X.n8 X.t13 22.7032
R243 X.n7 X.t10 22.7032
R244 X.n7 X.t11 22.7032
R245 X X.n13 15.1183
R246 X X.n6 7.60245
C0 X VGND 0.448736f
C1 VPB A 0.043072f
C2 VPB VPWR 0.214316f
C3 A VPWR 0.012727f
C4 VPB X 0.0255f
C5 VPB VGND 0.012108f
C6 A X 1.15e-19
C7 VPWR X 0.842854f
C8 A VGND 0.012208f
C9 VPWR VGND 0.120325f
C10 VGND VNB 0.889006f
C11 X VNB 0.064122f
C12 VPWR VNB 0.695827f
C13 A VNB 0.157043f
C14 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__bufinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__bufinv_8 VNB VPB VPWR VGND Y A
X0 VPWR.t11 A.t0 a_27_368.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_183_48.t2 a_27_368.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X2 Y.t15 a_183_48.t6 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3 Y.t14 a_183_48.t7 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 Y.t7 a_183_48.t8 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2408 pd=1.55 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t4 a_183_48.t9 Y.t6 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t5 a_183_48.t10 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VGND.t11 A.t1 a_27_368.t1 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 a_183_48.t5 a_27_368.t3 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 VGND.t5 a_183_48.t11 Y.t13 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 VPWR.t6 a_183_48.t12 Y.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t3 a_183_48.t13 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_183_48.t1 a_27_368.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X13 VGND.t4 a_183_48.t14 Y.t12 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VPWR.t8 a_183_48.t15 Y.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 VPWR.t0 a_27_368.t5 a_183_48.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VGND.t3 a_183_48.t16 Y.t11 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.111 ps=1.04 w=0.74 l=0.15
X17 Y.t1 a_183_48.t17 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X18 Y.t10 a_183_48.t18 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X19 VGND.t9 a_27_368.t6 a_183_48.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.10915 ps=1.035 w=0.74 l=0.15
X20 VPWR.t10 a_183_48.t19 Y.t0 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2408 ps=1.55 w=1.12 l=0.15
X21 VGND.t1 a_183_48.t20 Y.t9 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 Y.t8 a_183_48.t21 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1221 ps=1.07 w=0.74 l=0.15
X23 a_183_48.t3 a_27_368.t7 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.1295 ps=1.09 w=0.74 l=0.15
R0 A.n0 A.t0 248.017
R1 A.n0 A.t1 217.221
R2 A A.n0 158.847
R3 a_27_368.n7 a_27_368.n6 338.291
R4 a_27_368.n7 a_27_368.t1 263.87
R5 a_27_368.t0 a_27_368.n7 253.291
R6 a_27_368.n4 a_27_368.t4 237.642
R7 a_27_368.n0 a_27_368.t2 235.537
R8 a_27_368.n3 a_27_368.t5 234.841
R9 a_27_368.n0 a_27_368.t3 188.538
R10 a_27_368.n4 a_27_368.t7 186.374
R11 a_27_368.n2 a_27_368.t6 186.374
R12 a_27_368.n6 a_27_368.n1 158.696
R13 a_27_368.n6 a_27_368.n5 152
R14 a_27_368.n5 a_27_368.n4 48.9308
R15 a_27_368.n1 a_27_368.n0 37.2697
R16 a_27_368.n2 a_27_368.n1 33.5944
R17 a_27_368.n5 a_27_368.n3 14.6066
R18 a_27_368.n3 a_27_368.n2 1.46111
R19 VPWR.n11 VPWR.n10 617.255
R20 VPWR.n22 VPWR.n1 607.692
R21 VPWR.n20 VPWR.n3 607.692
R22 VPWR.n5 VPWR.n4 607.692
R23 VPWR.n14 VPWR.n7 607.692
R24 VPWR.n9 VPWR.n8 607.692
R25 VPWR.n1 VPWR.t11 35.1791
R26 VPWR.n8 VPWR.t1 35.1791
R27 VPWR.n10 VPWR.t0 35.1791
R28 VPWR.n14 VPWR.n13 32.7534
R29 VPWR.n15 VPWR.n5 28.2358
R30 VPWR.n1 VPWR.t9 26.3844
R31 VPWR.n3 VPWR.t7 26.3844
R32 VPWR.n3 VPWR.t8 26.3844
R33 VPWR.n4 VPWR.t5 26.3844
R34 VPWR.n4 VPWR.t6 26.3844
R35 VPWR.n7 VPWR.t3 26.3844
R36 VPWR.n7 VPWR.t4 26.3844
R37 VPWR.n8 VPWR.t10 26.3844
R38 VPWR.n10 VPWR.t2 26.3844
R39 VPWR.n21 VPWR.n20 23.7181
R40 VPWR.n20 VPWR.n19 23.7181
R41 VPWR.n13 VPWR.n9 19.9534
R42 VPWR.n22 VPWR.n21 19.2005
R43 VPWR.n19 VPWR.n5 19.2005
R44 VPWR.n15 VPWR.n14 14.6829
R45 VPWR.n13 VPWR.n12 9.3005
R46 VPWR.n14 VPWR.n6 9.3005
R47 VPWR.n16 VPWR.n15 9.3005
R48 VPWR.n17 VPWR.n5 9.3005
R49 VPWR.n19 VPWR.n18 9.3005
R50 VPWR.n20 VPWR.n2 9.3005
R51 VPWR.n21 VPWR.n0 9.3005
R52 VPWR.n23 VPWR.n22 7.43488
R53 VPWR.n11 VPWR.n9 6.94321
R54 VPWR.n12 VPWR.n11 0.516733
R55 VPWR VPWR.n23 0.160103
R56 VPWR.n23 VPWR.n0 0.1477
R57 VPWR.n12 VPWR.n6 0.122949
R58 VPWR.n16 VPWR.n6 0.122949
R59 VPWR.n17 VPWR.n16 0.122949
R60 VPWR.n18 VPWR.n17 0.122949
R61 VPWR.n18 VPWR.n2 0.122949
R62 VPWR.n2 VPWR.n0 0.122949
R63 VPB.t3 VPB.t10 296.238
R64 VPB VPB.t11 257.93
R65 VPB.t0 VPB.t2 255.376
R66 VPB.t10 VPB.t1 255.376
R67 VPB.t11 VPB.t9 255.376
R68 VPB.t1 VPB.t0 229.839
R69 VPB.t4 VPB.t3 229.839
R70 VPB.t5 VPB.t4 229.839
R71 VPB.t6 VPB.t5 229.839
R72 VPB.t7 VPB.t6 229.839
R73 VPB.t8 VPB.t7 229.839
R74 VPB.t9 VPB.t8 229.839
R75 a_183_48.n33 a_183_48.n32 350.305
R76 a_183_48.n2 a_183_48.t19 240.197
R77 a_183_48.n25 a_183_48.t8 240.197
R78 a_183_48.n5 a_183_48.t9 240.197
R79 a_183_48.n18 a_183_48.t10 240.197
R80 a_183_48.n11 a_183_48.t12 240.197
R81 a_183_48.n12 a_183_48.t13 240.197
R82 a_183_48.n9 a_183_48.t15 240.197
R83 a_183_48.n7 a_183_48.t17 240.197
R84 a_183_48.t2 a_183_48.n33 224.606
R85 a_183_48.n7 a_183_48.t21 182.138
R86 a_183_48.n2 a_183_48.t11 182.138
R87 a_183_48.n8 a_183_48.t16 179.947
R88 a_183_48.n13 a_183_48.t7 179.947
R89 a_183_48.n6 a_183_48.t14 179.947
R90 a_183_48.n20 a_183_48.t6 179.947
R91 a_183_48.n3 a_183_48.t20 179.947
R92 a_183_48.n26 a_183_48.t18 179.947
R93 a_183_48.n15 a_183_48.n10 165.189
R94 a_183_48.n15 a_183_48.n14 152
R95 a_183_48.n17 a_183_48.n16 152
R96 a_183_48.n19 a_183_48.n4 152
R97 a_183_48.n22 a_183_48.n21 152
R98 a_183_48.n24 a_183_48.n23 152
R99 a_183_48.n27 a_183_48.n1 152
R100 a_183_48.n29 a_183_48.n28 152
R101 a_183_48.n31 a_183_48.t5 145.654
R102 a_183_48.n30 a_183_48.n0 97.8675
R103 a_183_48.n8 a_183_48.n7 63.5369
R104 a_183_48.n10 a_183_48.n9 54.7732
R105 a_183_48.n28 a_183_48.n27 49.6611
R106 a_183_48.n30 a_183_48.n29 47.7561
R107 a_183_48.n21 a_183_48.n20 46.7399
R108 a_183_48.n33 a_183_48.n31 44.0715
R109 a_183_48.n18 a_183_48.n17 43.0884
R110 a_183_48.n31 a_183_48.n30 39.6805
R111 a_183_48.n24 a_183_48.n3 33.5944
R112 a_183_48.n14 a_183_48.n13 33.5944
R113 a_183_48.n14 a_183_48.n11 27.0217
R114 a_183_48.n32 a_183_48.t0 26.3844
R115 a_183_48.n32 a_183_48.t1 26.3844
R116 a_183_48.n25 a_183_48.n24 25.5611
R117 a_183_48.n0 a_183_48.t4 24.3248
R118 a_183_48.n0 a_183_48.t3 23.514
R119 a_183_48.n17 a_183_48.n6 20.449
R120 a_183_48.n26 a_183_48.n25 13.8763
R121 a_183_48.n29 a_183_48.n1 13.1884
R122 a_183_48.n23 a_183_48.n1 13.1884
R123 a_183_48.n23 a_183_48.n22 13.1884
R124 a_183_48.n22 a_183_48.n4 13.1884
R125 a_183_48.n16 a_183_48.n4 13.1884
R126 a_183_48.n16 a_183_48.n15 13.1884
R127 a_183_48.n28 a_183_48.n2 10.955
R128 a_183_48.n12 a_183_48.n10 10.955
R129 a_183_48.n27 a_183_48.n26 10.2247
R130 a_183_48.n21 a_183_48.n5 9.49444
R131 a_183_48.n5 a_183_48.n3 6.57323
R132 a_183_48.n19 a_183_48.n18 6.57323
R133 a_183_48.n13 a_183_48.n12 5.11262
R134 a_183_48.n20 a_183_48.n19 2.92171
R135 a_183_48.n11 a_183_48.n6 2.19141
R136 a_183_48.n9 a_183_48.n8 2.19141
R137 VGND.n9 VGND.n6 211.632
R138 VGND.n12 VGND.n5 209.243
R139 VGND.n22 VGND.n21 208.079
R140 VGND.n19 VGND.n2 207.109
R141 VGND.n8 VGND.n7 206.139
R142 VGND.n15 VGND.n14 206.139
R143 VGND.n6 VGND.t10 34.0546
R144 VGND.n7 VGND.t5 34.0546
R145 VGND.n5 VGND.t1 34.0546
R146 VGND.n14 VGND.t7 34.0546
R147 VGND.n2 VGND.t3 34.0546
R148 VGND.n21 VGND.t0 30.8113
R149 VGND.n15 VGND.n13 27.8593
R150 VGND.n20 VGND.n19 27.1064
R151 VGND.n8 VGND.n4 25.6005
R152 VGND.n12 VGND.n4 24.8476
R153 VGND.n22 VGND.n20 23.3417
R154 VGND.n6 VGND.t9 22.7032
R155 VGND.n7 VGND.t8 22.7032
R156 VGND.n5 VGND.t2 22.7032
R157 VGND.n14 VGND.t4 22.7032
R158 VGND.n2 VGND.t6 22.7032
R159 VGND.n21 VGND.t11 22.7032
R160 VGND.n13 VGND.n12 22.5887
R161 VGND.n19 VGND.n1 20.3299
R162 VGND.n15 VGND.n1 19.577
R163 VGND.n10 VGND.n4 9.3005
R164 VGND.n12 VGND.n11 9.3005
R165 VGND.n13 VGND.n3 9.3005
R166 VGND.n16 VGND.n15 9.3005
R167 VGND.n17 VGND.n1 9.3005
R168 VGND.n19 VGND.n18 9.3005
R169 VGND.n20 VGND.n0 9.3005
R170 VGND.n23 VGND.n22 7.25439
R171 VGND.n9 VGND.n8 6.52845
R172 VGND.n10 VGND.n9 0.629588
R173 VGND VGND.n23 0.157727
R174 VGND.n23 VGND.n0 0.150046
R175 VGND.n11 VGND.n10 0.122949
R176 VGND.n11 VGND.n3 0.122949
R177 VGND.n16 VGND.n3 0.122949
R178 VGND.n17 VGND.n16 0.122949
R179 VGND.n18 VGND.n17 0.122949
R180 VGND.n18 VGND.n0 0.122949
R181 Y.n2 Y.n0 630.749
R182 Y.n6 Y.n5 586.939
R183 Y.n2 Y.n1 585
R184 Y.n4 Y.n3 585
R185 Y.n14 Y.n13 185
R186 Y.n13 Y.n12 185
R187 Y.n10 Y.n8 151.77
R188 Y.n11 Y.n7 98.2648
R189 Y.n10 Y.n9 98.2201
R190 Y.n4 Y.n2 42.6672
R191 Y.n11 Y.n10 39.1685
R192 Y.n15 Y.n11 39.1685
R193 Y.n0 Y.t0 37.8175
R194 Y.n0 Y.t7 37.8175
R195 Y.n6 Y.n4 35.082
R196 Y.n8 Y.t10 34.0546
R197 Y.n5 Y.t2 26.3844
R198 Y.n5 Y.t1 26.3844
R199 Y.n3 Y.t4 26.3844
R200 Y.n3 Y.t3 26.3844
R201 Y.n1 Y.t6 26.3844
R202 Y.n1 Y.t5 26.3844
R203 Y.n13 Y.t8 25.9464
R204 Y.n13 Y.t11 22.7032
R205 Y.n7 Y.t12 22.7032
R206 Y.n7 Y.t14 22.7032
R207 Y.n9 Y.t9 22.7032
R208 Y.n9 Y.t15 22.7032
R209 Y.n8 Y.t13 22.7032
R210 Y Y.n6 13.7702
R211 Y.n12 Y 12.6066
R212 Y Y.n15 7.95202
R213 Y.n14 Y 4.84898
R214 Y.n12 Y 1.74595
R215 Y.n15 Y.n14 1.55202
R216 VNB VNB.t11 1177.95
R217 VNB.t9 VNB.t10 1154.86
R218 VNB.t5 VNB.t8 1154.86
R219 VNB.t2 VNB.t5 1154.86
R220 VNB.t1 VNB.t2 1154.86
R221 VNB.t4 VNB.t7 1154.86
R222 VNB.t3 VNB.t6 1154.86
R223 VNB.t11 VNB.t0 1108.66
R224 VNB.t0 VNB.t3 1039.37
R225 VNB.t8 VNB.t9 1027.82
R226 VNB.t7 VNB.t1 993.177
R227 VNB.t6 VNB.t4 993.177
C0 VPB A 0.03923f
C1 VPB VPWR 0.163802f
C2 VPB Y 0.012587f
C3 A VPWR 0.015202f
C4 A Y 7.67e-19
C5 VPB VGND 0.008268f
C6 VPWR Y 0.084206f
C7 A VGND 0.017679f
C8 VPWR VGND 0.1033f
C9 Y VGND 0.55494f
C10 VGND VNB 0.731944f
C11 Y VNB 0.02775f
C12 VPWR VNB 0.57501f
C13 A VNB 0.157515f
C14 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkbuf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkbuf_1 VNB VPB VPWR VGND A X
X0 VGND.t1 A.t0 a_27_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1 X.t1 a_27_74.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2 X.t0 a_27_74.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X3 VPWR.t1 A.t1 a_27_74.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 A.n0 A.t1 251.151
R1 A.n1 A.t0 231.361
R2 A.n2 A.n1 177.561
R3 A.n0 A 152.667
R4 A.n1 A.n0 24.1005
R5 A.n2 A 8.4005
R6 A A.n2 4.4005
R7 a_27_74.t1 a_27_74.n3 292.627
R8 a_27_74.n0 a_27_74.t0 287.827
R9 a_27_74.n2 a_27_74.t2 258.479
R10 a_27_74.n3 a_27_74.n2 152
R11 a_27_74.n1 a_27_74.n0 152
R12 a_27_74.n1 a_27_74.t3 140.389
R13 a_27_74.n2 a_27_74.n1 37.6741
R14 a_27_74.n3 a_27_74.n0 11.1595
R15 VGND.n0 VGND.t0 100.353
R16 VGND.n0 VGND.t1 100.343
R17 VGND VGND.n0 76.7841
R18 VNB.t1 VNB.t0 2148.03
R19 VNB VNB.t1 1143.31
R20 VPWR VPWR.n0 322.301
R21 VPWR.n0 VPWR.t0 35.1791
R22 VPWR.n0 VPWR.t1 35.1791
R23 X.n1 X 588.479
R24 X.n1 X.n0 585
R25 X.n2 X.n1 585
R26 X.n3 X.t0 216.073
R27 X.n1 X.t1 26.3844
R28 X X.n3 11.2005
R29 X.n2 X 9.32224
R30 X.n0 X 8.07007
R31 X.n3 X 3.87929
R32 X.n0 X 2.22659
R33 X X.n2 0.974413
R34 VPB VPB.t1 375.404
R35 VPB.t1 VPB.t0 280.914
C0 VPWR VGND 0.032165f
C1 X VGND 0.067618f
C2 A VPB 0.060059f
C3 VPWR VPB 0.060213f
C4 X VPB 0.019632f
C5 VGND VPB 0.006869f
C6 A VPWR 0.019428f
C7 A X 0.00109f
C8 A VGND 0.017997f
C9 VPWR X 0.110867f
C10 VGND VNB 0.280599f
C11 X VNB 0.114659f
C12 VPWR VNB 0.229932f
C13 A VNB 0.224803f
C14 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkbuf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkbuf_2 VNB VPB VPWR VGND X A
X0 a_43_192.t0 A.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3528 pd=2.87 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t1 a_43_192.t2 X.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 X.t0 a_43_192.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X3 a_43_192.t1 A.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X4 X.t1 a_43_192.t4 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5 VGND.t0 a_43_192.t5 X.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A.n1 A.t0 250.909
R1 A.n0 A.t1 162.274
R2 A.n0 A 153.094
R3 A.n2 A.n1 152
R4 A.n1 A.n0 49.6611
R5 A.n2 A 9.52245
R6 A A.n2 2.02977
R7 VPWR.n1 VPWR.t2 875.543
R8 VPWR.n1 VPWR.n0 611.904
R9 VPWR.n0 VPWR.t0 26.3844
R10 VPWR.n0 VPWR.t1 26.3844
R11 VPWR VPWR.n1 0.538891
R12 a_43_192.n3 a_43_192.t1 350.5
R13 a_43_192.t0 a_43_192.n3 324.954
R14 a_43_192.n1 a_43_192.t4 240.197
R15 a_43_192.n1 a_43_192.t2 240.197
R16 a_43_192.n3 a_43_192.n2 225.81
R17 a_43_192.n0 a_43_192.t5 122.108
R18 a_43_192.n0 a_43_192.t3 122.108
R19 a_43_192.n2 a_43_192.n0 19.491
R20 a_43_192.n2 a_43_192.n1 18.7093
R21 VPB VPB.t0 252.823
R22 VPB.t1 VPB.t2 229.839
R23 VPB.t0 VPB.t1 229.839
R24 X.n2 X.n0 677.236
R25 X.n2 X.n1 185
R26 X.n1 X.t3 40.0005
R27 X.n1 X.t0 40.0005
R28 X.n0 X.t2 26.3844
R29 X.n0 X.t1 26.3844
R30 X X.n2 3.76521
R31 VGND.n1 VGND.t1 261.106
R32 VGND.n1 VGND.n0 220.577
R33 VGND.n0 VGND.t2 60.0005
R34 VGND.n0 VGND.t0 40.0005
R35 VGND VGND.n1 0.447384
R36 VNB.t0 VNB.t2 1154.86
R37 VNB VNB.t1 1143.31
R38 VNB.t1 VNB.t0 993.177
C0 VPB A 0.036208f
C1 VPB VPWR 0.059632f
C2 VPB X 0.002461f
C3 A VPWR 0.022768f
C4 VGND VPB 0.004922f
C5 A X 0.08642f
C6 VGND A 0.040504f
C7 VPWR X 0.013217f
C8 VGND VPWR 0.034238f
C9 VGND X 0.110719f
C10 VGND VNB 0.305552f
C11 X VNB 0.012652f
C12 VPWR VNB 0.238361f
C13 A VNB 0.17296f
C14 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkbuf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkbuf_4 VNB VPB VPWR VGND A X
X0 X.t7 a_83_270.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 X.t3 a_83_270.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X2 a_83_270.t1 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X3 a_83_270.t0 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.126 pd=1.44 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 VPWR.t3 a_83_270.t4 X.t6 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5 X.t5 a_83_270.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t1 a_83_270.t6 X.t4 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VGND.t3 a_83_270.t7 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND.t2 a_83_270.t8 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.0672 ps=0.74 w=0.42 l=0.15
X9 X.t0 a_83_270.t9 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 a_83_270.n11 a_83_270.t0 292.901
R1 a_83_270.n2 a_83_270.t3 247.428
R2 a_83_270.n3 a_83_270.t7 247.428
R3 a_83_270.n6 a_83_270.t9 247.428
R4 a_83_270.n1 a_83_270.t8 247.428
R5 a_83_270.t1 a_83_270.n11 239.762
R6 a_83_270.n1 a_83_270.t4 229
R7 a_83_270.n2 a_83_270.t2 227.538
R8 a_83_270.n8 a_83_270.t5 226.809
R9 a_83_270.n4 a_83_270.t6 226.809
R10 a_83_270.n5 a_83_270.n0 162.881
R11 a_83_270.n7 a_83_270.n0 152
R12 a_83_270.n10 a_83_270.n9 152
R13 a_83_270.n3 a_83_270.n2 62.8066
R14 a_83_270.n6 a_83_270.n5 48.2005
R15 a_83_270.n9 a_83_270.n8 46.0096
R16 a_83_270.n11 a_83_270.n10 45.1864
R17 a_83_270.n9 a_83_270.n1 17.5278
R18 a_83_270.n5 a_83_270.n4 12.4157
R19 a_83_270.n10 a_83_270.n0 10.8805
R20 a_83_270.n8 a_83_270.n7 3.65202
R21 a_83_270.n4 a_83_270.n3 2.19141
R22 a_83_270.n7 a_83_270.n6 1.46111
R23 VPWR.n4 VPWR.n3 323.777
R24 VPWR.n6 VPWR.t4 259.171
R25 VPWR.n2 VPWR.n1 237.343
R26 VPWR.n1 VPWR.t0 35.1791
R27 VPWR.n6 VPWR.n5 26.7299
R28 VPWR.n3 VPWR.t2 26.3844
R29 VPWR.n3 VPWR.t1 26.3844
R30 VPWR.n1 VPWR.t3 26.3844
R31 VPWR.n5 VPWR.n4 22.2123
R32 VPWR.n5 VPWR.n0 9.3005
R33 VPWR.n7 VPWR.n6 9.3005
R34 VPWR.n4 VPWR.n2 7.12969
R35 VPWR.n2 VPWR.n0 0.486971
R36 VPWR.n7 VPWR.n0 0.122949
R37 VPWR VPWR.n7 0.0617245
R38 X.n3 X.n1 254.738
R39 X.n4 X.n0 243.719
R40 X.n3 X.n2 207.689
R41 X.n7 X.n6 185
R42 X.n4 X.n3 64.9275
R43 X.n0 X.t1 51.4291
R44 X.n6 X.t2 40.0005
R45 X.n6 X.t3 40.0005
R46 X.n0 X.t0 40.0005
R47 X.n2 X.t4 26.3844
R48 X.n2 X.t7 26.3844
R49 X.n1 X.t6 26.3844
R50 X.n1 X.t5 26.3844
R51 X X.n7 10.0853
R52 X X.n5 5.4308
R53 X.n5 X 5.04839
R54 X.n7 X 4.26717
R55 X.n5 X.n4 3.06529
R56 VPB VPB.t4 257.93
R57 VPB.t3 VPB.t0 255.376
R58 VPB.t2 VPB.t3 229.839
R59 VPB.t1 VPB.t2 229.839
R60 VPB.t4 VPB.t1 229.839
R61 VGND.n6 VGND.t4 254.696
R62 VGND.n4 VGND.n1 222.272
R63 VGND.n3 VGND.n2 213.114
R64 VGND.n2 VGND.t0 60.0005
R65 VGND.n2 VGND.t2 48.5719
R66 VGND.n1 VGND.t1 40.0005
R67 VGND.n1 VGND.t3 40.0005
R68 VGND.n5 VGND.n4 32.7534
R69 VGND.n6 VGND.n5 25.6005
R70 VGND.n4 VGND.n3 10.657
R71 VGND.n7 VGND.n6 9.3005
R72 VGND.n5 VGND.n0 9.3005
R73 VGND.n3 VGND.n0 0.504912
R74 VGND.n7 VGND.n0 0.122949
R75 VGND VGND.n7 0.0617245
R76 VNB.t2 VNB.t0 1224.15
R77 VNB VNB.t4 1177.95
R78 VNB.t1 VNB.t2 1085.56
R79 VNB.t3 VNB.t1 993.177
R80 VNB.t4 VNB.t3 993.177
R81 A.n0 A.t0 323.209
R82 A.n0 A.t1 184.768
R83 A A.n0 161.504
C0 VPB X 0.010279f
C1 A VPWR 0.021828f
C2 VPB VGND 0.005954f
C3 A X 0.00864f
C4 A VGND 0.03462f
C5 VPWR X 0.399795f
C6 VPWR VGND 0.056142f
C7 X VGND 0.250325f
C8 VPB A 0.032094f
C9 VPB VPWR 0.091009f
C10 VGND VNB 0.422577f
C11 X VNB 0.06623f
C12 VPWR VNB 0.353137f
C13 A VNB 0.173268f
C14 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__buf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__buf_16 VNB VPB VPWR X VGND A
X0 X.t29 a_83_260# VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 X.t15 a_83_260# VPWR.t21 VPB.t21 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t20 a_83_260# X.t14 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X.t13 a_83_260# VPWR.t19 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 X.t28 a_83_260# VGND.t16 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VGND.t15 a_83_260# X.t27 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VGND.t1 A.t0 a_83_260# VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X8 VPWR.t18 a_83_260# X.t12 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_83_260# A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_83_260# A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 X.t11 a_83_260# VPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VPWR.t2 A.t3 a_83_260# VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VPWR.t16 a_83_260# X.t10 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 X.t26 a_83_260# VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 X.t25 a_83_260# VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_83_260# A.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 X.t9 a_83_260# VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X18 VPWR.t4 A.t5 a_83_260# VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_83_260# A.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_83_260# A.t7 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X21 VGND.t12 a_83_260# X.t24 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 a_83_260# A.t8 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.11655 ps=1.055 w=0.74 l=0.15
X23 VGND.t11 a_83_260# X.t23 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 X.t22 a_83_260# VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X25 VGND.t9 a_83_260# X.t21 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 X.t20 a_83_260# VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X27 VPWR.t14 a_83_260# X.t8 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X28 X.t7 a_83_260# VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 VPWR.t12 a_83_260# X.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 VPWR.t11 a_83_260# X.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X32 X.t4 a_83_260# VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X33 VGND.t7 a_83_260# X.t19 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X34 VPWR.t9 a_83_260# X.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X35 X.t2 a_83_260# VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X36 X.t1 a_83_260# VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X37 VGND.t6 a_83_260# X.t18 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X38 VPWR.t6 a_83_260# X.t0 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X39 X.t17 a_83_260# VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X40 VPWR.t0 A.t9 a_83_260# VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X41 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1036 ps=1.02 w=0.74 l=0.15
X42 X.t16 a_83_260# VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X43 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 VGND.n12 VGND.t0 239.56
R1 VGND.n16 VGND.t2 233.886
R2 VGND.n10 VGND.t3 233.886
R3 VGND.n48 VGND.t14 171.77
R4 VGND.n13 VGND.t1 170.745
R5 VGND.n22 VGND.t10 149.756
R6 VGND.n32 VGND.n31 131.446
R7 VGND.n41 VGND.n40 130.206
R8 VGND.n38 VGND.n4 129.603
R9 VGND.n30 VGND.n29 120.704
R10 VGND.n46 VGND.n2 118.811
R11 VGND.n8 VGND.n7 115.2
R12 VGND.n24 VGND.n23 36.1417
R13 VGND.n37 VGND.n5 36.1417
R14 VGND.n42 VGND.n39 36.1417
R15 VGND.n33 VGND.n30 35.7652
R16 VGND.n21 VGND.n10 35.3887
R17 VGND.n28 VGND.n8 34.6358
R18 VGND.n7 VGND.t4 34.0546
R19 VGND.n7 VGND.t15 34.0546
R20 VGND.n29 VGND.t8 34.0546
R21 VGND.n29 VGND.t6 34.0546
R22 VGND.n46 VGND.n1 29.7417
R23 VGND.n17 VGND.n16 27.8593
R24 VGND.n33 VGND.n32 25.977
R25 VGND.n48 VGND.n47 25.6005
R26 VGND.n31 VGND.t17 22.7032
R27 VGND.n31 VGND.t12 22.7032
R28 VGND.n4 VGND.t16 22.7032
R29 VGND.n4 VGND.t11 22.7032
R30 VGND.n40 VGND.t13 22.7032
R31 VGND.n40 VGND.t9 22.7032
R32 VGND.n2 VGND.t5 22.7032
R33 VGND.n2 VGND.t7 22.7032
R34 VGND.n15 VGND.n12 20.3299
R35 VGND.n47 VGND.n46 20.3299
R36 VGND.n16 VGND.n15 19.577
R37 VGND.n38 VGND.n37 18.4476
R38 VGND.n39 VGND.n38 17.6946
R39 VGND.n41 VGND.n1 16.1887
R40 VGND.n30 VGND.n28 15.8123
R41 VGND.n24 VGND.n8 12.8005
R42 VGND.n17 VGND.n10 12.0476
R43 VGND.n32 VGND.n5 10.1652
R44 VGND.n22 VGND.n21 9.78874
R45 VGND.n49 VGND.n48 9.3005
R46 VGND.n15 VGND.n14 9.3005
R47 VGND.n16 VGND.n11 9.3005
R48 VGND.n18 VGND.n17 9.3005
R49 VGND.n19 VGND.n10 9.3005
R50 VGND.n21 VGND.n20 9.3005
R51 VGND.n23 VGND.n9 9.3005
R52 VGND.n25 VGND.n24 9.3005
R53 VGND.n26 VGND.n8 9.3005
R54 VGND.n28 VGND.n27 9.3005
R55 VGND.n30 VGND.n6 9.3005
R56 VGND.n34 VGND.n33 9.3005
R57 VGND.n35 VGND.n5 9.3005
R58 VGND.n37 VGND.n36 9.3005
R59 VGND.n39 VGND.n3 9.3005
R60 VGND.n43 VGND.n42 9.3005
R61 VGND.n44 VGND.n1 9.3005
R62 VGND.n46 VGND.n45 9.3005
R63 VGND.n47 VGND.n0 9.3005
R64 VGND.n13 VGND.n12 6.81903
R65 VGND.n42 VGND.n41 4.51815
R66 VGND.n23 VGND.n22 1.50638
R67 VGND.n14 VGND.n13 0.623326
R68 VGND.n14 VGND.n11 0.122949
R69 VGND.n18 VGND.n11 0.122949
R70 VGND.n19 VGND.n18 0.122949
R71 VGND.n20 VGND.n19 0.122949
R72 VGND.n20 VGND.n9 0.122949
R73 VGND.n25 VGND.n9 0.122949
R74 VGND.n26 VGND.n25 0.122949
R75 VGND.n27 VGND.n26 0.122949
R76 VGND.n27 VGND.n6 0.122949
R77 VGND.n34 VGND.n6 0.122949
R78 VGND.n35 VGND.n34 0.122949
R79 VGND.n36 VGND.n35 0.122949
R80 VGND.n36 VGND.n3 0.122949
R81 VGND.n43 VGND.n3 0.122949
R82 VGND.n44 VGND.n43 0.122949
R83 VGND.n45 VGND.n44 0.122949
R84 VGND.n45 VGND.n0 0.122949
R85 VGND.n49 VGND.n0 0.122949
R86 VGND VGND.n49 0.0617245
R87 X.n27 X.n25 204.577
R88 X.n23 X.n22 204.577
R89 X.n15 X.n14 204.577
R90 X.n19 X.n18 204.399
R91 X.n1 X.n0 204.227
R92 X.n3 X.n2 204.061
R93 X.n7 X.n6 203.315
R94 X.n11 X.n10 202.457
R95 X.n1 X.t22 197.91
R96 X.n3 X.t16 193.419
R97 X.n15 X.n13 167.712
R98 X.n11 X.n9 164.12
R99 X.n27 X.n26 150.649
R100 X.n23 X.n21 150.649
R101 X.n19 X.n17 147.464
R102 X.n7 X.n5 141.232
R103 X.n25 X.t5 26.3844
R104 X.n25 X.t15 26.3844
R105 X.n22 X.t8 26.3844
R106 X.n22 X.t7 26.3844
R107 X.n18 X.t10 26.3844
R108 X.n18 X.t9 26.3844
R109 X.n14 X.t12 26.3844
R110 X.n14 X.t11 26.3844
R111 X.n10 X.t14 26.3844
R112 X.n10 X.t13 26.3844
R113 X.n6 X.t0 26.3844
R114 X.n6 X.t2 26.3844
R115 X.n2 X.t3 26.3844
R116 X.n2 X.t1 26.3844
R117 X.n0 X.t6 26.3844
R118 X.n0 X.t4 26.3844
R119 X.n26 X.t19 22.7032
R120 X.n26 X.t26 22.7032
R121 X.n21 X.t21 22.7032
R122 X.n21 X.t17 22.7032
R123 X.n17 X.t23 22.7032
R124 X.n17 X.t25 22.7032
R125 X.n13 X.t24 22.7032
R126 X.n13 X.t28 22.7032
R127 X.n9 X.t18 22.7032
R128 X.n9 X.t29 22.7032
R129 X.n5 X.t27 22.7032
R130 X.n5 X.t20 22.7032
R131 X.n4 X.n1 10.6496
R132 X.n28 X.n27 10.1787
R133 X.n24 X.n23 10.1787
R134 X.n16 X.n15 10.1787
R135 X.n20 X.n19 10.1611
R136 X.n4 X.n3 10.1278
R137 X.n8 X.n7 10.055
R138 X.n12 X.n11 9.97218
R139 X.n24 X.n20 0.519522
R140 X.n16 X.n12 0.51137
R141 X.n8 X.n4 0.48963
R142 X.n12 X.n8 0.486913
R143 X.n20 X.n16 0.484196
R144 X.n28 X.n24 0.478761
R145 X X.n28 0.0793043
R146 VNB.t4 VNB.t10 2309.71
R147 VNB.t2 VNB.t0 2067.19
R148 VNB.t3 VNB.t2 1986.35
R149 VNB.t10 VNB.t3 1986.35
R150 VNB.t15 VNB.t4 1316.54
R151 VNB.t6 VNB.t8 1316.54
R152 VNB VNB.t14 1177.95
R153 VNB.t0 VNB.t1 1154.86
R154 VNB.t8 VNB.t15 993.177
R155 VNB.t17 VNB.t6 993.177
R156 VNB.t12 VNB.t17 993.177
R157 VNB.t16 VNB.t12 993.177
R158 VNB.t11 VNB.t16 993.177
R159 VNB.t13 VNB.t11 993.177
R160 VNB.t9 VNB.t13 993.177
R161 VNB.t5 VNB.t9 993.177
R162 VNB.t7 VNB.t5 993.177
R163 VNB.t14 VNB.t7 993.177
R164 VPWR.n22 VPWR.n14 331.5
R165 VPWR.n17 VPWR.n16 331.5
R166 VPWR.n25 VPWR.n24 323.406
R167 VPWR.n18 VPWR.t0 262.974
R168 VPWR.n58 VPWR.t21 259.171
R169 VPWR.n56 VPWR.n1 241.419
R170 VPWR.n43 VPWR.n42 241.419
R171 VPWR.n34 VPWR.n33 241.419
R172 VPWR.n40 VPWR.n8 241.2
R173 VPWR.n31 VPWR.n11 241.2
R174 VPWR.n49 VPWR.n5 241.081
R175 VPWR.n51 VPWR.n4 231.036
R176 VPWR.n18 VPWR.n17 40.1055
R177 VPWR.n55 VPWR.n2 36.1417
R178 VPWR.n30 VPWR.n12 36.1417
R179 VPWR.n35 VPWR.n32 36.1417
R180 VPWR.n39 VPWR.n9 36.1417
R181 VPWR.n44 VPWR.n41 36.1417
R182 VPWR.n48 VPWR.n6 36.1417
R183 VPWR.n21 VPWR.n15 36.1417
R184 VPWR.n26 VPWR.n23 36.1417
R185 VPWR.n4 VPWR.t14 35.1791
R186 VPWR.n24 VPWR.t5 35.1791
R187 VPWR.n57 VPWR.n56 34.6358
R188 VPWR.n51 VPWR.n50 32.0005
R189 VPWR.n22 VPWR.n21 30.1181
R190 VPWR.n50 VPWR.n49 29.3652
R191 VPWR.n58 VPWR.n57 26.7299
R192 VPWR.n1 VPWR.t13 26.3844
R193 VPWR.n1 VPWR.t11 26.3844
R194 VPWR.n4 VPWR.t15 26.3844
R195 VPWR.n5 VPWR.t17 26.3844
R196 VPWR.n5 VPWR.t16 26.3844
R197 VPWR.n42 VPWR.t19 26.3844
R198 VPWR.n42 VPWR.t18 26.3844
R199 VPWR.n8 VPWR.t8 26.3844
R200 VPWR.n8 VPWR.t20 26.3844
R201 VPWR.n33 VPWR.t7 26.3844
R202 VPWR.n33 VPWR.t6 26.3844
R203 VPWR.n11 VPWR.t10 26.3844
R204 VPWR.n11 VPWR.t9 26.3844
R205 VPWR.n24 VPWR.t12 26.3844
R206 VPWR.n14 VPWR.t3 26.3844
R207 VPWR.n14 VPWR.t4 26.3844
R208 VPWR.n16 VPWR.t1 26.3844
R209 VPWR.n16 VPWR.t2 26.3844
R210 VPWR.n31 VPWR.n30 24.8476
R211 VPWR.n43 VPWR.n6 24.8476
R212 VPWR.n51 VPWR.n2 21.4593
R213 VPWR.n35 VPWR.n34 20.3299
R214 VPWR.n41 VPWR.n40 20.3299
R215 VPWR.n26 VPWR.n25 16.9417
R216 VPWR.n34 VPWR.n9 15.8123
R217 VPWR.n40 VPWR.n39 15.8123
R218 VPWR.n32 VPWR.n31 11.2946
R219 VPWR.n44 VPWR.n43 11.2946
R220 VPWR.n19 VPWR.n15 9.3005
R221 VPWR.n21 VPWR.n20 9.3005
R222 VPWR.n23 VPWR.n13 9.3005
R223 VPWR.n27 VPWR.n26 9.3005
R224 VPWR.n28 VPWR.n12 9.3005
R225 VPWR.n30 VPWR.n29 9.3005
R226 VPWR.n32 VPWR.n10 9.3005
R227 VPWR.n36 VPWR.n35 9.3005
R228 VPWR.n37 VPWR.n9 9.3005
R229 VPWR.n39 VPWR.n38 9.3005
R230 VPWR.n41 VPWR.n7 9.3005
R231 VPWR.n45 VPWR.n44 9.3005
R232 VPWR.n46 VPWR.n6 9.3005
R233 VPWR.n48 VPWR.n47 9.3005
R234 VPWR.n50 VPWR.n3 9.3005
R235 VPWR.n52 VPWR.n51 9.3005
R236 VPWR.n53 VPWR.n2 9.3005
R237 VPWR.n55 VPWR.n54 9.3005
R238 VPWR.n57 VPWR.n0 9.3005
R239 VPWR.n59 VPWR.n58 9.3005
R240 VPWR.n49 VPWR.n48 6.77697
R241 VPWR.n23 VPWR.n22 6.02403
R242 VPWR.n19 VPWR.n18 2.0514
R243 VPWR.n56 VPWR.n55 1.50638
R244 VPWR.n17 VPWR.n15 1.50638
R245 VPWR.n25 VPWR.n12 0.376971
R246 VPWR.n20 VPWR.n19 0.122949
R247 VPWR.n20 VPWR.n13 0.122949
R248 VPWR.n27 VPWR.n13 0.122949
R249 VPWR.n28 VPWR.n27 0.122949
R250 VPWR.n29 VPWR.n28 0.122949
R251 VPWR.n29 VPWR.n10 0.122949
R252 VPWR.n36 VPWR.n10 0.122949
R253 VPWR.n37 VPWR.n36 0.122949
R254 VPWR.n38 VPWR.n37 0.122949
R255 VPWR.n38 VPWR.n7 0.122949
R256 VPWR.n45 VPWR.n7 0.122949
R257 VPWR.n46 VPWR.n45 0.122949
R258 VPWR.n47 VPWR.n46 0.122949
R259 VPWR.n47 VPWR.n3 0.122949
R260 VPWR.n52 VPWR.n3 0.122949
R261 VPWR.n53 VPWR.n52 0.122949
R262 VPWR.n54 VPWR.n53 0.122949
R263 VPWR.n54 VPWR.n0 0.122949
R264 VPWR.n59 VPWR.n0 0.122949
R265 VPWR VPWR.n59 0.0617245
R266 VPB VPB.t21 257.93
R267 VPB.t12 VPB.t5 255.376
R268 VPB.t14 VPB.t15 255.376
R269 VPB.t1 VPB.t0 229.839
R270 VPB.t2 VPB.t1 229.839
R271 VPB.t3 VPB.t2 229.839
R272 VPB.t4 VPB.t3 229.839
R273 VPB.t5 VPB.t4 229.839
R274 VPB.t10 VPB.t12 229.839
R275 VPB.t9 VPB.t10 229.839
R276 VPB.t7 VPB.t9 229.839
R277 VPB.t6 VPB.t7 229.839
R278 VPB.t8 VPB.t6 229.839
R279 VPB.t20 VPB.t8 229.839
R280 VPB.t19 VPB.t20 229.839
R281 VPB.t18 VPB.t19 229.839
R282 VPB.t17 VPB.t18 229.839
R283 VPB.t16 VPB.t17 229.839
R284 VPB.t15 VPB.t16 229.839
R285 VPB.t13 VPB.t14 229.839
R286 VPB.t11 VPB.t13 229.839
R287 VPB.t21 VPB.t11 229.839
R288 A.n9 A.t7 227.538
R289 A.n0 A.t9 226.809
R290 A.n1 A.t1 226.809
R291 A.n18 A.t3 226.809
R292 A.n4 A.t4 226.809
R293 A.n6 A.t5 226.809
R294 A.n0 A.t0 197.475
R295 A.n9 A.t6 196.013
R296 A.n8 A.n7 196.013
R297 A.n5 A.t2 196.013
R298 A.n17 A.n3 196.013
R299 A.n2 A.t8 196.013
R300 A.n11 A.n10 162.121
R301 A.n24 A.n23 152
R302 A.n22 A.n21 152
R303 A.n20 A.n19 152
R304 A.n16 A.n15 152
R305 A.n14 A.n13 152
R306 A.n12 A.n11 152
R307 A.n23 A.n22 49.6611
R308 A.n13 A.n12 49.6611
R309 A.n10 A.n8 43.8187
R310 A.n19 A.n2 38.7066
R311 A.n16 A.n4 37.246
R312 A.n19 A.n18 21.1793
R313 A.n17 A.n16 20.449
R314 A.n10 A.n9 18.9884
R315 A.n23 A.n0 10.955
R316 A.n21 A.n20 10.1214
R317 A.n15 A 9.37724
R318 A.n14 A 9.07957
R319 A.n18 A.n17 8.03383
R320 A A.n24 7.5912
R321 A.n13 A.n5 7.30353
R322 A.n24 A 6.69817
R323 A.n2 A.n1 5.84292
R324 A A.n14 5.2098
R325 A.n22 A.n1 5.11262
R326 A.n5 A.n4 5.11262
R327 A.n15 A 4.91213
R328 A.n12 A.n6 3.65202
R329 A.n21 A 3.42376
R330 A.n8 A.n6 2.19141
R331 A.n11 A 1.04236
R332 A.n20 A 0.744686
C0 X VGND 1.21826f
C1 a_83_260# VPB 0.585055f
C2 a_83_260# A 0.667664f
C3 a_83_260# VPWR 0.959495f
C4 a_83_260# X 2.24501f
C5 VPB A 0.212026f
C6 VPB VPWR 0.293064f
C7 a_83_260# VGND 1.10591f
C8 VPB X 0.042225f
C9 A VPWR 0.125552f
C10 VPB VGND 0.008047f
C11 A X 0.001474f
C12 A VGND 0.1397f
C13 VPWR X 1.79026f
C14 VPWR VGND 0.089074f
C15 VGND VNB 1.29846f
C16 X VNB 0.073381f
C17 VPWR VNB 1.07018f
C18 A VNB 0.646991f
C19 VPB VNB 2.44181f
C20 a_83_260# VNB 1.69982f
C21 X.t22 VNB 0.048105f
C22 X.t6 VNB 0.015992f
C23 X.t4 VNB 0.015992f
C24 X.n0 VNB 0.034723f
C25 X.n1 VNB 0.116307f
C26 X.t16 VNB 0.050748f
C27 X.t3 VNB 0.015992f
C28 X.t1 VNB 0.015992f
C29 X.n2 VNB 0.034727f
C30 X.n3 VNB 0.126199f
C31 X.n4 VNB 0.073014f
C32 X.t27 VNB 0.009861f
C33 X.t20 VNB 0.009861f
C34 X.n5 VNB 0.041867f
C35 X.t0 VNB 0.015992f
C36 X.t2 VNB 0.015992f
C37 X.n6 VNB 0.034744f
C38 X.n7 VNB 0.121497f
C39 X.n8 VNB 0.043178f
C40 X.t18 VNB 0.009861f
C41 X.t29 VNB 0.009861f
C42 X.n9 VNB 0.049668f
C43 X.t14 VNB 0.015992f
C44 X.t13 VNB 0.015992f
C45 X.n10 VNB 0.034764f
C46 X.n11 VNB 0.113291f
C47 X.n12 VNB 0.044091f
C48 X.t24 VNB 0.009861f
C49 X.t28 VNB 0.009861f
C50 X.n13 VNB 0.041904f
C51 X.t12 VNB 0.015992f
C52 X.t11 VNB 0.015992f
C53 X.n14 VNB 0.034715f
C54 X.n15 VNB 0.088498f
C55 X.n16 VNB 0.043891f
C56 X.t23 VNB 0.009861f
C57 X.t25 VNB 0.009861f
C58 X.n17 VNB 0.041158f
C59 X.t10 VNB 0.015992f
C60 X.t9 VNB 0.015992f
C61 X.n18 VNB 0.034719f
C62 X.n19 VNB 0.105232f
C63 X.n20 VNB 0.044227f
C64 X.t21 VNB 0.009861f
C65 X.t17 VNB 0.009861f
C66 X.n21 VNB 0.040491f
C67 X.t8 VNB 0.015992f
C68 X.t7 VNB 0.015992f
C69 X.n22 VNB 0.034715f
C70 X.n23 VNB 0.100339f
C71 X.n24 VNB 0.044f
C72 X.t5 VNB 0.015992f
C73 X.t15 VNB 0.015992f
C74 X.n25 VNB 0.034715f
C75 X.t19 VNB 0.009861f
C76 X.t26 VNB 0.009861f
C77 X.n26 VNB 0.040491f
C78 X.n27 VNB 0.100339f
C79 X.n28 VNB 0.026267f
.ends

* NGSPICE file created from sky130_fd_sc_hs__bufbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__bufbuf_16 VNB VPB VPWR X VGND A
X0 X.t25 a_588_74.t12 VGND.t18 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 VPWR.t16 A.t0 a_27_368.t0 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t20 a_203_74.t6 a_588_74.t8 VPB.t20 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VPWR.t10 a_588_74.t13 X.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VGND.t22 a_203_74.t7 a_588_74.t9 VNB.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_588_74.t10 a_203_74.t8 VGND.t23 VNB.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X6 VPWR.t9 a_588_74.t14 X.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 X.t8 a_588_74.t15 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t24 a_588_74.t16 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X9 VGND.t16 a_588_74.t17 X.t23 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VGND.t1 A.t1 a_27_368.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 VGND.t24 a_203_74.t9 a_588_74.t11 VNB.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VGND.t15 a_588_74.t18 X.t22 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VGND.t14 a_588_74.t19 X.t21 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1332 pd=1.1 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VGND.t13 a_588_74.t20 X.t20 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VGND.t12 a_588_74.t21 X.t19 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VPWR.t7 a_588_74.t22 X.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X17 X.t6 a_588_74.t23 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_203_74.t5 a_27_368.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.10545 ps=1.025 w=0.74 l=0.15
X19 a_588_74.t0 a_203_74.t10 VGND.t19 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X20 a_203_74.t2 a_27_368.t3 VPWR.t19 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X21 X.t18 a_588_74.t24 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 X.t5 a_588_74.t25 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 VPWR.t18 a_27_368.t4 a_203_74.t1 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_203_74.t0 a_27_368.t5 VPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 a_203_74.t4 a_27_368.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 VGND.t10 a_588_74.t26 X.t17 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 X.t16 a_588_74.t27 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X28 VPWR.t11 a_203_74.t11 a_588_74.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X29 X.t4 a_588_74.t28 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X30 X.t15 a_588_74.t29 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 VGND.t7 a_588_74.t30 X.t14 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 X.t3 a_588_74.t31 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X33 a_588_74.t2 a_203_74.t12 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X34 X.t2 a_588_74.t32 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X35 VPWR.t13 a_203_74.t13 a_588_74.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X36 VPWR.t1 a_588_74.t33 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X37 VGND.t20 a_203_74.t14 a_588_74.t4 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X38 X.t13 a_588_74.t34 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X39 a_588_74.t5 a_203_74.t15 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X40 X.t0 a_588_74.t35 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X41 VGND.t3 a_27_368.t7 a_203_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1036 ps=1.02 w=0.74 l=0.15
X42 X.t12 a_588_74.t36 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X43 VGND.t4 a_588_74.t37 X.t11 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X44 a_588_74.t6 a_203_74.t16 VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X45 a_588_74.t7 a_203_74.t17 VGND.t21 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
R0 a_588_74.n54 a_588_74.n2 249.742
R1 a_588_74.n15 a_588_74.t22 242.875
R2 a_588_74.n17 a_588_74.t31 234.841
R3 a_588_74.n20 a_588_74.t33 234.841
R4 a_588_74.n18 a_588_74.t35 234.841
R5 a_588_74.n23 a_588_74.t14 234.841
R6 a_588_74.n25 a_588_74.t15 234.841
R7 a_588_74.n28 a_588_74.n12 234.841
R8 a_588_74.n30 a_588_74.t23 234.841
R9 a_588_74.n35 a_588_74.n32 234.841
R10 a_588_74.n33 a_588_74.t25 234.841
R11 a_588_74.n38 a_588_74.n10 234.841
R12 a_588_74.n40 a_588_74.t28 234.841
R13 a_588_74.n43 a_588_74.n9 234.841
R14 a_588_74.n45 a_588_74.t32 234.841
R15 a_588_74.n50 a_588_74.t13 234.841
R16 a_588_74.n48 a_588_74.n47 234.841
R17 a_588_74.n53 a_588_74.n3 206.823
R18 a_588_74.n55 a_588_74.n54 206.822
R19 a_588_74.n48 a_588_74.t34 188.565
R20 a_588_74.n49 a_588_74.t37 186.374
R21 a_588_74.n46 a_588_74.t29 186.374
R22 a_588_74.n44 a_588_74.t20 186.374
R23 a_588_74.n41 a_588_74.t24 186.374
R24 a_588_74.n39 a_588_74.t18 186.374
R25 a_588_74.n11 a_588_74.t12 186.374
R26 a_588_74.n34 a_588_74.t17 186.374
R27 a_588_74.n31 a_588_74.t36 186.374
R28 a_588_74.n29 a_588_74.t26 186.374
R29 a_588_74.n26 a_588_74.t27 186.374
R30 a_588_74.n24 a_588_74.t21 186.374
R31 a_588_74.n13 a_588_74.t16 186.374
R32 a_588_74.n19 a_588_74.t19 186.374
R33 a_588_74.n16 a_588_74.n14 186.374
R34 a_588_74.n15 a_588_74.t30 186.374
R35 a_588_74.n37 a_588_74.n1 169.994
R36 a_588_74.n42 a_588_74.n1 169.994
R37 a_588_74.n0 a_588_74.n36 169.111
R38 a_588_74.n1 a_588_74.n51 168.732
R39 a_588_74.n27 a_588_74.n0 168.389
R40 a_588_74.n0 a_588_74.n21 167.637
R41 a_588_74.n22 a_588_74.n0 167.445
R42 a_588_74.n7 a_588_74.n5 154.244
R43 a_588_74.n7 a_588_74.n6 103.043
R44 a_588_74.n8 a_588_74.n4 98.6918
R45 a_588_74.n16 a_588_74.n15 62.8066
R46 a_588_74.n49 a_588_74.n48 60.6157
R47 a_588_74.n8 a_588_74.n7 60.6123
R48 a_588_74.n19 a_588_74.n18 59.155
R49 a_588_74.n25 a_588_74.n24 54.7732
R50 a_588_74.n30 a_588_74.n29 50.3914
R51 a_588_74.n45 a_588_74.n44 47.4702
R52 a_588_74.n34 a_588_74.n33 46.0096
R53 a_588_74.n54 a_588_74.n53 43.6711
R54 a_588_74.n40 a_588_74.n39 41.6278
R55 a_588_74.n27 a_588_74.n26 40.8975
R56 a_588_74.n21 a_588_74.n17 38.7066
R57 a_588_74.n22 a_588_74.n13 38.7066
R58 a_588_74.n36 a_588_74.n31 37.9763
R59 a_588_74.n37 a_588_74.n11 36.5157
R60 a_588_74.n51 a_588_74.n46 34.3247
R61 a_588_74.n42 a_588_74.n41 32.1338
R62 a_588_74.n21 a_588_74.n20 27.0217
R63 a_588_74.n3 a_588_74.t8 26.3844
R64 a_588_74.n3 a_588_74.t6 26.3844
R65 a_588_74.n2 a_588_74.t3 26.3844
R66 a_588_74.n2 a_588_74.t5 26.3844
R67 a_588_74.t1 a_588_74.n55 26.3844
R68 a_588_74.n55 a_588_74.t2 26.3844
R69 a_588_74.n39 a_588_74.n38 24.1005
R70 a_588_74.n23 a_588_74.n22 23.3702
R71 a_588_74.n51 a_588_74.n50 23.3702
R72 a_588_74.n5 a_588_74.t4 22.7032
R73 a_588_74.n5 a_588_74.t10 22.7032
R74 a_588_74.n6 a_588_74.t11 22.7032
R75 a_588_74.n6 a_588_74.t0 22.7032
R76 a_588_74.n4 a_588_74.t9 22.7032
R77 a_588_74.n4 a_588_74.t7 22.7032
R78 a_588_74.n52 a_588_74.n8 21.9025
R79 a_588_74.n41 a_588_74.n40 21.1793
R80 a_588_74.n35 a_588_74.n34 19.7187
R81 a_588_74.n44 a_588_74.n43 18.2581
R82 a_588_74.n28 a_588_74.n27 16.7975
R83 a_588_74.n33 a_588_74.n11 16.7975
R84 a_588_74.n29 a_588_74.n28 15.3369
R85 a_588_74.n36 a_588_74.n35 15.3369
R86 a_588_74.n46 a_588_74.n45 15.3369
R87 a_588_74.n31 a_588_74.n30 12.4157
R88 a_588_74.n38 a_588_74.n37 12.4157
R89 a_588_74.n43 a_588_74.n42 12.4157
R90 a_588_74.n24 a_588_74.n23 10.955
R91 a_588_74.n52 a_588_74.n1 9.81409
R92 a_588_74.n53 a_588_74.n52 8.89504
R93 a_588_74.n26 a_588_74.n25 8.03383
R94 a_588_74.n20 a_588_74.n19 6.57323
R95 a_588_74.n50 a_588_74.n49 5.11262
R96 a_588_74.n18 a_588_74.n13 3.65202
R97 a_588_74.n1 a_588_74.n0 2.47333
R98 a_588_74.n17 a_588_74.n16 2.19141
R99 VGND.n57 VGND.n56 217
R100 VGND.n45 VGND.n44 210.018
R101 VGND.n49 VGND.n4 210.018
R102 VGND.n60 VGND.n59 209.243
R103 VGND.n15 VGND.t7 161.441
R104 VGND.n51 VGND.t23 154.727
R105 VGND.n14 VGND.t14 154.2
R106 VGND.n42 VGND.n41 140.118
R107 VGND.n33 VGND.n32 129.406
R108 VGND.n35 VGND.n34 124.29
R109 VGND.n9 VGND.n8 122.508
R110 VGND.n26 VGND.n25 119.483
R111 VGND.n12 VGND.n11 118.189
R112 VGND.n19 VGND.n18 116.644
R113 VGND.n36 VGND.n33 36.1417
R114 VGND.n40 VGND.n6 36.1417
R115 VGND.n55 VGND.n1 36.1417
R116 VGND.n18 VGND.t17 34.0546
R117 VGND.n11 VGND.t9 34.0546
R118 VGND.n25 VGND.t5 34.0546
R119 VGND.n8 VGND.t18 34.0546
R120 VGND.n44 VGND.t21 34.0546
R121 VGND.n4 VGND.t19 34.0546
R122 VGND.n45 VGND.n43 32.7534
R123 VGND.n31 VGND.n9 30.8711
R124 VGND.n49 VGND.n3 30.4946
R125 VGND.n19 VGND.n17 28.2358
R126 VGND.n51 VGND.n50 28.2358
R127 VGND.n27 VGND.n26 26.3534
R128 VGND.n20 VGND.n12 25.977
R129 VGND.n26 VGND.n24 23.7181
R130 VGND.n56 VGND.t0 23.514
R131 VGND.n60 VGND.n58 23.3417
R132 VGND.n24 VGND.n12 22.9652
R133 VGND.n18 VGND.t12 22.7032
R134 VGND.n11 VGND.t10 22.7032
R135 VGND.n25 VGND.t16 22.7032
R136 VGND.n8 VGND.t15 22.7032
R137 VGND.n32 VGND.t11 22.7032
R138 VGND.n32 VGND.t13 22.7032
R139 VGND.n34 VGND.t8 22.7032
R140 VGND.n34 VGND.t4 22.7032
R141 VGND.n41 VGND.t6 22.7032
R142 VGND.n41 VGND.t22 22.7032
R143 VGND.n44 VGND.t24 22.7032
R144 VGND.n4 VGND.t20 22.7032
R145 VGND.n56 VGND.t3 22.7032
R146 VGND.n59 VGND.t2 22.7032
R147 VGND.n59 VGND.t1 22.7032
R148 VGND.n27 VGND.n9 21.4593
R149 VGND.n33 VGND.n31 19.9534
R150 VGND.n20 VGND.n19 19.2005
R151 VGND.n51 VGND.n1 19.2005
R152 VGND.n43 VGND.n42 17.6946
R153 VGND.n17 VGND.n14 16.9417
R154 VGND.n50 VGND.n49 16.9417
R155 VGND.n58 VGND.n57 16.5652
R156 VGND.n45 VGND.n3 14.6829
R157 VGND.n36 VGND.n35 12.424
R158 VGND.n58 VGND.n0 9.3005
R159 VGND.n55 VGND.n54 9.3005
R160 VGND.n53 VGND.n1 9.3005
R161 VGND.n52 VGND.n51 9.3005
R162 VGND.n17 VGND.n16 9.3005
R163 VGND.n19 VGND.n13 9.3005
R164 VGND.n21 VGND.n20 9.3005
R165 VGND.n22 VGND.n12 9.3005
R166 VGND.n24 VGND.n23 9.3005
R167 VGND.n26 VGND.n10 9.3005
R168 VGND.n28 VGND.n27 9.3005
R169 VGND.n29 VGND.n9 9.3005
R170 VGND.n31 VGND.n30 9.3005
R171 VGND.n33 VGND.n7 9.3005
R172 VGND.n37 VGND.n36 9.3005
R173 VGND.n38 VGND.n6 9.3005
R174 VGND.n40 VGND.n39 9.3005
R175 VGND.n43 VGND.n5 9.3005
R176 VGND.n46 VGND.n45 9.3005
R177 VGND.n47 VGND.n3 9.3005
R178 VGND.n49 VGND.n48 9.3005
R179 VGND.n50 VGND.n2 9.3005
R180 VGND.n61 VGND.n60 7.25439
R181 VGND.n15 VGND.n14 6.99787
R182 VGND.n35 VGND.n6 4.89462
R183 VGND.n42 VGND.n40 4.89462
R184 VGND.n57 VGND.n55 0.753441
R185 VGND.n16 VGND.n15 0.587308
R186 VGND VGND.n61 0.157727
R187 VGND.n61 VGND.n0 0.150046
R188 VGND.n16 VGND.n13 0.122949
R189 VGND.n21 VGND.n13 0.122949
R190 VGND.n22 VGND.n21 0.122949
R191 VGND.n23 VGND.n22 0.122949
R192 VGND.n23 VGND.n10 0.122949
R193 VGND.n28 VGND.n10 0.122949
R194 VGND.n29 VGND.n28 0.122949
R195 VGND.n30 VGND.n29 0.122949
R196 VGND.n30 VGND.n7 0.122949
R197 VGND.n37 VGND.n7 0.122949
R198 VGND.n38 VGND.n37 0.122949
R199 VGND.n39 VGND.n38 0.122949
R200 VGND.n39 VGND.n5 0.122949
R201 VGND.n46 VGND.n5 0.122949
R202 VGND.n47 VGND.n46 0.122949
R203 VGND.n48 VGND.n47 0.122949
R204 VGND.n48 VGND.n2 0.122949
R205 VGND.n52 VGND.n2 0.122949
R206 VGND.n53 VGND.n52 0.122949
R207 VGND.n54 VGND.n53 0.122949
R208 VGND.n54 VGND.n0 0.122949
R209 X.n23 X.t10 229.06
R210 X.n20 X.t2 229.016
R211 X.n17 X.t4 229.016
R212 X.n14 X.t5 229.016
R213 X.n11 X.t6 229.016
R214 X.n8 X.n7 202.631
R215 X.n4 X.n3 202.631
R216 X.n1 X.n0 202.409
R217 X.n1 X.t14 191.03
R218 X.n4 X.n2 159.66
R219 X.n20 X.n19 158.202
R220 X.n8 X.n6 155.733
R221 X.n11 X.n10 155.107
R222 X.n17 X.n16 151.246
R223 X.n14 X.n13 151.246
R224 X.n23 X.n22 151.058
R225 X.n0 X.t3 35.1791
R226 X.n7 X.t9 26.3844
R227 X.n7 X.t8 26.3844
R228 X.n3 X.t1 26.3844
R229 X.n3 X.t0 26.3844
R230 X.n0 X.t7 26.3844
R231 X.n22 X.t11 22.7032
R232 X.n22 X.t13 22.7032
R233 X.n19 X.t20 22.7032
R234 X.n19 X.t15 22.7032
R235 X.n16 X.t22 22.7032
R236 X.n16 X.t18 22.7032
R237 X.n13 X.t23 22.7032
R238 X.n13 X.t25 22.7032
R239 X.n10 X.t17 22.7032
R240 X.n10 X.t12 22.7032
R241 X.n6 X.t19 22.7032
R242 X.n6 X.t16 22.7032
R243 X.n2 X.t21 22.7032
R244 X.n2 X.t24 22.7032
R245 X.n5 X.n1 10.5462
R246 X.n21 X.n20 9.70406
R247 X.n18 X.n17 9.70406
R248 X.n15 X.n14 9.70406
R249 X.n12 X.n11 9.70406
R250 X.n9 X.n8 9.70406
R251 X.n5 X.n4 9.70406
R252 X.n24 X.n23 9.63695
R253 X.n15 X.n12 0.5005
R254 X.n21 X.n18 0.5005
R255 X.n24 X.n21 0.497783
R256 X.n9 X.n5 0.48963
R257 X.n12 X.n9 0.484196
R258 X.n18 X.n15 0.484196
R259 X X.n24 0.0793043
R260 VNB.t0 VNB.t23 2448.29
R261 VNB.t14 VNB.t7 2171.13
R262 VNB VNB.t1 1177.95
R263 VNB.t12 VNB.t17 1154.86
R264 VNB.t10 VNB.t9 1154.86
R265 VNB.t16 VNB.t5 1154.86
R266 VNB.t15 VNB.t18 1154.86
R267 VNB.t24 VNB.t21 1154.86
R268 VNB.t20 VNB.t19 1154.86
R269 VNB.t3 VNB.t0 1004.72
R270 VNB.t17 VNB.t14 993.177
R271 VNB.t9 VNB.t12 993.177
R272 VNB.t5 VNB.t10 993.177
R273 VNB.t18 VNB.t16 993.177
R274 VNB.t11 VNB.t15 993.177
R275 VNB.t13 VNB.t11 993.177
R276 VNB.t8 VNB.t13 993.177
R277 VNB.t4 VNB.t8 993.177
R278 VNB.t6 VNB.t4 993.177
R279 VNB.t22 VNB.t6 993.177
R280 VNB.t21 VNB.t22 993.177
R281 VNB.t19 VNB.t24 993.177
R282 VNB.t23 VNB.t20 993.177
R283 VNB.t2 VNB.t3 993.177
R284 VNB.t1 VNB.t2 993.177
R285 A.n0 A.t0 259.132
R286 A.n0 A.t1 198.882
R287 A A.n0 156.934
R288 a_27_368.t0 a_27_368.n8 279.683
R289 a_27_368.n1 a_27_368.t3 247.5
R290 a_27_368.n3 a_27_368.t4 240.197
R291 a_27_368.n5 a_27_368.t5 240.197
R292 a_27_368.n8 a_27_368.t1 190.91
R293 a_27_368.n5 a_27_368.t6 182.138
R294 a_27_368.n4 a_27_368.t7 179.947
R295 a_27_368.n1 a_27_368.t2 179.947
R296 a_27_368.n2 a_27_368.n0 165.189
R297 a_27_368.n7 a_27_368.n6 152
R298 a_27_368.n4 a_27_368.n0 152
R299 a_27_368.n6 a_27_368.n4 49.6611
R300 a_27_368.n3 a_27_368.n2 44.549
R301 a_27_368.n2 a_27_368.n1 13.8763
R302 a_27_368.n7 a_27_368.n0 13.1884
R303 a_27_368.n6 a_27_368.n5 10.955
R304 a_27_368.n8 a_27_368.n7 10.4732
R305 a_27_368.n4 a_27_368.n3 5.11262
R306 VPWR.n36 VPWR.t4 360.204
R307 VPWR.n61 VPWR.n2 334.173
R308 VPWR.n54 VPWR.n5 333.82
R309 VPWR.n48 VPWR.n47 333.82
R310 VPWR.n63 VPWR.n1 331.5
R311 VPWR.n39 VPWR.n38 325.01
R312 VPWR.n45 VPWR.t20 268.825
R313 VPWR.n30 VPWR.t5 268.825
R314 VPWR.n28 VPWR.t6 268.825
R315 VPWR.n22 VPWR.t8 268.825
R316 VPWR.n17 VPWR.t7 266.204
R317 VPWR.n56 VPWR.t14 259.171
R318 VPWR.n20 VPWR.n14 242.44
R319 VPWR.n16 VPWR.n15 231.752
R320 VPWR.n60 VPWR.n3 36.1417
R321 VPWR.n44 VPWR.n8 36.1417
R322 VPWR.n49 VPWR.n46 36.1417
R323 VPWR.n53 VPWR.n6 36.1417
R324 VPWR.n23 VPWR.n21 36.1417
R325 VPWR.n27 VPWR.n12 36.1417
R326 VPWR.n31 VPWR.n29 36.1417
R327 VPWR.n35 VPWR.n10 36.1417
R328 VPWR.n40 VPWR.n37 36.1417
R329 VPWR.n63 VPWR.n62 35.3887
R330 VPWR.n38 VPWR.t10 35.1791
R331 VPWR.n20 VPWR.n19 34.2593
R332 VPWR.n55 VPWR.n54 32.7534
R333 VPWR.n62 VPWR.n61 32.377
R334 VPWR.n23 VPWR.n22 29.7417
R335 VPWR.n56 VPWR.n55 28.6123
R336 VPWR.n48 VPWR.n6 28.2358
R337 VPWR.n47 VPWR.t15 28.1434
R338 VPWR.n19 VPWR.n16 27.1064
R339 VPWR.n1 VPWR.t17 26.3844
R340 VPWR.n1 VPWR.t16 26.3844
R341 VPWR.n2 VPWR.t19 26.3844
R342 VPWR.n2 VPWR.t18 26.3844
R343 VPWR.n5 VPWR.t12 26.3844
R344 VPWR.n5 VPWR.t13 26.3844
R345 VPWR.n47 VPWR.t11 26.3844
R346 VPWR.n38 VPWR.t2 26.3844
R347 VPWR.n14 VPWR.t0 26.3844
R348 VPWR.n14 VPWR.t9 26.3844
R349 VPWR.n15 VPWR.t3 26.3844
R350 VPWR.n15 VPWR.t1 26.3844
R351 VPWR.n28 VPWR.n27 25.224
R352 VPWR.n56 VPWR.n3 24.8476
R353 VPWR.n46 VPWR.n45 24.4711
R354 VPWR.n31 VPWR.n30 20.7064
R355 VPWR.n37 VPWR.n36 19.9534
R356 VPWR.n36 VPWR.n35 16.1887
R357 VPWR.n30 VPWR.n10 15.4358
R358 VPWR.n39 VPWR.n8 12.0476
R359 VPWR.n45 VPWR.n44 11.6711
R360 VPWR.n29 VPWR.n28 10.9181
R361 VPWR.n19 VPWR.n18 9.3005
R362 VPWR.n21 VPWR.n13 9.3005
R363 VPWR.n24 VPWR.n23 9.3005
R364 VPWR.n25 VPWR.n12 9.3005
R365 VPWR.n27 VPWR.n26 9.3005
R366 VPWR.n29 VPWR.n11 9.3005
R367 VPWR.n32 VPWR.n31 9.3005
R368 VPWR.n33 VPWR.n10 9.3005
R369 VPWR.n35 VPWR.n34 9.3005
R370 VPWR.n37 VPWR.n9 9.3005
R371 VPWR.n41 VPWR.n40 9.3005
R372 VPWR.n42 VPWR.n8 9.3005
R373 VPWR.n44 VPWR.n43 9.3005
R374 VPWR.n46 VPWR.n7 9.3005
R375 VPWR.n50 VPWR.n49 9.3005
R376 VPWR.n51 VPWR.n6 9.3005
R377 VPWR.n53 VPWR.n52 9.3005
R378 VPWR.n55 VPWR.n4 9.3005
R379 VPWR.n57 VPWR.n56 9.3005
R380 VPWR.n58 VPWR.n3 9.3005
R381 VPWR.n60 VPWR.n59 9.3005
R382 VPWR.n62 VPWR.n0 9.3005
R383 VPWR.n64 VPWR.n63 8.45673
R384 VPWR.n49 VPWR.n48 7.90638
R385 VPWR.n17 VPWR.n16 6.85153
R386 VPWR.n22 VPWR.n12 6.4005
R387 VPWR.n40 VPWR.n39 5.27109
R388 VPWR.n61 VPWR.n60 3.76521
R389 VPWR.n54 VPWR.n53 3.38874
R390 VPWR.n21 VPWR.n20 1.88285
R391 VPWR.n18 VPWR.n17 0.568865
R392 VPWR VPWR.n64 0.163644
R393 VPWR.n64 VPWR.n0 0.144205
R394 VPWR.n18 VPWR.n13 0.122949
R395 VPWR.n24 VPWR.n13 0.122949
R396 VPWR.n25 VPWR.n24 0.122949
R397 VPWR.n26 VPWR.n25 0.122949
R398 VPWR.n26 VPWR.n11 0.122949
R399 VPWR.n32 VPWR.n11 0.122949
R400 VPWR.n33 VPWR.n32 0.122949
R401 VPWR.n34 VPWR.n33 0.122949
R402 VPWR.n34 VPWR.n9 0.122949
R403 VPWR.n41 VPWR.n9 0.122949
R404 VPWR.n42 VPWR.n41 0.122949
R405 VPWR.n43 VPWR.n42 0.122949
R406 VPWR.n43 VPWR.n7 0.122949
R407 VPWR.n50 VPWR.n7 0.122949
R408 VPWR.n51 VPWR.n50 0.122949
R409 VPWR.n52 VPWR.n51 0.122949
R410 VPWR.n52 VPWR.n4 0.122949
R411 VPWR.n57 VPWR.n4 0.122949
R412 VPWR.n58 VPWR.n57 0.122949
R413 VPWR.n59 VPWR.n58 0.122949
R414 VPWR.n59 VPWR.n0 0.122949
R415 VPB.t19 VPB.t14 523.521
R416 VPB.t20 VPB.t10 464.786
R417 VPB.t6 VPB.t8 459.678
R418 VPB.t5 VPB.t6 459.678
R419 VPB.t4 VPB.t5 459.678
R420 VPB.t2 VPB.t4 459.678
R421 VPB VPB.t16 257.93
R422 VPB.t3 VPB.t7 255.376
R423 VPB.t10 VPB.t2 255.376
R424 VPB.t11 VPB.t15 234.946
R425 VPB.t1 VPB.t3 229.839
R426 VPB.t0 VPB.t1 229.839
R427 VPB.t9 VPB.t0 229.839
R428 VPB.t8 VPB.t9 229.839
R429 VPB.t15 VPB.t20 229.839
R430 VPB.t12 VPB.t11 229.839
R431 VPB.t13 VPB.t12 229.839
R432 VPB.t14 VPB.t13 229.839
R433 VPB.t18 VPB.t19 229.839
R434 VPB.t17 VPB.t18 229.839
R435 VPB.t16 VPB.t17 229.839
R436 a_203_74.n22 a_203_74.n0 250.518
R437 a_203_74.n3 a_203_74.t6 234.841
R438 a_203_74.n5 a_203_74.t16 234.841
R439 a_203_74.n7 a_203_74.t11 234.841
R440 a_203_74.n2 a_203_74.t12 234.841
R441 a_203_74.n14 a_203_74.t13 234.841
R442 a_203_74.n16 a_203_74.t15 234.841
R443 a_203_74.t2 a_203_74.n22 233.983
R444 a_203_74.n16 a_203_74.t8 188.565
R445 a_203_74.n3 a_203_74.t7 188.565
R446 a_203_74.n15 a_203_74.t14 186.374
R447 a_203_74.n9 a_203_74.t10 186.374
R448 a_203_74.n8 a_203_74.t9 186.374
R449 a_203_74.n4 a_203_74.t17 186.374
R450 a_203_74.n11 a_203_74.n6 165.189
R451 a_203_74.n20 a_203_74.n19 152.887
R452 a_203_74.n18 a_203_74.n17 152
R453 a_203_74.n15 a_203_74.n1 152
R454 a_203_74.n13 a_203_74.n12 152
R455 a_203_74.n11 a_203_74.n10 152
R456 a_203_74.n20 a_203_74.t5 146.603
R457 a_203_74.n4 a_203_74.n3 60.6157
R458 a_203_74.n6 a_203_74.n5 54.7732
R459 a_203_74.n17 a_203_74.n15 49.6611
R460 a_203_74.n14 a_203_74.n13 44.549
R461 a_203_74.n10 a_203_74.n8 36.5157
R462 a_203_74.n21 a_203_74.n18 31.4187
R463 a_203_74.n0 a_203_74.t1 26.3844
R464 a_203_74.n0 a_203_74.t0 26.3844
R465 a_203_74.n10 a_203_74.n9 26.2914
R466 a_203_74.n19 a_203_74.t3 22.7032
R467 a_203_74.n19 a_203_74.t4 22.7032
R468 a_203_74.n13 a_203_74.n2 21.1793
R469 a_203_74.n21 a_203_74.n20 17.9104
R470 a_203_74.n12 a_203_74.n11 13.1884
R471 a_203_74.n12 a_203_74.n1 13.1884
R472 a_203_74.n18 a_203_74.n1 13.1884
R473 a_203_74.n22 a_203_74.n21 12.8975
R474 a_203_74.n7 a_203_74.n6 12.4157
R475 a_203_74.n17 a_203_74.n16 10.955
R476 a_203_74.n5 a_203_74.n4 5.11262
R477 a_203_74.n15 a_203_74.n14 5.11262
R478 a_203_74.n9 a_203_74.n2 2.19141
R479 a_203_74.n8 a_203_74.n7 0.730803
C0 VPB A 0.0398f
C1 VPB VPWR 0.364852f
C2 VPB X 0.048826f
C3 A VPWR 0.015092f
C4 VPB VGND 0.014386f
C5 A X 1.01e-20
C6 VPWR X 1.99879f
C7 A VGND 0.01733f
C8 VPWR VGND 0.125633f
C9 X VGND 1.27215f
C10 VGND VNB 1.51429f
C11 X VNB 0.071257f
C12 VPWR VNB 1.22322f
C13 A VNB 0.162747f
C14 VPB VNB 2.97749f
C15 X.t14 VNB 0.046494f
C16 X.t7 VNB 0.014782f
C17 X.t3 VNB 0.01971f
C18 X.n0 VNB 0.037063f
C19 X.n1 VNB 0.130662f
C20 X.t21 VNB 0.009116f
C21 X.t24 VNB 0.009116f
C22 X.n2 VNB 0.035693f
C23 X.t1 VNB 0.014782f
C24 X.t0 VNB 0.014782f
C25 X.n3 VNB 0.032136f
C26 X.n4 VNB 0.09871f
C27 X.n5 VNB 0.067517f
C28 X.t19 VNB 0.009116f
C29 X.t16 VNB 0.009116f
C30 X.n6 VNB 0.0381f
C31 X.t9 VNB 0.014782f
C32 X.t8 VNB 0.014782f
C33 X.n7 VNB 0.032136f
C34 X.n8 VNB 0.102889f
C35 X.n9 VNB 0.038437f
C36 X.t17 VNB 0.009116f
C37 X.t12 VNB 0.009116f
C38 X.n10 VNB 0.039312f
C39 X.t6 VNB 0.056295f
C40 X.n11 VNB 0.109797f
C41 X.n12 VNB 0.038842f
C42 X.t23 VNB 0.009116f
C43 X.t25 VNB 0.009116f
C44 X.n13 VNB 0.040964f
C45 X.t5 VNB 0.056295f
C46 X.n14 VNB 0.115008f
C47 X.n15 VNB 0.038842f
C48 X.t22 VNB 0.009116f
C49 X.t18 VNB 0.009116f
C50 X.n16 VNB 0.040964f
C51 X.t4 VNB 0.056295f
C52 X.n17 VNB 0.115008f
C53 X.n18 VNB 0.038842f
C54 X.t20 VNB 0.009116f
C55 X.t15 VNB 0.009116f
C56 X.n19 VNB 0.038189f
C57 X.t2 VNB 0.056295f
C58 X.n20 VNB 0.106344f
C59 X.n21 VNB 0.039347f
C60 X.t10 VNB 0.056296f
C61 X.t11 VNB 0.009116f
C62 X.t13 VNB 0.009116f
C63 X.n22 VNB 0.037041f
C64 X.n23 VNB 0.112712f
C65 X.n24 VNB 0.023303f
C66 a_588_74.n0 VNB 0.202114f
C67 a_588_74.n1 VNB 0.165932f
C68 a_588_74.t2 VNB 0.012782f
C69 a_588_74.t3 VNB 0.012782f
C70 a_588_74.t5 VNB 0.012782f
C71 a_588_74.n2 VNB 0.039535f
C72 a_588_74.t8 VNB 0.012782f
C73 a_588_74.t6 VNB 0.012782f
C74 a_588_74.n3 VNB 0.028817f
C75 a_588_74.t9 VNB 0.007882f
C76 a_588_74.t7 VNB 0.007882f
C77 a_588_74.n4 VNB 0.017579f
C78 a_588_74.t4 VNB 0.007882f
C79 a_588_74.t10 VNB 0.007882f
C80 a_588_74.n5 VNB 0.030668f
C81 a_588_74.t11 VNB 0.007882f
C82 a_588_74.t0 VNB 0.007882f
C83 a_588_74.n6 VNB 0.018583f
C84 a_588_74.n7 VNB 0.071145f
C85 a_588_74.n8 VNB 0.045747f
C86 a_588_74.t29 VNB 0.012097f
C87 a_588_74.t32 VNB 0.018218f
C88 a_588_74.t20 VNB 0.012097f
C89 a_588_74.n9 VNB 0.018218f
C90 a_588_74.t24 VNB 0.012097f
C91 a_588_74.t28 VNB 0.018218f
C92 a_588_74.t18 VNB 0.012097f
C93 a_588_74.n10 VNB 0.018218f
C94 a_588_74.t12 VNB 0.012097f
C95 a_588_74.n11 VNB 0.015783f
C96 a_588_74.t36 VNB 0.012097f
C97 a_588_74.t23 VNB 0.018218f
C98 a_588_74.t26 VNB 0.012097f
C99 a_588_74.n12 VNB 0.018218f
C100 a_588_74.t27 VNB 0.012097f
C101 a_588_74.t15 VNB 0.018218f
C102 a_588_74.t21 VNB 0.012097f
C103 a_588_74.t14 VNB 0.018218f
C104 a_588_74.t16 VNB 0.012097f
C105 a_588_74.n13 VNB 0.0139f
C106 a_588_74.t31 VNB 0.018218f
C107 a_588_74.n14 VNB 0.012097f
C108 a_588_74.t30 VNB 0.012097f
C109 a_588_74.t22 VNB 0.018719f
C110 a_588_74.n15 VNB 0.033435f
C111 a_588_74.n16 VNB 0.017792f
C112 a_588_74.n17 VNB 0.01627f
C113 a_588_74.t33 VNB 0.018218f
C114 a_588_74.t19 VNB 0.012097f
C115 a_588_74.t35 VNB 0.018218f
C116 a_588_74.n18 VNB 0.020036f
C117 a_588_74.n19 VNB 0.017917f
C118 a_588_74.n20 VNB 0.015014f
C119 a_588_74.n21 VNB 0.013407f
C120 a_588_74.n22 VNB 0.012567f
C121 a_588_74.n23 VNB 0.01514f
C122 a_588_74.n24 VNB 0.017917f
C123 a_588_74.n25 VNB 0.020036f
C124 a_588_74.n26 VNB 0.01503f
C125 a_588_74.n27 VNB 0.011623f
C126 a_588_74.n28 VNB 0.014763f
C127 a_588_74.n29 VNB 0.017917f
C128 a_588_74.n30 VNB 0.020036f
C129 a_588_74.n31 VNB 0.015281f
C130 a_588_74.n32 VNB 0.018218f
C131 a_588_74.t17 VNB 0.012097f
C132 a_588_74.t25 VNB 0.018218f
C133 a_588_74.n33 VNB 0.020036f
C134 a_588_74.n34 VNB 0.017917f
C135 a_588_74.n35 VNB 0.015266f
C136 a_588_74.n36 VNB 0.010754f
C137 a_588_74.n37 VNB 0.009885f
C138 a_588_74.n38 VNB 0.015516f
C139 a_588_74.n39 VNB 0.017917f
C140 a_588_74.n40 VNB 0.020036f
C141 a_588_74.n41 VNB 0.015783f
C142 a_588_74.n42 VNB 0.009132f
C143 a_588_74.n43 VNB 0.014512f
C144 a_588_74.n44 VNB 0.017917f
C145 a_588_74.n45 VNB 0.020036f
C146 a_588_74.n46 VNB 0.015156f
C147 a_588_74.t13 VNB 0.018218f
C148 a_588_74.t37 VNB 0.012097f
C149 a_588_74.n47 VNB 0.018218f
C150 a_588_74.t34 VNB 0.012222f
C151 a_588_74.n48 VNB 0.030672f
C152 a_588_74.n49 VNB 0.017917f
C153 a_588_74.n50 VNB 0.014136f
C154 a_588_74.n51 VNB 0.011565f
C155 a_588_74.n52 VNB 0.038286f
C156 a_588_74.n53 VNB 0.06359f
C157 a_588_74.n54 VNB 0.121518f
C158 a_588_74.n55 VNB 0.028817f
C159 a_588_74.t1 VNB 0.012782f
.ends

* NGSPICE file created from sky130_fd_sc_hs__bufinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__bufinv_16 VNB VPB VPWR Y VGND A
X0 VGND.t20 A.t0 a_27_74.t2 VNB.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 Y.t24 a_384_74.t12 VGND.t21 VNB.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2 VPWR.t9 a_384_74.t13 Y.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1904 ps=1.46 w=1.12 l=0.15
X3 a_384_74.t11 a_27_74.t6 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 Y.t23 a_384_74.t14 VGND.t22 VNB.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 Y.t8 a_384_74.t15 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t15 a_27_74.t7 a_384_74.t5 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VPWR.t18 A.t1 a_27_74.t5 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8 a_384_74.t4 a_27_74.t8 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t22 a_384_74.t16 VGND.t23 VNB.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X10 VPWR.t13 a_27_74.t9 a_384_74.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VGND.t16 a_27_74.t10 a_384_74.t10 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 Y.t7 a_384_74.t17 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X13 VGND.t19 A.t2 a_27_74.t1 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.1258 pd=1.08 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 a_384_74.t2 a_27_74.t11 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 VGND.t15 a_27_74.t12 a_384_74.t9 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 Y.t21 a_384_74.t18 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t1 a_384_74.t19 Y.t20 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VPWR.t11 a_27_74.t13 a_384_74.t1 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X19 VPWR.t6 a_384_74.t20 Y.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X20 VGND.t14 a_27_74.t14 a_384_74.t8 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VGND.t2 a_384_74.t21 Y.t19 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 VGND.t3 a_384_74.t22 Y.t18 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 VPWR.t5 a_384_74.t23 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_384_74.t7 a_27_74.t15 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 Y.t17 a_384_74.t24 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X26 VPWR.t4 a_384_74.t25 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 Y.t3 a_384_74.t26 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.1736 ps=1.43 w=1.12 l=0.15
X28 Y.t16 a_384_74.t27 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X29 a_384_74.t0 a_27_74.t16 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_384_74.t6 a_27_74.t17 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 VGND.t6 a_384_74.t28 Y.t15 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 VPWR.t17 A.t3 a_27_74.t4 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X33 VPWR.t2 a_384_74.t29 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X34 VGND.t7 a_384_74.t30 Y.t14 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X35 Y.t13 a_384_74.t31 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X36 a_27_74.t3 A.t4 VPWR.t16 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X37 VPWR.t1 a_384_74.t32 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X38 a_27_74.t0 A.t5 VGND.t18 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1258 ps=1.08 w=0.74 l=0.15
X39 VPWR.t0 a_384_74.t33 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X40 VGND.t9 a_384_74.t34 Y.t12 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X41 VGND.t10 a_384_74.t35 Y.t11 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X42 VGND.t11 a_384_74.t36 Y.t10 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A.n0 A.t3 226.809
R1 A.n3 A.t4 226.809
R2 A.n4 A.t1 226.809
R3 A.n4 A.t2 198.204
R4 A.n0 A.t0 196.744
R5 A.n2 A.t5 196.013
R6 A A.n1 156.465
R7 A.n8 A.n7 152
R8 A.n6 A.n5 152
R9 A.n7 A.n6 49.6611
R10 A.n2 A.n1 40.8975
R11 A.n1 A.n0 21.1793
R12 A.n5 A 12.8005
R13 A.n6 A.n4 10.955
R14 A.n8 A 8.63306
R15 A A.n8 5.65631
R16 A.n7 A.n3 5.11262
R17 A.n3 A.n2 3.65202
R18 A.n5 A 1.48887
R19 a_27_74.n4 a_27_74.t7 309.284
R20 a_27_74.n21 a_27_74.t5 274.788
R21 a_27_74.n5 a_27_74.t8 240.197
R22 a_27_74.n8 a_27_74.t9 240.197
R23 a_27_74.n10 a_27_74.t11 240.197
R24 a_27_74.n15 a_27_74.t13 240.197
R25 a_27_74.n17 a_27_74.t16 240.197
R26 a_27_74.n1 a_27_74.t1 214.929
R27 a_27_74.n22 a_27_74.n21 205.486
R28 a_27_74.n17 a_27_74.t17 182.138
R29 a_27_74.n16 a_27_74.t14 179.947
R30 a_27_74.n4 a_27_74.t10 179.947
R31 a_27_74.n3 a_27_74.t15 179.947
R32 a_27_74.n9 a_27_74.t12 179.947
R33 a_27_74.n6 a_27_74.t6 179.947
R34 a_27_74.n12 a_27_74.n7 165.189
R35 a_27_74.n19 a_27_74.n18 152
R36 a_27_74.n16 a_27_74.n2 152
R37 a_27_74.n14 a_27_74.n13 152
R38 a_27_74.n12 a_27_74.n11 152
R39 a_27_74.n5 a_27_74.n4 107.939
R40 a_27_74.n1 a_27_74.n0 103.65
R41 a_27_74.n7 a_27_74.n6 49.6611
R42 a_27_74.n18 a_27_74.n16 49.6611
R43 a_27_74.n21 a_27_74.n20 49.3181
R44 a_27_74.n20 a_27_74.n1 45.5534
R45 a_27_74.n15 a_27_74.n14 41.6278
R46 a_27_74.n22 a_27_74.t4 26.3844
R47 a_27_74.t3 a_27_74.n22 26.3844
R48 a_27_74.n11 a_27_74.n9 26.2914
R49 a_27_74.n11 a_27_74.n10 25.5611
R50 a_27_74.n0 a_27_74.t2 22.7032
R51 a_27_74.n0 a_27_74.t0 22.7032
R52 a_27_74.n9 a_27_74.n8 13.8763
R53 a_27_74.n13 a_27_74.n12 13.1884
R54 a_27_74.n13 a_27_74.n2 13.1884
R55 a_27_74.n19 a_27_74.n2 13.1884
R56 a_27_74.n14 a_27_74.n3 13.146
R57 a_27_74.n10 a_27_74.n3 10.955
R58 a_27_74.n18 a_27_74.n17 10.955
R59 a_27_74.n20 a_27_74.n19 9.69747
R60 a_27_74.n8 a_27_74.n7 9.49444
R61 a_27_74.n16 a_27_74.n15 8.03383
R62 a_27_74.n6 a_27_74.n5 6.57323
R63 VGND.n49 VGND.n48 217
R64 VGND.n54 VGND.n2 211.183
R65 VGND.n57 VGND.n56 211.183
R66 VGND.n46 VGND.n45 209.243
R67 VGND.n14 VGND.t2 161.433
R68 VGND.n15 VGND.t11 152.998
R69 VGND.n36 VGND.n35 124.007
R70 VGND.n39 VGND.n38 116.644
R71 VGND.n13 VGND.n12 116.421
R72 VGND.n22 VGND.n21 116.421
R73 VGND.n10 VGND.n9 116.421
R74 VGND.n29 VGND.n28 116.421
R75 VGND.n7 VGND.n6 116.421
R76 VGND.n40 VGND.n37 36.1417
R77 VGND.n44 VGND.n4 36.1417
R78 VGND.n50 VGND.n47 36.1417
R79 VGND.n12 VGND.t8 34.0546
R80 VGND.n21 VGND.t22 34.0546
R81 VGND.n9 VGND.t4 34.0546
R82 VGND.n28 VGND.t5 34.0546
R83 VGND.n6 VGND.t23 34.0546
R84 VGND.n38 VGND.t21 34.0546
R85 VGND.n45 VGND.t17 34.0546
R86 VGND.n56 VGND.t18 32.4329
R87 VGND.n34 VGND.n7 28.9887
R88 VGND.n16 VGND.n13 27.4829
R89 VGND.n54 VGND.n1 27.4829
R90 VGND.n30 VGND.n29 26.7299
R91 VGND.n22 VGND.n20 25.224
R92 VGND.n27 VGND.n10 24.4711
R93 VGND.n57 VGND.n55 24.4711
R94 VGND.n23 VGND.n10 22.9652
R95 VGND.n12 VGND.t7 22.7032
R96 VGND.n21 VGND.t1 22.7032
R97 VGND.n9 VGND.t9 22.7032
R98 VGND.n28 VGND.t10 22.7032
R99 VGND.n6 VGND.t3 22.7032
R100 VGND.n35 VGND.t0 22.7032
R101 VGND.n35 VGND.t6 22.7032
R102 VGND.n38 VGND.t16 22.7032
R103 VGND.n45 VGND.t15 22.7032
R104 VGND.n48 VGND.t13 22.7032
R105 VGND.n48 VGND.t14 22.7032
R106 VGND.n2 VGND.t12 22.7032
R107 VGND.n2 VGND.t20 22.7032
R108 VGND.n56 VGND.t19 22.7032
R109 VGND.n23 VGND.n22 22.2123
R110 VGND.n29 VGND.n27 20.7064
R111 VGND.n20 VGND.n13 19.9534
R112 VGND.n55 VGND.n54 19.9534
R113 VGND.n30 VGND.n7 18.4476
R114 VGND.n16 VGND.n15 17.6946
R115 VGND.n36 VGND.n34 16.9417
R116 VGND.n49 VGND.n1 12.424
R117 VGND.n55 VGND.n0 9.3005
R118 VGND.n54 VGND.n53 9.3005
R119 VGND.n52 VGND.n1 9.3005
R120 VGND.n51 VGND.n50 9.3005
R121 VGND.n47 VGND.n3 9.3005
R122 VGND.n44 VGND.n43 9.3005
R123 VGND.n42 VGND.n4 9.3005
R124 VGND.n17 VGND.n16 9.3005
R125 VGND.n18 VGND.n13 9.3005
R126 VGND.n20 VGND.n19 9.3005
R127 VGND.n22 VGND.n11 9.3005
R128 VGND.n24 VGND.n23 9.3005
R129 VGND.n25 VGND.n10 9.3005
R130 VGND.n27 VGND.n26 9.3005
R131 VGND.n29 VGND.n8 9.3005
R132 VGND.n31 VGND.n30 9.3005
R133 VGND.n32 VGND.n7 9.3005
R134 VGND.n34 VGND.n33 9.3005
R135 VGND.n37 VGND.n5 9.3005
R136 VGND.n41 VGND.n40 9.3005
R137 VGND.n40 VGND.n39 8.65932
R138 VGND.n58 VGND.n57 7.19894
R139 VGND.n15 VGND.n14 6.96039
R140 VGND.n46 VGND.n44 6.4005
R141 VGND.n47 VGND.n46 4.89462
R142 VGND.n50 VGND.n49 4.89462
R143 VGND.n39 VGND.n4 2.63579
R144 VGND.n17 VGND.n14 0.594857
R145 VGND.n37 VGND.n36 0.376971
R146 VGND VGND.n58 0.156997
R147 VGND.n58 VGND.n0 0.150766
R148 VGND.n18 VGND.n17 0.122949
R149 VGND.n19 VGND.n18 0.122949
R150 VGND.n19 VGND.n11 0.122949
R151 VGND.n24 VGND.n11 0.122949
R152 VGND.n25 VGND.n24 0.122949
R153 VGND.n26 VGND.n25 0.122949
R154 VGND.n26 VGND.n8 0.122949
R155 VGND.n31 VGND.n8 0.122949
R156 VGND.n32 VGND.n31 0.122949
R157 VGND.n33 VGND.n32 0.122949
R158 VGND.n33 VGND.n5 0.122949
R159 VGND.n41 VGND.n5 0.122949
R160 VGND.n42 VGND.n41 0.122949
R161 VGND.n43 VGND.n42 0.122949
R162 VGND.n43 VGND.n3 0.122949
R163 VGND.n51 VGND.n3 0.122949
R164 VGND.n52 VGND.n51 0.122949
R165 VGND.n53 VGND.n52 0.122949
R166 VGND.n53 VGND.n0 0.122949
R167 VNB.t11 VNB.t2 2148.03
R168 VNB.t7 VNB.t8 1154.86
R169 VNB.t1 VNB.t22 1154.86
R170 VNB.t9 VNB.t4 1154.86
R171 VNB.t10 VNB.t5 1154.86
R172 VNB.t3 VNB.t23 1154.86
R173 VNB.t16 VNB.t21 1154.86
R174 VNB.t15 VNB.t17 1154.86
R175 VNB VNB.t19 1143.31
R176 VNB.t19 VNB.t18 1131.76
R177 VNB.t8 VNB.t11 993.177
R178 VNB.t22 VNB.t7 993.177
R179 VNB.t4 VNB.t1 993.177
R180 VNB.t5 VNB.t9 993.177
R181 VNB.t23 VNB.t10 993.177
R182 VNB.t0 VNB.t3 993.177
R183 VNB.t6 VNB.t0 993.177
R184 VNB.t21 VNB.t6 993.177
R185 VNB.t17 VNB.t16 993.177
R186 VNB.t13 VNB.t15 993.177
R187 VNB.t14 VNB.t13 993.177
R188 VNB.t12 VNB.t14 993.177
R189 VNB.t20 VNB.t12 993.177
R190 VNB.t18 VNB.t20 993.177
R191 a_384_74.n5 a_384_74.n3 250.518
R192 a_384_74.n18 a_384_74.t13 246.769
R193 a_384_74.n20 a_384_74.t26 240.197
R194 a_384_74.n24 a_384_74.t20 240.197
R195 a_384_74.n22 a_384_74.n21 240.197
R196 a_384_74.n28 a_384_74.n15 240.197
R197 a_384_74.n31 a_384_74.t17 240.197
R198 a_384_74.n34 a_384_74.t23 240.197
R199 a_384_74.n36 a_384_74.n14 240.197
R200 a_384_74.n39 a_384_74.t25 240.197
R201 a_384_74.n12 a_384_74.n11 240.197
R202 a_384_74.n44 a_384_74.t29 240.197
R203 a_384_74.n46 a_384_74.n10 240.197
R204 a_384_74.n49 a_384_74.t32 240.197
R205 a_384_74.n51 a_384_74.n9 240.197
R206 a_384_74.n55 a_384_74.t33 240.197
R207 a_384_74.n53 a_384_74.t15 240.197
R208 a_384_74.n5 a_384_74.n4 207.6
R209 a_384_74.n7 a_384_74.n6 207.6
R210 a_384_74.n53 a_384_74.t12 182.138
R211 a_384_74.n54 a_384_74.t28 179.947
R212 a_384_74.n52 a_384_74.t18 179.947
R213 a_384_74.n50 a_384_74.t22 179.947
R214 a_384_74.n47 a_384_74.t16 179.947
R215 a_384_74.n45 a_384_74.t35 179.947
R216 a_384_74.n37 a_384_74.t27 179.947
R217 a_384_74.n38 a_384_74.t34 179.947
R218 a_384_74.n35 a_384_74.t24 179.947
R219 a_384_74.n33 a_384_74.t19 179.947
R220 a_384_74.n30 a_384_74.t14 179.947
R221 a_384_74.n29 a_384_74.t30 179.947
R222 a_384_74.n16 a_384_74.t31 179.947
R223 a_384_74.n23 a_384_74.t36 179.947
R224 a_384_74.n19 a_384_74.n17 179.947
R225 a_384_74.n18 a_384_74.t21 179.947
R226 a_384_74.n57 a_384_74.n56 170.781
R227 a_384_74.n26 a_384_74.n25 169.566
R228 a_384_74.n27 a_384_74.n26 169.059
R229 a_384_74.n32 a_384_74.n13 169.059
R230 a_384_74.n41 a_384_74.n40 169.059
R231 a_384_74.n43 a_384_74.n42 169.059
R232 a_384_74.n48 a_384_74.n8 169.059
R233 a_384_74.n2 a_384_74.n0 152.511
R234 a_384_74.n2 a_384_74.n1 102.019
R235 a_384_74.n60 a_384_74.n59 102.019
R236 a_384_74.n19 a_384_74.n18 62.8066
R237 a_384_74.n30 a_384_74.n29 62.8066
R238 a_384_74.n38 a_384_74.n37 62.8066
R239 a_384_74.n23 a_384_74.n22 62.0763
R240 a_384_74.n35 a_384_74.n34 60.6157
R241 a_384_74.n54 a_384_74.n53 60.6157
R242 a_384_74.n46 a_384_74.n45 59.155
R243 a_384_74.n51 a_384_74.n50 54.7732
R244 a_384_74.n59 a_384_74.n2 51.2005
R245 a_384_74.n27 a_384_74.n16 43.0884
R246 a_384_74.n7 a_384_74.n5 42.9181
R247 a_384_74.n48 a_384_74.n47 42.3581
R248 a_384_74.n25 a_384_74.n20 40.8975
R249 a_384_74.n32 a_384_74.n31 40.8975
R250 a_384_74.n43 a_384_74.n12 40.1672
R251 a_384_74.n40 a_384_74.n36 37.246
R252 a_384_74.n56 a_384_74.n52 36.5157
R253 a_384_74.n33 a_384_74.n32 29.9429
R254 a_384_74.n3 a_384_74.t0 29.9023
R255 a_384_74.n28 a_384_74.n27 29.2126
R256 a_384_74.n40 a_384_74.n39 28.4823
R257 a_384_74.n6 a_384_74.t5 26.3844
R258 a_384_74.n6 a_384_74.t4 26.3844
R259 a_384_74.n3 a_384_74.t1 26.3844
R260 a_384_74.n4 a_384_74.t3 26.3844
R261 a_384_74.n4 a_384_74.t2 26.3844
R262 a_384_74.n25 a_384_74.n24 26.2914
R263 a_384_74.n44 a_384_74.n43 25.5611
R264 a_384_74.n0 a_384_74.t8 22.7032
R265 a_384_74.n0 a_384_74.t6 22.7032
R266 a_384_74.n1 a_384_74.t9 22.7032
R267 a_384_74.n1 a_384_74.t7 22.7032
R268 a_384_74.n60 a_384_74.t10 22.7032
R269 a_384_74.t11 a_384_74.n60 22.7032
R270 a_384_74.n58 a_384_74.n57 21.2906
R271 a_384_74.n56 a_384_74.n55 21.1793
R272 a_384_74.n49 a_384_74.n48 19.7187
R273 a_384_74.n59 a_384_74.n58 15.0476
R274 a_384_74.n50 a_384_74.n49 10.955
R275 a_384_74.n52 a_384_74.n51 8.03383
R276 a_384_74.n45 a_384_74.n44 6.57323
R277 a_384_74.n58 a_384_74.n7 5.23686
R278 a_384_74.n36 a_384_74.n35 5.11262
R279 a_384_74.n55 a_384_74.n54 5.11262
R280 a_384_74.n24 a_384_74.n23 3.65202
R281 a_384_74.n47 a_384_74.n46 3.65202
R282 a_384_74.n20 a_384_74.n19 2.19141
R283 a_384_74.n31 a_384_74.n30 2.19141
R284 a_384_74.n34 a_384_74.n33 2.19141
R285 a_384_74.n39 a_384_74.n38 2.19141
R286 a_384_74.n22 a_384_74.n16 0.730803
R287 a_384_74.n29 a_384_74.n28 0.730803
R288 a_384_74.n37 a_384_74.n12 0.730803
R289 a_384_74.n42 a_384_74.n8 0.51137
R290 a_384_74.n41 a_384_74.n13 0.505935
R291 a_384_74.n26 a_384_74.n13 0.503217
R292 a_384_74.n42 a_384_74.n41 0.497783
R293 a_384_74.n57 a_384_74.n8 0.484196
R294 Y.n18 Y.t1 229.026
R295 Y.n15 Y.t2 229.024
R296 Y.n3 Y.t6 229.022
R297 Y.n12 Y.t4 229.016
R298 Y.n6 Y.t7 228.835
R299 Y.n9 Y.t5 228.815
R300 Y.n22 Y.n20 202.641
R301 Y.n1 Y.n0 202.486
R302 Y.n1 Y.t19 184.966
R303 Y.n18 Y.n17 159.352
R304 Y.n15 Y.n14 154.112
R305 Y.n12 Y.n11 151.978
R306 Y.n9 Y.n8 150.885
R307 Y.n3 Y.n2 150.716
R308 Y.n6 Y.n5 150.657
R309 Y.n22 Y.n21 150.618
R310 Y.n0 Y.t3 33.4201
R311 Y.n20 Y.t0 26.3844
R312 Y.n20 Y.t8 26.3844
R313 Y.n0 Y.t9 26.3844
R314 Y.n21 Y.t15 22.7032
R315 Y.n21 Y.t24 22.7032
R316 Y.n17 Y.t18 22.7032
R317 Y.n17 Y.t21 22.7032
R318 Y.n14 Y.t11 22.7032
R319 Y.n14 Y.t22 22.7032
R320 Y.n11 Y.t12 22.7032
R321 Y.n11 Y.t16 22.7032
R322 Y.n8 Y.t20 22.7032
R323 Y.n8 Y.t17 22.7032
R324 Y.n5 Y.t14 22.7032
R325 Y.n5 Y.t23 22.7032
R326 Y.n2 Y.t10 22.7032
R327 Y.n2 Y.t13 22.7032
R328 Y.n4 Y.n1 10.4435
R329 Y.n10 Y.n9 10.0106
R330 Y.n7 Y.n6 9.97939
R331 Y.n13 Y.n12 9.70406
R332 Y.n4 Y.n3 9.69531
R333 Y.n16 Y.n15 9.69256
R334 Y.n23 Y.n22 9.68988
R335 Y.n19 Y.n18 9.68728
R336 Y.n7 Y.n4 0.516804
R337 Y.n10 Y.n7 0.516804
R338 Y.n13 Y.n10 0.48963
R339 Y.n16 Y.n13 0.48963
R340 Y.n19 Y.n16 0.48963
R341 Y.n23 Y.n19 0.484196
R342 Y Y.n23 0.0847391
R343 VPWR.n49 VPWR.n48 334.173
R344 VPWR.n46 VPWR.n5 334.173
R345 VPWR.n55 VPWR.n2 331.5
R346 VPWR.n57 VPWR.n1 331.5
R347 VPWR.n37 VPWR.t0 268.509
R348 VPWR.n31 VPWR.t1 268.509
R349 VPWR.n29 VPWR.t2 268.509
R350 VPWR.n23 VPWR.t4 268.509
R351 VPWR.n14 VPWR.t9 266.2
R352 VPWR.n40 VPWR.n39 242.125
R353 VPWR.n16 VPWR.n15 237.425
R354 VPWR.n22 VPWR.n12 235.556
R355 VPWR.n28 VPWR.n10 36.1417
R356 VPWR.n32 VPWR.n30 36.1417
R357 VPWR.n36 VPWR.n8 36.1417
R358 VPWR.n41 VPWR.n38 36.1417
R359 VPWR.n45 VPWR.n6 36.1417
R360 VPWR.n50 VPWR.n47 36.1417
R361 VPWR.n54 VPWR.n3 36.1417
R362 VPWR.n12 VPWR.t7 35.1791
R363 VPWR.n57 VPWR.n56 35.0123
R364 VPWR.n24 VPWR.n23 33.5064
R365 VPWR.n56 VPWR.n55 32.7534
R366 VPWR.n49 VPWR.n3 29.7417
R367 VPWR.n29 VPWR.n28 28.9887
R368 VPWR.n15 VPWR.t3 28.1434
R369 VPWR.n24 VPWR.n22 27.8593
R370 VPWR.n22 VPWR.n21 27.4829
R371 VPWR.n17 VPWR.n13 27.4829
R372 VPWR.n21 VPWR.n13 27.1064
R373 VPWR.n1 VPWR.t16 26.3844
R374 VPWR.n1 VPWR.t18 26.3844
R375 VPWR.n2 VPWR.t10 26.3844
R376 VPWR.n2 VPWR.t17 26.3844
R377 VPWR.n48 VPWR.t12 26.3844
R378 VPWR.n48 VPWR.t11 26.3844
R379 VPWR.n5 VPWR.t14 26.3844
R380 VPWR.n5 VPWR.t13 26.3844
R381 VPWR.n39 VPWR.t8 26.3844
R382 VPWR.n39 VPWR.t15 26.3844
R383 VPWR.n12 VPWR.t5 26.3844
R384 VPWR.n15 VPWR.t6 26.3844
R385 VPWR.n17 VPWR.n16 26.3534
R386 VPWR.n47 VPWR.n46 25.224
R387 VPWR.n32 VPWR.n31 24.4711
R388 VPWR.n40 VPWR.n6 20.7064
R389 VPWR.n37 VPWR.n36 19.9534
R390 VPWR.n38 VPWR.n37 16.1887
R391 VPWR.n41 VPWR.n40 15.4358
R392 VPWR.n31 VPWR.n8 11.6711
R393 VPWR.n46 VPWR.n45 10.9181
R394 VPWR.n18 VPWR.n17 9.3005
R395 VPWR.n19 VPWR.n13 9.3005
R396 VPWR.n21 VPWR.n20 9.3005
R397 VPWR.n22 VPWR.n11 9.3005
R398 VPWR.n25 VPWR.n24 9.3005
R399 VPWR.n26 VPWR.n10 9.3005
R400 VPWR.n28 VPWR.n27 9.3005
R401 VPWR.n30 VPWR.n9 9.3005
R402 VPWR.n33 VPWR.n32 9.3005
R403 VPWR.n34 VPWR.n8 9.3005
R404 VPWR.n36 VPWR.n35 9.3005
R405 VPWR.n38 VPWR.n7 9.3005
R406 VPWR.n42 VPWR.n41 9.3005
R407 VPWR.n43 VPWR.n6 9.3005
R408 VPWR.n45 VPWR.n44 9.3005
R409 VPWR.n47 VPWR.n4 9.3005
R410 VPWR.n51 VPWR.n50 9.3005
R411 VPWR.n52 VPWR.n3 9.3005
R412 VPWR.n54 VPWR.n53 9.3005
R413 VPWR.n56 VPWR.n0 9.3005
R414 VPWR.n58 VPWR.n57 8.8332
R415 VPWR.n30 VPWR.n29 7.15344
R416 VPWR.n16 VPWR.n14 7.02164
R417 VPWR.n50 VPWR.n49 6.4005
R418 VPWR.n55 VPWR.n54 3.38874
R419 VPWR.n23 VPWR.n10 2.63579
R420 VPWR.n18 VPWR.n14 0.543334
R421 VPWR VPWR.n58 0.163644
R422 VPWR.n58 VPWR.n0 0.144205
R423 VPWR.n19 VPWR.n18 0.122949
R424 VPWR.n20 VPWR.n19 0.122949
R425 VPWR.n20 VPWR.n11 0.122949
R426 VPWR.n25 VPWR.n11 0.122949
R427 VPWR.n26 VPWR.n25 0.122949
R428 VPWR.n27 VPWR.n26 0.122949
R429 VPWR.n27 VPWR.n9 0.122949
R430 VPWR.n33 VPWR.n9 0.122949
R431 VPWR.n34 VPWR.n33 0.122949
R432 VPWR.n35 VPWR.n34 0.122949
R433 VPWR.n35 VPWR.n7 0.122949
R434 VPWR.n42 VPWR.n7 0.122949
R435 VPWR.n43 VPWR.n42 0.122949
R436 VPWR.n44 VPWR.n43 0.122949
R437 VPWR.n44 VPWR.n4 0.122949
R438 VPWR.n51 VPWR.n4 0.122949
R439 VPWR.n52 VPWR.n51 0.122949
R440 VPWR.n53 VPWR.n52 0.122949
R441 VPWR.n53 VPWR.n0 0.122949
R442 VPB.t7 VPB.t6 715.054
R443 VPB.t4 VPB.t5 459.678
R444 VPB.t2 VPB.t4 459.678
R445 VPB.t1 VPB.t2 459.678
R446 VPB.t0 VPB.t1 459.678
R447 VPB VPB.t18 260.485
R448 VPB.t5 VPB.t7 255.376
R449 VPB.t3 VPB.t9 250.269
R450 VPB.t10 VPB.t11 240.054
R451 VPB.t6 VPB.t3 234.946
R452 VPB.t8 VPB.t0 229.839
R453 VPB.t15 VPB.t8 229.839
R454 VPB.t14 VPB.t15 229.839
R455 VPB.t13 VPB.t14 229.839
R456 VPB.t12 VPB.t13 229.839
R457 VPB.t11 VPB.t12 229.839
R458 VPB.t17 VPB.t10 229.839
R459 VPB.t16 VPB.t17 229.839
R460 VPB.t18 VPB.t16 229.839
C0 VPB VPWR 0.324458f
C1 A VPWR 0.047431f
C2 VPB Y 0.047977f
C3 A Y 5.85e-20
C4 VPB VGND 0.010846f
C5 VPWR Y 1.9952f
C6 A VGND 0.054906f
C7 VPWR VGND 0.111478f
C8 Y VGND 1.24531f
C9 VPB A 0.101906f
C10 VGND VNB 1.39278f
C11 Y VNB 0.069213f
C12 VPWR VNB 1.13625f
C13 A VNB 0.342428f
C14 VPB VNB 2.76322f
C15 Y.t19 VNB 0.045159f
C16 Y.t9 VNB 0.014784f
C17 Y.t3 VNB 0.018726f
C18 Y.n0 VNB 0.036081f
C19 Y.n1 VNB 0.140904f
C20 Y.t6 VNB 0.056301f
C21 Y.t10 VNB 0.009117f
C22 Y.t13 VNB 0.009117f
C23 Y.n2 VNB 0.036933f
C24 Y.n3 VNB 0.112867f
C25 Y.n4 VNB 0.067707f
C26 Y.t7 VNB 0.056297f
C27 Y.t14 VNB 0.009117f
C28 Y.t23 VNB 0.009117f
C29 Y.n5 VNB 0.036905f
C30 Y.n6 VNB 0.111056f
C31 Y.n7 VNB 0.042113f
C32 Y.t5 VNB 0.056296f
C33 Y.t20 VNB 0.009117f
C34 Y.t17 VNB 0.009117f
C35 Y.n8 VNB 0.036979f
C36 Y.n9 VNB 0.110476f
C37 Y.n10 VNB 0.041255f
C38 Y.t12 VNB 0.009117f
C39 Y.t16 VNB 0.009117f
C40 Y.n11 VNB 0.03681f
C41 Y.t4 VNB 0.056301f
C42 Y.n12 VNB 0.111303f
C43 Y.n13 VNB 0.038643f
C44 Y.t2 VNB 0.056301f
C45 Y.t11 VNB 0.009117f
C46 Y.t22 VNB 0.009117f
C47 Y.n14 VNB 0.03639f
C48 Y.n15 VNB 0.109372f
C49 Y.n16 VNB 0.038583f
C50 Y.t1 VNB 0.056301f
C51 Y.t18 VNB 0.009117f
C52 Y.t21 VNB 0.009117f
C53 Y.n17 VNB 0.035617f
C54 Y.n18 VNB 0.104822f
C55 Y.n19 VNB 0.038353f
C56 Y.t0 VNB 0.014784f
C57 Y.t8 VNB 0.014784f
C58 Y.n20 VNB 0.032139f
C59 Y.t15 VNB 0.009117f
C60 Y.t24 VNB 0.009117f
C61 Y.n21 VNB 0.0369f
C62 Y.n22 VNB 0.107699f
C63 Y.n23 VNB 0.023288f
C64 a_384_74.t10 VNB 0.007836f
C65 a_384_74.t8 VNB 0.007836f
C66 a_384_74.t6 VNB 0.007836f
C67 a_384_74.n0 VNB 0.025874f
C68 a_384_74.t9 VNB 0.007836f
C69 a_384_74.t7 VNB 0.007836f
C70 a_384_74.n1 VNB 0.018234f
C71 a_384_74.n2 VNB 0.061222f
C72 a_384_74.t1 VNB 0.012707f
C73 a_384_74.t0 VNB 0.014401f
C74 a_384_74.n3 VNB 0.041293f
C75 a_384_74.t3 VNB 0.012707f
C76 a_384_74.t2 VNB 0.012707f
C77 a_384_74.n4 VNB 0.028839f
C78 a_384_74.n5 VNB 0.122187f
C79 a_384_74.t5 VNB 0.012707f
C80 a_384_74.t4 VNB 0.012707f
C81 a_384_74.n6 VNB 0.028839f
C82 a_384_74.n7 VNB 0.061936f
C83 a_384_74.n8 VNB 0.052456f
C84 a_384_74.t18 VNB 0.011799f
C85 a_384_74.n9 VNB 0.018322f
C86 a_384_74.t22 VNB 0.011799f
C87 a_384_74.t32 VNB 0.018322f
C88 a_384_74.t16 VNB 0.011799f
C89 a_384_74.n10 VNB 0.018322f
C90 a_384_74.t35 VNB 0.011799f
C91 a_384_74.t29 VNB 0.018322f
C92 a_384_74.n11 VNB 0.018322f
C93 a_384_74.n12 VNB 0.016508f
C94 a_384_74.n13 VNB 0.052891f
C95 a_384_74.n14 VNB 0.018322f
C96 a_384_74.t24 VNB 0.011799f
C97 a_384_74.t23 VNB 0.018322f
C98 a_384_74.t19 VNB 0.011799f
C99 a_384_74.t17 VNB 0.018322f
C100 a_384_74.t14 VNB 0.011799f
C101 a_384_74.t30 VNB 0.011799f
C102 a_384_74.n15 VNB 0.018322f
C103 a_384_74.t31 VNB 0.011799f
C104 a_384_74.n16 VNB 0.013841f
C105 a_384_74.t26 VNB 0.018322f
C106 a_384_74.n17 VNB 0.011799f
C107 a_384_74.t21 VNB 0.011799f
C108 a_384_74.t13 VNB 0.018725f
C109 a_384_74.n18 VNB 0.032941f
C110 a_384_74.n19 VNB 0.017461f
C111 a_384_74.n20 VNB 0.016882f
C112 a_384_74.t20 VNB 0.018322f
C113 a_384_74.t36 VNB 0.011799f
C114 a_384_74.n21 VNB 0.018322f
C115 a_384_74.n22 VNB 0.020252f
C116 a_384_74.n23 VNB 0.017585f
C117 a_384_74.n24 VNB 0.014636f
C118 a_384_74.n25 VNB 0.01345f
C119 a_384_74.n26 VNB 0.094784f
C120 a_384_74.n27 VNB 0.014198f
C121 a_384_74.n28 VNB 0.014636f
C122 a_384_74.n29 VNB 0.017211f
C123 a_384_74.n30 VNB 0.017461f
C124 a_384_74.n31 VNB 0.016882f
C125 a_384_74.n32 VNB 0.013948f
C126 a_384_74.n33 VNB 0.011844f
C127 a_384_74.n34 VNB 0.020252f
C128 a_384_74.n35 VNB 0.017585f
C129 a_384_74.n36 VNB 0.016758f
C130 a_384_74.t25 VNB 0.018322f
C131 a_384_74.t34 VNB 0.011799f
C132 a_384_74.t27 VNB 0.011799f
C133 a_384_74.n37 VNB 0.017211f
C134 a_384_74.n38 VNB 0.017461f
C135 a_384_74.n39 VNB 0.014761f
C136 a_384_74.n40 VNB 0.013075f
C137 a_384_74.n41 VNB 0.052717f
C138 a_384_74.n42 VNB 0.052891f
C139 a_384_74.n43 VNB 0.013075f
C140 a_384_74.n44 VNB 0.01501f
C141 a_384_74.n45 VNB 0.017585f
C142 a_384_74.n46 VNB 0.020252f
C143 a_384_74.n47 VNB 0.014216f
C144 a_384_74.n48 VNB 0.012451f
C145 a_384_74.n49 VNB 0.014761f
C146 a_384_74.n50 VNB 0.017585f
C147 a_384_74.n51 VNB 0.020252f
C148 a_384_74.n52 VNB 0.013966f
C149 a_384_74.t33 VNB 0.018322f
C150 a_384_74.t28 VNB 0.011799f
C151 a_384_74.t15 VNB 0.018322f
C152 a_384_74.t12 VNB 0.011925f
C153 a_384_74.n53 VNB 0.030598f
C154 a_384_74.n54 VNB 0.017585f
C155 a_384_74.n55 VNB 0.014012f
C156 a_384_74.n56 VNB 0.011461f
C157 a_384_74.n57 VNB 0.07936f
C158 a_384_74.n58 VNB 0.042081f
C159 a_384_74.n59 VNB 0.039095f
C160 a_384_74.n60 VNB 0.018234f
C161 a_384_74.t11 VNB 0.007836f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkbuf_8 VNB VPB VPWR VGND X A
X0 X.t15 a_125_368.t4 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0882 ps=0.84 w=0.42 l=0.15
X1 VGND.t6 a_125_368.t5 X.t14 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND.t5 a_125_368.t6 X.t13 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0882 pd=0.84 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 X.t5 a_125_368.t7 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.196 ps=1.47 w=1.12 l=0.15
X4 a_125_368.t3 A.t0 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1491 ps=1.55 w=0.42 l=0.15
X5 X.t12 a_125_368.t8 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR.t9 A.t1 a_125_368.t2 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.1708 ps=1.425 w=1.12 l=0.15
X7 X.t11 a_125_368.t9 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 a_125_368.t1 A.t2 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1708 pd=1.425 as=0.3808 ps=2.92 w=1.12 l=0.15
X9 VPWR.t6 a_125_368.t10 X.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VGND.t2 a_125_368.t11 X.t10 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 X.t7 a_125_368.t12 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VPWR.t4 a_125_368.t13 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 X.t2 a_125_368.t14 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 X.t9 a_125_368.t15 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.06405 pd=0.725 as=0.08295 ps=0.815 w=0.42 l=0.15
X15 VGND.t8 a_125_368.t16 X.t8 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VGND.t0 A.t3 a_125_368.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.08295 pd=0.815 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR.t2 a_125_368.t17 X.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VPWR.t1 a_125_368.t18 X.t4 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X19 X.t1 a_125_368.t19 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
R0 a_125_368.n8 a_125_368.t18 269.652
R1 a_125_368.n9 a_125_368.t7 269.652
R2 a_125_368.n12 a_125_368.t10 269.652
R3 a_125_368.n7 a_125_368.t12 269.652
R4 a_125_368.n18 a_125_368.t13 269.652
R5 a_125_368.n6 a_125_368.t14 269.652
R6 a_125_368.n24 a_125_368.t17 269.652
R7 a_125_368.n27 a_125_368.t19 269.652
R8 a_125_368.n31 a_125_368.n30 269.111
R9 a_125_368.n30 a_125_368.n4 238.071
R10 a_125_368.n27 a_125_368.t15 198.204
R11 a_125_368.n8 a_125_368.t5 198.204
R12 a_125_368.n25 a_125_368.t6 196.013
R13 a_125_368.n19 a_125_368.t4 196.013
R14 a_125_368.n3 a_125_368.t16 196.013
R15 a_125_368.n13 a_125_368.t9 196.013
R16 a_125_368.n11 a_125_368.t11 196.013
R17 a_125_368.n1 a_125_368.t8 196.013
R18 a_125_368.n1 a_125_368.n0 165.189
R19 a_125_368.n29 a_125_368.n28 152
R20 a_125_368.n26 a_125_368.n5 152
R21 a_125_368.n23 a_125_368.n22 152
R22 a_125_368.n21 a_125_368.n20 152
R23 a_125_368.n3 a_125_368.n2 152
R24 a_125_368.n17 a_125_368.n16 152
R25 a_125_368.n15 a_125_368.n14 152
R26 a_125_368.n10 a_125_368.n0 152
R27 a_125_368.n1 a_125_368.n8 60.6157
R28 a_125_368.n28 a_125_368.n26 49.6611
R29 a_125_368.n3 a_125_368.n17 48.9308
R30 a_125_368.n24 a_125_368.n23 44.549
R31 a_125_368.n10 a_125_368.n9 43.0884
R32 a_125_368.n4 a_125_368.t0 40.0005
R33 a_125_368.n4 a_125_368.t3 40.0005
R34 a_125_368.n20 a_125_368.n18 37.246
R35 a_125_368.n14 a_125_368.n13 35.7853
R36 a_125_368.t1 a_125_368.n31 27.2639
R37 a_125_368.n31 a_125_368.t2 26.3844
R38 a_125_368.n11 a_125_368.n10 22.6399
R39 a_125_368.n23 a_125_368.n6 21.1793
R40 a_125_368.n14 a_125_368.n12 19.7187
R41 a_125_368.n19 a_125_368.n6 16.0672
R42 a_125_368.n15 a_125_368.n0 13.1884
R43 a_125_368.n16 a_125_368.n15 13.1884
R44 a_125_368.n16 a_125_368.n2 13.1884
R45 a_125_368.n21 a_125_368.n2 13.1884
R46 a_125_368.n22 a_125_368.n21 13.1884
R47 a_125_368.n22 a_125_368.n5 13.1884
R48 a_125_368.n29 a_125_368.n5 13.1884
R49 a_125_368.n18 a_125_368.n3 13.146
R50 a_125_368.n20 a_125_368.n19 12.4157
R51 a_125_368.n28 a_125_368.n27 10.955
R52 a_125_368.n30 a_125_368.n29 10.4732
R53 a_125_368.n13 a_125_368.n7 10.2247
R54 a_125_368.n12 a_125_368.n11 7.30353
R55 a_125_368.n9 a_125_368.n1 7.30353
R56 a_125_368.n17 a_125_368.n7 3.65202
R57 a_125_368.n26 a_125_368.n25 3.65202
R58 a_125_368.n25 a_125_368.n24 1.46111
R59 VGND.n20 VGND.t9 267.498
R60 VGND.n8 VGND.t6 251.506
R61 VGND.n18 VGND.n2 207.498
R62 VGND.n11 VGND.n5 204.976
R63 VGND.n14 VGND.n13 204.976
R64 VGND.n7 VGND.n6 201.481
R65 VGND.n13 VGND.t7 60.0005
R66 VGND.n13 VGND.t5 60.0005
R67 VGND.n2 VGND.t0 60.0005
R68 VGND.n2 VGND.t1 52.8576
R69 VGND.n6 VGND.t4 50.0005
R70 VGND.n6 VGND.t2 50.0005
R71 VGND.n5 VGND.t3 40.0005
R72 VGND.n5 VGND.t8 40.0005
R73 VGND.n14 VGND.n1 32.7534
R74 VGND.n12 VGND.n11 30.4946
R75 VGND.n19 VGND.n18 29.7417
R76 VGND.n7 VGND.n4 22.9652
R77 VGND.n20 VGND.n19 20.7064
R78 VGND.n18 VGND.n1 17.6946
R79 VGND.n11 VGND.n4 16.9417
R80 VGND.n14 VGND.n12 14.6829
R81 VGND.n21 VGND.n20 9.3005
R82 VGND.n9 VGND.n4 9.3005
R83 VGND.n11 VGND.n10 9.3005
R84 VGND.n12 VGND.n3 9.3005
R85 VGND.n15 VGND.n14 9.3005
R86 VGND.n16 VGND.n1 9.3005
R87 VGND.n18 VGND.n17 9.3005
R88 VGND.n19 VGND.n0 9.3005
R89 VGND.n8 VGND.n7 6.26985
R90 VGND.n9 VGND.n8 0.733933
R91 VGND.n10 VGND.n9 0.122949
R92 VGND.n10 VGND.n3 0.122949
R93 VGND.n15 VGND.n3 0.122949
R94 VGND.n16 VGND.n15 0.122949
R95 VGND.n17 VGND.n16 0.122949
R96 VGND.n17 VGND.n0 0.122949
R97 VGND.n21 VGND.n0 0.122949
R98 VGND VGND.n21 0.0617245
R99 X.n2 X.n0 269.019
R100 X.n11 X.n9 249.218
R101 X.n2 X.n1 216.333
R102 X.n6 X.n5 216.333
R103 X.n4 X.n3 215.936
R104 X.n12 X.n8 205.329
R105 X.n13 X.n7 205.329
R106 X.n11 X.n10 203.177
R107 X.n13 X.n12 70.024
R108 X.n12 X.n11 58.3534
R109 X.n6 X.n4 53.0829
R110 X.n9 X.t9 47.1434
R111 X.n4 X.n2 42.9181
R112 X.n9 X.t13 40.0005
R113 X.n10 X.t8 40.0005
R114 X.n10 X.t15 40.0005
R115 X.n8 X.t10 40.0005
R116 X.n8 X.t11 40.0005
R117 X.n7 X.t14 40.0005
R118 X.n7 X.t12 40.0005
R119 X X.n13 29.8517
R120 X.n5 X.t4 28.1434
R121 X.n5 X.t5 27.2639
R122 X.n0 X.t0 26.3844
R123 X.n0 X.t1 26.3844
R124 X.n1 X.t3 26.3844
R125 X.n1 X.t2 26.3844
R126 X.n3 X.t6 26.3844
R127 X.n3 X.t7 26.3844
R128 X X.n6 10.5036
R129 VNB.t6 VNB.t8 1316.54
R130 VNB VNB.t9 1304.99
R131 VNB.t0 VNB.t2 1258.79
R132 VNB.t3 VNB.t5 1154.86
R133 VNB.t2 VNB.t6 1050.92
R134 VNB.t5 VNB.t7 993.177
R135 VNB.t4 VNB.t3 993.177
R136 VNB.t1 VNB.t4 993.177
R137 VNB.t8 VNB.t1 993.177
R138 VNB.t9 VNB.t0 993.177
R139 VPWR.n12 VPWR.n6 336.101
R140 VPWR.n19 VPWR.n2 315.928
R141 VPWR.n21 VPWR.t8 256.659
R142 VPWR.n9 VPWR.t1 255.514
R143 VPWR.n4 VPWR.n3 222.486
R144 VPWR.n8 VPWR.n7 222.486
R145 VPWR.n14 VPWR.n13 36.1417
R146 VPWR.n12 VPWR.n11 35.3887
R147 VPWR.n2 VPWR.t0 35.1791
R148 VPWR.n2 VPWR.t9 35.1791
R149 VPWR.n7 VPWR.t7 35.1791
R150 VPWR.n20 VPWR.n19 29.7417
R151 VPWR.n18 VPWR.n4 28.9887
R152 VPWR.n3 VPWR.t3 26.3844
R153 VPWR.n3 VPWR.t2 26.3844
R154 VPWR.n6 VPWR.t5 26.3844
R155 VPWR.n6 VPWR.t4 26.3844
R156 VPWR.n7 VPWR.t6 26.3844
R157 VPWR.n21 VPWR.n20 20.7064
R158 VPWR.n11 VPWR.n8 19.9534
R159 VPWR.n14 VPWR.n4 18.4476
R160 VPWR.n19 VPWR.n18 17.6946
R161 VPWR.n11 VPWR.n10 9.3005
R162 VPWR.n13 VPWR.n5 9.3005
R163 VPWR.n15 VPWR.n14 9.3005
R164 VPWR.n16 VPWR.n4 9.3005
R165 VPWR.n18 VPWR.n17 9.3005
R166 VPWR.n19 VPWR.n1 9.3005
R167 VPWR.n20 VPWR.n0 9.3005
R168 VPWR.n22 VPWR.n21 9.3005
R169 VPWR.n9 VPWR.n8 6.83455
R170 VPWR.n13 VPWR.n12 0.753441
R171 VPWR.n10 VPWR.n9 0.623818
R172 VPWR.n10 VPWR.n5 0.122949
R173 VPWR.n15 VPWR.n5 0.122949
R174 VPWR.n16 VPWR.n15 0.122949
R175 VPWR.n17 VPWR.n16 0.122949
R176 VPWR.n17 VPWR.n1 0.122949
R177 VPWR.n1 VPWR.n0 0.122949
R178 VPWR.n22 VPWR.n0 0.122949
R179 VPWR VPWR.n22 0.0617245
R180 VPB.t9 VPB.t0 280.914
R181 VPB VPB.t8 280.914
R182 VPB.t6 VPB.t7 255.376
R183 VPB.t7 VPB.t1 237.5
R184 VPB.t8 VPB.t9 232.393
R185 VPB.t5 VPB.t6 229.839
R186 VPB.t4 VPB.t5 229.839
R187 VPB.t3 VPB.t4 229.839
R188 VPB.t2 VPB.t3 229.839
R189 VPB.t0 VPB.t2 229.839
R190 A.n2 A.t0 247.428
R191 A.n0 A.t3 247.428
R192 A.n2 A.t2 229
R193 A.n0 A.t1 228.268
R194 A A.n1 160.781
R195 A.n4 A.n3 152
R196 A.n3 A.n1 49.6611
R197 A.n4 A 12.9493
R198 A.n1 A.n0 9.49444
R199 A.n3 A.n2 3.65202
R200 A A.n4 1.34003
C0 VPWR X 0.852784f
C1 A VGND 0.049326f
C2 VPWR VGND 0.090671f
C3 X VGND 0.498722f
C4 VPB A 0.070217f
C5 VPB VPWR 0.154593f
C6 A VPWR 0.072656f
C7 VPB X 0.026065f
C8 A X 0.001199f
C9 VPB VGND 0.006067f
C10 VGND VNB 0.687486f
C11 X VNB 0.110387f
C12 VPWR VNB 0.569777f
C13 A VNB 0.298135f
C14 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkbuf_16 VNB VPB VPWR VGND X A
X0 VPWR.t11 a_114_74.t8 X.t27 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 X.t26 a_114_74.t9 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X2 VGND.t15 a_114_74.t10 X.t13 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X.t12 a_114_74.t11 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 X.t11 a_114_74.t12 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5 X.t10 a_114_74.t13 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 a_114_74.t7 A.t0 VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 VPWR.t9 a_114_74.t14 X.t25 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_114_74.t0 A.t1 VGND.t16 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X9 a_114_74.t2 A.t2 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X10 VPWR.t8 a_114_74.t15 X.t24 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VGND.t11 a_114_74.t16 X.t9 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 VPWR.t7 a_114_74.t17 X.t23 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t19 A.t3 a_114_74.t5 VNB.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 X.t8 a_114_74.t18 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X15 X.t22 a_114_74.t19 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 X.t7 a_114_74.t20 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR.t5 a_114_74.t21 X.t21 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VPWR.t4 a_114_74.t22 X.t20 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 X.t6 a_114_74.t23 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X20 VPWR.t13 A.t4 a_114_74.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X21 VGND.t18 A.t5 a_114_74.t4 VNB.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 VGND.t7 a_114_74.t24 X.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 X.t4 a_114_74.t25 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X24 a_114_74.t1 A.t6 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 VGND.t5 a_114_74.t26 X.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 VPWR.t14 A.t7 a_114_74.t6 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 X.t2 a_114_74.t27 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X28 VGND.t3 a_114_74.t28 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X.t19 a_114_74.t29 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X30 VPWR.t2 a_114_74.t30 X.t18 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X31 VGND.t2 a_114_74.t31 X.t16 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 VPWR.t1 a_114_74.t32 X.t17 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X33 VGND.t1 a_114_74.t33 X.t15 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 X.t0 a_114_74.t34 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X35 VGND.t0 a_114_74.t35 X.t14 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 a_114_74.n14 a_114_74.t30 269.652
R1 a_114_74.n16 a_114_74.n13 269.652
R2 a_114_74.n2 a_114_74.t14 269.652
R3 a_114_74.n12 a_114_74.n11 269.652
R4 a_114_74.n20 a_114_74.t15 269.652
R5 a_114_74.n3 a_114_74.n10 269.652
R6 a_114_74.n23 a_114_74.t17 269.652
R7 a_114_74.n25 a_114_74.n9 269.652
R8 a_114_74.n29 a_114_74.t22 269.652
R9 a_114_74.n27 a_114_74.t19 269.652
R10 a_114_74.n32 a_114_74.t21 269.652
R11 a_114_74.n34 a_114_74.t29 269.652
R12 a_114_74.n37 a_114_74.t32 269.652
R13 a_114_74.n39 a_114_74.t34 269.652
R14 a_114_74.n43 a_114_74.t8 269.652
R15 a_114_74.n41 a_114_74.t9 269.652
R16 a_114_74.n7 a_114_74.n5 257.267
R17 a_114_74.n46 a_114_74.n4 248.405
R18 a_114_74.n7 a_114_74.n6 209.833
R19 a_114_74.n47 a_114_74.n46 205.486
R20 a_114_74.n41 a_114_74.t12 198.204
R21 a_114_74.n14 a_114_74.t28 198.204
R22 a_114_74.n42 a_114_74.t33 196.013
R23 a_114_74.n40 a_114_74.t11 196.013
R24 a_114_74.n38 a_114_74.t26 196.013
R25 a_114_74.n35 a_114_74.t20 196.013
R26 a_114_74.n33 a_114_74.t24 196.013
R27 a_114_74.n8 a_114_74.t18 196.013
R28 a_114_74.n28 a_114_74.t10 196.013
R29 a_114_74.n26 a_114_74.t27 196.013
R30 a_114_74.n24 a_114_74.t35 196.013
R31 a_114_74.n3 a_114_74.t25 196.013
R32 a_114_74.n21 a_114_74.t16 196.013
R33 a_114_74.n17 a_114_74.t13 196.013
R34 a_114_74.n2 a_114_74.t31 196.013
R35 a_114_74.n15 a_114_74.t23 196.013
R36 a_114_74.n1 a_114_74.n44 164.144
R37 a_114_74.n0 a_114_74.n18 164.133
R38 a_114_74.n19 a_114_74.n0 163.627
R39 a_114_74.n22 a_114_74.n0 163.627
R40 a_114_74.n1 a_114_74.n30 163.627
R41 a_114_74.n31 a_114_74.n1 163.627
R42 a_114_74.n36 a_114_74.n1 163.627
R43 a_114_74.n46 a_114_74.n45 65.491
R44 a_114_74.n2 a_114_74.n17 62.0763
R45 a_114_74.n3 a_114_74.n21 62.0763
R46 a_114_74.n15 a_114_74.n14 60.6157
R47 a_114_74.n42 a_114_74.n41 60.6157
R48 a_114_74.n25 a_114_74.n24 57.6944
R49 a_114_74.n39 a_114_74.n38 54.7732
R50 a_114_74.n28 a_114_74.n27 53.3126
R51 a_114_74.n34 a_114_74.n33 48.9308
R52 a_114_74.n30 a_114_74.n26 43.0884
R53 a_114_74.n22 a_114_74.n3 42.3581
R54 a_114_74.n31 a_114_74.n8 40.8975
R55 a_114_74.n5 a_114_74.t4 40.0005
R56 a_114_74.n5 a_114_74.t0 40.0005
R57 a_114_74.n6 a_114_74.t5 40.0005
R58 a_114_74.n6 a_114_74.t2 40.0005
R59 a_114_74.n19 a_114_74.n12 37.9763
R60 a_114_74.n18 a_114_74.n16 36.5157
R61 a_114_74.n45 a_114_74.n7 36.5028
R62 a_114_74.n18 a_114_74.n2 32.1338
R63 a_114_74.n44 a_114_74.n43 29.9429
R64 a_114_74.n20 a_114_74.n19 27.752
R65 a_114_74.n36 a_114_74.n35 27.752
R66 a_114_74.n44 a_114_74.n40 27.752
R67 a_114_74.n4 a_114_74.t6 26.3844
R68 a_114_74.n4 a_114_74.t7 26.3844
R69 a_114_74.n47 a_114_74.t3 26.3844
R70 a_114_74.t1 a_114_74.n47 26.3844
R71 a_114_74.n37 a_114_74.n36 24.1005
R72 a_114_74.n23 a_114_74.n22 23.3702
R73 a_114_74.n30 a_114_74.n29 17.5278
R74 a_114_74.n33 a_114_74.n32 16.7975
R75 a_114_74.n32 a_114_74.n31 15.3369
R76 a_114_74.n35 a_114_74.n34 13.8763
R77 a_114_74.n29 a_114_74.n28 12.4157
R78 a_114_74.n38 a_114_74.n37 10.955
R79 a_114_74.n45 a_114_74.n1 9.77876
R80 a_114_74.n27 a_114_74.n8 9.49444
R81 a_114_74.n24 a_114_74.n23 8.03383
R82 a_114_74.n40 a_114_74.n39 8.03383
R83 a_114_74.n16 a_114_74.n15 5.11262
R84 a_114_74.n26 a_114_74.n25 5.11262
R85 a_114_74.n43 a_114_74.n42 5.11262
R86 a_114_74.n17 a_114_74.n12 3.65202
R87 a_114_74.n21 a_114_74.n20 3.65202
R88 a_114_74.n1 a_114_74.n0 2.438
R89 X.n17 X.n15 282.548
R90 X.n21 X.n19 266.019
R91 X.n13 X.n11 263.05
R92 X.n3 X.n2 259.947
R93 X.n1 X.n0 259.716
R94 X.n6 X.n5 259.281
R95 X.n9 X.n8 258.664
R96 X.n25 X.n24 253.141
R97 X.n9 X.t23 233.202
R98 X.n6 X.t24 233.202
R99 X.n3 X.t25 232.933
R100 X.n1 X.t18 232.428
R101 X.n17 X.n16 207.101
R102 X.n21 X.n20 206.819
R103 X.n13 X.n12 206.548
R104 X.n25 X.n23 205.381
R105 X.n24 X.t15 40.0005
R106 X.n24 X.t11 40.0005
R107 X.n19 X.t3 40.0005
R108 X.n19 X.t12 40.0005
R109 X.n15 X.t5 40.0005
R110 X.n15 X.t7 40.0005
R111 X.n11 X.t13 40.0005
R112 X.n11 X.t8 40.0005
R113 X.n8 X.t14 40.0005
R114 X.n8 X.t2 40.0005
R115 X.n5 X.t9 40.0005
R116 X.n5 X.t4 40.0005
R117 X.n2 X.t16 40.0005
R118 X.n2 X.t10 40.0005
R119 X.n0 X.t1 40.0005
R120 X.n0 X.t6 40.0005
R121 X.n23 X.t27 26.3844
R122 X.n23 X.t26 26.3844
R123 X.n20 X.t17 26.3844
R124 X.n20 X.t0 26.3844
R125 X.n16 X.t21 26.3844
R126 X.n16 X.t19 26.3844
R127 X.n12 X.t20 26.3844
R128 X.n12 X.t22 26.3844
R129 X.n4 X.n1 10.8256
R130 X.n18 X.n17 10.4339
R131 X.n22 X.n21 10.4047
R132 X.n10 X.n9 10.4047
R133 X.n7 X.n6 10.4047
R134 X.n14 X.n13 10.377
R135 X.n4 X.n3 10.377
R136 X.n26 X.n25 10.1332
R137 X.n18 X.n14 0.497783
R138 X.n7 X.n4 0.48963
R139 X.n10 X.n7 0.48963
R140 X.n14 X.n10 0.48963
R141 X.n26 X.n22 0.48963
R142 X.n22 X.n18 0.481478
R143 X X.n26 0.0847391
R144 VPWR.n41 VPWR.n1 331.5
R145 VPWR.n36 VPWR.n4 323.406
R146 VPWR.n43 VPWR.t15 257.433
R147 VPWR.n14 VPWR.t2 255.337
R148 VPWR.n22 VPWR.t4 248.744
R149 VPWR.n21 VPWR.t7 248.744
R150 VPWR.n13 VPWR.t8 248.744
R151 VPWR.n15 VPWR.t9 248.744
R152 VPWR.n34 VPWR.n6 222.486
R153 VPWR.n8 VPWR.n7 222.361
R154 VPWR.n28 VPWR.n10 222.361
R155 VPWR.n40 VPWR.n2 36.1417
R156 VPWR.n30 VPWR.n29 36.1417
R157 VPWR.n27 VPWR.n11 36.1417
R158 VPWR.n42 VPWR.n41 35.0123
R159 VPWR.n34 VPWR.n33 33.1299
R160 VPWR.n23 VPWR.n21 32.377
R161 VPWR.n36 VPWR.n35 29.3652
R162 VPWR.n4 VPWR.t10 28.1434
R163 VPWR.n20 VPWR.n13 27.8593
R164 VPWR.n1 VPWR.t12 26.3844
R165 VPWR.n1 VPWR.t14 26.3844
R166 VPWR.n4 VPWR.t13 26.3844
R167 VPWR.n6 VPWR.t0 26.3844
R168 VPWR.n6 VPWR.t11 26.3844
R169 VPWR.n7 VPWR.t3 26.3844
R170 VPWR.n7 VPWR.t1 26.3844
R171 VPWR.n10 VPWR.t6 26.3844
R172 VPWR.n10 VPWR.t5 26.3844
R173 VPWR.n43 VPWR.n42 26.3534
R174 VPWR.n36 VPWR.n2 24.0946
R175 VPWR.n16 VPWR.n15 23.3417
R176 VPWR.n16 VPWR.n13 19.577
R177 VPWR.n21 VPWR.n20 15.0593
R178 VPWR.n35 VPWR.n34 14.3064
R179 VPWR.n23 VPWR.n22 10.5417
R180 VPWR.n33 VPWR.n8 9.78874
R181 VPWR.n17 VPWR.n16 9.3005
R182 VPWR.n18 VPWR.n13 9.3005
R183 VPWR.n20 VPWR.n19 9.3005
R184 VPWR.n21 VPWR.n12 9.3005
R185 VPWR.n24 VPWR.n23 9.3005
R186 VPWR.n25 VPWR.n11 9.3005
R187 VPWR.n27 VPWR.n26 9.3005
R188 VPWR.n29 VPWR.n9 9.3005
R189 VPWR.n31 VPWR.n30 9.3005
R190 VPWR.n33 VPWR.n32 9.3005
R191 VPWR.n34 VPWR.n5 9.3005
R192 VPWR.n35 VPWR.n3 9.3005
R193 VPWR.n37 VPWR.n36 9.3005
R194 VPWR.n38 VPWR.n2 9.3005
R195 VPWR.n40 VPWR.n39 9.3005
R196 VPWR.n42 VPWR.n0 9.3005
R197 VPWR.n44 VPWR.n43 9.3005
R198 VPWR.n15 VPWR.n14 6.62873
R199 VPWR.n28 VPWR.n27 6.02403
R200 VPWR.n29 VPWR.n28 5.27109
R201 VPWR.n30 VPWR.n8 1.50638
R202 VPWR.n41 VPWR.n40 1.12991
R203 VPWR.n22 VPWR.n11 0.753441
R204 VPWR.n17 VPWR.n14 0.665573
R205 VPWR.n18 VPWR.n17 0.122949
R206 VPWR.n19 VPWR.n18 0.122949
R207 VPWR.n19 VPWR.n12 0.122949
R208 VPWR.n24 VPWR.n12 0.122949
R209 VPWR.n25 VPWR.n24 0.122949
R210 VPWR.n26 VPWR.n25 0.122949
R211 VPWR.n26 VPWR.n9 0.122949
R212 VPWR.n31 VPWR.n9 0.122949
R213 VPWR.n32 VPWR.n31 0.122949
R214 VPWR.n32 VPWR.n5 0.122949
R215 VPWR.n5 VPWR.n3 0.122949
R216 VPWR.n37 VPWR.n3 0.122949
R217 VPWR.n38 VPWR.n37 0.122949
R218 VPWR.n39 VPWR.n38 0.122949
R219 VPWR.n39 VPWR.n0 0.122949
R220 VPWR.n44 VPWR.n0 0.122949
R221 VPWR VPWR.n44 0.0617245
R222 VPB.t9 VPB.t2 469.892
R223 VPB.t8 VPB.t9 459.678
R224 VPB.t7 VPB.t8 459.678
R225 VPB.t4 VPB.t7 459.678
R226 VPB VPB.t15 260.485
R227 VPB.t13 VPB.t10 234.946
R228 VPB.t6 VPB.t4 229.839
R229 VPB.t5 VPB.t6 229.839
R230 VPB.t3 VPB.t5 229.839
R231 VPB.t1 VPB.t3 229.839
R232 VPB.t0 VPB.t1 229.839
R233 VPB.t11 VPB.t0 229.839
R234 VPB.t10 VPB.t11 229.839
R235 VPB.t12 VPB.t13 229.839
R236 VPB.t14 VPB.t12 229.839
R237 VPB.t15 VPB.t14 229.839
R238 VGND.n45 VGND.t16 254.696
R239 VGND.n12 VGND.t3 254.125
R240 VGND.n36 VGND.n4 217.376
R241 VGND.n30 VGND.n29 216.858
R242 VGND.n43 VGND.n2 214.696
R243 VGND.n28 VGND.n27 207.647
R244 VGND.n39 VGND.n38 207.498
R245 VGND.n14 VGND.n13 204.976
R246 VGND.n11 VGND.n10 204.976
R247 VGND.n21 VGND.n20 204.976
R248 VGND.n8 VGND.n7 204.976
R249 VGND.n13 VGND.t8 60.0005
R250 VGND.n10 VGND.t12 60.0005
R251 VGND.n20 VGND.t6 60.0005
R252 VGND.n7 VGND.t4 60.0005
R253 VGND.n27 VGND.t10 60.0005
R254 VGND.n38 VGND.t13 60.0005
R255 VGND.n2 VGND.t17 45.7148
R256 VGND.n13 VGND.t2 40.0005
R257 VGND.n10 VGND.t11 40.0005
R258 VGND.n20 VGND.t0 40.0005
R259 VGND.n7 VGND.t15 40.0005
R260 VGND.n27 VGND.t7 40.0005
R261 VGND.n29 VGND.t9 40.0005
R262 VGND.n29 VGND.t5 40.0005
R263 VGND.n4 VGND.t14 40.0005
R264 VGND.n4 VGND.t1 40.0005
R265 VGND.n38 VGND.t19 40.0005
R266 VGND.n2 VGND.t18 40.0005
R267 VGND.n35 VGND.n5 36.1417
R268 VGND.n39 VGND.n37 34.2593
R269 VGND.n43 VGND.n1 34.2593
R270 VGND.n31 VGND.n28 32.377
R271 VGND.n26 VGND.n8 29.7417
R272 VGND.n22 VGND.n21 27.4829
R273 VGND.n45 VGND.n44 26.7299
R274 VGND.n19 VGND.n11 25.224
R275 VGND.n37 VGND.n36 23.3417
R276 VGND.n15 VGND.n14 22.9652
R277 VGND.n15 VGND.n11 22.2123
R278 VGND.n21 VGND.n19 19.9534
R279 VGND.n44 VGND.n43 19.2005
R280 VGND.n22 VGND.n8 17.6946
R281 VGND.n28 VGND.n26 15.4358
R282 VGND.n31 VGND.n30 13.9299
R283 VGND.n39 VGND.n1 13.177
R284 VGND.n36 VGND.n35 12.8005
R285 VGND.n46 VGND.n45 9.3005
R286 VGND.n16 VGND.n15 9.3005
R287 VGND.n17 VGND.n11 9.3005
R288 VGND.n19 VGND.n18 9.3005
R289 VGND.n21 VGND.n9 9.3005
R290 VGND.n23 VGND.n22 9.3005
R291 VGND.n24 VGND.n8 9.3005
R292 VGND.n26 VGND.n25 9.3005
R293 VGND.n28 VGND.n6 9.3005
R294 VGND.n32 VGND.n31 9.3005
R295 VGND.n33 VGND.n5 9.3005
R296 VGND.n35 VGND.n34 9.3005
R297 VGND.n37 VGND.n3 9.3005
R298 VGND.n40 VGND.n39 9.3005
R299 VGND.n41 VGND.n1 9.3005
R300 VGND.n43 VGND.n42 9.3005
R301 VGND.n44 VGND.n0 9.3005
R302 VGND.n14 VGND.n12 6.6595
R303 VGND.n30 VGND.n5 5.27109
R304 VGND.n16 VGND.n12 0.655456
R305 VGND.n17 VGND.n16 0.122949
R306 VGND.n18 VGND.n17 0.122949
R307 VGND.n18 VGND.n9 0.122949
R308 VGND.n23 VGND.n9 0.122949
R309 VGND.n24 VGND.n23 0.122949
R310 VGND.n25 VGND.n24 0.122949
R311 VGND.n25 VGND.n6 0.122949
R312 VGND.n32 VGND.n6 0.122949
R313 VGND.n33 VGND.n32 0.122949
R314 VGND.n34 VGND.n33 0.122949
R315 VGND.n34 VGND.n3 0.122949
R316 VGND.n40 VGND.n3 0.122949
R317 VGND.n41 VGND.n40 0.122949
R318 VGND.n42 VGND.n41 0.122949
R319 VGND.n42 VGND.n0 0.122949
R320 VGND.n46 VGND.n0 0.122949
R321 VGND VGND.n46 0.0617245
R322 VNB.t2 VNB.t8 1154.86
R323 VNB.t11 VNB.t12 1154.86
R324 VNB.t0 VNB.t6 1154.86
R325 VNB.t15 VNB.t4 1154.86
R326 VNB.t7 VNB.t10 1154.86
R327 VNB.t19 VNB.t13 1154.86
R328 VNB VNB.t16 1143.31
R329 VNB.t18 VNB.t17 1039.37
R330 VNB.t8 VNB.t3 993.177
R331 VNB.t12 VNB.t2 993.177
R332 VNB.t6 VNB.t11 993.177
R333 VNB.t4 VNB.t0 993.177
R334 VNB.t10 VNB.t15 993.177
R335 VNB.t9 VNB.t7 993.177
R336 VNB.t5 VNB.t9 993.177
R337 VNB.t14 VNB.t5 993.177
R338 VNB.t1 VNB.t14 993.177
R339 VNB.t13 VNB.t1 993.177
R340 VNB.t17 VNB.t19 993.177
R341 VNB.t16 VNB.t18 993.177
R342 A.n4 A.t1 249.619
R343 A.n8 A.t5 247.428
R344 A.n3 A.t2 247.428
R345 A.n0 A.t3 247.428
R346 A.n0 A.t4 234.841
R347 A.n2 A.t6 226.809
R348 A.n9 A.t7 226.809
R349 A.n4 A.t0 226.809
R350 A A.n1 152.298
R351 A.n11 A.n10 152
R352 A.n8 A.n7 152
R353 A.n6 A.n5 152
R354 A.n8 A.n5 49.6611
R355 A.n10 A.n9 44.549
R356 A.n1 A.n0 29.2126
R357 A.n2 A.n1 28.4823
R358 A.n10 A.n3 16.0672
R359 A.n6 A 12.8005
R360 A.n5 A.n4 10.955
R361 A A.n11 9.82376
R362 A.n7 A 8.63306
R363 A.n7 A 5.65631
R364 A.n3 A.n2 5.11262
R365 A.n9 A.n8 5.11262
R366 A.n11 A 4.46562
R367 A A.n6 1.48887
C0 VPB A 0.138577f
C1 VPB VPWR 0.261252f
C2 A VPWR 0.09178f
C3 VPB X 0.052418f
C4 A X 0.002012f
C5 VPB VGND 0.007898f
C6 VPWR X 1.85268f
C7 A VGND 0.079105f
C8 VPWR VGND 0.071786f
C9 X VGND 0.700464f
C10 VGND VNB 1.1887f
C11 X VNB 0.148395f
C12 VPWR VNB 0.949526f
C13 A VNB 0.527453f
C14 VPB VNB 2.22754f
.ends

* NGSPICE file created from sky130_fd_sc_hs__clkdlyinv3sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkdlyinv3sd1_1 VNB VPB VPWR VGND A Y
X0 Y.t0 a_285_392.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 Y.t1 a_285_392.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.308 ps=2.79 w=1.12 l=0.15
X2 VGND.t1 A.t0 a_28_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.15435 pd=1.155 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 VPWR.t1 A.t1 a_28_74.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3684 pd=1.825 as=0.3136 ps=2.8 w=1.12 l=0.15
X4 a_285_392.t1 a_28_74.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.28 pd=2.56 as=0.3684 ps=1.825 w=1 l=0.15
X5 a_285_392.t0 a_28_74.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0.15435 ps=1.155 w=0.42 l=0.15
R0 a_285_392.n0 a_285_392.t3 265.637
R1 a_285_392.n1 a_285_392.t0 262.938
R2 a_285_392.t1 a_285_392.n1 257.397
R3 a_285_392.n0 a_285_392.t2 253.853
R4 a_285_392.n1 a_285_392.n0 177.794
R5 VGND.n1 VGND.t0 253.761
R6 VGND.n1 VGND.n0 212.68
R7 VGND.n0 VGND.t2 154.286
R8 VGND.n0 VGND.t1 55.7148
R9 VGND VGND.n1 0.263065
R10 Y.n1 Y 589.268
R11 Y.n1 Y.n0 585
R12 Y.n2 Y.n1 585
R13 Y.n3 Y.t0 225
R14 Y.n1 Y.t1 27.2639
R15 Y.n2 Y 11.9116
R16 Y Y.n3 9.97283
R17 Y.n0 Y 9.24494
R18 Y.n3 Y 4.26717
R19 Y.n0 Y 3.91161
R20 Y Y.n2 1.24494
R21 VNB.t2 VNB.t0 2194.23
R22 VNB.t1 VNB.t2 2044.09
R23 VNB VNB.t1 1108.66
R24 VPWR.n1 VPWR.n0 321.021
R25 VPWR.n1 VPWR.t0 256.077
R26 VPWR.n0 VPWR.t2 105.395
R27 VPWR.n0 VPWR.t1 31.6309
R28 VPWR VPWR.n1 0.260042
R29 VPB.t2 VPB.t0 497.985
R30 VPB.t1 VPB.t2 436.695
R31 VPB VPB.t1 252.823
R32 A.n0 A.t1 293.752
R33 A.n0 A.t0 220.113
R34 A A.n0 159.929
R35 a_28_74.t0 a_28_74.n1 448.507
R36 a_28_74.n0 a_28_74.t2 338.438
R37 a_28_74.n1 a_28_74.t1 289.522
R38 a_28_74.n0 a_28_74.t3 193.838
R39 a_28_74.n1 a_28_74.n0 152
C0 VPWR VGND 0.050205f
C1 Y VGND 0.073742f
C2 VPB A 0.041909f
C3 VPB VPWR 0.094064f
C4 A VPWR 0.021276f
C5 VPB Y 0.019107f
C6 VPB VGND 0.006931f
C7 VPWR Y 0.14736f
C8 A VGND 0.017461f
C9 VGND VNB 0.394438f
C10 Y VNB 0.124951f
C11 VPWR VNB 0.311738f
C12 A VNB 0.209054f
C13 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a31o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31o_2 VNB VPB VPWR VGND A1 A2 A3 B1 X
X0 VPWR.t1 a_97_296.t3 X.t3 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3064 pd=1.68 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t2 A2.t0 a_362_368.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.245 pd=1.49 as=0.15 ps=1.3 w=1 l=0.15
X2 X.t1 a_97_296.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2627 ps=2.19 w=0.74 l=0.15
X3 X.t2 a_97_296.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4 a_362_368.t1 A3.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.3064 ps=1.68 w=1 l=0.15
X5 a_97_296.t0 B1.t0 a_362_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.175 ps=1.35 w=1 l=0.15
X6 a_449_74.t1 A2.t1 a_371_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X7 a_371_74.t0 A3.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.23495 ps=1.375 w=0.74 l=0.15
X8 VGND.t2 B1.t1 a_97_296.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 VGND.t0 a_97_296.t6 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.23495 pd=1.375 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_362_368.t2 A1.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.245 ps=1.49 w=1 l=0.15
X11 a_97_296.t2 A1.t1 a_449_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
R0 a_97_296.t0 a_97_296.n4 415.406
R1 a_97_296.n4 a_97_296.n0 247.09
R2 a_97_296.n1 a_97_296.t5 240.98
R3 a_97_296.n3 a_97_296.t3 240.197
R4 a_97_296.n1 a_97_296.t4 181.387
R5 a_97_296.n2 a_97_296.t6 179.947
R6 a_97_296.n4 a_97_296.n3 165.876
R7 a_97_296.n2 a_97_296.n1 61.3654
R8 a_97_296.n0 a_97_296.t1 35.6762
R9 a_97_296.n0 a_97_296.t2 32.4329
R10 a_97_296.n3 a_97_296.n2 4.38232
R11 X.n2 X 590.08
R12 X.n2 X.n0 585
R13 X.n3 X.n2 585
R14 X X.n1 162.373
R15 X.n2 X.t3 26.3844
R16 X.n2 X.t2 26.3844
R17 X.n1 X.t0 22.7032
R18 X.n1 X.t1 22.7032
R19 X X.n3 13.6132
R20 X X.n0 11.7846
R21 X X.n0 3.25129
R22 X.n3 X 1.42272
R23 VPWR.n2 VPWR.n1 620.36
R24 VPWR.n6 VPWR.t0 259.171
R25 VPWR.n4 VPWR.n3 202.155
R26 VPWR.n3 VPWR.t3 60.2627
R27 VPWR.n1 VPWR.t2 50.2355
R28 VPWR.n1 VPWR.t4 46.2955
R29 VPWR.n3 VPWR.t1 39.876
R30 VPWR.n5 VPWR.n4 27.8593
R31 VPWR.n6 VPWR.n5 21.4593
R32 VPWR.n5 VPWR.n0 9.3005
R33 VPWR.n7 VPWR.n6 9.3005
R34 VPWR.n4 VPWR.n2 4.97951
R35 VPWR.n2 VPWR.n0 0.366107
R36 VPWR.n7 VPWR.n0 0.122949
R37 VPWR VPWR.n7 0.0617245
R38 VPB.t1 VPB.t4 362.635
R39 VPB.t2 VPB.t5 326.882
R40 VPB VPB.t0 293.683
R41 VPB.t5 VPB.t3 255.376
R42 VPB.t4 VPB.t2 229.839
R43 VPB.t0 VPB.t1 229.839
R44 A2.n0 A2.t0 266.44
R45 A2.n0 A2.t1 178.34
R46 A2 A2.n0 158.4
R47 a_362_368.n1 a_362_368.n0 653.878
R48 a_362_368.t0 a_362_368.n1 39.4005
R49 a_362_368.n0 a_362_368.t3 29.5505
R50 a_362_368.n0 a_362_368.t1 29.5505
R51 a_362_368.n1 a_362_368.t2 29.5505
R52 VGND.n2 VGND.n1 185
R53 VGND.n4 VGND.n3 185
R54 VGND.n9 VGND.t1 154.727
R55 VGND.n5 VGND.t2 145.576
R56 VGND.n3 VGND.n2 55.1356
R57 VGND.n8 VGND.n7 28.2166
R58 VGND.n2 VGND.t0 25.1356
R59 VGND.n3 VGND.t3 22.7032
R60 VGND.n9 VGND.n8 20.7064
R61 VGND.n5 VGND.n4 9.69319
R62 VGND.n10 VGND.n9 9.3005
R63 VGND.n7 VGND.n6 9.3005
R64 VGND.n8 VGND.n0 9.3005
R65 VGND.n4 VGND.n1 6.35378
R66 VGND.n7 VGND.n1 0.467653
R67 VGND.n6 VGND.n5 0.164396
R68 VGND.n6 VGND.n0 0.122949
R69 VGND.n10 VGND.n0 0.122949
R70 VGND VGND.n10 0.0617245
R71 VNB.t0 VNB.t4 1813.12
R72 VNB.t3 VNB.t2 1316.54
R73 VNB.t5 VNB.t3 1316.54
R74 VNB VNB.t1 1304.99
R75 VNB.t1 VNB.t0 993.177
R76 VNB.t4 VNB.t5 900.788
R77 A3.n0 A3.t0 266.44
R78 A3.n0 A3.t1 178.34
R79 A3 A3.n0 158.788
R80 B1.n0 B1.t0 258.245
R81 B1.n0 B1.t1 170.147
R82 B1 B1.n0 158.788
R83 a_371_74.t0 a_371_74.t1 38.9194
R84 a_449_74.t0 a_449_74.t1 68.1086
R85 A1.n0 A1.t0 266.44
R86 A1.n0 A1.t1 178.34
R87 A1 A1.n0 159.093
C0 VPWR X 0.213692f
C1 VPB A3 0.03453f
C2 X B1 6.68e-20
C3 VPWR A3 0.016693f
C4 VPB A2 0.031947f
C5 A2 A1 0.070301f
C6 X VGND 0.122704f
C7 VPB A1 0.032964f
C8 VPWR A2 0.011945f
C9 A3 VGND 0.015608f
C10 VPB VPWR 0.127345f
C11 VPB B1 0.041127f
C12 VPWR A1 0.014224f
C13 A1 B1 0.088108f
C14 A2 VGND 0.008971f
C15 VPB VGND 0.009683f
C16 VPWR B1 0.010209f
C17 A1 VGND 0.012007f
C18 VPWR VGND 0.077066f
C19 B1 VGND 0.05074f
C20 X A3 0.001363f
C21 X A2 5.67e-19
C22 VPB X 0.005782f
C23 A3 A2 0.090744f
C24 X A1 2.85e-19
C25 VGND VNB 0.555518f
C26 B1 VNB 0.16948f
C27 A1 VNB 0.110722f
C28 A2 VNB 0.106125f
C29 A3 VNB 0.108479f
C30 X VNB 0.029057f
C31 VPWR VNB 0.429929f
C32 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a31o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31o_4 VNB VPB VPWR VGND A1 A2 A3 B1 X
X0 VGND.t5 a_83_274.t6 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.11285 ps=1.045 w=0.74 l=0.15
X1 X.t3 a_83_274.t7 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VPWR.t5 a_83_274.t8 X.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VGND.t0 B1.t0 a_83_274.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.1824 ps=1.85 w=0.64 l=0.15
X4 X.t1 a_83_274.t9 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X5 a_529_392.t1 A3.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X6 X.t6 a_83_274.t10 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.2294 ps=2.1 w=0.74 l=0.15
X7 a_83_274.t5 A1.t0 a_775_74.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2272 pd=1.99 as=0.112 ps=0.99 w=0.64 l=0.15
X8 a_1000_74.t0 A3.t1 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 VPWR.t9 A3.t2 a_529_392.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X10 VPWR.t8 A1.t1 a_529_392.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.225 ps=1.45 w=1 l=0.15
X11 a_1000_74.t2 A2.t0 a_775_74.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X12 X.t5 a_83_274.t11 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_775_74.t1 A1.t2 a_83_274.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X14 a_83_274.t1 B1.t1 a_529_392.t4 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.185 pd=1.37 as=0.295 ps=2.59 w=1 l=0.15
X15 VPWR.t3 a_83_274.t12 X.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_529_392.t6 A2.t1 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.205 ps=1.41 w=1 l=0.15
X17 a_775_74.t0 A2.t2 a_1000_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X18 VGND.t2 a_83_274.t13 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X19 a_83_274.t2 B1.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.112 ps=0.99 w=0.64 l=0.15
X20 a_529_392.t5 A1.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X21 VPWR.t1 A2.t3 a_529_392.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.205 pd=1.41 as=0.15 ps=1.3 w=1 l=0.15
X22 a_529_392.t3 B1.t3 a_83_274.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
R0 a_83_274.n17 a_83_274.n16 349.212
R1 a_83_274.n1 a_83_274.t5 295.774
R2 a_83_274.n4 a_83_274.t7 264.413
R3 a_83_274.n13 a_83_274.t8 261.62
R4 a_83_274.n10 a_83_274.t9 261.62
R5 a_83_274.n5 a_83_274.t12 261.62
R6 a_83_274.n14 a_83_274.n13 183.404
R7 a_83_274.n8 a_83_274.n7 165.189
R8 a_83_274.n4 a_83_274.t10 154.24
R9 a_83_274.n6 a_83_274.t13 154.24
R10 a_83_274.n3 a_83_274.t11 154.24
R11 a_83_274.n12 a_83_274.t6 154.24
R12 a_83_274.n9 a_83_274.n8 152
R13 a_83_274.n11 a_83_274.n2 152
R14 a_83_274.n15 a_83_274.t0 151.594
R15 a_83_274.n1 a_83_274.n0 108.046
R16 a_83_274.n5 a_83_274.n4 63.5369
R17 a_83_274.n16 a_83_274.n15 56.4711
R18 a_83_274.n11 a_83_274.n10 47.4702
R19 a_83_274.t1 a_83_274.n17 41.3705
R20 a_83_274.n7 a_83_274.n3 40.1672
R21 a_83_274.n17 a_83_274.t3 31.5205
R22 a_83_274.n0 a_83_274.t4 26.2505
R23 a_83_274.n0 a_83_274.t2 26.2505
R24 a_83_274.n7 a_83_274.n6 22.6399
R25 a_83_274.n15 a_83_274.n14 16.6997
R26 a_83_274.n8 a_83_274.n2 13.1884
R27 a_83_274.n13 a_83_274.n12 10.955
R28 a_83_274.n14 a_83_274.n2 10.9027
R29 a_83_274.n9 a_83_274.n3 9.49444
R30 a_83_274.n12 a_83_274.n11 7.30353
R31 a_83_274.n6 a_83_274.n5 5.84292
R32 a_83_274.n16 a_83_274.n1 3.54021
R33 a_83_274.n10 a_83_274.n9 2.19141
R34 X.n6 X 589.85
R35 X.n6 X.n0 585
R36 X.n7 X.n6 585
R37 X.n5 X.n1 261.149
R38 X.n4 X.n3 158.095
R39 X.n4 X.n2 96.7184
R40 X X.n4 32.3216
R41 X.n2 X.t6 30.0005
R42 X.n3 X.t7 26.7573
R43 X.n6 X.t0 26.3844
R44 X.n6 X.t3 26.3844
R45 X.n1 X.t2 26.3844
R46 X.n1 X.t1 26.3844
R47 X.n2 X.t4 22.7032
R48 X.n3 X.t5 22.7032
R49 X X.n7 12.9944
R50 X X.n0 11.249
R51 X.n5 X 8.72777
R52 X X.n5 5.62474
R53 X X.n0 3.10353
R54 X.n7 X 1.35808
R55 VGND.n12 VGND.n2 206.916
R56 VGND.n14 VGND.t4 160.254
R57 VGND.n4 VGND.t6 158.029
R58 VGND.n8 VGND.t5 138.363
R59 VGND.n6 VGND.n5 114.883
R60 VGND.n5 VGND.t1 39.3755
R61 VGND.n8 VGND.n7 28.6123
R62 VGND.n5 VGND.t0 26.2505
R63 VGND.n13 VGND.n12 24.4711
R64 VGND.n12 VGND.n1 22.9652
R65 VGND.n2 VGND.t3 22.7032
R66 VGND.n2 VGND.t2 22.7032
R67 VGND.n7 VGND.n6 21.0829
R68 VGND.n14 VGND.n13 20.7064
R69 VGND.n8 VGND.n1 18.824
R70 VGND.n15 VGND.n14 9.3005
R71 VGND.n7 VGND.n3 9.3005
R72 VGND.n9 VGND.n8 9.3005
R73 VGND.n10 VGND.n1 9.3005
R74 VGND.n12 VGND.n11 9.3005
R75 VGND.n13 VGND.n0 9.3005
R76 VGND.n6 VGND.n4 7.27857
R77 VGND.n4 VGND.n3 0.155399
R78 VGND.n9 VGND.n3 0.122949
R79 VGND.n10 VGND.n9 0.122949
R80 VGND.n11 VGND.n10 0.122949
R81 VGND.n11 VGND.n0 0.122949
R82 VGND.n15 VGND.n0 0.122949
R83 VGND VGND.n15 0.0617245
R84 VNB.t8 VNB.t0 2448.29
R85 VNB.t7 VNB.t1 2286.61
R86 VNB.t9 VNB.t10 1986.35
R87 VNB VNB.t6 1201.05
R88 VNB.t3 VNB.t8 1154.86
R89 VNB.t1 VNB.t2 1154.86
R90 VNB.t6 VNB.t4 1097.11
R91 VNB.t5 VNB.t7 1050.92
R92 VNB.t0 VNB.t9 993.177
R93 VNB.t2 VNB.t3 993.177
R94 VNB.t4 VNB.t5 993.177
R95 VPWR.n9 VPWR.n8 321.834
R96 VPWR.n13 VPWR.n7 316.211
R97 VPWR.n11 VPWR.n10 316.211
R98 VPWR.n26 VPWR.t6 259.171
R99 VPWR.n3 VPWR.t5 258.875
R100 VPWR.n24 VPWR.n2 221.766
R101 VPWR.n10 VPWR.t7 41.3705
R102 VPWR.n7 VPWR.t2 39.4005
R103 VPWR.n7 VPWR.t8 39.4005
R104 VPWR.n10 VPWR.t1 39.4005
R105 VPWR.n8 VPWR.t0 39.4005
R106 VPWR.n17 VPWR.n5 36.1417
R107 VPWR.n18 VPWR.n17 36.1417
R108 VPWR.n19 VPWR.n18 36.1417
R109 VPWR.n2 VPWR.t4 35.1791
R110 VPWR.n2 VPWR.t3 35.1791
R111 VPWR.n13 VPWR.n12 35.0123
R112 VPWR.n8 VPWR.t9 29.5505
R113 VPWR.n23 VPWR.n3 28.9887
R114 VPWR.n26 VPWR.n25 26.7299
R115 VPWR.n25 VPWR.n24 25.977
R116 VPWR.n24 VPWR.n23 21.4593
R117 VPWR.n19 VPWR.n3 18.4476
R118 VPWR.n12 VPWR.n11 15.4358
R119 VPWR.n13 VPWR.n5 12.424
R120 VPWR.n12 VPWR.n6 9.3005
R121 VPWR.n14 VPWR.n13 9.3005
R122 VPWR.n15 VPWR.n5 9.3005
R123 VPWR.n17 VPWR.n16 9.3005
R124 VPWR.n18 VPWR.n4 9.3005
R125 VPWR.n20 VPWR.n19 9.3005
R126 VPWR.n21 VPWR.n3 9.3005
R127 VPWR.n23 VPWR.n22 9.3005
R128 VPWR.n24 VPWR.n1 9.3005
R129 VPWR.n25 VPWR.n0 9.3005
R130 VPWR.n27 VPWR.n26 9.3005
R131 VPWR.n11 VPWR.n9 7.11161
R132 VPWR.n9 VPWR.n6 0.52313
R133 VPWR.n14 VPWR.n6 0.122949
R134 VPWR.n15 VPWR.n14 0.122949
R135 VPWR.n16 VPWR.n15 0.122949
R136 VPWR.n16 VPWR.n4 0.122949
R137 VPWR.n20 VPWR.n4 0.122949
R138 VPWR.n21 VPWR.n20 0.122949
R139 VPWR.n22 VPWR.n21 0.122949
R140 VPWR.n22 VPWR.n1 0.122949
R141 VPWR.n1 VPWR.n0 0.122949
R142 VPWR.n27 VPWR.n0 0.122949
R143 VPWR VPWR.n27 0.0617245
R144 VPB.t7 VPB.t2 541.399
R145 VPB.t3 VPB.t10 306.452
R146 VPB.t1 VPB.t9 286.022
R147 VPB.t10 VPB.t4 280.914
R148 VPB.t5 VPB.t6 280.914
R149 VPB.t2 VPB.t3 265.591
R150 VPB VPB.t8 257.93
R151 VPB.t11 VPB.t0 255.376
R152 VPB.t9 VPB.t11 255.376
R153 VPB.t4 VPB.t1 229.839
R154 VPB.t6 VPB.t7 229.839
R155 VPB.t8 VPB.t5 229.839
R156 B1.n3 B1.t0 250.641
R157 B1.n0 B1.t2 250.641
R158 B1.n0 B1.t3 238.566
R159 B1.n2 B1.t1 207.529
R160 B1 B1.n3 184.28
R161 B1 B1.n1 153.358
R162 B1.n1 B1.n0 43.8187
R163 B1.n3 B1.n2 21.1793
R164 B1.n2 B1.n1 8.03383
R165 A3.n2 A3.n1 244.214
R166 A3.n0 A3.t1 244.214
R167 A3.n0 A3.t0 219.457
R168 A3.n2 A3.t2 216.536
R169 A3.n3 A3 156.462
R170 A3.n5 A3.n4 152
R171 A3.n4 A3.n3 49.6611
R172 A3 A3.n5 9.89141
R173 A3.n3 A3.n2 8.76414
R174 A3.n5 A3 8.72777
R175 A3.n4 A3.n0 4.38232
R176 a_529_392.n1 a_529_392.t4 310.685
R177 a_529_392.t1 a_529_392.n5 285.483
R178 a_529_392.n3 a_529_392.n2 205.487
R179 a_529_392.n5 a_529_392.n4 205.487
R180 a_529_392.n1 a_529_392.n0 189.115
R181 a_529_392.n3 a_529_392.n1 66.8196
R182 a_529_392.n0 a_529_392.t3 59.1005
R183 a_529_392.n5 a_529_392.n3 51.2005
R184 a_529_392.n4 a_529_392.t0 39.4005
R185 a_529_392.n0 a_529_392.t7 29.5505
R186 a_529_392.n2 a_529_392.t2 29.5505
R187 a_529_392.n2 a_529_392.t5 29.5505
R188 a_529_392.n4 a_529_392.t6 29.5505
R189 A1.n0 A1.t3 232.602
R190 A1.n2 A1.t1 223.839
R191 A1.n1 A1.t2 205.654
R192 A1 A1.n0 154.91
R193 A1.n3 A1.n2 152
R194 A1.n1 A1.t0 137.881
R195 A1.n2 A1.n0 49.6611
R196 A1.n2 A1.n1 42.3581
R197 A1 A1.n3 10.2793
R198 A1.n3 A1 8.33989
R199 a_775_74.n1 a_775_74.n0 290.733
R200 a_775_74.n1 a_775_74.t1 39.3755
R201 a_775_74.n0 a_775_74.t3 26.2505
R202 a_775_74.n0 a_775_74.t0 26.2505
R203 a_775_74.t2 a_775_74.n1 26.2505
R204 a_1000_74.n0 a_1000_74.t1 291.875
R205 a_1000_74.t0 a_1000_74.n0 208.923
R206 a_1000_74.n0 a_1000_74.t2 154.72
R207 A2.n2 A2.t2 263.493
R208 A2.n0 A2.t0 257.36
R209 A2.n2 A2.t3 214.793
R210 A2.n1 A2.t1 212.883
R211 A2 A2.n0 162.28
R212 A2.n4 A2.n3 152
R213 A2.n3 A2.n1 48.9308
R214 A2.n3 A2.n2 30.6732
R215 A2.n4 A2 15.7096
R216 A2 A2.n4 2.90959
R217 A2.n1 A2.n0 0.730803
C0 VPB VGND 0.014257f
C1 B1 X 0.005358f
C2 A2 A3 0.090939f
C3 A1 VPWR 0.035463f
C4 B1 VGND 0.037789f
C5 A2 VPWR 0.037867f
C6 A1 VGND 0.017488f
C7 A3 VPWR 0.039915f
C8 A2 VGND 0.016902f
C9 VPWR X 0.45636f
C10 A3 VGND 0.038938f
C11 VPB B1 0.113838f
C12 VPWR VGND 0.128251f
C13 VPB A1 0.09203f
C14 X VGND 0.26885f
C15 VPB A2 0.088393f
C16 B1 A1 0.048304f
C17 VPB A3 0.085293f
C18 VPB VPWR 0.21512f
C19 A1 A2 0.072276f
C20 B1 VPWR 0.016428f
C21 VPB X 0.013667f
C22 VGND VNB 0.882957f
C23 X VNB 0.040656f
C24 VPWR VNB 0.704893f
C25 A3 VNB 0.257176f
C26 A2 VNB 0.240735f
C27 A1 VNB 0.246288f
C28 B1 VNB 0.25459f
C29 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a31oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31oi_1 VNB VPB VPWR VGND Y A3 B1 A2 A1
X0 VGND.t0 B1.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X1 VPWR.t1 A2.t0 a_136_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2744 pd=1.61 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_136_368.t0 A3.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.4312 ps=3.01 w=1.12 l=0.15
X3 a_145_74.t1 A3.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.3182 ps=2.34 w=0.74 l=0.15
X4 Y.t1 B1.t1 a_136_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.196 ps=1.47 w=1.12 l=0.15
X5 Y.t2 A1.t0 a_223_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X6 a_136_368.t3 A1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2744 ps=1.61 w=1.12 l=0.15
X7 a_223_74.t1 A2.t1 a_145_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
R0 B1.n0 B1.t1 261.62
R1 B1.n0 B1.t0 156.431
R2 B1.n1 B1.n0 95.6291
R3 B1 B1.n1 10.8481
R4 B1.n1 B1 5.49334
R5 Y.n2 Y 588.201
R6 Y.n2 Y.n0 585
R7 Y.n3 Y.n2 585
R8 Y Y.n1 386.252
R9 Y.n1 Y.t0 34.0546
R10 Y.n1 Y.t2 34.0546
R11 Y.n2 Y.t1 26.3844
R12 Y Y.n3 8.5765
R13 Y Y.n0 7.4245
R14 Y Y.n0 2.0485
R15 Y.n3 Y 0.8965
R16 VGND.n0 VGND.t1 169.07
R17 VGND.n0 VGND.t0 162.303
R18 VGND VGND.n0 0.106149
R19 VNB VNB.t1 1501.31
R20 VNB.t2 VNB.t0 1316.54
R21 VNB.t3 VNB.t2 1316.54
R22 VNB.t1 VNB.t3 900.788
R23 A2.n0 A2.t0 285.719
R24 A2.n0 A2.t1 178.34
R25 A2 A2.n0 158.4
R26 a_136_368.n1 a_136_368.n0 461.577
R27 a_136_368.n0 a_136_368.t2 35.1791
R28 a_136_368.n0 a_136_368.t3 26.3844
R29 a_136_368.n1 a_136_368.t1 26.3844
R30 a_136_368.t0 a_136_368.n1 26.3844
R31 VPWR.n1 VPWR.n0 320.866
R32 VPWR.n1 VPWR.t0 272.56
R33 VPWR.n0 VPWR.t2 43.9737
R34 VPWR.n0 VPWR.t1 42.2148
R35 VPWR VPWR.n1 0.375167
R36 VPB.t1 VPB.t3 326.882
R37 VPB VPB.t0 309.005
R38 VPB.t3 VPB.t2 255.376
R39 VPB.t0 VPB.t1 229.839
R40 A3.n0 A3.t0 261.62
R41 A3 A3.n0 204.798
R42 A3.n0 A3.t1 160.814
R43 a_145_74.t0 a_145_74.t1 38.9194
R44 A1.n0 A1.t1 285.719
R45 A1.n0 A1.t0 178.34
R46 A1 A1.n0 158.788
R47 a_223_74.t0 a_223_74.t1 68.1086
C0 VPB A3 0.044691f
C1 VPWR VGND 0.051362f
C2 VPB A2 0.031266f
C3 Y VGND 0.247518f
C4 A3 A2 0.061674f
C5 VPB A1 0.032043f
C6 VPB B1 0.048771f
C7 VPB VPWR 0.089445f
C8 A2 A1 0.074813f
C9 A3 VPWR 0.046862f
C10 A2 B1 4.35e-19
C11 VPB Y 0.031012f
C12 VPB VGND 0.006145f
C13 A1 B1 0.081468f
C14 A2 VPWR 0.017374f
C15 A3 Y 0.057401f
C16 A1 VPWR 0.012652f
C17 A2 Y 0.142573f
C18 A3 VGND 0.045152f
C19 A1 Y 0.070812f
C20 B1 VPWR 0.008698f
C21 A2 VGND 0.01037f
C22 A1 VGND 0.007459f
C23 B1 Y 0.095838f
C24 VPWR Y 0.076544f
C25 B1 VGND 0.058399f
C26 VGND VNB 0.447546f
C27 Y VNB 0.085331f
C28 VPWR VNB 0.349927f
C29 B1 VNB 0.193391f
C30 A1 VNB 0.108173f
C31 A2 VNB 0.111134f
C32 A3 VNB 0.176999f
C33 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a31oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31oi_2 VNB VPB VPWR VGND A2 A1 A3 Y B1
X0 VPWR.t2 A1.t0 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1 Y.t4 B1.t0 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.1554 ps=1.16 w=0.74 l=0.15
X2 VPWR.t4 A3.t0 a_27_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_27_368.t7 A3.t1 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.196 ps=1.47 w=1.12 l=0.15
X4 VGND.t0 A3.t2 a_114_74.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1295 ps=1.09 w=0.74 l=0.15
X5 Y.t0 A1.t1 a_200_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.10915 ps=1.035 w=0.74 l=0.15
X6 a_114_74.t1 A3.t3 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7 VPWR.t3 A2.t0 a_27_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1904 ps=1.46 w=1.12 l=0.15
X8 a_27_368.t4 B1.t1 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t2 B1.t2 a_27_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X10 a_114_74.t0 A2.t1 a_200_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X11 a_200_74.t1 A1.t2 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.24605 ps=1.405 w=0.74 l=0.15
X12 a_200_74.t3 A2.t2 a_114_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_27_368.t0 A2.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1904 pd=1.46 as=0.1736 ps=1.43 w=1.12 l=0.15
X14 a_27_368.t1 A1.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A1.n0 A1.t3 235.571
R1 A1.n1 A1.t0 226.809
R2 A1.n1 A1.t2 205.796
R3 A1.n0 A1.t1 196.013
R4 A1 A1.n2 161.327
R5 A1.n2 A1.n1 54.7732
R6 A1.n2 A1.n0 2.19141
R7 a_27_368.n2 a_27_368.t1 297.808
R8 a_27_368.n4 a_27_368.t6 284.75
R9 a_27_368.n5 a_27_368.n4 203.381
R10 a_27_368.n2 a_27_368.n1 188.19
R11 a_27_368.n3 a_27_368.n0 187.786
R12 a_27_368.n3 a_27_368.n2 101.097
R13 a_27_368.n4 a_27_368.n3 66.8953
R14 a_27_368.n1 a_27_368.t4 35.1791
R15 a_27_368.t0 a_27_368.n5 33.4201
R16 a_27_368.n0 a_27_368.t5 27.2639
R17 a_27_368.n0 a_27_368.t7 27.2639
R18 a_27_368.n1 a_27_368.t2 26.3844
R19 a_27_368.n5 a_27_368.t3 26.3844
R20 VPWR.n5 VPWR.n4 323.406
R21 VPWR.n3 VPWR.n2 321.248
R22 VPWR.n7 VPWR.n1 316.351
R23 VPWR.n4 VPWR.t5 35.1791
R24 VPWR.n6 VPWR.n5 29.7417
R25 VPWR.n1 VPWR.t0 28.1434
R26 VPWR.n1 VPWR.t4 26.3844
R27 VPWR.n4 VPWR.t3 26.3844
R28 VPWR.n2 VPWR.t1 26.3844
R29 VPWR.n2 VPWR.t2 26.3844
R30 VPWR.n7 VPWR.n6 22.9652
R31 VPWR.n6 VPWR.n0 9.3005
R32 VPWR.n8 VPWR.n7 7.27223
R33 VPWR.n5 VPWR.n3 7.13599
R34 VPWR.n3 VPWR.n0 0.169443
R35 VPWR VPWR.n8 0.157962
R36 VPWR.n8 VPWR.n0 0.149814
R37 VPB VPB.t6 257.93
R38 VPB.t4 VPB.t2 255.376
R39 VPB.t3 VPB.t7 255.376
R40 VPB.t0 VPB.t3 250.269
R41 VPB.t7 VPB.t5 234.946
R42 VPB.t6 VPB.t0 234.946
R43 VPB.t2 VPB.t1 229.839
R44 VPB.t5 VPB.t4 229.839
R45 B1.n2 B1.t2 272.574
R46 B1.n0 B1.t1 266.731
R47 B1 B1.n0 161.514
R48 B1 B1.n2 154.25
R49 B1.n1 B1.t0 154.24
R50 B1.n1 B1.n0 48.9308
R51 B1.n2 B1.n1 0.730803
R52 VGND.n1 VGND.t1 252.109
R53 VGND.n1 VGND.n0 210.419
R54 VGND.n0 VGND.t2 34.0546
R55 VGND.n0 VGND.t0 34.0546
R56 VGND VGND.n1 0.103468
R57 Y.n1 Y.n0 331.729
R58 Y.t0 Y.n1 261.057
R59 Y.n2 Y.t0 261.057
R60 Y Y.n3 140.579
R61 Y.n3 Y.t4 50.6233
R62 Y.n3 Y.t1 48.5083
R63 Y.n0 Y.t3 26.3844
R64 Y.n0 Y.t2 26.3844
R65 Y.n2 Y 12.6066
R66 Y.n1 Y 4.84898
R67 Y Y.n2 1.74595
R68 VNB.t6 VNB.t1 1882.41
R69 VNB.t3 VNB.t6 1316.54
R70 VNB.t0 VNB.t3 1154.86
R71 VNB.t5 VNB.t0 1154.86
R72 VNB VNB.t4 1143.31
R73 VNB.t1 VNB.t2 1027.82
R74 VNB.t4 VNB.t5 993.177
R75 A3.n0 A3.t1 285.719
R76 A3.n1 A3.t0 277.849
R77 A3.n2 A3.n0 266.385
R78 A3.n0 A3.t2 178.34
R79 A3.n1 A3.t3 170.471
R80 A3.n2 A3.n1 152
R81 A3 A3.n2 3.2005
R82 a_114_74.n1 a_114_74.n0 343.642
R83 a_114_74.n1 a_114_74.t0 34.0546
R84 a_114_74.n0 a_114_74.t3 22.7032
R85 a_114_74.n0 a_114_74.t1 22.7032
R86 a_114_74.t2 a_114_74.n1 22.7032
R87 a_200_74.n1 a_200_74.n0 536.861
R88 a_200_74.n0 a_200_74.t3 34.0546
R89 a_200_74.n1 a_200_74.t1 25.1356
R90 a_200_74.n0 a_200_74.t0 22.7032
R91 a_200_74.t2 a_200_74.n1 22.7032
R92 A2.n0 A2.t0 231.19
R93 A2.n2 A2.t3 226.809
R94 A2.n2 A2.t2 203.141
R95 A2.n0 A2.t1 196.013
R96 A2 A2.n1 161.691
R97 A2.n4 A2.n3 152
R98 A2.n3 A2.n1 49.6611
R99 A2.n4 A2 14.8119
R100 A2.n3 A2.n2 10.955
R101 A2.n1 A2.n0 6.57323
R102 A2 A2.n4 2.74336
C0 VPB A2 0.068469f
C1 Y VGND 0.226305f
C2 VPB B1 0.058571f
C3 A3 A2 0.238387f
C4 VPB A1 0.06733f
C5 A3 B1 0.085002f
C6 VPB VPWR 0.111587f
C7 A2 B1 9.37e-19
C8 VPB Y 0.007683f
C9 A3 VPWR 0.039345f
C10 VPB VGND 0.006625f
C11 A2 VPWR 0.036357f
C12 A3 Y 0.003914f
C13 B1 A1 0.047722f
C14 B1 VPWR 0.011415f
C15 A3 VGND 0.063966f
C16 A2 Y 0.004564f
C17 B1 Y 0.121237f
C18 A1 VPWR 0.038543f
C19 A2 VGND 0.012588f
C20 A1 Y 0.15139f
C21 B1 VGND 0.01693f
C22 VPWR Y 0.015905f
C23 A1 VGND 0.012151f
C24 VPB A3 0.070674f
C25 VPWR VGND 0.069787f
C26 VGND VNB 0.54353f
C27 Y VNB 0.0781f
C28 VPWR VNB 0.4206f
C29 A1 VNB 0.242102f
C30 B1 VNB 0.170521f
C31 A2 VNB 0.208169f
C32 A3 VNB 0.290253f
C33 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a31oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31oi_4 VNB VPB VPWR VGND B1 A3 A2 A1 Y
X0 VPWR.t11 A3.t0 a_27_368.t15 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t3 A1.t0 a_27_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.4648 ps=1.95 w=1.12 l=0.15
X2 a_27_368.t10 B1.t0 Y.t5 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_475_74# A2.t0 a_30_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 Y A1 a_475_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=1.31 w=0.74 l=0.15
X5 Y.t4 B1.t1 a_27_368.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_27_368.t4 B1.t2 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X7 VPWR.t7 A2.t1 a_27_368.t11 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_27_368.t1 A2.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X9 VGND.t5 A3.t1 a_30_74.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 a_27_368.t6 A1.t1 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.4648 pd=1.95 as=0.196 ps=1.47 w=1.12 l=0.15
X11 a_475_74# A2.t3 a_30_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VGND.t1 B1.t3 Y.t7 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.40885 pd=1.845 as=0.1295 ps=1.09 w=0.74 l=0.15
X13 a_30_74.t1 A2.t4 a_475_74# VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.202325 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X14 a_27_368.t7 A1.t2 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.224 ps=1.52 w=1.12 l=0.15
X15 VPWR.t1 A2.t5 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X16 Y.t2 B1.t4 a_27_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.1848 ps=1.45 w=1.12 l=0.15
X17 a_27_368.t14 A3.t2 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_30_74.t6 A3.t3 VGND.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X19 Y.t1 A1.t3 a_475_74# VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VPWR.t6 A1.t4 a_27_368.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X21 Y.t6 B1.t5 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.40885 ps=1.845 w=0.74 l=0.15
X22 VPWR.t9 A3.t4 a_27_368.t13 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 a_27_368.t12 A3.t5 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_30_74.t5 A3.t6 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 VGND.t2 A3.t7 a_30_74.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 a_475_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X27 a_27_368.t3 A2.t6 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X28 a_475_74# A1.t5 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=1.31 as=0.19805 ps=2.07 w=0.74 l=0.15
X29 a_30_74.t0 A2.t7 a_475_74# VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1073 ps=1.03 w=0.74 l=0.15
R0 A3.n7 A3.t0 227.538
R1 A3.n1 A3.t2 226.809
R2 A3.n3 A3.t4 226.809
R3 A3.n6 A3.t5 226.809
R4 A3.n1 A3.t3 198.204
R5 A3.n10 A3.t6 196.013
R6 A3.n7 A3.t1 196.013
R7 A3.n4 A3.t7 196.013
R8 A3.n2 A3.n0 162.121
R9 A3.n5 A3.n0 152
R10 A3.n11 A3.n10 152
R11 A3.n9 A3.n8 152
R12 A3.n10 A3.n9 49.6611
R13 A3.n6 A3.n5 47.4702
R14 A3.n2 A3.n1 34.3247
R15 A3.n3 A3.n2 31.4035
R16 A3.n8 A3 13.247
R17 A3.n5 A3.n4 13.146
R18 A3.n9 A3.n7 13.146
R19 A3.n11 A3 9.07957
R20 A3 A3.n11 5.2098
R21 A3.n4 A3.n3 5.11262
R22 A3 A3.n0 4.91213
R23 A3.n10 A3.n6 2.19141
R24 A3.n8 A3 1.04236
R25 a_27_368.n13 a_27_368.n12 309.351
R26 a_27_368.n9 a_27_368.n8 292.5
R27 a_27_368.n11 a_27_368.n10 292.5
R28 a_27_368.n13 a_27_368.t10 289.711
R29 a_27_368.n15 a_27_368.n14 288.108
R30 a_27_368.n2 a_27_368.t15 281.61
R31 a_27_368.n2 a_27_368.n1 205.96
R32 a_27_368.n5 a_27_368.n4 203.014
R33 a_27_368.n3 a_27_368.n0 202.71
R34 a_27_368.n7 a_27_368.n6 194.792
R35 a_27_368.n10 a_27_368.n9 92.3443
R36 a_27_368.n3 a_27_368.n2 67.7835
R37 a_27_368.n14 a_27_368.n13 67.5062
R38 a_27_368.n14 a_27_368.n11 62.5353
R39 a_27_368.n7 a_27_368.n5 59.4308
R40 a_27_368.n8 a_27_368.n7 57.2393
R41 a_27_368.n5 a_27_368.n3 46.2829
R42 a_27_368.n6 a_27_368.t3 35.1791
R43 a_27_368.t0 a_27_368.n15 31.6612
R44 a_27_368.n9 a_27_368.t6 27.2639
R45 a_27_368.n10 a_27_368.t5 26.3844
R46 a_27_368.n4 a_27_368.t11 26.3844
R47 a_27_368.n4 a_27_368.t1 26.3844
R48 a_27_368.n0 a_27_368.t2 26.3844
R49 a_27_368.n0 a_27_368.t14 26.3844
R50 a_27_368.n1 a_27_368.t13 26.3844
R51 a_27_368.n1 a_27_368.t12 26.3844
R52 a_27_368.n6 a_27_368.t8 26.3844
R53 a_27_368.n12 a_27_368.t9 26.3844
R54 a_27_368.n12 a_27_368.t4 26.3844
R55 a_27_368.n15 a_27_368.t7 26.3844
R56 a_27_368.n11 a_27_368.n8 10.5005
R57 VPWR.n11 VPWR.n10 612.984
R58 VPWR.n9 VPWR.n8 606.915
R59 VPWR.n20 VPWR.n3 316.096
R60 VPWR.n14 VPWR.n7 316.096
R61 VPWR.n22 VPWR.n1 316.094
R62 VPWR.n5 VPWR.n4 315.812
R63 VPWR.n4 VPWR.t0 35.1791
R64 VPWR.n7 VPWR.t7 35.1791
R65 VPWR.n8 VPWR.t6 35.1791
R66 VPWR.n10 VPWR.t5 35.1791
R67 VPWR.n10 VPWR.t3 35.1791
R68 VPWR.n15 VPWR.n5 32.0005
R69 VPWR.n14 VPWR.n13 28.9887
R70 VPWR.n20 VPWR.n19 27.4829
R71 VPWR.n1 VPWR.t8 26.3844
R72 VPWR.n1 VPWR.t11 26.3844
R73 VPWR.n3 VPWR.t10 26.3844
R74 VPWR.n3 VPWR.t9 26.3844
R75 VPWR.n4 VPWR.t1 26.3844
R76 VPWR.n7 VPWR.t2 26.3844
R77 VPWR.n8 VPWR.t4 26.3844
R78 VPWR.n22 VPWR.n21 22.9652
R79 VPWR.n13 VPWR.n9 21.4593
R80 VPWR.n21 VPWR.n20 19.9534
R81 VPWR.n15 VPWR.n14 18.4476
R82 VPWR.n19 VPWR.n5 15.4358
R83 VPWR.n13 VPWR.n12 9.3005
R84 VPWR.n14 VPWR.n6 9.3005
R85 VPWR.n16 VPWR.n15 9.3005
R86 VPWR.n17 VPWR.n5 9.3005
R87 VPWR.n19 VPWR.n18 9.3005
R88 VPWR.n20 VPWR.n2 9.3005
R89 VPWR.n21 VPWR.n0 9.3005
R90 VPWR.n23 VPWR.n22 7.27223
R91 VPWR.n11 VPWR.n9 7.19852
R92 VPWR.n12 VPWR.n11 0.217359
R93 VPWR VPWR.n23 0.157962
R94 VPWR.n23 VPWR.n0 0.149814
R95 VPWR.n12 VPWR.n6 0.122949
R96 VPWR.n16 VPWR.n6 0.122949
R97 VPWR.n17 VPWR.n16 0.122949
R98 VPWR.n18 VPWR.n17 0.122949
R99 VPWR.n18 VPWR.n2 0.122949
R100 VPWR.n2 VPWR.n0 0.122949
R101 VPB.t6 VPB.t5 500.538
R102 VPB.t5 VPB.t7 280.914
R103 VPB VPB.t15 257.93
R104 VPB.t8 VPB.t6 255.376
R105 VPB.t3 VPB.t8 255.376
R106 VPB.t11 VPB.t3 255.376
R107 VPB.t2 VPB.t1 255.376
R108 VPB.t7 VPB.t0 245.161
R109 VPB.t0 VPB.t4 240.054
R110 VPB.t9 VPB.t10 229.839
R111 VPB.t4 VPB.t9 229.839
R112 VPB.t1 VPB.t11 229.839
R113 VPB.t14 VPB.t2 229.839
R114 VPB.t13 VPB.t14 229.839
R115 VPB.t12 VPB.t13 229.839
R116 VPB.t15 VPB.t12 229.839
R117 A1.n5 A1.t4 335.793
R118 A1.n6 A1.t5 234.573
R119 A1.n2 A1.t2 226.809
R120 A1.n11 A1.t0 226.809
R121 A1.n5 A1.t1 224.131
R122 A1.n2 A1.t3 206.511
R123 A1.n9 A1.n4 186.374
R124 A1.n3 A1.n1 186.374
R125 A1.n13 A1.n12 152
R126 A1.n10 A1.n0 152
R127 A1.n8 A1.n7 152
R128 A1.n6 A1.n5 50.8783
R129 A1.n8 A1.n6 46.1922
R130 A1.n3 A1.n2 43.5144
R131 A1.n9 A1.n8 36.1505
R132 A1.n11 A1.n10 27.4477
R133 A1.n12 A1.n11 18.0755
R134 A1.n12 A1.n3 12.0505
R135 A1.n13 A1.n0 10.1214
R136 A1.n10 A1.n9 9.37272
R137 A1.n7 A1 7.29352
R138 A1.n7 A1 6.99585
R139 A1 A1.n0 2.82841
R140 A1 A1.n13 1.34003
R141 B1.n3 B1.t4 237.762
R142 B1.n1 B1.t1 226.809
R143 B1.n7 B1.t2 226.809
R144 B1.n0 B1.t0 206.87
R145 B1.n0 B1.t5 198.196
R146 B1.n2 B1.t3 196.013
R147 B1.n9 B1.n8 152
R148 B1.n6 B1.n5 152
R149 B1.n4 B1.n3 152
R150 B1.n1 B1.n0 65.0033
R151 B1.n6 B1.n2 42.3581
R152 B1.n8 B1.n7 41.6278
R153 B1.n8 B1.n1 24.1005
R154 B1.n4 B1 13.247
R155 B1 B1.n9 9.37724
R156 B1.n5 B1 9.07957
R157 B1.n7 B1.n6 8.03383
R158 B1.n3 B1.n2 7.30353
R159 B1.n5 B1 5.2098
R160 B1.n9 B1 4.91213
R161 B1 B1.n4 1.04236
R162 Y.n2 Y.n0 341.913
R163 Y.n2 Y.n1 298.997
R164 Y.n4 Y.t6 251.167
R165 Y.n5 Y.t0 218.552
R166 Y Y.n2 186.03
R167 Y.n4 Y.n3 101.71
R168 Y.n5 Y.n4 100.236
R169 Y.n3 Y.t1 34.0546
R170 Y.n1 Y.t2 29.9023
R171 Y.n0 Y.t5 26.3844
R172 Y.n0 Y.t4 26.3844
R173 Y.n1 Y.t3 26.3844
R174 Y.n3 Y.t7 22.7032
R175 Y Y.n5 7.31479
R176 A2.n1 A2.t6 228.47
R177 A2.n3 A2.t1 226.809
R178 A2.n4 A2.t2 225.47
R179 A2.n6 A2.t5 207.042
R180 A2.n6 A2.t3 197.445
R181 A2.n5 A2.t7 196.013
R182 A2.n1 A2.t4 196.013
R183 A2.n10 A2.t0 196.013
R184 A2 A2.n7 152.447
R185 A2.n2 A2.n0 152
R186 A2.n12 A2.n11 152
R187 A2.n9 A2.n8 152
R188 A2.n3 A2.n2 44.549
R189 A2.n10 A2.n9 42.3254
R190 A2.n7 A2.n6 33.0996
R191 A2.n7 A2.n5 28.7766
R192 A2.n2 A2.n1 26.2914
R193 A2.n0 A2 12.9493
R194 A2.n9 A2.n4 10.7915
R195 A2.n8 A2 9.67492
R196 A2.n5 A2.n4 9.35274
R197 A2 A2.n12 8.7819
R198 A2.n11 A2.n10 7.30353
R199 A2.n12 A2 5.50748
R200 A2.n11 A2.n3 5.11262
R201 A2.n8 A2 4.61445
R202 A2 A2.n0 1.34003
R203 a_30_74.n4 a_30_74.t1 272.349
R204 a_30_74.n1 a_30_74.t7 210.411
R205 a_30_74.n5 a_30_74.n4 199.536
R206 a_30_74.n3 a_30_74.n2 104.007
R207 a_30_74.n1 a_30_74.n0 103.65
R208 a_30_74.n3 a_30_74.n1 57.6005
R209 a_30_74.n4 a_30_74.n3 49.3181
R210 a_30_74.n0 a_30_74.t4 22.7032
R211 a_30_74.n0 a_30_74.t5 22.7032
R212 a_30_74.n2 a_30_74.t2 22.7032
R213 a_30_74.n2 a_30_74.t6 22.7032
R214 a_30_74.t3 a_30_74.n5 22.7032
R215 a_30_74.n5 a_30_74.t0 22.7032
R216 VNB.t0 VNB.t1 3811.02
R217 VNB.t3 VNB.t2 2898.69
R218 VNB.t5 VNB.t0 2309.71
R219 VNB.t7 VNB.t5 1316.54
R220 VNB VNB.t11 1177.95
R221 VNB.t1 VNB.t3 1154.86
R222 VNB.t8 VNB.t10 1154.86
R223 VNB.t6 VNB.t4 1016.27
R224 VNB.t4 VNB.t7 993.177
R225 VNB.t10 VNB.t6 993.177
R226 VNB.t9 VNB.t8 993.177
R227 VNB.t11 VNB.t9 993.177
R228 VGND.n33 VGND.n2 211.183
R229 VGND.n36 VGND.n35 211.183
R230 VGND.n11 VGND.n9 185.113
R231 VGND.n15 VGND.n14 185
R232 VGND.n13 VGND.n12 185
R233 VGND.n13 VGND.n9 67.2978
R234 VGND.n14 VGND.n13 66.487
R235 VGND.n17 VGND.n16 36.1417
R236 VGND.n17 VGND.n6 36.1417
R237 VGND.n21 VGND.n6 36.1417
R238 VGND.n22 VGND.n21 36.1417
R239 VGND.n23 VGND.n22 36.1417
R240 VGND.n23 VGND.n4 36.1417
R241 VGND.n27 VGND.n4 36.1417
R242 VGND.n28 VGND.n27 36.1417
R243 VGND.n29 VGND.n28 36.1417
R244 VGND.n29 VGND.n1 36.1417
R245 VGND.n2 VGND.t4 34.0546
R246 VGND.n33 VGND.n1 30.8711
R247 VGND.n36 VGND.n34 23.3417
R248 VGND.n9 VGND.t0 22.7032
R249 VGND.n14 VGND.t1 22.7032
R250 VGND.n2 VGND.t2 22.7032
R251 VGND.n35 VGND.t3 22.7032
R252 VGND.n35 VGND.t5 22.7032
R253 VGND.n34 VGND.n33 16.5652
R254 VGND.n10 VGND.n8 9.3005
R255 VGND.n16 VGND.n7 9.3005
R256 VGND.n18 VGND.n17 9.3005
R257 VGND.n19 VGND.n6 9.3005
R258 VGND.n21 VGND.n20 9.3005
R259 VGND.n22 VGND.n5 9.3005
R260 VGND.n24 VGND.n23 9.3005
R261 VGND.n25 VGND.n4 9.3005
R262 VGND.n27 VGND.n26 9.3005
R263 VGND.n28 VGND.n3 9.3005
R264 VGND.n30 VGND.n29 9.3005
R265 VGND.n31 VGND.n1 9.3005
R266 VGND.n33 VGND.n32 9.3005
R267 VGND.n34 VGND.n0 9.3005
R268 VGND.n11 VGND.n10 7.61028
R269 VGND.n37 VGND.n36 7.25439
R270 VGND.n12 VGND.n11 5.63191
R271 VGND.n16 VGND.n15 5.0798
R272 VGND.n15 VGND.n8 4.63618
R273 VGND.n12 VGND.n8 1.03834
R274 VGND VGND.n37 0.157727
R275 VGND.n37 VGND.n0 0.150046
R276 VGND.n10 VGND.n7 0.122949
R277 VGND.n18 VGND.n7 0.122949
R278 VGND.n19 VGND.n18 0.122949
R279 VGND.n20 VGND.n19 0.122949
R280 VGND.n20 VGND.n5 0.122949
R281 VGND.n24 VGND.n5 0.122949
R282 VGND.n25 VGND.n24 0.122949
R283 VGND.n26 VGND.n25 0.122949
R284 VGND.n26 VGND.n3 0.122949
R285 VGND.n30 VGND.n3 0.122949
R286 VGND.n31 VGND.n30 0.122949
R287 VGND.n32 VGND.n31 0.122949
R288 VGND.n32 VGND.n0 0.122949
C0 VPWR VGND 0.138271f
C1 a_475_74# B1 4.29e-19
C2 VPB A2 0.142989f
C3 Y VGND 0.296758f
C4 A3 A2 0.074713f
C5 a_475_74# VPWR 0.005124f
C6 VPB A1 0.183751f
C7 VPB B1 0.141962f
C8 a_475_74# Y 0.233998f
C9 VPB VPWR 0.210059f
C10 A2 A1 0.034666f
C11 a_475_74# VGND 0.452569f
C12 A3 VPWR 0.085014f
C13 VPB Y 0.007392f
C14 A1 B1 0.092122f
C15 A2 VPWR 0.081826f
C16 A3 Y 2.16e-19
C17 VPB VGND 0.008523f
C18 A3 VGND 0.072437f
C19 A1 VPWR 0.063408f
C20 A2 Y 0.031438f
C21 a_475_74# VPB 1.41e-20
C22 A1 Y 0.359318f
C23 A2 VGND 0.030283f
C24 B1 VPWR 0.025062f
C25 a_475_74# A3 3.86e-19
C26 A1 VGND 0.029451f
C27 B1 Y 0.420112f
C28 a_475_74# A2 0.051162f
C29 B1 VGND 0.045225f
C30 VPWR Y 0.046123f
C31 VPB A3 0.138459f
C32 a_475_74# A1 0.050197f
C33 VGND VNB 0.969379f
C34 Y VNB 0.077925f
C35 VPWR VNB 0.768727f
C36 B1 VNB 0.391669f
C37 A1 VNB 0.470896f
C38 A2 VNB 0.422829f
C39 A3 VNB 0.444444f
C40 VPB VNB 2.01326f
C41 a_475_74# VNB 0.034777f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a32o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32o_1 VNB VPB VPWR VGND X B2 B1 A2 A1 A3
X0 a_601_94.t1 B1.t0 a_84_48.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2016 ps=1.27 w=0.64 l=0.15
X1 a_337_94.t1 A2.t0 a_259_94.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
X2 a_84_48.t0 A1.t0 a_337_94.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2016 pd=1.27 as=0.1248 ps=1.03 w=0.64 l=0.15
X3 VGND.t2 a_84_48.t4 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.209 pd=1.315 as=0.2109 ps=2.05 w=0.74 l=0.15
X4 VPWR.t0 a_84_48.t5 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2607 pd=1.6 as=0.3304 ps=2.83 w=1.12 l=0.15
X5 VPWR.t2 A2.t1 a_244_368.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=1.59 as=0.15 ps=1.3 w=1 l=0.15
X6 a_84_48.t1 B1.t1 a_244_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X7 a_244_368.t0 A3.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2607 ps=1.6 w=1 l=0.15
X8 a_244_368.t3 A1.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=1.59 w=1 l=0.15
X9 a_259_94.t0 A3.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.209 ps=1.315 w=0.64 l=0.15
X10 a_244_368.t4 B2.t0 a_84_48.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2 ps=1.4 w=1 l=0.15
X11 VGND.t0 B2.t1 a_601_94.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0768 ps=0.88 w=0.64 l=0.15
R0 B1.n0 B1.t1 266.44
R1 B1.n0 B1.t0 162.274
R2 B1 B1.n0 162.133
R3 a_84_48.n3 a_84_48.n2 385.579
R4 a_84_48.n1 a_84_48.t5 263.938
R5 a_84_48.n1 a_84_48.t4 203.688
R6 a_84_48.n2 a_84_48.n0 178.416
R7 a_84_48.n2 a_84_48.n1 152
R8 a_84_48.n0 a_84_48.t2 51.6892
R9 a_84_48.n0 a_84_48.t0 49.7595
R10 a_84_48.n3 a_84_48.t3 39.4005
R11 a_84_48.t1 a_84_48.n3 39.4005
R12 a_601_94.t0 a_601_94.t1 45.0005
R13 VNB.t2 VNB.t5 1801.57
R14 VNB.t3 VNB.t1 1674.54
R15 VNB.t4 VNB.t2 1247.24
R16 VNB VNB.t3 1143.31
R17 VNB.t5 VNB.t0 900.788
R18 VNB.t1 VNB.t4 900.788
R19 A2.n0 A2.t1 266.44
R20 A2.n0 A2.t0 162.274
R21 A2 A2.n0 158.788
R22 a_259_94.t0 a_259_94.t1 45.0005
R23 a_337_94.t0 a_337_94.t1 73.1255
R24 A1.n0 A1.t1 263.269
R25 A1.n0 A1.t0 159.102
R26 A1 A1.n0 158.788
R27 X.n0 X.t0 292.712
R28 X.t1 X.n0 279.738
R29 X.n1 X.t1 279.738
R30 X.n1 X 11.5561
R31 X.n0 X 4.44494
R32 X X.n1 1.6005
R33 VGND.n1 VGND.n0 207.796
R34 VGND.n1 VGND.t0 162.93
R35 VGND.n0 VGND.t1 55.313
R36 VGND.n0 VGND.t2 32.825
R37 VGND VGND.n1 0.211269
R38 VPWR.n2 VPWR.n0 621
R39 VPWR.n2 VPWR.n1 316.601
R40 VPWR.n0 VPWR.t3 58.1155
R41 VPWR.n0 VPWR.t2 58.1155
R42 VPWR.n1 VPWR.t1 49.2881
R43 VPWR.n1 VPWR.t0 41.2186
R44 VPWR VPWR.n2 0.355379
R45 VPB.t3 VPB.t4 377.957
R46 VPB.t0 VPB.t1 321.774
R47 VPB.t2 VPB.t5 280.914
R48 VPB VPB.t0 263.038
R49 VPB.t4 VPB.t2 229.839
R50 VPB.t1 VPB.t3 229.839
R51 a_244_368.n2 a_244_368.n1 374.7
R52 a_244_368.n1 a_244_368.t4 315.19
R53 a_244_368.n1 a_244_368.n0 287.591
R54 a_244_368.n0 a_244_368.t1 29.5505
R55 a_244_368.n0 a_244_368.t3 29.5505
R56 a_244_368.n2 a_244_368.t2 29.5505
R57 a_244_368.t0 a_244_368.n2 29.5505
R58 A3.n0 A3.t0 266.44
R59 A3.n0 A3.t1 162.274
R60 A3 A3.n0 158.4
R61 B2.n0 B2.t0 263.548
R62 B2.n0 B2.t1 159.381
R63 B2 B2.n0 157.272
C0 VPB A3 0.033564f
C1 X VPWR 0.12111f
C2 B1 VGND 0.015909f
C3 VPB A2 0.032916f
C4 X A3 0.001814f
C5 B2 VGND 0.051211f
C6 VPB A1 0.034919f
C7 VPWR A3 0.016018f
C8 X A2 5.57e-19
C9 VPWR A2 0.012357f
C10 X A1 2.36e-19
C11 VPB B1 0.030911f
C12 VPWR A1 0.013531f
C13 VPB B2 0.037221f
C14 X B1 7.83e-20
C15 A3 A2 0.092848f
C16 VPWR B1 0.005627f
C17 VPB VGND 0.006249f
C18 VPWR B2 0.005974f
C19 A2 A1 0.073038f
C20 X VGND 0.067926f
C21 VPWR VGND 0.063521f
C22 A1 B1 0.082829f
C23 A3 VGND 0.011437f
C24 VPB X 0.014306f
C25 A2 VGND 0.008636f
C26 VPB VPWR 0.104254f
C27 B1 B2 0.076799f
C28 A1 VGND 0.006793f
C29 VGND VNB 0.534482f
C30 B2 VNB 0.155282f
C31 B1 VNB 0.109451f
C32 A1 VNB 0.113463f
C33 A2 VNB 0.103819f
C34 A3 VNB 0.109254f
C35 VPWR VNB 0.384026f
C36 X VNB 0.112145f
C37 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a41oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a41oi_4 VNB VPB VPWR VGND Y A1 A2 A3 A4 B1
X0 VPWR.t3 A1.t0 a_27_368# VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_27_368# A4.t0 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_27_368# B1.t0 Y.t9 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5 Y.t8 B1.t1 a_27_368# VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6 a_325_74.t7 A1.t1 Y.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2294 pd=1.36 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 a_852_74.t7 A3.t0 a_1235_74.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 Y.t7 B1.t2 a_27_368# VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.336 ps=2.84 w=1.12 l=0.15
X9 VPWR.t8 A2.t0 a_27_368# VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_325_74.t6 A1.t2 Y.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_27_368# A1.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1988 ps=1.475 w=1.12 l=0.15
X12 a_1235_74.t3 A3.t1 a_852_74.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_27_368# A2.t1 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2016 ps=1.48 w=1.12 l=0.15
X14 Y.t5 B1.t3 VGND.t5 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 VPWR.t10 A2.t2 a_27_368# VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X16 Y.t1 A1.t4 a_325_74.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X17 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X18 a_27_368# B1.t4 Y.t6 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1932 ps=1.465 w=1.12 l=0.15
X19 VPWR.t1 A1.t5 a_27_368# VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.475 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_27_368# A1.t6 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
X21 Y.t0 A1.t7 a_325_74.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2294 ps=1.36 w=0.74 l=0.15
X22 a_325_74.t3 A2.t3 a_852_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_1235_74.t7 A4.t1 VGND.t3 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X25 a_27_368# A4.t2 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X26 a_27_368# A3.t2 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X27 a_1235_74.t1 A3.t3 a_852_74.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 a_1235_74.t6 A4.t3 VGND.t2 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X29 a_325_74.t2 A2.t4 a_852_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X30 VGND.t1 A4.t4 a_1235_74.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X31 VGND.t4 B1.t5 Y.t4 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X32 a_852_74.t1 A2.t5 a_325_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X33 VGND.t0 A4.t5 a_1235_74.t4 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X34 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X35 VPWR.t5 A3.t4 a_27_368# VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X36 a_852_74.t0 A2.t6 a_325_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1295 ps=1.09 w=0.74 l=0.15
X37 a_852_74.t4 A3.t5 a_1235_74.t0 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A1.n5 A1.t4 256.531
R1 A1.n0 A1.t3 255.46
R2 A1.n1 A1.t5 209.403
R3 A1.n4 A1.t6 209.403
R4 A1.n5 A1.t0 209.403
R5 A1.n6 A1 155.126
R6 A1 A1.n3 154.828
R7 A1.n9 A1.n8 152
R8 A1.n7 A1.t1 149.421
R9 A1.n2 A1.t7 149.421
R10 A1.n0 A1.t2 149.421
R11 A1.n8 A1.n7 27.2246
R12 A1.n1 A1.n0 24.9931
R13 A1.n4 A1.n3 15.6209
R14 A1.n8 A1.n4 14.7283
R15 A1.n2 A1.n1 13.3894
R16 A1.n3 A1.n2 11.1579
R17 A1 A1.n9 7.29352
R18 A1.n9 A1 6.99585
R19 A1.n6 A1.n5 4.01717
R20 A1.n7 A1.n6 3.12457
R21 VPWR.n26 VPWR.n3 612.393
R22 VPWR.n28 VPWR.n1 608.08
R23 VPWR.n11 VPWR.t7 365.046
R24 VPWR.n20 VPWR.t10 349.789
R25 VPWR.n10 VPWR.t6 349.789
R26 VPWR.n5 VPWR.n4 323.793
R27 VPWR.n8 VPWR.n7 323.406
R28 VPWR.n4 VPWR.t9 36.938
R29 VPWR.n3 VPWR.t2 36.0585
R30 VPWR.n1 VPWR.t0 35.1791
R31 VPWR.n1 VPWR.t3 35.1791
R32 VPWR.n7 VPWR.t4 35.1791
R33 VPWR.n27 VPWR.n26 32.0005
R34 VPWR.n25 VPWR.n5 31.624
R35 VPWR.n21 VPWR.n20 31.624
R36 VPWR.n19 VPWR.n8 30.8711
R37 VPWR.n15 VPWR.n14 30.1181
R38 VPWR.n13 VPWR.n10 27.1064
R39 VPWR.n3 VPWR.t1 26.3844
R40 VPWR.n4 VPWR.t8 26.3844
R41 VPWR.n7 VPWR.t5 26.3844
R42 VPWR.n14 VPWR.n13 23.3417
R43 VPWR.n15 VPWR.n8 22.5887
R44 VPWR.n21 VPWR.n5 21.8358
R45 VPWR.n20 VPWR.n19 21.8358
R46 VPWR.n26 VPWR.n25 21.4593
R47 VPWR.n28 VPWR.n27 20.7064
R48 VPWR.n13 VPWR.n12 9.3005
R49 VPWR.n14 VPWR.n9 9.3005
R50 VPWR.n16 VPWR.n15 9.3005
R51 VPWR.n17 VPWR.n8 9.3005
R52 VPWR.n19 VPWR.n18 9.3005
R53 VPWR.n20 VPWR.n6 9.3005
R54 VPWR.n22 VPWR.n21 9.3005
R55 VPWR.n23 VPWR.n5 9.3005
R56 VPWR.n25 VPWR.n24 9.3005
R57 VPWR.n26 VPWR.n2 9.3005
R58 VPWR.n27 VPWR.n0 9.3005
R59 VPWR.n29 VPWR.n28 7.29602
R60 VPWR.n11 VPWR.n10 6.94902
R61 VPWR VPWR.n29 0.644871
R62 VPWR.n12 VPWR.n11 0.485017
R63 VPWR.n29 VPWR.n0 0.155053
R64 VPWR.n12 VPWR.n9 0.122949
R65 VPWR.n16 VPWR.n9 0.122949
R66 VPWR.n17 VPWR.n16 0.122949
R67 VPWR.n18 VPWR.n17 0.122949
R68 VPWR.n18 VPWR.n6 0.122949
R69 VPWR.n22 VPWR.n6 0.122949
R70 VPWR.n23 VPWR.n22 0.122949
R71 VPWR.n24 VPWR.n23 0.122949
R72 VPWR.n24 VPWR.n2 0.122949
R73 VPWR.n2 VPWR.n0 0.122949
R74 VPB.t7 VPB.t9 970.431
R75 VPB.t14 VPB.t8 485.216
R76 VPB.t9 VPB.t10 459.678
R77 VPB.t3 VPB.t0 280.914
R78 VPB.t11 VPB.t12 260.485
R79 VPB VPB.t5 260.485
R80 VPB.t1 VPB.t2 257.93
R81 VPB.t8 VPB.t7 255.376
R82 VPB.t4 VPB.t13 255.376
R83 VPB.t5 VPB.t4 252.823
R84 VPB.t12 VPB.t14 229.839
R85 VPB.t2 VPB.t11 229.839
R86 VPB.t0 VPB.t1 229.839
R87 VPB.t6 VPB.t3 229.839
R88 VPB.t13 VPB.t6 229.839
R89 A4.n6 A4.n5 231.921
R90 A4.n0 A4.t2 226.809
R91 A4.n2 A4.n1 226.809
R92 A4.n8 A4.t0 226.809
R93 A4.n0 A4.t3 198.204
R94 A4.n6 A4.t5 196.013
R95 A4.n9 A4.t1 196.013
R96 A4.n4 A4.t4 196.013
R97 A4.n15 A4.n14 152
R98 A4.n13 A4.n12 152
R99 A4.n11 A4.n10 152
R100 A4.n7 A4.n3 152
R101 A4.n14 A4.n13 49.6611
R102 A4.n10 A4.n4 47.4702
R103 A4.n8 A4.n7 32.1338
R104 A4.n7 A4.n6 28.4823
R105 A4.n10 A4.n9 15.3369
R106 A4.n14 A4.n0 14.6066
R107 A4.n11 A4.n3 10.1214
R108 A4.n12 A4 9.97259
R109 A4 A4.n15 8.48422
R110 A4.n15 A4 5.80515
R111 A4.n12 A4 4.31678
R112 A4.n3 A4 4.0191
R113 A4.n9 A4.n8 2.19141
R114 A4.n13 A4.n2 1.46111
R115 A4.n4 A4.n2 0.730803
R116 A4 A4.n11 0.149337
R117 B1.n0 B1.t0 336.164
R118 B1.n0 B1.t1 217.436
R119 B1.n2 B1.t4 217.436
R120 B1.n4 B1.t2 217.436
R121 B1.n4 B1.t3 197.994
R122 B1.n3 B1.t5 196.013
R123 B1 B1.n1 156.465
R124 B1.n8 B1.n7 152
R125 B1.n6 B1.n5 152
R126 B1.n7 B1.n6 44.8991
R127 B1.n2 B1.n1 34.3347
R128 B1.n1 B1.n0 31.6936
R129 B1.n5 B1 12.8005
R130 B1.n6 B1.n4 9.90461
R131 B1.n7 B1.n3 9.24434
R132 B1.n8 B1 8.63306
R133 B1 B1.n8 5.65631
R134 B1.n5 B1 1.48887
R135 B1.n3 B1.n2 1.32105
R136 Y.n5 Y.n4 355.483
R137 Y.n5 Y.n3 300.733
R138 Y Y.n7 236.287
R139 Y.n2 Y.n1 197.994
R140 Y.n2 Y.n0 172.488
R141 Y Y.n6 131.883
R142 Y.n4 Y.t7 34.2996
R143 Y.n1 Y.t1 34.0546
R144 Y.n0 Y.t4 34.0546
R145 Y.n6 Y.n2 32.0005
R146 Y.n3 Y.t9 26.3844
R147 Y.n3 Y.t8 26.3844
R148 Y.n4 Y.t6 26.3844
R149 Y.n1 Y.t3 22.7032
R150 Y.n0 Y.t5 22.7032
R151 Y.n7 Y.t2 22.7032
R152 Y.n7 Y.t0 22.7032
R153 Y.n6 Y.n5 9.81383
R154 A2.n2 A2.n1 298.396
R155 A2.n4 A2.t2 234.841
R156 A2.n0 A2.t1 234.841
R157 A2.n10 A2.t0 234.841
R158 A2.n10 A2.t6 186.482
R159 A2.n6 A2.n3 165.189
R160 A2.n6 A2.n5 152
R161 A2.n8 A2.n7 152
R162 A2.n12 A2.n11 152
R163 A2.n5 A2.t5 149.421
R164 A2.n9 A2.t4 149.421
R165 A2.n2 A2.t3 149.421
R166 A2.n11 A2.n9 27.0792
R167 A2.n5 A2.n0 26.5376
R168 A2.n5 A2.n4 22.205
R169 A2.n4 A2.n3 14.623
R170 A2.n7 A2.n6 13.1884
R171 A2 A2.n12 12.244
R172 A2.n8 A2.n0 10.2904
R173 A2.n3 A2.n2 9.74881
R174 A2.n9 A2.n8 9.74881
R175 A2.n7 A2 9.44451
R176 A2.n11 A2.n10 8.1241
R177 A2.n12 A2 1.11354
R178 a_325_74.n1 a_325_74.t3 309.897
R179 a_325_74.n7 a_325_74.t5 270.368
R180 a_325_74.n4 a_325_74.n2 185
R181 a_325_74.n3 a_325_74.n2 185
R182 a_325_74.n1 a_325_74.n0 185
R183 a_325_74.n9 a_325_74.n8 95.7292
R184 a_325_74.n6 a_325_74.n5 80.5048
R185 a_325_74.n8 a_325_74.n7 56.2339
R186 a_325_74.t6 a_325_74.n9 34.0546
R187 a_325_74.n8 a_325_74.n1 32.6142
R188 a_325_74.n5 a_325_74.n4 23.9934
R189 a_325_74.n5 a_325_74.n3 23.9934
R190 a_325_74.n0 a_325_74.t1 22.7032
R191 a_325_74.n0 a_325_74.t2 22.7032
R192 a_325_74.n3 a_325_74.t4 22.7032
R193 a_325_74.n4 a_325_74.t7 22.7032
R194 a_325_74.n9 a_325_74.t0 22.7032
R195 a_325_74.n6 a_325_74.n2 10.8684
R196 a_325_74.n7 a_325_74.n6 4.22692
R197 VNB.t3 VNB.t8 2286.61
R198 VNB.t16 VNB.t5 2286.61
R199 VNB.t7 VNB.t4 1778.48
R200 VNB.t0 VNB.t2 1154.86
R201 VNB.t6 VNB.t0 1154.86
R202 VNB.t5 VNB.t7 1154.86
R203 VNB.t17 VNB.t16 1154.86
R204 VNB VNB.t17 1143.31
R205 VNB.t13 VNB.t14 1085.56
R206 VNB.t15 VNB.t13 993.177
R207 VNB.t12 VNB.t15 993.177
R208 VNB.t10 VNB.t12 993.177
R209 VNB.t11 VNB.t10 993.177
R210 VNB.t9 VNB.t11 993.177
R211 VNB.t8 VNB.t9 993.177
R212 VNB.t1 VNB.t3 993.177
R213 VNB.t2 VNB.t1 993.177
R214 VNB.t4 VNB.t6 993.177
R215 A3.n7 A3.t4 237.762
R216 A3.n2 A3.n1 226.809
R217 A3.n13 A3.n3 226.809
R218 A3.n5 A3.t2 226.809
R219 A3.n2 A3.t3 211.351
R220 A3.n8 A3.t0 196.013
R221 A3.n4 A3.t1 196.013
R222 A3.n15 A3.t5 196.013
R223 A3.n17 A3.n16 152
R224 A3.n14 A3.n0 152
R225 A3.n12 A3.n11 152
R226 A3.n10 A3.n9 152
R227 A3.n7 A3.n6 152
R228 A3.n16 A3.n15 45.2793
R229 A3.n13 A3.n12 28.4823
R230 A3.n5 A3.n4 28.4823
R231 A3.n8 A3.n7 27.752
R232 A3.n9 A3.n8 21.9096
R233 A3.n14 A3.n13 21.1793
R234 A3.n6 A3 12.8005
R235 A3.n9 A3.n5 12.4157
R236 A3.n17 A3.n0 10.1214
R237 A3.n11 A3 9.82376
R238 A3.n12 A3.n4 8.76414
R239 A3.n10 A3 8.63306
R240 A3 A3.n10 5.65631
R241 A3.n11 A3 4.46562
R242 A3.n15 A3.n14 4.38232
R243 A3 A3.n17 3.87027
R244 A3.n16 A3.n2 2.19141
R245 A3.n6 A3 1.48887
R246 A3 A3.n0 0.298174
R247 a_1235_74.n4 a_1235_74.t2 318.933
R248 a_1235_74.n1 a_1235_74.t6 213.423
R249 a_1235_74.n5 a_1235_74.n4 185
R250 a_1235_74.n1 a_1235_74.n0 103.65
R251 a_1235_74.n3 a_1235_74.n2 86.1054
R252 a_1235_74.n3 a_1235_74.n1 80.9333
R253 a_1235_74.n4 a_1235_74.n3 56.8241
R254 a_1235_74.n2 a_1235_74.t4 22.7032
R255 a_1235_74.n2 a_1235_74.t1 22.7032
R256 a_1235_74.n0 a_1235_74.t5 22.7032
R257 a_1235_74.n0 a_1235_74.t7 22.7032
R258 a_1235_74.t0 a_1235_74.n5 22.7032
R259 a_1235_74.n5 a_1235_74.t3 22.7032
R260 a_852_74.n2 a_852_74.n0 217.376
R261 a_852_74.n4 a_852_74.n3 217.376
R262 a_852_74.n2 a_852_74.n1 185
R263 a_852_74.n5 a_852_74.n4 185
R264 a_852_74.n4 a_852_74.n2 53.4593
R265 a_852_74.n3 a_852_74.t0 34.0546
R266 a_852_74.n3 a_852_74.t2 22.7032
R267 a_852_74.n1 a_852_74.t6 22.7032
R268 a_852_74.n1 a_852_74.t7 22.7032
R269 a_852_74.n0 a_852_74.t5 22.7032
R270 a_852_74.n0 a_852_74.t4 22.7032
R271 a_852_74.t3 a_852_74.n5 22.7032
R272 a_852_74.n5 a_852_74.t1 22.7032
R273 VGND.n34 VGND.t4 233.886
R274 VGND.n9 VGND.n8 216.702
R275 VGND.n11 VGND.n10 211.183
R276 VGND.n36 VGND.t5 171.77
R277 VGND.n12 VGND.n7 36.1417
R278 VGND.n16 VGND.n7 36.1417
R279 VGND.n17 VGND.n16 36.1417
R280 VGND.n18 VGND.n17 36.1417
R281 VGND.n18 VGND.n5 36.1417
R282 VGND.n22 VGND.n5 36.1417
R283 VGND.n23 VGND.n22 36.1417
R284 VGND.n24 VGND.n23 36.1417
R285 VGND.n24 VGND.n3 36.1417
R286 VGND.n28 VGND.n3 36.1417
R287 VGND.n29 VGND.n28 36.1417
R288 VGND.n30 VGND.n29 36.1417
R289 VGND.n30 VGND.n1 36.1417
R290 VGND.n8 VGND.t2 29.1897
R291 VGND.n12 VGND.n11 28.9887
R292 VGND.n36 VGND.n35 26.7299
R293 VGND.n35 VGND.n34 24.4711
R294 VGND.n34 VGND.n1 22.9652
R295 VGND.n8 VGND.t1 22.7032
R296 VGND.n10 VGND.t3 22.7032
R297 VGND.n10 VGND.t0 22.7032
R298 VGND.n37 VGND.n36 9.3005
R299 VGND.n13 VGND.n12 9.3005
R300 VGND.n14 VGND.n7 9.3005
R301 VGND.n16 VGND.n15 9.3005
R302 VGND.n17 VGND.n6 9.3005
R303 VGND.n19 VGND.n18 9.3005
R304 VGND.n20 VGND.n5 9.3005
R305 VGND.n22 VGND.n21 9.3005
R306 VGND.n23 VGND.n4 9.3005
R307 VGND.n25 VGND.n24 9.3005
R308 VGND.n26 VGND.n3 9.3005
R309 VGND.n28 VGND.n27 9.3005
R310 VGND.n29 VGND.n2 9.3005
R311 VGND.n31 VGND.n30 9.3005
R312 VGND.n32 VGND.n1 9.3005
R313 VGND.n34 VGND.n33 9.3005
R314 VGND.n35 VGND.n0 9.3005
R315 VGND.n11 VGND.n9 6.30563
R316 VGND.n13 VGND.n9 0.64124
R317 VGND.n14 VGND.n13 0.122949
R318 VGND.n15 VGND.n14 0.122949
R319 VGND.n15 VGND.n6 0.122949
R320 VGND.n19 VGND.n6 0.122949
R321 VGND.n20 VGND.n19 0.122949
R322 VGND.n21 VGND.n20 0.122949
R323 VGND.n21 VGND.n4 0.122949
R324 VGND.n25 VGND.n4 0.122949
R325 VGND.n26 VGND.n25 0.122949
R326 VGND.n27 VGND.n26 0.122949
R327 VGND.n27 VGND.n2 0.122949
R328 VGND.n31 VGND.n2 0.122949
R329 VGND.n32 VGND.n31 0.122949
R330 VGND.n33 VGND.n32 0.122949
R331 VGND.n33 VGND.n0 0.122949
R332 VGND.n37 VGND.n0 0.122949
R333 VGND VGND.n37 0.0617245
C0 a_27_368# A1 0.070829f
C1 A2 A3 0.067753f
C2 VPB VPWR 0.24705f
C3 B1 Y 0.275649f
C4 a_27_368# A2 0.210769f
C5 A2 A4 3.03e-20
C6 VPB VGND 0.009815f
C7 A1 Y 0.288291f
C8 B1 VPWR 0.023412f
C9 a_27_368# A3 0.259385f
C10 A2 Y 0.031289f
C11 B1 VGND 0.062917f
C12 A1 VPWR 0.060361f
C13 A3 A4 0.091367f
C14 a_27_368# A4 0.219398f
C15 A1 VGND 0.028784f
C16 A2 VPWR 0.07221f
C17 A3 Y 2.05e-19
C18 a_27_368# Y 0.451269f
C19 A2 VGND 0.024265f
C20 A3 VPWR 0.073668f
C21 A4 Y 6.97e-20
C22 a_27_368# VPWR 1.66753f
C23 VPB B1 0.142853f
C24 A3 VGND 0.02732f
C25 A4 VPWR 0.069748f
C26 a_27_368# VGND 0.02033f
C27 VPB A1 0.147876f
C28 A4 VGND 0.074068f
C29 Y VPWR 0.043413f
C30 VPB A2 0.146626f
C31 B1 A1 0.046606f
C32 Y VGND 0.208152f
C33 VPB A3 0.149261f
C34 VPWR VGND 0.161116f
C35 a_27_368# VPB 0.056953f
C36 VPB A4 0.138914f
C37 A1 A2 0.053874f
C38 a_27_368# B1 0.100734f
C39 VPB Y 0.010239f
C40 VGND VNB 1.16511f
C41 VPWR VNB 0.893245f
C42 Y VNB 0.047925f
C43 A4 VNB 0.441505f
C44 A3 VNB 0.42311f
C45 A2 VNB 0.42466f
C46 A1 VNB 0.452175f
C47 B1 VNB 0.374535f
C48 VPB VNB 2.33467f
C49 a_27_368# VNB 0.085002f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a41oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a41oi_2 VNB VPB VPWR VGND A1 Y A2 A3 A4 B1
X0 Y.t1 B1.t0 a_27_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y.t2 B1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2 VPWR.t1 A1.t0 a_27_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=1.71 as=0.196 ps=1.47 w=1.12 l=0.15
X3 a_512_74.t1 A2.t0 a_239_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4 VPWR.t5 A4.t0 a_27_368.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2156 ps=1.505 w=1.12 l=0.15
X5 a_27_368.t3 A4.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3584 pd=2.88 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_27_368.t8 A3.t0 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.2156 pd=1.505 as=0.224 ps=1.52 w=1.12 l=0.15
X7 a_239_74.t0 A2.t1 a_512_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_239_74.t3 A1.t1 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VPWR.t4 A2.t2 a_27_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_27_368.t0 B1.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X11 a_27_368.t4 A1.t2 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=1.71 w=1.12 l=0.15
X12 a_709_74.t1 A4.t2 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2257 pd=2.09 as=0.1221 ps=1.07 w=0.74 l=0.15
X13 a_709_74.t3 A3.t1 a_512_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 Y.t3 A1.t3 a_239_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X15 VGND.t2 A4.t3 a_709_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VPWR.t7 A3.t2 a_27_368.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_512_74.t2 A3.t3 a_709_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X18 a_27_368.t2 A2.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.224 ps=1.52 w=1.12 l=0.15
R0 B1.n0 B1.t2 239.224
R1 B1.n1 B1.t0 235.571
R2 B1.n1 B1.t1 179.947
R3 B1 B1.n0 160.484
R4 B1.n3 B1.n2 152
R5 B1.n2 B1.n0 49.6611
R6 B1.n3 B1 12.6517
R7 B1.n2 B1.n1 2.19141
R8 B1 B1.n3 1.63771
R9 a_27_368.n6 a_27_368.t1 301.221
R10 a_27_368.n7 a_27_368.n6 288.625
R11 a_27_368.n2 a_27_368.t3 282.741
R12 a_27_368.n4 a_27_368.n3 205.487
R13 a_27_368.n2 a_27_368.n1 202.68
R14 a_27_368.n5 a_27_368.n0 194.504
R15 a_27_368.n6 a_27_368.n5 78.2327
R16 a_27_368.n5 a_27_368.n4 59.0719
R17 a_27_368.n4 a_27_368.n2 50.4476
R18 a_27_368.n1 a_27_368.t7 38.6969
R19 a_27_368.t0 a_27_368.n7 35.1791
R20 a_27_368.n1 a_27_368.t8 29.0228
R21 a_27_368.n0 a_27_368.t6 26.3844
R22 a_27_368.n0 a_27_368.t4 26.3844
R23 a_27_368.n3 a_27_368.t9 26.3844
R24 a_27_368.n3 a_27_368.t2 26.3844
R25 a_27_368.n7 a_27_368.t5 26.3844
R26 Y Y.n0 424.284
R27 Y.n2 Y.t2 202.923
R28 Y.n2 Y.n1 202.153
R29 Y.n0 Y.t1 35.1791
R30 Y.n0 Y.t0 26.3844
R31 Y.n1 Y.t4 22.7032
R32 Y.n1 Y.t3 22.7032
R33 Y Y.n2 7.80048
R34 VPB.t5 VPB.t4 377.957
R35 VPB.t9 VPB.t8 280.914
R36 VPB.t6 VPB.t2 280.914
R37 VPB.t8 VPB.t7 273.253
R38 VPB VPB.t1 257.93
R39 VPB.t0 VPB.t5 255.376
R40 VPB.t1 VPB.t0 255.376
R41 VPB.t7 VPB.t3 229.839
R42 VPB.t2 VPB.t9 229.839
R43 VPB.t4 VPB.t6 229.839
R44 VGND.n1 VGND.n0 218.155
R45 VGND.n1 VGND.t0 163.643
R46 VGND.n0 VGND.t1 30.8113
R47 VGND.n0 VGND.t2 22.7032
R48 VGND VGND.n1 0.0988719
R49 VNB.t0 VNB.t6 2286.61
R50 VNB.t1 VNB.t4 2286.61
R51 VNB VNB.t1 1304.99
R52 VNB.t5 VNB.t2 1154.86
R53 VNB.t8 VNB.t3 1108.66
R54 VNB.t7 VNB.t8 993.177
R55 VNB.t6 VNB.t7 993.177
R56 VNB.t2 VNB.t0 993.177
R57 VNB.t4 VNB.t5 993.177
R58 A1.n0 A1.t2 275.009
R59 A1.n1 A1.t0 221.185
R60 A1.n1 A1.t3 196.013
R61 A1.n0 A1.t1 196.013
R62 A1 A1.n2 154.19
R63 A1.n2 A1.n0 52.0565
R64 A1.n2 A1.n1 3.21383
R65 VPWR.n14 VPWR.n1 598.538
R66 VPWR.n5 VPWR.n4 321.45
R67 VPWR.n3 VPWR.n2 316.353
R68 VPWR.n7 VPWR.n6 316.353
R69 VPWR.n1 VPWR.t0 51.8889
R70 VPWR.n1 VPWR.t1 51.8889
R71 VPWR.n13 VPWR.n12 36.1417
R72 VPWR.n2 VPWR.t2 35.1791
R73 VPWR.n2 VPWR.t4 35.1791
R74 VPWR.n6 VPWR.t6 35.1791
R75 VPWR.n6 VPWR.t7 35.1791
R76 VPWR.n8 VPWR.n3 35.0123
R77 VPWR.n4 VPWR.t3 26.3844
R78 VPWR.n4 VPWR.t5 26.3844
R79 VPWR.n8 VPWR.n7 15.4358
R80 VPWR.n12 VPWR.n3 12.424
R81 VPWR.n9 VPWR.n8 9.3005
R82 VPWR.n10 VPWR.n3 9.3005
R83 VPWR.n12 VPWR.n11 9.3005
R84 VPWR.n13 VPWR.n0 9.3005
R85 VPWR.n15 VPWR.n14 7.4836
R86 VPWR.n7 VPWR.n5 7.13828
R87 VPWR.n14 VPWR.n13 1.88285
R88 VPWR.n9 VPWR.n5 0.500685
R89 VPWR VPWR.n15 0.401983
R90 VPWR.n15 VPWR.n0 0.151923
R91 VPWR.n10 VPWR.n9 0.122949
R92 VPWR.n11 VPWR.n10 0.122949
R93 VPWR.n11 VPWR.n0 0.122949
R94 A2.n1 A2.t3 248.321
R95 A2.n3 A2.t2 240.197
R96 A2.n3 A2.t0 191.303
R97 A2 A2.n4 159.589
R98 A2.n1 A2.n0 152
R99 A2.n2 A2.t1 142.994
R100 A2.n2 A2.n1 27.6207
R101 A2.n4 A2.n3 14.623
R102 A2.n4 A2.n2 9.20724
R103 A2.n0 A2 9.2005
R104 A2 A2.n0 3.6005
R105 a_239_74.n1 a_239_74.t0 319.327
R106 a_239_74.t2 a_239_74.n1 282.123
R107 a_239_74.n1 a_239_74.n0 88.3446
R108 a_239_74.n0 a_239_74.t3 34.0546
R109 a_239_74.n0 a_239_74.t1 22.7032
R110 a_512_74.n1 a_512_74.n0 440.291
R111 a_512_74.n0 a_512_74.t3 22.7032
R112 a_512_74.n0 a_512_74.t2 22.7032
R113 a_512_74.n1 a_512_74.t0 22.7032
R114 a_512_74.t1 a_512_74.n1 22.7032
R115 A4.n0 A4.t1 226.809
R116 A4.n1 A4.t0 226.809
R117 A4.n1 A4.t3 198.204
R118 A4.n0 A4.t2 198.204
R119 A4.n3 A4.n2 152
R120 A4.n2 A4.n1 45.2793
R121 A4.n2 A4.n0 20.449
R122 A4 A4.n3 10.2703
R123 A4.n3 A4 4.0191
R124 A3.n0 A3.t2 333.651
R125 A3.n2 A3.t0 250.909
R126 A3.n1 A3.t1 206.969
R127 A3.n0 A3.t3 196.013
R128 A3.n3 A3.n2 152
R129 A3.n1 A3.n0 56.2338
R130 A3.n2 A3.n1 13.146
R131 A3.n3 A3 7.44236
R132 A3 A3.n3 6.84701
R133 a_709_74.n1 a_709_74.t2 308.851
R134 a_709_74.t1 a_709_74.n1 205.141
R135 a_709_74.n1 a_709_74.n0 102.144
R136 a_709_74.n0 a_709_74.t0 22.7032
R137 a_709_74.n0 a_709_74.t3 22.7032
C0 A1 A2 0.046131f
C1 VPB A4 0.066712f
C2 VPB Y 0.007655f
C3 B1 Y 0.119314f
C4 VPB VPWR 0.142749f
C5 A2 A3 0.086119f
C6 A2 A4 1.45e-19
C7 B1 VPWR 0.012258f
C8 A1 Y 0.160211f
C9 VPB VGND 0.00764f
C10 A2 Y 0.029599f
C11 A3 A4 0.089307f
C12 B1 VGND 0.052542f
C13 A1 VPWR 0.029435f
C14 A3 Y 3.12e-19
C15 A2 VPWR 0.037972f
C16 A1 VGND 0.012133f
C17 A2 VGND 0.019312f
C18 A3 VPWR 0.037484f
C19 A4 Y 1.09e-19
C20 VPB B1 0.070968f
C21 A4 VPWR 0.041727f
C22 A3 VGND 0.016944f
C23 VPB A1 0.080675f
C24 A4 VGND 0.036371f
C25 Y VPWR 0.029132f
C26 B1 A1 0.055657f
C27 VPB A2 0.074504f
C28 Y VGND 0.114882f
C29 VPB A3 0.070574f
C30 VPWR VGND 0.093124f
C31 VGND VNB 0.721858f
C32 VPWR VNB 0.534802f
C33 Y VNB 0.041324f
C34 A4 VNB 0.240908f
C35 A3 VNB 0.21805f
C36 A2 VNB 0.238073f
C37 A1 VNB 0.222536f
C38 B1 VNB 0.213309f
C39 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a41oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a41oi_1 VNB VPB VPWR VGND Y A2 A1 B1 A4 A3
X0 a_116_368.t4 B1.t0 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t3 A2.t0 a_116_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2296 pd=1.53 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_355_74.t1 A3.t0 a_277_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X3 a_116_368.t1 A3.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=1.81 w=1.12 l=0.15
X4 Y.t0 A1.t0 a_469_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 VGND.t1 B1.t1 Y.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VPWR.t2 A4.t0 a_116_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=1.81 as=0.196 ps=1.47 w=1.12 l=0.15
X7 a_277_74.t0 A4.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.24605 ps=1.405 w=0.74 l=0.15
X8 a_469_74.t1 A2.t1 a_355_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 a_116_368.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2296 ps=1.53 w=1.12 l=0.15
R0 B1.n0 B1.t0 256.428
R1 B1.n0 B1.t1 196.178
R2 B1 B1.n0 155.067
R3 Y.n0 Y.t0 301.933
R4 Y Y.t2 287.738
R5 Y.n0 Y.t1 159.251
R6 Y Y.n0 9.18311
R7 a_116_368.n2 a_116_368.n1 585
R8 a_116_368.n2 a_116_368.n0 348.284
R9 a_116_368.t0 a_116_368.n2 263.293
R10 a_116_368.n0 a_116_368.t4 35.1791
R11 a_116_368.n1 a_116_368.t3 26.3844
R12 a_116_368.n1 a_116_368.t1 26.3844
R13 a_116_368.n0 a_116_368.t2 26.3844
R14 VPB.t2 VPB.t1 429.033
R15 VPB.t3 VPB.t0 286.022
R16 VPB VPB.t4 257.93
R17 VPB.t4 VPB.t2 255.376
R18 VPB.t1 VPB.t3 229.839
R19 A2.n0 A2.t0 250.909
R20 A2.n0 A2.t1 220.113
R21 A2 A2.n0 157.805
R22 VPWR.n2 VPWR.n1 617.351
R23 VPWR.n2 VPWR.n0 292.151
R24 VPWR.n0 VPWR.t2 63.5898
R25 VPWR.n0 VPWR.t1 54.874
R26 VPWR.n1 VPWR.t0 36.0585
R27 VPWR.n1 VPWR.t3 36.0585
R28 VPWR VPWR.n2 0.575046
R29 A3.n0 A3.t1 250.909
R30 A3.n0 A3.t0 220.113
R31 A3 A3.n0 157.805
R32 a_277_74.t0 a_277_74.t1 38.9194
R33 a_355_74.t0 a_355_74.t1 68.1086
R34 VNB.t4 VNB.t1 1882.41
R35 VNB.t2 VNB.t0 1316.54
R36 VNB.t3 VNB.t2 1316.54
R37 VNB VNB.t4 1143.31
R38 VNB.t1 VNB.t3 900.788
R39 A1.n0 A1.t1 256.428
R40 A1.n0 A1.t0 196.178
R41 A1 A1.n0 156.462
R42 a_469_74.t0 a_469_74.t1 68.1086
R43 VGND VGND.n0 83.5068
R44 VGND.n0 VGND.t0 49.4909
R45 VGND.n0 VGND.t1 49.4328
R46 A4.n0 A4.t0 243.73
R47 A4.n0 A4.t1 212.935
R48 A4 A4.n0 154.522
C0 A2 A1 0.090455f
C1 A4 VPWR 0.01823f
C2 A3 Y 0.039897f
C3 B1 VGND 0.016103f
C4 A3 VPWR 0.021449f
C5 A2 Y 0.052818f
C6 A4 VGND 0.017575f
C7 A2 VPWR 0.021568f
C8 A3 VGND 0.009392f
C9 A1 Y 0.047013f
C10 VPB B1 0.043842f
C11 A2 VGND 0.010736f
C12 A1 VPWR 0.016804f
C13 VPB A4 0.043519f
C14 Y VPWR 0.047072f
C15 A1 VGND 0.011721f
C16 B1 A4 0.039071f
C17 VPB A3 0.036168f
C18 Y VGND 0.217057f
C19 VPB A2 0.033983f
C20 VPWR VGND 0.055301f
C21 A4 A3 0.085155f
C22 VPB A1 0.044556f
C23 VPB Y 0.015261f
C24 VPB VPWR 0.089952f
C25 A4 A1 4.56e-20
C26 B1 Y 0.151622f
C27 A3 A2 0.081004f
C28 A3 A1 7.39e-20
C29 B1 VPWR 0.011625f
C30 VPB VGND 0.005987f
C31 A4 Y 0.083799f
C32 VGND VNB 0.429218f
C33 VPWR VNB 0.339151f
C34 Y VNB 0.149193f
C35 A1 VNB 0.172202f
C36 A2 VNB 0.109192f
C37 A3 VNB 0.104191f
C38 A4 VNB 0.120376f
C39 B1 VNB 0.175169f
C40 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a41o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a41o_4 VNB VPB VPWR VGND X A3 A4 A1 A2 B1
X0 VPWR.t6 a_113_98.t6 X.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2009 pd=1.49 as=0.168 ps=1.42 w=1.12 l=0.15
X1 X.t2 a_113_98.t7 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_113_98.t3 B1.t0 a_27_392.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X3 a_113_98.t2 B1.t1 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2072 ps=2.04 w=0.74 l=0.15
X4 VPWR.t4 a_113_98.t8 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t1 A4.t0 a_27_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X6 X.t0 a_113_98.t9 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7 VPWR.t10 A1.t0 a_27_392.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.2625 pd=1.525 as=0.2475 ps=1.495 w=1 l=0.15
X8 a_27_392.t2 A4.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X9 a_751_74.t1 A1.t1 a_113_98.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 X.t7 a_113_98.t10 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1955 ps=1.43 w=0.74 l=0.15
X11 VPWR.t9 A2.t0 a_27_392.t5 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X12 a_27_392.t4 A2.t1 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2625 ps=1.525 w=1 l=0.15
X13 VGND.t3 a_113_98.t11 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.3495 pd=2.81 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_27_392.t8 B1.t2 a_113_98.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X15 a_27_392.t0 A1.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2475 pd=1.495 as=0.2009 ps=1.49 w=1 l=0.15
X16 a_113_98.t0 A1.t3 a_751_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X17 VPWR.t7 A3.t0 a_27_392.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X18 VGND A4 a_1205_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 X.t5 a_113_98.t12 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.193 ps=1.425 w=0.74 l=0.15
X20 a_1205_74# A4.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 a_27_392.t7 A3.t1 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.2 ps=1.4 w=1 l=0.15
X22 a_1205_74# A3.t2 a_1010_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_1010_74.t1 A2.t2 a_751_74.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VGND.t1 a_113_98.t13 X.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.193 pd=1.425 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 a_751_74.t3 A2.t3 a_1010_74.t0 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=2.03 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 VGND.t5 B1.t3 a_113_98.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1955 pd=1.43 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 a_113_98.n2 a_113_98.n0 433.993
R1 a_113_98.n15 a_113_98.n14 331.493
R2 a_113_98.n4 a_113_98.t6 292.293
R3 a_113_98.n5 a_113_98.t7 229.487
R4 a_113_98.n7 a_113_98.t8 229.487
R5 a_113_98.n9 a_113_98.t9 229.487
R6 a_113_98.n8 a_113_98.n3 165.189
R7 a_113_98.n12 a_113_98.t10 160.083
R8 a_113_98.n10 a_113_98.t13 154.24
R9 a_113_98.n6 a_113_98.t12 154.24
R10 a_113_98.n4 a_113_98.t11 154.24
R11 a_113_98.n13 a_113_98.n12 152
R12 a_113_98.n11 a_113_98.n3 152
R13 a_113_98.n2 a_113_98.n1 91.5745
R14 a_113_98.n6 a_113_98.n5 59.8853
R15 a_113_98.n12 a_113_98.n11 49.6611
R16 a_113_98.n15 a_113_98.t3 39.4005
R17 a_113_98.n8 a_113_98.n7 35.7853
R18 a_113_98.n9 a_113_98.n8 29.9429
R19 a_113_98.t1 a_113_98.n15 29.5505
R20 a_113_98.n0 a_113_98.t5 22.7032
R21 a_113_98.n0 a_113_98.t0 22.7032
R22 a_113_98.n1 a_113_98.t4 22.7032
R23 a_113_98.n1 a_113_98.t2 22.7032
R24 a_113_98.n14 a_113_98.n13 19.9901
R25 a_113_98.n13 a_113_98.n3 13.1884
R26 a_113_98.n10 a_113_98.n9 12.4157
R27 a_113_98.n11 a_113_98.n10 7.30353
R28 a_113_98.n14 a_113_98.n2 6.18615
R29 a_113_98.n7 a_113_98.n6 5.84292
R30 a_113_98.n5 a_113_98.n4 2.92171
R31 X.n2 X.n0 599.4
R32 X.n2 X.n1 585.513
R33 X.n5 X.n3 248.248
R34 X.n5 X.n4 185
R35 X.n1 X.t3 26.3844
R36 X.n1 X.t2 26.3844
R37 X.n0 X.t1 26.3844
R38 X.n0 X.t0 26.3844
R39 X.n4 X.t6 22.7032
R40 X.n4 X.t5 22.7032
R41 X.n3 X.t4 22.7032
R42 X.n3 X.t7 22.7032
R43 X X.n5 2.13383
R44 X X.n2 0.5125
R45 VPWR.n27 VPWR.t3 844.371
R46 VPWR.n25 VPWR.n2 607.303
R47 VPWR.n4 VPWR.n3 605.663
R48 VPWR.n9 VPWR.n8 316.305
R49 VPWR.n12 VPWR.n11 316.305
R50 VPWR.n18 VPWR.n7 309.861
R51 VPWR.n10 VPWR.t1 267.649
R52 VPWR.n7 VPWR.t8 52.2055
R53 VPWR.n7 VPWR.t10 51.2205
R54 VPWR.n3 VPWR.t0 41.3705
R55 VPWR.n8 VPWR.t11 39.4005
R56 VPWR.n8 VPWR.t9 39.4005
R57 VPWR.n11 VPWR.t2 39.4005
R58 VPWR.n20 VPWR.n19 36.1417
R59 VPWR.n18 VPWR.n17 32.0005
R60 VPWR.n3 VPWR.t6 29.6609
R61 VPWR.n11 VPWR.t7 29.5505
R62 VPWR.n13 VPWR.n9 28.9887
R63 VPWR.n26 VPWR.n25 27.4829
R64 VPWR.n2 VPWR.t5 26.3844
R65 VPWR.n2 VPWR.t4 26.3844
R66 VPWR.n24 VPWR.n4 22.9652
R67 VPWR.n20 VPWR.n4 22.9652
R68 VPWR.n13 VPWR.n12 21.4593
R69 VPWR.n25 VPWR.n24 19.9534
R70 VPWR.n17 VPWR.n9 18.4476
R71 VPWR.n27 VPWR.n26 15.4358
R72 VPWR.n14 VPWR.n13 9.3005
R73 VPWR.n15 VPWR.n9 9.3005
R74 VPWR.n17 VPWR.n16 9.3005
R75 VPWR.n18 VPWR.n6 9.3005
R76 VPWR.n19 VPWR.n5 9.3005
R77 VPWR.n21 VPWR.n20 9.3005
R78 VPWR.n22 VPWR.n4 9.3005
R79 VPWR.n24 VPWR.n23 9.3005
R80 VPWR.n25 VPWR.n1 9.3005
R81 VPWR.n26 VPWR.n0 9.3005
R82 VPWR.n28 VPWR.n27 7.51147
R83 VPWR.n12 VPWR.n10 6.8344
R84 VPWR.n19 VPWR.n18 5.64756
R85 VPWR.n14 VPWR.n10 0.569119
R86 VPWR VPWR.n28 0.402426
R87 VPWR.n28 VPWR.n0 0.151487
R88 VPWR.n15 VPWR.n14 0.122949
R89 VPWR.n16 VPWR.n15 0.122949
R90 VPWR.n16 VPWR.n6 0.122949
R91 VPWR.n6 VPWR.n5 0.122949
R92 VPWR.n21 VPWR.n5 0.122949
R93 VPWR.n22 VPWR.n21 0.122949
R94 VPWR.n23 VPWR.n22 0.122949
R95 VPWR.n23 VPWR.n1 0.122949
R96 VPWR.n1 VPWR.n0 0.122949
R97 VPB.t7 VPB.t3 515.861
R98 VPB.t12 VPB.t10 344.759
R99 VPB.t0 VPB.t12 329.435
R100 VPB.t11 VPB.t13 280.914
R101 VPB.t6 VPB.t0 265.591
R102 VPB VPB.t9 257.93
R103 VPB.t8 VPB.t2 255.376
R104 VPB.t13 VPB.t8 255.376
R105 VPB.t9 VPB.t7 255.376
R106 VPB.t2 VPB.t1 229.839
R107 VPB.t10 VPB.t11 229.839
R108 VPB.t5 VPB.t6 229.839
R109 VPB.t4 VPB.t5 229.839
R110 VPB.t3 VPB.t4 229.839
R111 B1.n2 B1.t0 234.091
R112 B1.n0 B1.t2 233.012
R113 B1.n1 B1.t1 208.868
R114 B1.n0 B1.t3 189.588
R115 B1 B1.n2 160.922
R116 B1.n1 B1.n0 51.3612
R117 B1.n2 B1.n1 1.9285
R118 a_27_392.n7 a_27_392.t9 302.262
R119 a_27_392.n2 a_27_392.n0 255.934
R120 a_27_392.t8 a_27_392.n7 221.968
R121 a_27_392.n7 a_27_392.n6 209.627
R122 a_27_392.n2 a_27_392.n1 205.487
R123 a_27_392.n4 a_27_392.n3 205.487
R124 a_27_392.n6 a_27_392.n5 195.66
R125 a_27_392.n6 a_27_392.n4 76.7139
R126 a_27_392.n4 a_27_392.n2 50.4476
R127 a_27_392.n5 a_27_392.t0 49.2505
R128 a_27_392.n5 a_27_392.t6 48.2655
R129 a_27_392.n1 a_27_392.t3 39.4005
R130 a_27_392.n0 a_27_392.t1 29.5505
R131 a_27_392.n0 a_27_392.t2 29.5505
R132 a_27_392.n1 a_27_392.t7 29.5505
R133 a_27_392.n3 a_27_392.t5 29.5505
R134 a_27_392.n3 a_27_392.t4 29.5505
R135 VGND.n5 VGND.t3 397.425
R136 VGND.n8 VGND.n7 249.727
R137 VGND.n12 VGND.n2 248.832
R138 VGND.n14 VGND.t6 178.762
R139 VGND.n4 VGND.t0 144.507
R140 VGND.n7 VGND.t2 34.8654
R141 VGND.n2 VGND.t4 34.8654
R142 VGND.n2 VGND.t5 34.8654
R143 VGND.n7 VGND.t1 34.0546
R144 VGND.n6 VGND.n5 31.2476
R145 VGND.n8 VGND.n1 28.2358
R146 VGND.n14 VGND.n13 27.1064
R147 VGND.n13 VGND.n12 24.4711
R148 VGND.n12 VGND.n1 22.9652
R149 VGND.n8 VGND.n6 19.2005
R150 VGND.n15 VGND.n14 9.3005
R151 VGND.n6 VGND.n3 9.3005
R152 VGND.n9 VGND.n8 9.3005
R153 VGND.n10 VGND.n1 9.3005
R154 VGND.n12 VGND.n11 9.3005
R155 VGND.n13 VGND.n0 9.3005
R156 VGND.n5 VGND.n4 7.06559
R157 VGND.n4 VGND.n3 0.158694
R158 VGND.n9 VGND.n3 0.122949
R159 VGND.n10 VGND.n9 0.122949
R160 VGND.n11 VGND.n10 0.122949
R161 VGND.n11 VGND.n0 0.122949
R162 VGND.n15 VGND.n0 0.122949
R163 VGND VGND.n15 0.0617245
R164 VNB.t8 VNB.t6 3245.14
R165 VNB.t4 VNB.t0 2725.46
R166 VNB.t6 VNB.t1 1986.35
R167 VNB.t10 VNB.t5 1339.63
R168 VNB.t2 VNB.t3 1328.08
R169 VNB VNB.t11 1131.76
R170 VNB.t7 VNB.t8 993.177
R171 VNB.t9 VNB.t7 993.177
R172 VNB.t0 VNB.t9 993.177
R173 VNB.t3 VNB.t4 993.177
R174 VNB.t5 VNB.t2 993.177
R175 VNB.t11 VNB.t10 993.177
R176 A4.n0 A4.t2 230.339
R177 A4.n2 A4.n1 228.148
R178 A4.n2 A4.t1 217.995
R179 A4.n0 A4.t0 212.883
R180 A4.n4 A4.n3 152
R181 A4.n3 A4.n2 36.5157
R182 A4.n3 A4.n0 24.1005
R183 A4 A4.n4 13.3823
R184 A4.n4 A4 5.23686
R185 A1.n2 A1.t2 234.062
R186 A1.n0 A1.t1 230.339
R187 A1.n1 A1.t3 228.148
R188 A1.n0 A1.t0 212.883
R189 A1 A1.n2 153.358
R190 A1.n1 A1.n0 60.6157
R191 A1.n2 A1.n1 12.4157
R192 a_751_74.n0 a_751_74.t0 242.858
R193 a_751_74.n0 a_751_74.t3 159.46
R194 a_751_74.n1 a_751_74.n0 89.408
R195 a_751_74.n1 a_751_74.t2 22.7032
R196 a_751_74.t1 a_751_74.n1 22.7032
R197 A2.n0 A2.t0 271.236
R198 A2.n2 A2.t2 241.292
R199 A2.n0 A2.t3 228.148
R200 A2.n1 A2.t1 212.883
R201 A2.n3 A2.n2 152
R202 A2.n1 A2.n0 29.2126
R203 A2.n2 A2.n1 20.449
R204 A2 A2.n3 14.352
R205 A2.n3 A2 4.26717
R206 A3.n0 A3.t2 243.483
R207 A3.n4 A3.n1 228.148
R208 A3.n3 A3.t1 223.839
R209 A3.n0 A3.t0 212.883
R210 A3.n6 A3.n5 152
R211 A3.n3 A3.n2 152
R212 A3.n5 A3.n4 35.055
R213 A3.n4 A3.n3 14.6066
R214 A3.n2 A3 14.1581
R215 A3.n5 A3.n0 12.4157
R216 A3 A3.n6 9.89141
R217 A3.n6 A3 8.72777
R218 A3.n2 A3 4.46111
R219 a_1010_74.n0 a_1010_74.t2 528.61
R220 a_1010_74.n0 a_1010_74.t0 22.7032
R221 a_1010_74.t1 a_1010_74.n0 22.7032
C0 VGND VPWR 0.133384f
C1 VPB A3 0.087469f
C2 a_1205_74# VPWR 0.003957f
C3 VGND X 0.03343f
C4 VPB A4 0.080334f
C5 A1 A2 0.070107f
C6 VPB VPWR 0.223517f
C7 VGND a_1205_74# 0.306315f
C8 A2 A3 0.057242f
C9 VPB X 0.012259f
C10 B1 VPWR 0.012583f
C11 B1 X 9.09e-19
C12 A1 VPWR 0.036283f
C13 VGND VPB 0.013763f
C14 a_1205_74# VPB 4.44e-19
C15 A1 X 0.031328f
C16 A2 VPWR 0.038122f
C17 A3 A4 0.091748f
C18 VGND B1 0.047249f
C19 A2 X 5.51e-19
C20 A3 VPWR 0.039649f
C21 VGND A1 0.013261f
C22 a_1205_74# A1 6.96e-20
C23 A4 VPWR 0.060489f
C24 A3 X 1.82e-19
C25 VGND A2 0.012351f
C26 a_1205_74# A2 8.72e-19
C27 VPB B1 0.102248f
C28 A4 X 1.1e-19
C29 VGND A3 0.013273f
C30 a_1205_74# A3 0.056908f
C31 VPB A1 0.097999f
C32 VPWR X 0.041449f
C33 VGND A4 0.03824f
C34 VPB A2 0.090389f
C35 a_1205_74# A4 0.097524f
C36 B1 A1 7.06e-19
C37 VGND VNB 0.990643f
C38 X VNB 0.016836f
C39 VPWR VNB 0.770831f
C40 A4 VNB 0.236438f
C41 A3 VNB 0.215564f
C42 A2 VNB 0.214694f
C43 A1 VNB 0.224644f
C44 B1 VNB 0.242371f
C45 VPB VNB 1.90613f
C46 a_1205_74# VNB 0.063896f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a41o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a41o_2 VNB VPB VPWR VGND A1 A2 A3 A4 B1 X
X0 a_441_74.t0 B1.t0 a_27_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.15 ps=1.3 w=1 l=0.15
X1 VPWR.t5 A4.t0 a_27_392.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.295 ps=2.59 w=1 l=0.15
X2 a_27_392.t1 A1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.29 ps=1.58 w=1 l=0.15
X3 VPWR.t1 A2.t0 a_27_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=1.58 as=0.15 ps=1.3 w=1 l=0.15
X4 a_27_392.t3 A3.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2 ps=1.4 w=1 l=0.15
X5 VPWR.t2 a_441_74.t3 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_199_74.t0 A3.t1 a_121_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X7 X.t1 a_441_74.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X8 VGND.t0 B1.t1 a_441_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1591 pd=1.17 as=0.1443 ps=1.13 w=0.74 l=0.15
X9 VGND.t2 a_441_74.t5 X.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.5772 pd=3.04 as=0.1517 ps=1.15 w=0.74 l=0.15
X10 a_313_74.t0 A2.t1 a_199_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1813 pd=1.23 as=0.1554 ps=1.16 w=0.74 l=0.15
X11 a_121_74.t1 A4.t1 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X12 X.t0 a_441_74.t6 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1517 pd=1.15 as=0.1591 ps=1.17 w=0.74 l=0.15
X13 a_441_74.t2 A1.t1 a_313_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1813 ps=1.23 w=0.74 l=0.15
R0 B1.n0 B1.t1 252.248
R1 B1.n0 B1.t0 236.983
R2 B1 B1.n0 159.952
R3 a_27_392.n1 a_27_392.t4 303.043
R4 a_27_392.n2 a_27_392.n1 269.486
R5 a_27_392.n1 a_27_392.n0 205.202
R6 a_27_392.n0 a_27_392.t2 29.5505
R7 a_27_392.n0 a_27_392.t3 29.5505
R8 a_27_392.t0 a_27_392.n2 29.5505
R9 a_27_392.n2 a_27_392.t1 29.5505
R10 a_441_74.n0 a_441_74.t3 325.156
R11 a_441_74.t0 a_441_74.n4 288.384
R12 a_441_74.n1 a_441_74.t4 261.62
R13 a_441_74.n2 a_441_74.t6 188.149
R14 a_441_74.n0 a_441_74.t5 154.24
R15 a_441_74.n4 a_441_74.n3 148.345
R16 a_441_74.n4 a_441_74.n2 72.3417
R17 a_441_74.n2 a_441_74.n1 38.912
R18 a_441_74.n3 a_441_74.t1 32.4329
R19 a_441_74.n3 a_441_74.t2 30.8113
R20 a_441_74.n1 a_441_74.n0 2.19141
R21 VPB.t0 VPB.t3 566.936
R22 VPB.t2 VPB.t1 372.849
R23 VPB.t6 VPB.t5 280.914
R24 VPB VPB.t6 257.93
R25 VPB.t3 VPB.t4 229.839
R26 VPB.t1 VPB.t0 229.839
R27 VPB.t5 VPB.t2 229.839
R28 A4.n0 A4.t0 291.041
R29 A4.n0 A4.t1 170.81
R30 A4 A4.n0 158.788
R31 VPWR.n6 VPWR.t3 351.815
R32 VPWR.n12 VPWR.n3 308.161
R33 VPWR.n5 VPWR.t2 265.579
R34 VPWR.n14 VPWR.n1 221.764
R35 VPWR.n3 VPWR.t0 57.1305
R36 VPWR.n3 VPWR.t1 57.1305
R37 VPWR.n1 VPWR.t4 39.4005
R38 VPWR.n1 VPWR.t5 39.4005
R39 VPWR.n7 VPWR.n4 36.1417
R40 VPWR.n11 VPWR.n4 36.1417
R41 VPWR.n13 VPWR.n12 31.2476
R42 VPWR.n14 VPWR.n13 19.2005
R43 VPWR.n7 VPWR.n6 17.6946
R44 VPWR.n8 VPWR.n7 9.3005
R45 VPWR.n9 VPWR.n4 9.3005
R46 VPWR.n11 VPWR.n10 9.3005
R47 VPWR.n12 VPWR.n2 9.3005
R48 VPWR.n13 VPWR.n0 9.3005
R49 VPWR.n15 VPWR.n14 7.43488
R50 VPWR.n6 VPWR.n5 6.96039
R51 VPWR.n12 VPWR.n11 2.63579
R52 VPWR.n8 VPWR.n5 0.594857
R53 VPWR VPWR.n15 0.160103
R54 VPWR.n15 VPWR.n0 0.1477
R55 VPWR.n9 VPWR.n8 0.122949
R56 VPWR.n10 VPWR.n9 0.122949
R57 VPWR.n10 VPWR.n2 0.122949
R58 VPWR.n2 VPWR.n0 0.122949
R59 A1.n0 A1.t1 252.248
R60 A1.n0 A1.t0 236.983
R61 A1 A1.n0 156.462
R62 A2.n0 A2.t0 294.356
R63 A2.n0 A2.t1 174.123
R64 A2 A2.n0 158.788
R65 A3.n0 A3.t0 298.572
R66 A3.n0 A3.t1 178.34
R67 A3 A3.n0 156.767
R68 X.n2 X.n0 312.096
R69 X.n2 X.n1 89.137
R70 X.n1 X.t0 36.487
R71 X.n1 X.t3 30.0005
R72 X.n0 X.t2 26.3844
R73 X.n0 X.t1 26.3844
R74 X X.n2 7.69861
R75 a_121_74.t0 a_121_74.t1 38.9194
R76 a_199_74.t0 a_199_74.t1 68.1086
R77 VNB.t4 VNB.t5 1478.22
R78 VNB.t1 VNB.t2 1339.63
R79 VNB.t0 VNB.t4 1316.54
R80 VNB.t2 VNB.t3 1293.44
R81 VNB.t5 VNB.t1 1247.24
R82 VNB VNB.t6 1224.15
R83 VNB.t6 VNB.t0 900.788
R84 VGND.n13 VGND.t3 155.453
R85 VGND.n3 VGND.t2 131.436
R86 VGND.n5 VGND.n4 115.659
R87 VGND.n7 VGND.n6 36.1417
R88 VGND.n7 VGND.n1 36.1417
R89 VGND.n11 VGND.n1 36.1417
R90 VGND.n12 VGND.n11 36.1417
R91 VGND.n4 VGND.t1 35.6762
R92 VGND.n4 VGND.t0 34.0546
R93 VGND.n13 VGND.n12 18.0711
R94 VGND.n6 VGND.n5 11.2946
R95 VGND.n14 VGND.n13 9.3005
R96 VGND.n6 VGND.n2 9.3005
R97 VGND.n8 VGND.n7 9.3005
R98 VGND.n9 VGND.n1 9.3005
R99 VGND.n11 VGND.n10 9.3005
R100 VGND.n12 VGND.n0 9.3005
R101 VGND.n5 VGND.n3 7.42972
R102 VGND.n3 VGND.n2 0.354742
R103 VGND.n8 VGND.n2 0.122949
R104 VGND.n9 VGND.n8 0.122949
R105 VGND.n10 VGND.n9 0.122949
R106 VGND.n10 VGND.n0 0.122949
R107 VGND.n14 VGND.n0 0.122949
R108 VGND VGND.n14 0.0617245
R109 a_313_74.t0 a_313_74.t1 79.46
C0 VPB X 0.00831f
C1 A4 VPWR 0.020549f
C2 A2 A1 0.064145f
C3 A2 B1 4.43e-19
C4 VPB VGND 0.011509f
C5 A3 VPWR 0.021944f
C6 A1 B1 0.086188f
C7 A2 VPWR 0.020388f
C8 A4 VGND 0.051507f
C9 A3 VGND 0.077326f
C10 A1 VPWR 0.016836f
C11 A2 VGND 0.038089f
C12 B1 VPWR 0.012107f
C13 VPB A4 0.049028f
C14 B1 X 3.98e-19
C15 A1 VGND 0.011742f
C16 VPB A3 0.037556f
C17 VPWR X 0.197816f
C18 B1 VGND 0.015581f
C19 VPB A2 0.043518f
C20 A4 A3 0.085557f
C21 VPWR VGND 0.093037f
C22 VPB A1 0.044927f
C23 X VGND 0.147737f
C24 A3 A2 0.159876f
C25 VPB B1 0.049305f
C26 A4 A1 2.07e-19
C27 A3 A1 4.41e-19
C28 VPB VPWR 0.151052f
C29 VGND VNB 0.643465f
C30 X VNB 0.047015f
C31 VPWR VNB 0.506656f
C32 B1 VNB 0.108756f
C33 A1 VNB 0.108998f
C34 A2 VNB 0.119707f
C35 A3 VNB 0.115475f
C36 A4 VNB 0.17022f
C37 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a41o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a41o_1 VNB VPB VPWR VGND A4 A1 A2 A3 B1 X
X0 a_354_392.t1 B1.t0 a_83_244.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X1 VPWR.t3 a_83_244.t3 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3304 ps=2.83 w=1.12 l=0.15
X2 VGND.t2 a_83_244.t4 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.7104 ps=3.4 w=0.74 l=0.15
X3 VPWR.t1 A3.t0 a_354_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.15 ps=1.3 w=1 l=0.15
X4 a_354_392.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.215 ps=1.43 w=1 l=0.15
X5 a_354_392.t4 A4.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.21 ps=1.42 w=1 l=0.15
X6 a_657_74.t1 A3.t1 a_543_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X7 a_83_244.t1 B1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8 a_543_74.t0 A2.t1 a_449_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1184 ps=1.06 w=0.74 l=0.15
X9 a_449_74.t1 A1.t0 a_83_244.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VGND.t0 A4.t1 a_657_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X11 VPWR.t2 A1.t1 a_354_392.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.215 pd=1.43 as=0.175 ps=1.35 w=1 l=0.15
R0 B1.n0 B1.t1 252.248
R1 B1.n0 B1.t0 236.983
R2 B1 B1.n0 154.133
R3 a_83_244.n1 a_83_244.t3 318.058
R4 a_83_244.t0 a_83_244.n2 263.986
R5 a_83_244.n1 a_83_244.t4 188.149
R6 a_83_244.n2 a_83_244.n0 143.827
R7 a_83_244.n2 a_83_244.n1 72.0508
R8 a_83_244.n0 a_83_244.t2 22.7032
R9 a_83_244.n0 a_83_244.t1 22.7032
R10 a_354_392.n1 a_354_392.t4 304.548
R11 a_354_392.n1 a_354_392.n0 258.193
R12 a_354_392.n2 a_354_392.n1 205.202
R13 a_354_392.n0 a_354_392.t1 39.4005
R14 a_354_392.n0 a_354_392.t3 29.5505
R15 a_354_392.n2 a_354_392.t2 29.5505
R16 a_354_392.t0 a_354_392.n2 29.5505
R17 VPB.t4 VPB.t1 607.797
R18 VPB.t3 VPB.t0 296.238
R19 VPB.t2 VPB.t5 291.13
R20 VPB VPB.t4 257.93
R21 VPB.t1 VPB.t3 255.376
R22 VPB.t0 VPB.t2 229.839
R23 X.n0 X.t0 283.438
R24 X.n0 X.t1 93.0157
R25 X X.n0 1.57588
R26 VPWR.n4 VPWR.n3 315.928
R27 VPWR.n10 VPWR.t3 259.171
R28 VPWR.n5 VPWR.n2 227.293
R29 VPWR.n3 VPWR.t0 45.3105
R30 VPWR.n2 VPWR.t4 43.3405
R31 VPWR.n3 VPWR.t2 39.4005
R32 VPWR.n2 VPWR.t1 39.4005
R33 VPWR.n8 VPWR.n1 36.1417
R34 VPWR.n9 VPWR.n8 36.1417
R35 VPWR.n10 VPWR.n9 22.9652
R36 VPWR.n4 VPWR.n1 10.9181
R37 VPWR.n6 VPWR.n1 9.3005
R38 VPWR.n8 VPWR.n7 9.3005
R39 VPWR.n9 VPWR.n0 9.3005
R40 VPWR.n5 VPWR.n4 7.61686
R41 VPWR.n11 VPWR.n10 7.52053
R42 VPWR.n6 VPWR.n5 0.528998
R43 VPWR VPWR.n11 0.161231
R44 VPWR.n11 VPWR.n0 0.146587
R45 VPWR.n7 VPWR.n6 0.122949
R46 VPWR.n7 VPWR.n0 0.122949
R47 VGND.n1 VGND.t0 163.436
R48 VGND.n1 VGND.n0 122.219
R49 VGND.n0 VGND.t1 34.0546
R50 VGND.n0 VGND.t2 34.0546
R51 VGND VGND.n1 0.378187
R52 VNB VNB.t3 2702.36
R53 VNB.t4 VNB.t0 1316.54
R54 VNB.t1 VNB.t4 1316.54
R55 VNB.t3 VNB.t2 1316.54
R56 VNB.t5 VNB.t1 1085.56
R57 VNB.t2 VNB.t5 993.177
R58 A3.n0 A3.t0 298.572
R59 A3.n0 A3.t1 178.34
R60 A3 A3.n0 159.439
R61 A2.n0 A2.t0 298.572
R62 A2.n0 A2.t1 178.34
R63 A2 A2.n0 158.054
R64 A4.n0 A4.t0 290.067
R65 A4.n0 A4.t1 169.834
R66 A4 A4.n0 158.788
R67 a_543_74.t0 a_543_74.t1 68.1086
R68 a_657_74.t0 a_657_74.t1 68.1086
R69 a_449_74.t0 a_449_74.t1 51.8924
R70 A1.n0 A1.t0 252.248
R71 A1.n0 A1.t1 236.983
R72 A1 A1.n0 156.462
C0 A1 VPWR 0.015143f
C1 A3 A4 0.090316f
C2 B1 VGND 0.014434f
C3 A1 VGND 0.01125f
C4 A2 VPWR 0.018098f
C5 A3 VPWR 0.020637f
C6 A2 VGND 0.050792f
C7 VPB B1 0.049688f
C8 A3 VGND 0.026439f
C9 A4 VPWR 0.020923f
C10 VPB A1 0.043247f
C11 X VPWR 0.129987f
C12 A4 VGND 0.050277f
C13 B1 A1 0.090664f
C14 VPB A2 0.038303f
C15 X VGND 0.17725f
C16 VPB A3 0.038048f
C17 B1 A2 4.99e-19
C18 VPWR VGND 0.070431f
C19 A1 A2 0.069978f
C20 VPB A4 0.051454f
C21 A1 A3 5.19e-19
C22 VPB X 0.014085f
C23 A2 A3 0.092292f
C24 B1 X 3.37e-19
C25 A1 A4 2.28e-19
C26 VPB VPWR 0.135066f
C27 A2 A4 0.001621f
C28 B1 VPWR 0.010848f
C29 VPB VGND 0.010846f
C30 VGND VNB 0.571349f
C31 VPWR VNB 0.428602f
C32 X VNB 0.118279f
C33 A4 VNB 0.174417f
C34 A3 VNB 0.112421f
C35 A2 VNB 0.116693f
C36 A1 VNB 0.105163f
C37 B1 VNB 0.105357f
C38 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a32oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32oi_4 VNB VPB VPWR VGND B2 B1 A3 A2 A1 Y
X0 Y.t10 B1.t0 a_27_368.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X1 VPWR.t3 A3.t0 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2268 pd=1.525 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_1313_74.t3 A3.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3 a_27_74.t3 B1.t1 Y.t6 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_27_368.t9 B1.t2 Y.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.2744 pd=1.61 as=0.196 ps=1.47 w=1.12 l=0.15
X5 VGND.t2 A3.t2 a_1313_74.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_27_74.t2 B1.t3 Y.t5 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t11 A2.t0 a_27_368.t19 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1736 ps=1.43 w=1.12 l=0.15
X8 a_868_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VGND.t1 A3.t3 a_1313_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 Y.t13 B2.t0 a_27_368.t17 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.336 ps=2.84 w=1.12 l=0.15
X11 VPWR.t9 A2.t1 a_27_368.t15 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_27_368.t16 A2.t2 VPWR.t10 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2184 ps=1.51 w=1.12 l=0.15
X13 a_868_74# A1.t0 Y.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X14 a_27_368.t18 B2.t1 Y.t14 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X15 VGND.t7 B2.t2 a_27_74.t7 VNB.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X16 Y.t11 B2.t3 a_27_368.t11 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_27_368.t13 A3.t4 VPWR.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X18 a_27_368.t12 B2.t4 Y.t12 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1932 ps=1.465 w=1.12 l=0.15
X19 Y.t8 B1.t4 a_27_368.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X20 a_27_368.t3 A1.t1 VPWR.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X21 VPWR.t6 A1.t2 a_27_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.168 ps=1.42 w=1.12 l=0.15
X22 Y.t4 B1.t5 a_27_74.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_868_74# A2.t3 a_1313_74.t6 VNB.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 VGND.t4 B2.t5 a_27_74.t4 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.12765 pd=1.085 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 Y.t1 A1.t3 a_868_74# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X26 VPWR.t1 A3.t5 a_27_368.t14 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X27 a_27_368.t1 A3.t6 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2268 ps=1.525 w=1.12 l=0.15
X28 VPWR.t7 A1.t4 a_27_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2744 ps=1.61 w=1.12 l=0.15
X29 a_27_368.t7 B1.t6 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X30 a_27_74.t5 B2.t6 VGND.t5 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12765 ps=1.085 w=0.74 l=0.15
X31 a_1313_74.t4 A2.t4 a_868_74# VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.10545 ps=1.025 w=0.74 l=0.15
X32 a_27_74.t6 B2.t7 VGND.t6 VNB.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X33 a_27_368.t6 A1.t5 VPWR.t8 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.224 ps=1.52 w=1.12 l=0.15
X34 Y.t3 B1.t7 a_27_74.t0 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X35 a_1313_74.t5 A2.t5 a_868_74# VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X36 a_1313_74.t0 A3.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X37 a_27_368.t0 A2.t6 VPWR.t4 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X38 Y.t2 A1.t6 a_868_74# VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 B1.n13 B1.t2 242.144
R1 B1.n0 B1.t4 226.809
R2 B1.n7 B1.t6 226.809
R3 B1.n2 B1.t0 226.809
R4 B1.n2 B1.t5 204.048
R5 B1.n6 B1.t3 196.013
R6 B1.n1 B1.t7 196.013
R7 B1.n12 B1.t1 196.013
R8 B1.n14 B1.n13 152
R9 B1.n11 B1.n10 152
R10 B1.n9 B1.n8 152
R11 B1.n6 B1.n5 152
R12 B1.n4 B1.n3 152
R13 B1.n6 B1.n3 49.6611
R14 B1.n12 B1.n11 36.5157
R15 B1.n8 B1.n7 31.4035
R16 B1.n8 B1.n1 23.3702
R17 B1.n1 B1.n0 18.2581
R18 B1.n7 B1.n6 18.2581
R19 B1.n13 B1.n12 13.146
R20 B1.n4 B1 10.8656
R21 B1.n10 B1.n9 10.1214
R22 B1.n14 B1 8.48422
R23 B1.n11 B1.n0 8.03383
R24 B1.n5 B1 7.5912
R25 B1.n5 B1 6.69817
R26 B1 B1.n14 5.80515
R27 B1.n3 B1.n2 5.11262
R28 B1 B1.n4 3.42376
R29 B1.n9 B1 2.53073
R30 B1.n10 B1 1.63771
R31 a_27_368.n1 a_27_368.n0 305.901
R32 a_27_368.n3 a_27_368.n2 302.74
R33 a_27_368.n5 a_27_368.n4 302.74
R34 a_27_368.n9 a_27_368.n8 299.053
R35 a_27_368.n11 a_27_368.n10 299.053
R36 a_27_368.n1 a_27_368.t17 295.541
R37 a_27_368.n7 a_27_368.n6 289.051
R38 a_27_368.n15 a_27_368.t1 282.695
R39 a_27_368.n15 a_27_368.n14 205.487
R40 a_27_368.n17 a_27_368.n16 205.486
R41 a_27_368.n13 a_27_368.n12 195.787
R42 a_27_368.n9 a_27_368.n7 67.227
R43 a_27_368.n7 a_27_368.n5 64.1354
R44 a_27_368.n16 a_27_368.n13 60.1471
R45 a_27_368.n3 a_27_368.n1 59.1064
R46 a_27_368.n13 a_27_368.n11 53.8232
R47 a_27_368.n6 a_27_368.t5 51.0094
R48 a_27_368.n5 a_27_368.n3 50.4476
R49 a_27_368.n11 a_27_368.n9 50.4476
R50 a_27_368.n16 a_27_368.n15 50.4476
R51 a_27_368.n14 a_27_368.t13 35.1791
R52 a_27_368.n6 a_27_368.t9 35.1791
R53 a_27_368.n2 a_27_368.t18 35.1791
R54 a_27_368.n4 a_27_368.t7 35.1791
R55 a_27_368.t0 a_27_368.n17 35.1791
R56 a_27_368.n10 a_27_368.t19 28.1434
R57 a_27_368.n14 a_27_368.t2 26.3844
R58 a_27_368.n12 a_27_368.t15 26.3844
R59 a_27_368.n12 a_27_368.t16 26.3844
R60 a_27_368.n0 a_27_368.t11 26.3844
R61 a_27_368.n0 a_27_368.t12 26.3844
R62 a_27_368.n2 a_27_368.t10 26.3844
R63 a_27_368.n4 a_27_368.t8 26.3844
R64 a_27_368.n8 a_27_368.t4 26.3844
R65 a_27_368.n8 a_27_368.t3 26.3844
R66 a_27_368.n10 a_27_368.t6 26.3844
R67 a_27_368.n17 a_27_368.t14 26.3844
R68 Y.n2 Y.n0 342.868
R69 Y.n2 Y.n1 299.95
R70 Y.n4 Y.n3 299.95
R71 Y.n6 Y.n5 299.95
R72 Y.n7 Y.t2 275
R73 Y Y.n6 256.397
R74 Y.n10 Y.n8 224.234
R75 Y.n10 Y.n9 185
R76 Y.n12 Y.n11 185
R77 Y Y.n10 98.5963
R78 Y.n4 Y.n2 50.4476
R79 Y.n6 Y.n4 50.4476
R80 Y.n3 Y.t10 35.1791
R81 Y.n5 Y.t8 35.1791
R82 Y.n0 Y.t13 34.2996
R83 Y.n11 Y.t1 34.0546
R84 Y.n0 Y.t12 26.3844
R85 Y.n1 Y.t14 26.3844
R86 Y.n1 Y.t11 26.3844
R87 Y.n3 Y.t7 26.3844
R88 Y.n5 Y.t9 26.3844
R89 Y.n11 Y.t0 22.7032
R90 Y.n9 Y.t6 22.7032
R91 Y.n9 Y.t3 22.7032
R92 Y.n8 Y.t5 22.7032
R93 Y.n8 Y.t4 22.7032
R94 Y Y.n12 15.2851
R95 Y Y.n7 14.5783
R96 Y.n7 Y 2.48939
R97 Y.n12 Y 0.937085
R98 VPB.t9 VPB.t5 326.882
R99 VPB.t2 VPB.t1 283.469
R100 VPB.t4 VPB.t6 280.914
R101 VPB.t19 VPB.t16 275.807
R102 VPB VPB.t17 260.485
R103 VPB.t13 VPB.t2 255.376
R104 VPB.t14 VPB.t13 255.376
R105 VPB.t0 VPB.t14 255.376
R106 VPB.t15 VPB.t0 255.376
R107 VPB.t5 VPB.t3 255.376
R108 VPB.t8 VPB.t9 255.376
R109 VPB.t7 VPB.t8 255.376
R110 VPB.t10 VPB.t7 255.376
R111 VPB.t18 VPB.t10 255.376
R112 VPB.t17 VPB.t12 252.823
R113 VPB.t6 VPB.t19 234.946
R114 VPB.t16 VPB.t15 229.839
R115 VPB.t3 VPB.t4 229.839
R116 VPB.t11 VPB.t18 229.839
R117 VPB.t12 VPB.t11 229.839
R118 A3.n3 A3.t5 294.8
R119 A3.n0 A3.t6 226.809
R120 A3.n1 A3.t0 226.809
R121 A3.n5 A3.t4 226.809
R122 A3.n0 A3.t2 198.204
R123 A3.n3 A3.t1 196.013
R124 A3.n6 A3.t3 196.013
R125 A3.n11 A3.t7 196.013
R126 A3.n13 A3.n12 152
R127 A3.n10 A3.n9 152
R128 A3.n8 A3.n7 152
R129 A3.n4 A3.n2 152
R130 A3.n12 A3.n11 46.0096
R131 A3.n7 A3.n1 32.8641
R132 A3.n6 A3.n5 30.6732
R133 A3.n4 A3.n3 22.6399
R134 A3.n10 A3.n1 16.7975
R135 A3.n12 A3.n0 14.6066
R136 A3.n8 A3.n2 10.1214
R137 A3.n9 A3 9.97259
R138 A3.n7 A3.n6 9.49444
R139 A3.n5 A3.n4 9.49444
R140 A3 A3.n13 8.48422
R141 A3.n13 A3 5.80515
R142 A3.n9 A3 4.31678
R143 A3.n2 A3 4.0191
R144 A3.n11 A3.n10 3.65202
R145 A3 A3.n8 0.149337
R146 VPWR.n26 VPWR.n1 605.365
R147 VPWR.n3 VPWR.n2 605.365
R148 VPWR.n19 VPWR.n5 605.365
R149 VPWR.n10 VPWR.n9 321.521
R150 VPWR.n14 VPWR.n8 315.928
R151 VPWR.n12 VPWR.n11 315.928
R152 VPWR.n25 VPWR.n24 36.1417
R153 VPWR.n21 VPWR.n20 36.1417
R154 VPWR.n18 VPWR.n6 36.1417
R155 VPWR.n9 VPWR.t0 36.0585
R156 VPWR.n1 VPWR.t5 35.1791
R157 VPWR.n2 VPWR.t8 35.1791
R158 VPWR.n2 VPWR.t6 35.1791
R159 VPWR.n5 VPWR.t10 35.1791
R160 VPWR.n8 VPWR.t9 35.1791
R161 VPWR.n11 VPWR.t1 35.1791
R162 VPWR.n9 VPWR.t3 35.1791
R163 VPWR.n14 VPWR.n13 35.0123
R164 VPWR.n5 VPWR.t11 33.4201
R165 VPWR.n1 VPWR.t7 26.3844
R166 VPWR.n8 VPWR.t4 26.3844
R167 VPWR.n11 VPWR.t2 26.3844
R168 VPWR.n13 VPWR.n12 15.4358
R169 VPWR.n14 VPWR.n6 12.424
R170 VPWR.n27 VPWR.n26 11.0387
R171 VPWR.n20 VPWR.n19 9.41227
R172 VPWR.n13 VPWR.n7 9.3005
R173 VPWR.n15 VPWR.n14 9.3005
R174 VPWR.n16 VPWR.n6 9.3005
R175 VPWR.n18 VPWR.n17 9.3005
R176 VPWR.n20 VPWR.n4 9.3005
R177 VPWR.n22 VPWR.n21 9.3005
R178 VPWR.n24 VPWR.n23 9.3005
R179 VPWR.n25 VPWR.n0 9.3005
R180 VPWR.n26 VPWR.n25 7.90638
R181 VPWR.n12 VPWR.n10 7.10021
R182 VPWR.n24 VPWR.n3 6.4005
R183 VPWR.n21 VPWR.n3 4.89462
R184 VPWR.n19 VPWR.n18 1.88285
R185 VPWR VPWR.n27 1.14267
R186 VPWR.n10 VPWR.n7 0.532715
R187 VPWR.n27 VPWR.n0 0.149471
R188 VPWR.n15 VPWR.n7 0.122949
R189 VPWR.n16 VPWR.n15 0.122949
R190 VPWR.n17 VPWR.n16 0.122949
R191 VPWR.n17 VPWR.n4 0.122949
R192 VPWR.n22 VPWR.n4 0.122949
R193 VPWR.n23 VPWR.n22 0.122949
R194 VPWR.n23 VPWR.n0 0.122949
R195 VGND.n14 VGND.t3 269.132
R196 VGND.n12 VGND.n11 208.079
R197 VGND.n36 VGND.n2 208.079
R198 VGND.n39 VGND.n38 208.079
R199 VGND.n10 VGND.t2 170.607
R200 VGND.n18 VGND.n8 36.1417
R201 VGND.n19 VGND.n18 36.1417
R202 VGND.n20 VGND.n19 36.1417
R203 VGND.n20 VGND.n6 36.1417
R204 VGND.n24 VGND.n6 36.1417
R205 VGND.n25 VGND.n24 36.1417
R206 VGND.n26 VGND.n25 36.1417
R207 VGND.n26 VGND.n4 36.1417
R208 VGND.n30 VGND.n4 36.1417
R209 VGND.n31 VGND.n30 36.1417
R210 VGND.n32 VGND.n31 36.1417
R211 VGND.n32 VGND.n1 36.1417
R212 VGND.n14 VGND.n8 35.7652
R213 VGND.n38 VGND.t7 34.0546
R214 VGND.n2 VGND.t5 33.2437
R215 VGND.n13 VGND.n12 28.2358
R216 VGND.n36 VGND.n1 26.7299
R217 VGND.n11 VGND.t0 22.7032
R218 VGND.n11 VGND.t1 22.7032
R219 VGND.n2 VGND.t4 22.7032
R220 VGND.n38 VGND.t6 22.7032
R221 VGND.n37 VGND.n36 20.7064
R222 VGND.n39 VGND.n37 19.2005
R223 VGND.n14 VGND.n13 11.6711
R224 VGND.n37 VGND.n0 9.3005
R225 VGND.n36 VGND.n35 9.3005
R226 VGND.n34 VGND.n1 9.3005
R227 VGND.n33 VGND.n32 9.3005
R228 VGND.n31 VGND.n3 9.3005
R229 VGND.n30 VGND.n29 9.3005
R230 VGND.n28 VGND.n4 9.3005
R231 VGND.n27 VGND.n26 9.3005
R232 VGND.n25 VGND.n5 9.3005
R233 VGND.n24 VGND.n23 9.3005
R234 VGND.n22 VGND.n6 9.3005
R235 VGND.n21 VGND.n20 9.3005
R236 VGND.n19 VGND.n7 9.3005
R237 VGND.n18 VGND.n17 9.3005
R238 VGND.n16 VGND.n8 9.3005
R239 VGND.n15 VGND.n14 9.3005
R240 VGND.n13 VGND.n9 9.3005
R241 VGND.n40 VGND.n39 7.43488
R242 VGND.n12 VGND.n10 6.26985
R243 VGND.n10 VGND.n9 0.733933
R244 VGND VGND.n40 0.160103
R245 VGND.n40 VGND.n0 0.1477
R246 VGND.n15 VGND.n9 0.122949
R247 VGND.n16 VGND.n15 0.122949
R248 VGND.n17 VGND.n16 0.122949
R249 VGND.n17 VGND.n7 0.122949
R250 VGND.n21 VGND.n7 0.122949
R251 VGND.n22 VGND.n21 0.122949
R252 VGND.n23 VGND.n22 0.122949
R253 VGND.n23 VGND.n5 0.122949
R254 VGND.n27 VGND.n5 0.122949
R255 VGND.n28 VGND.n27 0.122949
R256 VGND.n29 VGND.n28 0.122949
R257 VGND.n29 VGND.n3 0.122949
R258 VGND.n33 VGND.n3 0.122949
R259 VGND.n34 VGND.n33 0.122949
R260 VGND.n35 VGND.n34 0.122949
R261 VGND.n35 VGND.n0 0.122949
R262 a_1313_74.n2 a_1313_74.t5 308.553
R263 a_1313_74.n2 a_1313_74.n1 185
R264 a_1313_74.n3 a_1313_74.n0 168.403
R265 a_1313_74.n4 a_1313_74.n3 103.65
R266 a_1313_74.n3 a_1313_74.n2 100.894
R267 a_1313_74.n1 a_1313_74.t6 22.7032
R268 a_1313_74.n1 a_1313_74.t4 22.7032
R269 a_1313_74.n0 a_1313_74.t2 22.7032
R270 a_1313_74.n0 a_1313_74.t0 22.7032
R271 a_1313_74.n4 a_1313_74.t1 22.7032
R272 a_1313_74.t3 a_1313_74.n4 22.7032
R273 VNB.t16 VNB.t3 2286.61
R274 VNB.t12 VNB.t7 2286.61
R275 VNB.t5 VNB.t4 1997.9
R276 VNB.t8 VNB.t5 1986.35
R277 VNB.t7 VNB.t6 1154.86
R278 VNB.t11 VNB.t9 1154.86
R279 VNB.t17 VNB.t15 1154.86
R280 VNB.t13 VNB.t14 1143.31
R281 VNB VNB.t17 1143.31
R282 VNB.t0 VNB.t2 993.177
R283 VNB.t1 VNB.t0 993.177
R284 VNB.t3 VNB.t1 993.177
R285 VNB.t4 VNB.t16 993.177
R286 VNB.t6 VNB.t8 993.177
R287 VNB.t9 VNB.t12 993.177
R288 VNB.t10 VNB.t11 993.177
R289 VNB.t14 VNB.t10 993.177
R290 VNB.t15 VNB.t13 993.177
R291 a_27_74.t3 a_27_74.n5 325.339
R292 a_27_74.n1 a_27_74.t7 206.744
R293 a_27_74.n5 a_27_74.n4 185
R294 a_27_74.n1 a_27_74.n0 103.65
R295 a_27_74.n3 a_27_74.n1 88.5562
R296 a_27_74.n3 a_27_74.n2 84.741
R297 a_27_74.n5 a_27_74.n3 84.5392
R298 a_27_74.n4 a_27_74.t2 34.0546
R299 a_27_74.n4 a_27_74.t0 22.7032
R300 a_27_74.n2 a_27_74.t1 22.7032
R301 a_27_74.n2 a_27_74.t5 22.7032
R302 a_27_74.n0 a_27_74.t4 22.7032
R303 a_27_74.n0 a_27_74.t6 22.7032
R304 A2.n1 A2.t6 237.762
R305 A2.n12 A2.t1 226.809
R306 A2.n3 A2.t2 226.809
R307 A2.n6 A2.t0 226.809
R308 A2.n6 A2.t5 198.204
R309 A2.n5 A2.n4 196.013
R310 A2.n11 A2.t4 196.013
R311 A2.n2 A2.t3 196.013
R312 A2.n1 A2.n0 152
R313 A2.n14 A2.n13 152
R314 A2.n10 A2.n9 152
R315 A2.n8 A2.n7 152
R316 A2.n7 A2.n6 57.6944
R317 A2.n13 A2.n2 29.9429
R318 A2.n10 A2.n3 28.4823
R319 A2.n12 A2.n11 20.449
R320 A2.n2 A2.n1 19.7187
R321 A2.n5 A2.n3 18.2581
R322 A2.n11 A2.n10 16.7975
R323 A2.n13 A2.n12 12.4157
R324 A2.n0 A2 11.7586
R325 A2.n9 A2.n8 10.1214
R326 A2 A2.n14 7.5912
R327 A2.n14 A2 6.69817
R328 A2.n9 A2 3.42376
R329 A2.n7 A2.n5 2.92171
R330 A2 A2.n0 2.53073
R331 A2.n8 A2 0.744686
R332 A1.n7 A1.t4 237.762
R333 A1.n1 A1.t5 226.809
R334 A1.n5 A1.t2 226.809
R335 A1.n10 A1.t1 226.809
R336 A1.n1 A1.n0 198.204
R337 A1.n8 A1.t3 196.013
R338 A1.n11 A1.t0 196.013
R339 A1.n4 A1.t6 196.013
R340 A1 A1.n2 158.102
R341 A1.n13 A1.n12 152
R342 A1.n9 A1.n3 152
R343 A1.n7 A1.n6 152
R344 A1.n2 A1.n1 59.155
R345 A1.n9 A1.n8 37.9763
R346 A1.n12 A1.n5 28.4823
R347 A1.n11 A1.n10 22.6399
R348 A1.n5 A1.n4 19.7187
R349 A1.n12 A1.n11 14.6066
R350 A1.n10 A1.n9 12.4157
R351 A1.n8 A1.n7 11.6853
R352 A1.n13 A1.n3 10.1214
R353 A1.n6 A1 9.97259
R354 A1.n6 A1 4.31678
R355 A1 A1.n13 4.0191
R356 A1.n4 A1.n2 1.46111
R357 A1 A1.n3 0.149337
R358 B2.n0 B2.t1 226.809
R359 B2.n2 B2.t3 226.809
R360 B2.n10 B2.t4 226.809
R361 B2.n4 B2.t0 226.809
R362 B2.n4 B2.t2 198.204
R363 B2.n0 B2.t6 198.204
R364 B2.n9 B2.t7 196.013
R365 B2.n3 B2.t5 196.013
R366 B2 B2.n1 152.298
R367 B2.n12 B2.n11 152
R368 B2.n8 B2.n7 152
R369 B2.n6 B2.n5 152
R370 B2.n8 B2.n5 49.6611
R371 B2.n1 B2.n0 43.8187
R372 B2.n11 B2.n10 37.9763
R373 B2.n11 B2.n3 23.3702
R374 B2.n2 B2.n1 21.9096
R375 B2.n6 B2 12.8005
R376 B2.n5 B2.n4 10.955
R377 B2.n9 B2.n8 10.2247
R378 B2 B2.n12 9.82376
R379 B2.n7 B2 8.63306
R380 B2.n7 B2 5.65631
R381 B2.n12 B2 4.46562
R382 B2.n3 B2.n2 4.38232
R383 B2 B2.n6 1.48887
R384 B2.n10 B2.n9 1.46111
C0 B2 B1 0.089308f
C1 VPB A1 0.147004f
C2 a_868_74# Y 0.200976f
C3 Y VGND 0.051711f
C4 VPB A2 0.145966f
C5 a_868_74# VPWR 0.004394f
C6 VPWR VGND 0.166751f
C7 a_868_74# VGND 0.368289f
C8 VPB A3 0.155155f
C9 B1 A1 0.058151f
C10 VPB Y 0.011693f
C11 VPB VPWR 0.240221f
C12 B2 Y 0.16311f
C13 A1 A2 0.055438f
C14 a_868_74# VPB 1.22e-19
C15 B1 Y 0.44352f
C16 VPB VGND 0.009595f
C17 B2 VPWR 0.025621f
C18 B2 VGND 0.072769f
C19 A1 Y 0.33816f
C20 B1 VPWR 0.025699f
C21 A2 A3 0.071996f
C22 a_868_74# B1 9.55e-19
C23 A1 VPWR 0.050354f
C24 A2 Y 0.041168f
C25 B1 VGND 0.026882f
C26 a_868_74# A1 0.033654f
C27 A1 VGND 0.025437f
C28 A2 VPWR 0.06732f
C29 A3 Y 4.27e-19
C30 VPB B2 0.142534f
C31 a_868_74# A2 0.036279f
C32 A3 VPWR 0.078562f
C33 A2 VGND 0.029688f
C34 VPB B1 0.15277f
C35 a_868_74# A3 6.98e-20
C36 A3 VGND 0.10329f
C37 Y VPWR 0.069939f
C38 VGND VNB 1.22098f
C39 VPWR VNB 0.935831f
C40 Y VNB 0.045894f
C41 A3 VNB 0.465262f
C42 A2 VNB 0.417445f
C43 A1 VNB 0.416217f
C44 B1 VNB 0.426749f
C45 B2 VNB 0.450244f
C46 VPB VNB 2.44181f
C47 a_868_74# VNB 0.025707f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a32oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32oi_2 VNB VPB VPWR VGND B2 B1 A3 A2 A1 Y
X0 Y.t2 B1.t0 a_27_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X1 a_27_368.t2 A3.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2 Y.t4 B1.t1 a_27_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_507_74.t2 A1.t0 Y.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.11285 pd=1.045 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t1 A3.t1 a_771_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 Y.t6 B2.t0 a_27_368.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.465 as=0.336 ps=2.84 w=1.12 l=0.15
X6 VPWR.t3 A2.t0 a_27_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2044 pd=1.485 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_27_368.t8 A1.t1 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=1.81 w=1.12 l=0.15
X8 VGND.t3 B2.t1 a_27_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_27_368.t0 B2.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.1932 ps=1.465 w=1.12 l=0.15
X10 Y.t5 A1.t2 a_507_74.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X11 VPWR.t4 A1.t3 a_27_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3864 pd=1.81 as=0.196 ps=1.47 w=1.12 l=0.15
X12 a_27_368.t1 A2.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.266 pd=1.595 as=0.2044 ps=1.485 w=1.12 l=0.15
X13 a_771_74.t0 A3.t2 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 VPWR.t1 A3.t3 a_27_368.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.266 ps=1.595 w=1.12 l=0.15
X15 a_507_74.t3 A2.t2 a_771_74.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.14615 ps=1.135 w=0.74 l=0.15
X16 a_771_74.t2 A2.t3 a_507_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.14615 pd=1.135 as=0.11285 ps=1.045 w=0.74 l=0.15
X17 a_27_368.t3 B1.t2 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X18 a_27_74.t0 B1.t3 Y.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_27_74.t2 B2.t3 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
R0 B1.n1 B1.t2 261.62
R1 B1.n3 B1.t0 261.62
R2 B1.n3 B1.t1 172.125
R3 B1.n2 B1.t3 154.24
R4 B1.n1 B1.n0 152.731
R5 B1.n5 B1.n4 152
R6 B1.n2 B1.n1 24.8308
R7 B1.n4 B1.n2 24.1005
R8 B1.n4 B1.n3 24.1005
R9 B1.n5 B1.n0 11.7627
R10 B1 B1.n5 2.59509
R11 B1.n0 B1 2.24915
R12 a_27_368.n3 a_27_368.n2 585
R13 a_27_368.n4 a_27_368.n1 305.659
R14 a_27_368.n9 a_27_368.n8 304.481
R15 a_27_368.n3 a_27_368.t2 297.7
R16 a_27_368.n8 a_27_368.t9 286.882
R17 a_27_368.n5 a_27_368.n0 204.643
R18 a_27_368.n7 a_27_368.n6 188.306
R19 a_27_368.n7 a_27_368.n5 106.484
R20 a_27_368.n8 a_27_368.n7 72.4324
R21 a_27_368.n5 a_27_368.n4 54.0471
R22 a_27_368.n1 a_27_368.t1 35.1791
R23 a_27_368.n6 a_27_368.t3 35.1791
R24 a_27_368.t0 a_27_368.n9 35.1791
R25 a_27_368.n0 a_27_368.t5 26.3844
R26 a_27_368.n0 a_27_368.t8 26.3844
R27 a_27_368.n2 a_27_368.t7 26.3844
R28 a_27_368.n6 a_27_368.t6 26.3844
R29 a_27_368.n9 a_27_368.t4 26.3844
R30 a_27_368.n2 a_27_368.n1 21.9871
R31 a_27_368.n4 a_27_368.n3 1.40709
R32 Y.n5 Y.n3 281.949
R33 Y.n2 Y.n0 255.727
R34 Y.n2 Y.n1 205.475
R35 Y.n5 Y.n4 195.829
R36 Y Y.n2 95.437
R37 Y Y.n5 39.0405
R38 Y.n1 Y.t2 35.1791
R39 Y.n0 Y.t6 34.2996
R40 Y.n1 Y.t1 26.3844
R41 Y.n0 Y.t0 26.3844
R42 Y.n3 Y.t3 22.7032
R43 Y.n3 Y.t4 22.7032
R44 Y.n4 Y.t7 22.7032
R45 Y.n4 Y.t5 22.7032
R46 VPB.t6 VPB.t8 429.033
R47 VPB.t1 VPB.t7 319.221
R48 VPB.t7 VPB.t2 280.914
R49 VPB.t5 VPB.t1 263.038
R50 VPB VPB.t9 260.485
R51 VPB.t3 VPB.t6 255.376
R52 VPB.t4 VPB.t3 255.376
R53 VPB.t0 VPB.t4 255.376
R54 VPB.t9 VPB.t0 252.823
R55 VPB.t8 VPB.t5 229.839
R56 A3.n0 A3.t3 317.123
R57 A3.n1 A3.t0 261.62
R58 A3 A3.n2 188.731
R59 A3.n0 A3.t2 154.24
R60 A3.n2 A3.t1 154.24
R61 A3.n2 A3.n1 37.9763
R62 A3.n1 A3.n0 24.8308
R63 VPWR.n3 VPWR.n1 585
R64 VPWR.n2 VPWR.n1 585
R65 VPWR.n9 VPWR.n8 315.634
R66 VPWR.n5 VPWR.n4 276.695
R67 VPWR.n7 VPWR.n6 226.929
R68 VPWR.n8 VPWR.t3 36.0585
R69 VPWR.n6 VPWR.t2 35.1791
R70 VPWR.n6 VPWR.t1 35.1791
R71 VPWR.n4 VPWR.n3 31.6146
R72 VPWR.n4 VPWR.n2 31.6146
R73 VPWR.n8 VPWR.t0 28.1434
R74 VPWR.n2 VPWR.t5 27.2639
R75 VPWR.n3 VPWR.t4 27.2639
R76 VPWR.n11 VPWR.n10 24.0946
R77 VPWR.n10 VPWR.n9 22.9652
R78 VPWR.n10 VPWR.n0 9.3005
R79 VPWR.n11 VPWR.n5 8.92444
R80 VPWR.n9 VPWR.n7 6.87305
R81 VPWR.n5 VPWR.n1 6.13008
R82 VPWR.n12 VPWR.n11 4.1063
R83 VPWR VPWR.n12 0.714876
R84 VPWR.n7 VPWR.n0 0.410331
R85 VPWR.n12 VPWR.n0 0.207182
R86 a_27_74.n0 a_27_74.t0 306.938
R87 a_27_74.n0 a_27_74.t3 226.978
R88 a_27_74.n1 a_27_74.n0 84.8201
R89 a_27_74.t1 a_27_74.n1 22.7032
R90 a_27_74.n1 a_27_74.t2 22.7032
R91 VNB.t0 VNB.t7 2448.29
R92 VNB.t8 VNB.t2 2286.61
R93 VNB.t4 VNB.t8 1258.79
R94 VNB VNB.t6 1143.31
R95 VNB.t6 VNB.t5 1108.66
R96 VNB.t9 VNB.t4 1050.92
R97 VNB.t2 VNB.t3 993.177
R98 VNB.t7 VNB.t9 993.177
R99 VNB.t1 VNB.t0 993.177
R100 VNB.t5 VNB.t1 993.177
R101 A1.n2 A1.t3 276.955
R102 A1.n0 A1.t1 264.541
R103 A1 A1.n2 158.788
R104 A1.n1 A1.t2 154.24
R105 A1.n0 A1.t0 154.24
R106 A1.n1 A1.n0 62.8066
R107 A1.n2 A1.n1 41.6278
R108 a_507_74.n0 a_507_74.t1 313.051
R109 a_507_74.n0 a_507_74.t3 271.144
R110 a_507_74.n1 a_507_74.n0 103.456
R111 a_507_74.n1 a_507_74.t0 26.7573
R112 a_507_74.t2 a_507_74.n1 22.7032
R113 a_771_74.n1 a_771_74.n0 389.914
R114 a_771_74.n0 a_771_74.t3 34.0546
R115 a_771_74.n0 a_771_74.t2 30.0005
R116 a_771_74.n1 a_771_74.t1 22.7032
R117 a_771_74.t0 a_771_74.n1 22.7032
R118 VGND.n5 VGND.t0 242.263
R119 VGND.n19 VGND.n18 209.243
R120 VGND.n4 VGND.t1 145.002
R121 VGND.n6 VGND.n3 36.1417
R122 VGND.n10 VGND.n3 36.1417
R123 VGND.n11 VGND.n10 36.1417
R124 VGND.n12 VGND.n11 36.1417
R125 VGND.n12 VGND.n1 36.1417
R126 VGND.n16 VGND.n1 36.1417
R127 VGND.n17 VGND.n16 36.1417
R128 VGND.n18 VGND.t2 30.8113
R129 VGND.n6 VGND.n5 28.2358
R130 VGND.n19 VGND.n17 24.4711
R131 VGND.n18 VGND.t3 22.7032
R132 VGND.n17 VGND.n0 9.3005
R133 VGND.n16 VGND.n15 9.3005
R134 VGND.n14 VGND.n1 9.3005
R135 VGND.n13 VGND.n12 9.3005
R136 VGND.n11 VGND.n2 9.3005
R137 VGND.n10 VGND.n9 9.3005
R138 VGND.n8 VGND.n3 9.3005
R139 VGND.n7 VGND.n6 9.3005
R140 VGND.n20 VGND.n19 7.19894
R141 VGND.n5 VGND.n4 6.70714
R142 VGND.n7 VGND.n4 0.645862
R143 VGND VGND.n20 0.156997
R144 VGND.n20 VGND.n0 0.150766
R145 VGND.n8 VGND.n7 0.122949
R146 VGND.n9 VGND.n8 0.122949
R147 VGND.n9 VGND.n2 0.122949
R148 VGND.n13 VGND.n2 0.122949
R149 VGND.n14 VGND.n13 0.122949
R150 VGND.n15 VGND.n14 0.122949
R151 VGND.n15 VGND.n0 0.122949
R152 B2.n1 B2.t2 244.579
R153 B2.n0 B2.t0 240.197
R154 B2.n0 B2.t1 182.138
R155 B2.n1 B2.t3 179.947
R156 B2.n3 B2.n2 81.8268
R157 B2.n2 B2.n0 31.5319
R158 B2.n2 B2.n1 29.6657
R159 B2 B2.n3 7.25383
R160 B2.n3 B2 3.29747
R161 A2.n0 A2.t1 226.809
R162 A2.n2 A2.t0 226.809
R163 A2.n2 A2.t3 198.204
R164 A2.n0 A2.t2 198.204
R165 A2 A2.n1 158.4
R166 A2.n4 A2.n3 152
R167 A2.n3 A2.n1 49.6611
R168 A2.n1 A2.n0 14.6066
R169 A2.n3 A2.n2 10.955
R170 A2.n4 A2 10.5679
R171 A2 A2.n4 3.72143
C0 VPB B1 0.066948f
C1 A3 VGND 0.07163f
C2 Y VPWR 0.030992f
C3 VPB A1 0.080883f
C4 B2 B1 0.066913f
C5 Y VGND 0.030073f
C6 B2 A1 1.69e-19
C7 VPB A2 0.069568f
C8 VPWR VGND 0.099811f
C9 B1 A1 0.078528f
C10 VPB A3 0.096981f
C11 VPB Y 0.014736f
C12 A1 A2 0.063064f
C13 B2 Y 0.073536f
C14 VPB VPWR 0.152364f
C15 VPB VGND 0.009646f
C16 A1 A3 9.04e-20
C17 B1 Y 0.192251f
C18 B2 VPWR 0.012712f
C19 A1 Y 0.146946f
C20 A2 A3 0.039161f
C21 B2 VGND 0.035533f
C22 B1 VPWR 0.012251f
C23 B1 VGND 0.014162f
C24 A1 VPWR 0.040262f
C25 A2 Y 0.030151f
C26 A3 Y 0.002125f
C27 A1 VGND 0.014049f
C28 A2 VPWR 0.04157f
C29 VPB B2 0.070357f
C30 A2 VGND 0.013939f
C31 A3 VPWR 0.043667f
C32 VGND VNB 0.765625f
C33 VPWR VNB 0.577412f
C34 Y VNB 0.031385f
C35 A3 VNB 0.314553f
C36 A2 VNB 0.214908f
C37 A1 VNB 0.239257f
C38 B1 VNB 0.225345f
C39 B2 VNB 0.252675f
C40 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a32oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32oi_1 VNB VPB VPWR VGND A3 B2 B1 A2 Y A1
X0 a_27_368.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3584 ps=1.76 w=1.12 l=0.15
X1 a_391_74.t1 A1.t0 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.3034 ps=1.56 w=0.74 l=0.15
X2 Y.t1 B2.t0 a_27_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X3 a_119_74.t0 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2294 ps=2.1 w=0.74 l=0.15
X4 VPWR.t2 A1.t1 a_27_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3584 pd=1.76 as=0.2576 ps=1.58 w=1.12 l=0.15
X5 VGND.t1 A3.t0 a_469_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X6 Y.t0 B1.t0 a_119_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3034 pd=1.56 as=0.0888 ps=0.98 w=0.74 l=0.15
X7 a_27_368.t4 B1.t1 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2576 pd=1.58 as=0.196 ps=1.47 w=1.12 l=0.15
X8 a_469_74.t1 A2.t1 a_391_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X9 VPWR.t1 A3.t1 a_27_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A2.n0 A2.t0 285.719
R1 A2.n0 A2.t1 178.34
R2 A2 A2.n0 156.667
R3 VPWR.n4 VPWR.n3 585
R4 VPWR.n6 VPWR.n5 585
R5 VPWR.n2 VPWR.t1 264.714
R6 VPWR.n5 VPWR.n4 59.8041
R7 VPWR.n3 VPWR.n2 30.4793
R8 VPWR.n4 VPWR.t0 26.3844
R9 VPWR.n5 VPWR.t2 26.3844
R10 VPWR.n7 VPWR.n6 10.3542
R11 VPWR.n1 VPWR.n0 9.3005
R12 VPWR.n6 VPWR.n1 5.42567
R13 VPWR.n2 VPWR.n0 2.0514
R14 VPWR VPWR.n7 0.404497
R15 VPWR.n3 VPWR.n1 0.339573
R16 VPWR.n7 VPWR.n0 0.149448
R17 a_27_368.n1 a_27_368.t2 301.925
R18 a_27_368.n1 a_27_368.n0 290.389
R19 a_27_368.n2 a_27_368.n1 283.553
R20 a_27_368.n0 a_27_368.t3 45.7326
R21 a_27_368.n0 a_27_368.t4 35.1791
R22 a_27_368.n2 a_27_368.t1 26.3844
R23 a_27_368.t0 a_27_368.n2 26.3844
R24 VPB.t3 VPB.t0 403.495
R25 VPB.t4 VPB.t3 311.56
R26 VPB VPB.t2 257.93
R27 VPB.t2 VPB.t4 255.376
R28 VPB.t0 VPB.t1 229.839
R29 A1.n0 A1.t1 280.115
R30 A1.n0 A1.t0 172.736
R31 A1 A1.n0 158.788
R32 Y.n2 Y.n0 305.048
R33 Y.n2 Y.n1 98.6516
R34 Y Y.n2 63.0024
R35 Y.n1 Y.t2 54.5616
R36 Y.n1 Y.t0 51.3215
R37 Y.n0 Y.t1 35.1791
R38 Y.n0 Y.t3 26.3844
R39 a_391_74.t0 a_391_74.t1 38.9194
R40 VNB.t2 VNB.t4 2240.42
R41 VNB.t3 VNB.t1 1316.54
R42 VNB VNB.t0 1201.05
R43 VNB.t4 VNB.t3 900.788
R44 VNB.t0 VNB.t2 900.788
R45 B2.n0 B2.t0 278.188
R46 B2.n0 B2.t1 170.81
R47 B2 B2.n0 158.788
R48 VGND.n0 VGND.t1 163.578
R49 VGND.n0 VGND.t0 149.754
R50 VGND VGND.n0 0.0994077
R51 a_119_74.t0 a_119_74.t1 38.9194
R52 A3.n0 A3.t1 285.719
R53 A3.n0 A3.t0 178.34
R54 A3 A3.n0 156.767
R55 a_469_74.t0 a_469_74.t1 68.1086
R56 B1.n0 B1.t1 279.293
R57 B1.n0 B1.t0 171.913
R58 B1 B1.n0 158.222
C0 A3 VGND 0.053373f
C1 Y VPWR 0.03022f
C2 B2 B1 0.058121f
C3 Y VGND 0.189267f
C4 VPWR VGND 0.055263f
C5 B1 A1 0.069314f
C6 VPB B2 0.039968f
C7 B1 A2 2.85e-19
C8 VPB B1 0.036444f
C9 A1 A2 0.086827f
C10 B2 Y 0.055459f
C11 VPB A1 0.038899f
C12 B1 Y 0.141936f
C13 B2 VPWR 0.006785f
C14 VPB A2 0.033058f
C15 B2 VGND 0.053897f
C16 B1 VPWR 0.006044f
C17 A2 A3 0.084593f
C18 A1 Y 0.082487f
C19 VPB A3 0.033654f
C20 B1 VGND 0.007474f
C21 A2 Y 0.071099f
C22 A1 VPWR 0.013851f
C23 VPB Y 0.012291f
C24 A1 VGND 0.012344f
C25 A2 VPWR 0.017478f
C26 A3 Y 7.38e-19
C27 VPB VPWR 0.093822f
C28 A3 VPWR 0.039212f
C29 A2 VGND 0.077508f
C30 VPB VGND 0.00623f
C31 VGND VNB 0.496703f
C32 VPWR VNB 0.38216f
C33 Y VNB 0.04121f
C34 A3 VNB 0.154826f
C35 A2 VNB 0.11749f
C36 A1 VNB 0.120095f
C37 B1 VNB 0.121329f
C38 B2 VNB 0.16526f
C39 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a32o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32o_4 VNB VPB VPWR VGND B1 A3 A1 X B2 A2
X0 X.t3 a_83_283.t7 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 VPWR.t0 A2.t0 a_509_392.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2325 pd=1.465 as=0.2725 ps=1.545 w=1 l=0.15
X2 VGND.t6 a_83_283.t8 X.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2557 pd=1.5 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_83_283.t2 B2.t0 a_509_392.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X4 a_509_392.t1 A3.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.175 ps=1.35 w=1 l=0.15
X5 a_509_392.t6 B2.t1 a_83_283.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2725 pd=1.545 as=0.175 ps=1.35 w=1 l=0.15
X6 a_1079_122.t1 A2.t1 a_992_122.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X7 VPWR.t7 a_83_283.t9 X.t2 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t1 a_83_283.t10 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X9 X.t6 a_83_283.t11 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.10915 pd=1.035 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 X.t5 a_83_283.t12 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1591 ps=1.17 w=0.74 l=0.15
X11 a_992_122.t0 A3.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.12 ps=1.015 w=0.64 l=0.15
X12 VPWR.t4 A1.t0 a_509_392.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.18 pd=1.36 as=0.16 ps=1.32 w=1 l=0.15
X13 VPWR.t2 A3.t2 a_509_392.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X14 a_587_110.t3 B1.t0 a_83_283.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.127875 ps=1.145 w=0.64 l=0.15
X15 a_509_392.t2 A2.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.18 ps=1.36 w=1 l=0.15
X16 a_83_283.t6 A1.t1 a_1079_122.t2 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X17 a_83_283.t1 B1.t1 a_509_392.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X18 VPWR.t5 a_83_283.t13 X.t0 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VGND.t3 a_83_283.t14 X.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1591 pd=1.17 as=0.10915 ps=1.035 w=0.74 l=0.15
X20 a_587_110.t1 B2.t2 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2557 ps=1.5 w=0.64 l=0.15
X21 VGND.t2 B2.t3 a_587_110.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.192025 pd=1.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X22 a_509_392.t9 A1.t2 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.32 as=0.2325 ps=1.465 w=1 l=0.15
X23 a_509_392.t8 B1.t2 a_83_283.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X24 a_992_122.t1 A2.t3 a_1079_122.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.096 pd=0.94 as=0.1152 ps=1 w=0.64 l=0.15
X25 a_83_283.t0 B1.t3 a_587_110.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.127875 pd=1.145 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 a_83_283.n1 a_83_283.t6 401.767
R1 a_83_283.n16 a_83_283.n15 313.74
R2 a_83_283.n14 a_83_283.n13 300.281
R3 a_83_283.n3 a_83_283.t9 226.809
R4 a_83_283.n8 a_83_283.t10 226.809
R5 a_83_283.n6 a_83_283.t13 225.709
R6 a_83_283.n1 a_83_283.n0 213.359
R7 a_83_283.n4 a_83_283.t7 204.048
R8 a_83_283.n3 a_83_283.t8 177.555
R9 a_83_283.n10 a_83_283.t12 170.308
R10 a_83_283.n7 a_83_283.n2 165.189
R11 a_83_283.n9 a_83_283.n2 152
R12 a_83_283.n12 a_83_283.n11 152
R13 a_83_283.n4 a_83_283.t11 144.155
R14 a_83_283.n5 a_83_283.t14 142.994
R15 a_83_283.n14 a_83_283.n12 100.45
R16 a_83_283.n5 a_83_283.n4 50.5234
R17 a_83_283.n15 a_83_283.n1 50.4476
R18 a_83_283.n15 a_83_283.n14 46.3064
R19 a_83_283.n11 a_83_283.n10 45.2793
R20 a_83_283.n0 a_83_283.t0 44.9092
R21 a_83_283.n8 a_83_283.n7 44.549
R22 a_83_283.n13 a_83_283.t2 39.4005
R23 a_83_283.t1 a_83_283.n16 39.4005
R24 a_83_283.n13 a_83_283.t4 29.5505
R25 a_83_283.n16 a_83_283.t3 29.5505
R26 a_83_283.n7 a_83_283.n6 25.4879
R27 a_83_283.n0 a_83_283.t5 22.9787
R28 a_83_283.n12 a_83_283.n2 13.1884
R29 a_83_283.n11 a_83_283.n3 10.955
R30 a_83_283.n9 a_83_283.n8 5.11262
R31 a_83_283.n10 a_83_283.n9 4.38232
R32 a_83_283.n6 a_83_283.n5 1.59292
R33 VPWR.n10 VPWR.n9 604.023
R34 VPWR.n15 VPWR.n8 603.173
R35 VPWR.n3 VPWR.t7 342.784
R36 VPWR.n12 VPWR.n11 325.146
R37 VPWR.n28 VPWR.n2 317.435
R38 VPWR.n30 VPWR.t8 259.171
R39 VPWR.n8 VPWR.t9 51.2205
R40 VPWR.n8 VPWR.t0 40.3855
R41 VPWR.n11 VPWR.t3 39.4005
R42 VPWR.n9 VPWR.t4 38.4155
R43 VPWR.n17 VPWR.n16 36.1417
R44 VPWR.n17 VPWR.n5 36.1417
R45 VPWR.n21 VPWR.n5 36.1417
R46 VPWR.n22 VPWR.n21 36.1417
R47 VPWR.n23 VPWR.n22 36.1417
R48 VPWR.n2 VPWR.t6 35.1791
R49 VPWR.n9 VPWR.t1 32.5055
R50 VPWR.n11 VPWR.t2 29.5505
R51 VPWR.n15 VPWR.n14 28.9887
R52 VPWR.n30 VPWR.n29 26.7299
R53 VPWR.n2 VPWR.t5 26.3844
R54 VPWR.n23 VPWR.n3 25.977
R55 VPWR.n28 VPWR.n27 25.224
R56 VPWR.n29 VPWR.n28 22.2123
R57 VPWR.n27 VPWR.n3 21.4593
R58 VPWR.n14 VPWR.n10 21.4593
R59 VPWR.n16 VPWR.n15 12.8005
R60 VPWR.n14 VPWR.n13 9.3005
R61 VPWR.n15 VPWR.n7 9.3005
R62 VPWR.n16 VPWR.n6 9.3005
R63 VPWR.n18 VPWR.n17 9.3005
R64 VPWR.n19 VPWR.n5 9.3005
R65 VPWR.n21 VPWR.n20 9.3005
R66 VPWR.n22 VPWR.n4 9.3005
R67 VPWR.n24 VPWR.n23 9.3005
R68 VPWR.n25 VPWR.n3 9.3005
R69 VPWR.n27 VPWR.n26 9.3005
R70 VPWR.n28 VPWR.n1 9.3005
R71 VPWR.n29 VPWR.n0 9.3005
R72 VPWR.n31 VPWR.n30 9.3005
R73 VPWR.n12 VPWR.n10 6.71627
R74 VPWR.n13 VPWR.n12 0.560449
R75 VPWR.n13 VPWR.n7 0.122949
R76 VPWR.n7 VPWR.n6 0.122949
R77 VPWR.n18 VPWR.n6 0.122949
R78 VPWR.n19 VPWR.n18 0.122949
R79 VPWR.n20 VPWR.n19 0.122949
R80 VPWR.n20 VPWR.n4 0.122949
R81 VPWR.n24 VPWR.n4 0.122949
R82 VPWR.n25 VPWR.n24 0.122949
R83 VPWR.n26 VPWR.n25 0.122949
R84 VPWR.n26 VPWR.n1 0.122949
R85 VPWR.n1 VPWR.n0 0.122949
R86 VPWR.n31 VPWR.n0 0.122949
R87 VPWR VPWR.n31 0.0617245
R88 X.n2 X.n0 261.183
R89 X.n2 X.n1 208.98
R90 X.n5 X.n4 141.73
R91 X.n5 X.n3 97.7287
R92 X X.n2 54.5128
R93 X.n1 X.t0 26.3844
R94 X.n1 X.t3 26.3844
R95 X.n0 X.t2 26.3844
R96 X.n0 X.t1 26.3844
R97 X X.n5 25.9901
R98 X.n3 X.t4 24.3248
R99 X.n3 X.t6 23.514
R100 X.n4 X.t7 22.7032
R101 X.n4 X.t5 22.7032
R102 VPB.n0 VPB 2500.13
R103 VPB VPB.n1 1692.53
R104 VPB.t5 VPB.t11 515.861
R105 VPB.t0 VPB.t13 314.113
R106 VPB.t4 VPB.t6 272.988
R107 VPB.t8 VPB.t4 272.988
R108 VPB.t6 VPB.n0 262.07
R109 VPB.t7 VPB.t1 260.485
R110 VPB.t12 VPB 257.93
R111 VPB.t2 VPB.t3 255.376
R112 VPB.t10 VPB.t9 255.376
R113 VPB.t13 VPB.t7 240.054
R114 VPB.t1 VPB.t2 229.839
R115 VPB.t11 VPB.t10 229.839
R116 VPB.t9 VPB.t12 229.839
R117 VPB.n1 VPB.t8 171.983
R118 VPB.n0 VPB.t0 109.812
R119 VPB.n1 VPB.t5 94.4898
R120 A2.n2 A2.n0 279.822
R121 A2.n0 A2.t2 239.661
R122 A2.n1 A2.t0 228.737
R123 A2.n1 A2.t1 194.728
R124 A2.n0 A2.t3 187.981
R125 A2.n2 A2.n1 152
R126 A2 A2.n2 9.2005
R127 a_509_392.n1 a_509_392.t5 383.207
R128 a_509_392.n1 a_509_392.n0 303.212
R129 a_509_392.n5 a_509_392.n4 296.705
R130 a_509_392.n3 a_509_392.t1 291
R131 a_509_392.n3 a_509_392.n2 195.901
R132 a_509_392.n7 a_509_392.n6 192.501
R133 a_509_392.n6 a_509_392.n1 72.8863
R134 a_509_392.n6 a_509_392.n5 71.1553
R135 a_509_392.t3 a_509_392.n7 54.1755
R136 a_509_392.n7 a_509_392.t6 53.1905
R137 a_509_392.n5 a_509_392.n3 52.709
R138 a_509_392.n0 a_509_392.t8 39.4005
R139 a_509_392.n4 a_509_392.t7 33.4905
R140 a_509_392.n0 a_509_392.t4 29.5505
R141 a_509_392.n2 a_509_392.t0 29.5505
R142 a_509_392.n2 a_509_392.t2 29.5505
R143 a_509_392.n4 a_509_392.t9 29.5505
R144 VGND.n7 VGND.t2 303.053
R145 VGND.n22 VGND.t5 302.817
R146 VGND.n6 VGND.t0 260.68
R147 VGND.n20 VGND.n2 203.577
R148 VGND.n16 VGND.n15 122.316
R149 VGND.n15 VGND.t1 103.126
R150 VGND.n2 VGND.t4 40.541
R151 VGND.n9 VGND.n8 36.1417
R152 VGND.n9 VGND.n4 36.1417
R153 VGND.n13 VGND.n4 36.1417
R154 VGND.n14 VGND.n13 36.1417
R155 VGND.n15 VGND.t6 35.7861
R156 VGND.n7 VGND.n6 35.5073
R157 VGND.n16 VGND.n1 29.3652
R158 VGND.n2 VGND.t3 29.1897
R159 VGND.n20 VGND.n1 21.0829
R160 VGND.n22 VGND.n21 20.7064
R161 VGND.n21 VGND.n20 20.3299
R162 VGND.n16 VGND.n14 18.0711
R163 VGND.n23 VGND.n22 9.3005
R164 VGND.n21 VGND.n0 9.3005
R165 VGND.n20 VGND.n19 9.3005
R166 VGND.n18 VGND.n1 9.3005
R167 VGND.n17 VGND.n16 9.3005
R168 VGND.n8 VGND.n5 9.3005
R169 VGND.n10 VGND.n9 9.3005
R170 VGND.n11 VGND.n4 9.3005
R171 VGND.n13 VGND.n12 9.3005
R172 VGND.n14 VGND.n3 9.3005
R173 VGND.n8 VGND.n7 8.28285
R174 VGND.n6 VGND.n5 0.151403
R175 VGND.n10 VGND.n5 0.122949
R176 VGND.n11 VGND.n10 0.122949
R177 VGND.n12 VGND.n11 0.122949
R178 VGND.n12 VGND.n3 0.122949
R179 VGND.n17 VGND.n3 0.122949
R180 VGND.n18 VGND.n17 0.122949
R181 VGND.n19 VGND.n18 0.122949
R182 VGND.n19 VGND.n0 0.122949
R183 VGND.n23 VGND.n0 0.122949
R184 VGND VGND.n23 0.0617245
R185 VNB.t5 VNB.t3 2517.59
R186 VNB.t2 VNB.t1 2251.97
R187 VNB.t11 VNB.t2 2171.13
R188 VNB.t9 VNB.t4 2101.84
R189 VNB.t6 VNB.t7 1339.63
R190 VNB.t0 VNB.t10 1177.95
R191 VNB VNB.t8 1143.31
R192 VNB.t8 VNB.t6 1027.82
R193 VNB.t3 VNB.t11 993.177
R194 VNB.t4 VNB.t0 993.177
R195 VNB.t7 VNB.t9 993.177
R196 VNB.t10 VNB.t5 993.177
R197 B2.n1 B2.t1 768.223
R198 B2 B2.n1 348.289
R199 B2.n0 B2.t0 228.79
R200 B2.n0 B2.t2 202.28
R201 B2 B2.n0 153.358
R202 B2.n1 B2.t3 141.095
R203 A3.n0 A3.t0 212.883
R204 A3.n2 A3.t2 212.883
R205 A3.n2 A3.n1 169.285
R206 A3.n0 A3.t1 168.554
R207 A3.n3 A3 156.849
R208 A3.n5 A3.n4 152
R209 A3.n4 A3.n3 61.346
R210 A3.n5 A3 11.4429
R211 A3.n3 A3.n2 10.955
R212 A3 A3.n5 7.17626
R213 A3.n4 A3.n0 0.730803
R214 a_992_122.n0 a_992_122.t2 422.844
R215 a_992_122.t0 a_992_122.n0 203.095
R216 a_992_122.n0 a_992_122.t1 123.174
R217 a_1079_122.n0 a_1079_122.t0 382.168
R218 a_1079_122.n0 a_1079_122.t2 26.2505
R219 a_1079_122.t1 a_1079_122.n0 26.2505
R220 A1.n2 A1.t2 216.536
R221 A1.n1 A1.t0 215.075
R222 A1.n2 A1.t1 167.094
R223 A1.n1 A1.n0 167.094
R224 A1 A1.n3 156.462
R225 A1.n3 A1.n1 55.5035
R226 A1.n3 A1.n2 7.30353
R227 B1.n1 B1.t3 210.975
R228 B1.n0 B1.t1 205.109
R229 B1.n1 B1.t2 192.8
R230 B1.n3 B1.n2 152
R231 B1.n0 B1.t0 139.78
R232 B1.n2 B1.n0 36.8943
R233 B1.n3 B1 17.649
R234 B1.n2 B1.n1 8.92643
R235 B1 B1.n3 0.970197
R236 a_587_110.n1 a_587_110.n0 339.147
R237 a_587_110.n0 a_587_110.t0 26.2505
R238 a_587_110.n0 a_587_110.t3 26.2505
R239 a_587_110.n1 a_587_110.t2 26.2505
R240 a_587_110.t1 a_587_110.n1 26.2505
C0 B2 X 0.003268f
C1 A2 A3 0.080085f
C2 B1 VPWR 0.012137f
C3 VPB VGND 0.014089f
C4 A2 VPWR 0.046284f
C5 B2 VGND 0.366728f
C6 B1 X 1.11e-19
C7 B1 VGND 0.011325f
C8 A1 VPWR 0.03043f
C9 A2 VGND 0.014061f
C10 A3 VPWR 0.03802f
C11 VPB B2 0.105543f
C12 A1 VGND 0.009434f
C13 VPB B1 0.068551f
C14 VPWR X 0.412897f
C15 A3 VGND 0.027351f
C16 B2 B1 0.142722f
C17 VPB A2 0.100675f
C18 VPWR VGND 0.132409f
C19 B2 A2 0.064179f
C20 VPB A1 0.076181f
C21 X VGND 0.303044f
C22 B1 A2 5.32e-19
C23 B2 A1 6.35e-20
C24 VPB A3 0.088075f
C25 VPB VPWR 0.221326f
C26 A2 A1 0.210104f
C27 VPB X 0.012906f
C28 B2 VPWR 0.015503f
C29 VGND VNB 0.993176f
C30 X VNB 0.058193f
C31 VPWR VNB 0.779373f
C32 A3 VNB 0.231344f
C33 A1 VNB 0.174858f
C34 A2 VNB 0.205387f
C35 B1 VNB 0.212635f
C36 B2 VNB 0.46567f
C37 VPB VNB 1.88028f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a32o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32o_2 VNB VPB VPWR VGND B2 B1 A3 A2 A1 X
X0 X.t3 a_45_264.t4 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 a_355_74.t1 A3.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2035 ps=1.29 w=0.74 l=0.15
X2 X.t1 a_45_264.t5 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1073 pd=1.03 as=0.259 ps=2.18 w=0.74 l=0.15
X3 a_45_264.t3 A1.t0 a_433_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X4 VGND.t0 B2.t0 a_661_74.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 a_45_264.t0 B1.t0 a_346_368.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X6 VPWR.t0 A2.t0 a_346_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.28 pd=1.56 as=0.15 ps=1.3 w=1 l=0.15
X7 a_346_368.t2 A3.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.3026 ps=1.67 w=1 l=0.15
X8 a_346_368.t1 A1.t1 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.28 ps=1.56 w=1 l=0.15
X9 a_433_74.t1 A2.t1 a_355_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X10 VPWR.t2 a_45_264.t6 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.3026 pd=1.67 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_661_74.t0 B1.t1 a_45_264.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1554 ps=1.16 w=0.74 l=0.15
X12 VGND.t2 a_45_264.t7 X.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2035 pd=1.29 as=0.1073 ps=1.03 w=0.74 l=0.15
X13 a_346_368.t4 B2.t1 a_45_264.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2 ps=1.4 w=1 l=0.15
R0 a_45_264.n5 a_45_264.n4 463.373
R1 a_45_264.n4 a_45_264.n2 306.962
R2 a_45_264.n4 a_45_264.n3 279.029
R3 a_45_264.n0 a_45_264.t6 234.841
R4 a_45_264.n2 a_45_264.t4 234.841
R5 a_45_264.n0 a_45_264.t7 193.963
R6 a_45_264.n1 a_45_264.t5 186.374
R7 a_45_264.n1 a_45_264.n0 57.6944
R8 a_45_264.n5 a_45_264.t1 39.4005
R9 a_45_264.t0 a_45_264.n5 39.4005
R10 a_45_264.n3 a_45_264.t2 34.8654
R11 a_45_264.n3 a_45_264.t3 33.2437
R12 a_45_264.n2 a_45_264.n1 8.03383
R13 VPWR.n6 VPWR.t3 860.096
R14 VPWR.n2 VPWR.n1 610.923
R15 VPWR.n4 VPWR.n3 600.766
R16 VPWR.n1 VPWR.t4 55.1605
R17 VPWR.n1 VPWR.t0 55.1605
R18 VPWR.n3 VPWR.t1 54.1755
R19 VPWR.n3 VPWR.t2 45.3924
R20 VPWR.n5 VPWR.n4 28.6123
R21 VPWR.n6 VPWR.n5 20.7064
R22 VPWR.n5 VPWR.n0 9.3005
R23 VPWR.n7 VPWR.n6 9.3005
R24 VPWR.n4 VPWR.n2 6.19401
R25 VPWR.n2 VPWR.n0 0.332068
R26 VPWR.n7 VPWR.n0 0.122949
R27 VPWR VPWR.n7 0.0617245
R28 X.n2 X.n1 585
R29 X.n2 X.n0 148.471
R30 X.n1 X.t2 26.3844
R31 X.n1 X.t3 26.3844
R32 X.n0 X.t0 23.514
R33 X.n0 X.t1 23.514
R34 X X.n2 3.68535
R35 VPB.t1 VPB.t6 362.635
R36 VPB.t4 VPB.t2 357.527
R37 VPB.t0 VPB.t3 280.914
R38 VPB VPB.t5 257.93
R39 VPB.t6 VPB.t0 229.839
R40 VPB.t2 VPB.t1 229.839
R41 VPB.t5 VPB.t4 229.839
R42 A3.n0 A3.t1 231.629
R43 A3.n0 A3.t0 220.113
R44 A3 A3.n0 154.522
R45 VGND.n3 VGND.n2 211.183
R46 VGND.n1 VGND.t0 171.583
R47 VGND.n5 VGND.t3 155.272
R48 VGND.n2 VGND.t1 44.5951
R49 VGND.n2 VGND.t2 44.5951
R50 VGND.n4 VGND.n3 35.0123
R51 VGND.n5 VGND.n4 20.7064
R52 VGND.n6 VGND.n5 9.3005
R53 VGND.n4 VGND.n0 9.3005
R54 VGND.n3 VGND.n1 6.32375
R55 VGND.n1 VGND.n0 0.171064
R56 VGND.n6 VGND.n0 0.122949
R57 VGND VGND.n6 0.0617245
R58 a_355_74.t0 a_355_74.t1 38.9194
R59 VNB.t3 VNB.t2 1616.8
R60 VNB.t5 VNB.t0 1316.54
R61 VNB.t6 VNB.t5 1316.54
R62 VNB.t1 VNB.t6 1316.54
R63 VNB VNB.t4 1293.44
R64 VNB.t4 VNB.t3 1016.27
R65 VNB.t2 VNB.t1 900.788
R66 A1.n0 A1.t1 231.629
R67 A1.n0 A1.t0 220.113
R68 A1 A1.n0 157.805
R69 a_433_74.t0 a_433_74.t1 68.1086
R70 B2.n0 B2.t1 237.148
R71 B2.n0 B2.t0 196.178
R72 B2 B2.n0 156.462
R73 a_661_74.t0 a_661_74.t1 68.1086
R74 B1.n0 B1.t0 231.629
R75 B1.n0 B1.t1 220.113
R76 B1 B1.n0 157.805
R77 a_346_368.n1 a_346_368.t4 482.736
R78 a_346_368.n2 a_346_368.n1 364.776
R79 a_346_368.n1 a_346_368.n0 289.24
R80 a_346_368.n0 a_346_368.t3 29.5505
R81 a_346_368.n0 a_346_368.t1 29.5505
R82 a_346_368.t0 a_346_368.n2 29.5505
R83 a_346_368.n2 a_346_368.t2 29.5505
R84 A2.n0 A2.t0 231.629
R85 A2.n0 A2.t1 220.113
R86 A2 A2.n0 155.126
C0 A3 VGND 0.013299f
C1 A2 B2 3.76e-20
C2 A1 B1 0.081004f
C3 VPB VPWR 0.121497f
C4 A1 B2 7.39e-20
C5 A2 VGND 0.010658f
C6 VPB X 0.002503f
C7 A1 VGND 0.008115f
C8 B1 B2 0.090732f
C9 VPB A3 0.037285f
C10 VPWR X 0.013686f
C11 B1 VGND 0.025125f
C12 VPB A2 0.035344f
C13 VPWR A3 0.011027f
C14 B2 VGND 0.052861f
C15 X A3 5.17e-19
C16 VPWR A2 0.010932f
C17 VPB A1 0.035679f
C18 X A2 2.77e-19
C19 VPB B1 0.034511f
C20 VPWR A1 0.012252f
C21 VPB B2 0.045077f
C22 A3 A2 0.091576f
C23 X A1 1.37e-19
C24 VPWR B1 0.006276f
C25 VPB VGND 0.008097f
C26 VPWR B2 0.006894f
C27 VPWR VGND 0.075239f
C28 A2 A1 0.079931f
C29 X VGND 0.142562f
C30 A3 B2 2.6e-20
C31 VGND VNB 0.616484f
C32 B2 VNB 0.171647f
C33 B1 VNB 0.110276f
C34 A1 VNB 0.106663f
C35 A2 VNB 0.102436f
C36 A3 VNB 0.107603f
C37 X VNB 0.012023f
C38 VPWR VNB 0.435282f
C39 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a221oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221oi_1 VNB VPB VPWR VGND C1 Y B2 B1 A1 A2
X0 VGND.t0 C1.t0 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.4477 ps=2.69 w=0.74 l=0.15
X1 a_351_74.t1 B2.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1443 ps=1.13 w=0.74 l=0.15
X2 a_118_368.t0 C1.t1 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X3 Y.t2 B1.t0 a_351_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=1.31 as=0.0777 ps=0.95 w=0.74 l=0.15
X4 a_567_74.t0 A1.t0 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.2109 ps=1.31 w=0.74 l=0.15
X5 a_263_368.t3 B1.t1 a_118_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t1 A1.t1 a_263_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1848 ps=1.45 w=1.12 l=0.15
X7 VGND.t2 A2.t0 a_567_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.0777 ps=0.95 w=0.74 l=0.15
X8 a_118_368.t2 B2.t1 a_263_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X9 a_263_368.t1 A2.t1 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.2184 ps=1.51 w=1.12 l=0.15
R0 C1.n0 C1.t0 261.317
R1 C1.n0 C1.t1 255.291
R2 C1 C1.n0 154.233
R3 Y.n7 Y 591.4
R4 Y.n7 Y.n0 585
R5 Y.n8 Y.n7 585
R6 Y.n5 Y.n4 185
R7 Y.n4 Y.n3 185
R8 Y.n3 Y.n2 182.633
R9 Y.t1 Y.n1 135.837
R10 Y.n2 Y.t3 50.2708
R11 Y.n4 Y.t1 44.6286
R12 Y.n2 Y.t2 42.1627
R13 Y.n7 Y.t0 26.3844
R14 Y Y.n8 17.1525
R15 Y Y.n0 14.8485
R16 Y.n6 Y.n5 5.16677
R17 Y Y.n0 4.0965
R18 Y.n3 Y.n1 2.58605
R19 Y.n5 Y.n1 2.58605
R20 Y.n8 Y 1.7925
R21 Y Y.n6 1.5365
R22 Y.n6 Y 1.46556
R23 VGND.n1 VGND.n0 214.185
R24 VGND.n1 VGND.t2 166.915
R25 VGND.n0 VGND.t0 37.2978
R26 VGND.n0 VGND.t1 25.9464
R27 VGND VGND.n1 0.386927
R28 VNB VNB.t0 2633.07
R29 VNB.t1 VNB.t3 1662.99
R30 VNB.t0 VNB.t2 1247.24
R31 VNB.t3 VNB.t4 831.496
R32 VNB.t2 VNB.t1 831.496
R33 B2.n0 B2.t1 250.909
R34 B2.n0 B2.t0 220.113
R35 B2.n1 B2.n0 152
R36 B2.n1 B2 14.14
R37 B2 B2.n1 0.149337
R38 a_351_74.t0 a_351_74.t1 34.0546
R39 a_118_368.t0 a_118_368.n0 599.968
R40 a_118_368.n0 a_118_368.t1 26.3844
R41 a_118_368.n0 a_118_368.t2 26.3844
R42 VPB.t0 VPB.t3 587.366
R43 VPB.t2 VPB.t4 275.807
R44 VPB VPB.t0 263.038
R45 VPB.t1 VPB.t2 245.161
R46 VPB.t3 VPB.t1 229.839
R47 B1.n0 B1.t1 250.909
R48 B1.n0 B1.t0 220.113
R49 B1 B1.n0 154.522
R50 A1.n0 A1.t1 250.909
R51 A1.n0 A1.t0 220.113
R52 A1 A1.n0 155.423
R53 a_567_74.t0 a_567_74.t1 34.0546
R54 a_263_368.t0 a_263_368.n1 446.045
R55 a_263_368.n1 a_263_368.t1 281.464
R56 a_263_368.n1 a_263_368.n0 205.998
R57 a_263_368.n0 a_263_368.t2 31.6612
R58 a_263_368.n0 a_263_368.t3 26.3844
R59 VPWR VPWR.n0 321.284
R60 VPWR.n0 VPWR.t0 36.938
R61 VPWR.n0 VPWR.t1 31.6612
R62 A2.n0 A2.t1 285.719
R63 A2.n0 A2.t0 178.34
R64 A2.n1 A2.n0 152
R65 A2.n1 A2 10.5519
R66 A2 A2.n1 6.05455
C0 C1 VPWR 0.013229f
C1 B2 Y 0.072683f
C2 B1 A2 3.7e-19
C3 VPB VGND 0.011411f
C4 A1 A2 0.085956f
C5 C1 VGND 0.015102f
C6 B1 Y 0.045627f
C7 B2 VPWR 0.006769f
C8 B2 VGND 0.016114f
C9 B1 VPWR 0.007299f
C10 A1 Y 0.016267f
C11 B1 VGND 0.013049f
C12 A1 VPWR 0.017608f
C13 A2 Y 0.00494f
C14 VPB C1 0.063683f
C15 A1 VGND 0.020039f
C16 A2 VPWR 0.017615f
C17 VPB B2 0.042941f
C18 A2 VGND 0.05605f
C19 Y VPWR 0.037255f
C20 VPB B1 0.031827f
C21 C1 B2 0.087609f
C22 Y VGND 0.289923f
C23 VPB A1 0.034595f
C24 VPWR VGND 0.060442f
C25 VPB A2 0.040137f
C26 B2 B1 0.105286f
C27 VPB Y 0.018843f
C28 C1 A2 1.19e-19
C29 B1 A1 0.08156f
C30 VPB VPWR 0.100339f
C31 B2 A2 2.2e-19
C32 C1 Y 0.107199f
C33 VGND VNB 0.523742f
C34 VPWR VNB 0.389732f
C35 Y VNB 0.149067f
C36 A2 VNB 0.159945f
C37 A1 VNB 0.110168f
C38 B1 VNB 0.103024f
C39 B2 VNB 0.103008f
C40 C1 VNB 0.178289f
C41 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a221o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221o_4 VNB VPB VPWR X VGND C1 B1 A2 B2 A1
X0 a_157_376.t4 A1.t0 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.275 ps=2.55 w=1 l=0.15
X1 a_71_135.t1 A2.t0 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X2 VGND.t0 a_154_135.t6 X.t7 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.25005 pd=1.48 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 VGND.t7 C1.t0 a_154_135.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.17 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 VGND.t8 B2.t0 a_1346_123.t1 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 a_154_135.t4 A1.t1 a_71_135.t3 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X6 VPWR.t6 A1.t2 a_157_376.t3 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.3725 pd=1.745 as=0.21 ps=1.42 w=1 l=0.15
X7 VPWR.t0 a_154_135.t7 X.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_1102_392.t0 B2.t1 a_157_376.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.295 pd=1.59 as=0.15 ps=1.3 w=1 l=0.15
X9 X.t2 a_154_135.t8 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 X.t6 a_154_135.t9 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12335 ps=1.095 w=0.74 l=0.15
X11 a_157_376.t5 B1.t0 a_1102_392.t2 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.17 pd=1.34 as=0.295 ps=1.59 w=1 l=0.15
X12 VPWR.t2 a_154_135.t10 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_1102_392.t1 C1.t1 a_154_135.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X14 VGND.t6 A2.t1 a_71_135.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.12335 pd=1.095 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 X.t0 a_154_135.t11 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2465 ps=1.58 w=1.12 l=0.15
X16 a_71_135.t2 A1.t3 a_154_135.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X17 a_1346_123.t3 B1.t1 a_154_135.t5 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.2144 pd=1.95 as=0.0896 ps=0.92 w=0.64 l=0.15
X18 VGND.t2 a_154_135.t12 X.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_154_135.t2 B1.t2 a_1346_123.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X20 X.t4 a_154_135.t13 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 VPWR.t4 A2.t2 a_157_376.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2465 pd=1.58 as=0.15 ps=1.3 w=1 l=0.15
X22 a_1346_123.t0 B2.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1648 ps=1.17 w=0.64 l=0.15
X23 a_157_376.t1 A2.t3 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.3725 ps=1.745 w=1 l=0.15
R0 A1.t3 A1.t2 432.462
R1 A1.t1 A1.t0 422.822
R2 A1 A1.n0 278.428
R3 A1.n0 A1.t1 276.348
R4 A1.n0 A1.t3 138.173
R5 A1.n1 A1 20.7064
R6 A1 A1.n1 7.15344
R7 A1.n1 A1 3.68535
R8 VPWR.n5 VPWR.t0 898.125
R9 VPWR.n4 VPWR.n3 605.558
R10 VPWR.n7 VPWR.n6 605.558
R11 VPWR.n14 VPWR.n1 585
R12 VPWR.n16 VPWR.n15 585
R13 VPWR.n22 VPWR.t7 350.329
R14 VPWR.n15 VPWR.n14 66.9805
R15 VPWR.n3 VPWR.t4 61.0705
R16 VPWR.n14 VPWR.t6 40.3855
R17 VPWR.n15 VPWR.t5 39.4005
R18 VPWR.n21 VPWR.n20 36.1417
R19 VPWR.n13 VPWR.n12 36.1417
R20 VPWR.n8 VPWR.n4 32.0005
R21 VPWR.n6 VPWR.t1 26.3844
R22 VPWR.n6 VPWR.t2 26.3844
R23 VPWR.n3 VPWR.t3 25.8649
R24 VPWR.n20 VPWR.n1 17.2743
R25 VPWR.n12 VPWR.n4 15.4358
R26 VPWR.n23 VPWR.n22 15.324
R27 VPWR.n8 VPWR.n7 10.9181
R28 VPWR.n16 VPWR.n13 9.74485
R29 VPWR.n9 VPWR.n8 9.3005
R30 VPWR.n10 VPWR.n4 9.3005
R31 VPWR.n12 VPWR.n11 9.3005
R32 VPWR.n13 VPWR.n2 9.3005
R33 VPWR.n18 VPWR.n17 9.3005
R34 VPWR.n20 VPWR.n19 9.3005
R35 VPWR.n21 VPWR.n0 9.3005
R36 VPWR.n7 VPWR.n5 7.24017
R37 VPWR.n22 VPWR.n21 5.27109
R38 VPWR.n17 VPWR.n16 3.45571
R39 VPWR.n17 VPWR.n1 1.88516
R40 VPWR.n9 VPWR.n5 0.891649
R41 VPWR.n10 VPWR.n9 0.122949
R42 VPWR.n11 VPWR.n10 0.122949
R43 VPWR.n11 VPWR.n2 0.122949
R44 VPWR.n18 VPWR.n2 0.122949
R45 VPWR.n19 VPWR.n18 0.122949
R46 VPWR.n19 VPWR.n0 0.122949
R47 VPWR.n23 VPWR.n0 0.122949
R48 VPWR VPWR.n23 0.0617245
R49 a_157_376.n0 a_157_376.t5 407.452
R50 a_157_376.n3 a_157_376.n2 374.762
R51 a_157_376.n2 a_157_376.n0 328.88
R52 a_157_376.n0 a_157_376.t2 320.067
R53 a_157_376.n2 a_157_376.n1 294.51
R54 a_157_376.t4 a_157_376.n3 53.1905
R55 a_157_376.n1 a_157_376.t0 29.5505
R56 a_157_376.n1 a_157_376.t1 29.5505
R57 a_157_376.n3 a_157_376.t3 29.5505
R58 VPB.t0 VPB.t6 881.048
R59 VPB.t6 VPB.t7 459.678
R60 VPB.t8 VPB.t5 457.125
R61 VPB.t7 VPB.t10 377.957
R62 VPB VPB.t9 362.635
R63 VPB.t4 VPB.t3 311.56
R64 VPB.t9 VPB.t8 291.13
R65 VPB.t1 VPB.t0 229.839
R66 VPB.t2 VPB.t1 229.839
R67 VPB.t3 VPB.t2 229.839
R68 VPB.t5 VPB.t4 229.839
R69 A2.n1 A2.t3 354.538
R70 A2 A2.t0 320.161
R71 A2.n0 A2.t2 291.878
R72 A2.n0 A2.t1 183.161
R73 A2.t0 A2.n1 126.927
R74 A2.n1 A2.n0 24.1005
R75 VGND.n6 VGND.t8 264.361
R76 VGND.n0 VGND.t5 262.966
R77 VGND.n16 VGND.n15 228.294
R78 VGND.n21 VGND.n3 218.792
R79 VGND.n13 VGND.t0 146.32
R80 VGND.n8 VGND.n7 136.667
R81 VGND.n7 VGND.t7 53.2739
R82 VGND.n7 VGND.t4 36.252
R83 VGND.n9 VGND.n5 36.1417
R84 VGND.n17 VGND.n14 36.1417
R85 VGND.n23 VGND.n22 36.1417
R86 VGND.n3 VGND.t6 35.0202
R87 VGND.n25 VGND.n0 33.2507
R88 VGND.n16 VGND.n2 32.0005
R89 VGND.n8 VGND.n6 27.2321
R90 VGND.n22 VGND.n21 27.1064
R91 VGND.n21 VGND.n2 26.3534
R92 VGND.n15 VGND.t3 22.7032
R93 VGND.n15 VGND.t2 22.7032
R94 VGND.n3 VGND.t1 22.1288
R95 VGND.n9 VGND.n8 16.1887
R96 VGND.n14 VGND.n13 12.0476
R97 VGND.n23 VGND.n0 10.5417
R98 VGND.n24 VGND.n23 9.3005
R99 VGND.n22 VGND.n1 9.3005
R100 VGND.n21 VGND.n20 9.3005
R101 VGND.n19 VGND.n2 9.3005
R102 VGND.n18 VGND.n17 9.3005
R103 VGND.n14 VGND.n4 9.3005
R104 VGND.n13 VGND.n12 9.3005
R105 VGND.n11 VGND.n5 9.3005
R106 VGND.n10 VGND.n9 9.3005
R107 VGND.n13 VGND.n5 6.02403
R108 VGND.n17 VGND.n16 4.14168
R109 VGND.n10 VGND.n6 0.497178
R110 VGND VGND.n25 0.404642
R111 VGND.n25 VGND.n24 0.149306
R112 VGND.n11 VGND.n10 0.122949
R113 VGND.n12 VGND.n11 0.122949
R114 VGND.n12 VGND.n4 0.122949
R115 VGND.n18 VGND.n4 0.122949
R116 VGND.n19 VGND.n18 0.122949
R117 VGND.n20 VGND.n19 0.122949
R118 VGND.n20 VGND.n1 0.122949
R119 VGND.n24 VGND.n1 0.122949
R120 a_71_135.n0 a_71_135.t3 330.923
R121 a_71_135.n1 a_71_135.n0 302.353
R122 a_71_135.n0 a_71_135.t2 211.25
R123 a_71_135.n1 a_71_135.t0 26.2505
R124 a_71_135.t1 a_71_135.n1 26.2505
R125 VNB.t10 VNB.t6 3083.46
R126 VNB.t0 VNB.t7 3048.82
R127 VNB.t9 VNB.t8 2263.52
R128 VNB VNB.t11 1605.25
R129 VNB.t7 VNB.t4 1535.96
R130 VNB.t5 VNB.t1 1131.76
R131 VNB.t8 VNB.t12 993.177
R132 VNB.t4 VNB.t9 993.177
R133 VNB.t3 VNB.t0 993.177
R134 VNB.t2 VNB.t3 993.177
R135 VNB.t1 VNB.t2 993.177
R136 VNB.t6 VNB.t5 993.177
R137 VNB.t11 VNB.t10 993.177
R138 a_154_135.n3 a_154_135.t1 834.409
R139 a_154_135.n15 a_154_135.n14 399.416
R140 a_154_135.n3 a_154_135.n2 361.303
R141 a_154_135.n11 a_154_135.t11 253.119
R142 a_154_135.n1 a_154_135.t7 224.131
R143 a_154_135.n8 a_154_135.t8 224.131
R144 a_154_135.n12 a_154_135.t10 224.131
R145 a_154_135.n1 a_154_135.t6 168.237
R146 a_154_135.n11 a_154_135.t9 154.24
R147 a_154_135.n10 a_154_135.t12 154.24
R148 a_154_135.n7 a_154_135.t13 154.24
R149 a_154_135.n14 a_154_135.n13 152
R150 a_154_135.n9 a_154_135.n0 152
R151 a_154_135.n6 a_154_135.n5 152
R152 a_154_135.n4 a_154_135.t0 134.667
R153 a_154_135.n5 a_154_135.n4 88.9134
R154 a_154_135.n12 a_154_135.n11 43.2387
R155 a_154_135.n4 a_154_135.n3 43.2034
R156 a_154_135.n10 a_154_135.n9 41.1123
R157 a_154_135.n7 a_154_135.n6 28.3534
R158 a_154_135.n2 a_154_135.t5 26.2505
R159 a_154_135.n2 a_154_135.t2 26.2505
R160 a_154_135.n15 a_154_135.t3 26.2505
R161 a_154_135.t4 a_154_135.n15 26.2505
R162 a_154_135.n6 a_154_135.n1 20.5564
R163 a_154_135.n8 a_154_135.n7 14.8858
R164 a_154_135.n5 a_154_135.n0 10.8805
R165 a_154_135.n14 a_154_135.n0 10.8805
R166 a_154_135.n13 a_154_135.n12 10.6329
R167 a_154_135.n13 a_154_135.n10 7.08874
R168 a_154_135.n9 a_154_135.n8 4.96226
R169 X.n5 X.n3 627.668
R170 X.n5 X.n4 585
R171 X X.n5 268.014
R172 X.n2 X.n0 141.008
R173 X.n2 X.n1 99.0584
R174 X X.n2 35.1595
R175 X.n4 X.t1 26.3844
R176 X.n4 X.t0 26.3844
R177 X.n3 X.t3 26.3844
R178 X.n3 X.t2 26.3844
R179 X.n0 X.t7 22.7032
R180 X.n0 X.t4 22.7032
R181 X.n1 X.t5 22.7032
R182 X.n1 X.t6 22.7032
R183 C1.n1 C1.t1 363.089
R184 C1.n2 C1.n0 207.529
R185 C1.n4 C1.n3 168.433
R186 C1.n1 C1.t0 163.825
R187 C1.n5 C1.n4 152
R188 C1.n4 C1.n2 38.8283
R189 C1.n2 C1.n1 23.3879
R190 C1.n5 C1 12.2187
R191 C1 C1.n5 2.13383
R192 B2.n3 B2.n2 769.155
R193 B2.n1 B2.n0 309.82
R194 B2.n1 B2.t0 221.72
R195 B2.n2 B2.t1 214.222
R196 B2 B2.n3 164.288
R197 B2.n3 B2.t2 162.274
R198 B2.n2 B2.n1 40.1672
R199 a_1346_123.n1 a_1346_123.n0 277.921
R200 a_1346_123.n0 a_1346_123.t3 205.339
R201 a_1346_123.n0 a_1346_123.t2 127.79
R202 a_1346_123.t1 a_1346_123.n1 26.2505
R203 a_1346_123.n1 a_1346_123.t0 26.2505
R204 a_1102_392.n0 a_1102_392.t1 1171.93
R205 a_1102_392.t0 a_1102_392.n0 60.0855
R206 a_1102_392.n0 a_1102_392.t2 56.1455
R207 B1.n1 B1.t0 248.762
R208 B1.n2 B1.n0 226.585
R209 B1.n1 B1.t2 218.507
R210 B1.n3 B1.t1 192.8
R211 B1.n4 B1.n3 114.766
R212 B1.n2 B1.n1 51.4893
R213 B1.n4 B1 9.48193
R214 B1.n3 B1.n2 6.19307
R215 B1 B1.n4 3.9385
C0 A1 C1 4.88e-20
C1 C1 VPWR 0.01411f
C2 A2 X 0.038252f
C3 A1 VGND 0.123249f
C4 VPWR VGND 0.101998f
C5 A2 C1 9.6e-19
C6 A2 VGND 0.145423f
C7 C1 X 0.007645f
C8 X VGND 0.390388f
C9 C1 VGND 0.027558f
C10 VPB B2 0.095489f
C11 B2 B1 0.05032f
C12 VPB B1 0.144157f
C13 A1 B2 1.73e-19
C14 B2 VPWR 0.011965f
C15 VPB A1 0.077294f
C16 A2 B2 8.88e-19
C17 VPB VPWR 0.270326f
C18 B2 X 4.6e-19
C19 B1 VPWR 0.025583f
C20 VPB A2 0.079653f
C21 VPB X 0.031645f
C22 C1 B2 0.040437f
C23 A1 VPWR 0.0254f
C24 B1 X 1.42e-19
C25 B2 VGND 0.213974f
C26 A1 A2 0.02581f
C27 VPB C1 0.111195f
C28 A1 X 0.04727f
C29 VPB VGND 0.01672f
C30 A2 VPWR 0.018578f
C31 VPWR X 0.193042f
C32 B1 VGND 0.028407f
C33 VGND VNB 1.14909f
C34 X VNB 0.094304f
C35 VPWR VNB 0.890257f
C36 B1 VNB 0.347863f
C37 B2 VNB 0.458593f
C38 C1 VNB 0.224087f
C39 A2 VNB 0.267866f
C40 A1 VNB 0.346999f
C41 VPB VNB 2.22754f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a221o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221o_2 VNB VPB VPWR VGND C1 B2 B1 A2 A1 X
X0 VPWR.t2 A1.t0 a_316_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X1 a_316_392.t2 A2.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.199 ps=1.485 w=1 l=0.15
X2 X.t1 a_89_260.t4 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X3 a_89_260.t2 C1.t0 a_515_392.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X4 a_515_392.t0 B2.t0 a_316_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X5 a_316_392.t3 B1.t0 a_515_392.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X6 X.t3 a_89_260.t5 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X7 a_603_74.t0 B1.t1 a_89_260.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.3034 ps=1.56 w=0.74 l=0.15
X8 a_337_74.t1 A2.t1 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.17575 ps=1.215 w=0.74 l=0.15
X9 VGND.t3 B2.t1 a_603_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X10 a_89_260.t3 C1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X11 VGND.t1 a_89_260.t6 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.17575 pd=1.215 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VPWR.t1 a_89_260.t7 X.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.199 pd=1.485 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_89_260.t1 A1.t1 a_337_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.3034 pd=1.56 as=0.0777 ps=0.95 w=0.74 l=0.15
R0 A1.n0 A1.t1 250.87
R1 A1.n0 A1.t0 235.821
R2 A1 A1.n0 153.319
R3 a_316_392.n1 a_316_392.n0 588.567
R4 a_316_392.n0 a_316_392.t1 29.5505
R5 a_316_392.n0 a_316_392.t2 29.5505
R6 a_316_392.t0 a_316_392.n1 29.5505
R7 a_316_392.n1 a_316_392.t3 29.5505
R8 VPWR.n1 VPWR.t2 351.842
R9 VPWR.n5 VPWR.t0 351.637
R10 VPWR.n3 VPWR.n2 231.049
R11 VPWR.n2 VPWR.t3 42.3555
R12 VPWR.n4 VPWR.n3 30.8711
R13 VPWR.n2 VPWR.t1 27.4811
R14 VPWR.n5 VPWR.n4 24.0946
R15 VPWR.n4 VPWR.n0 9.3005
R16 VPWR.n6 VPWR.n5 9.3005
R17 VPWR.n3 VPWR.n1 6.6864
R18 VPWR.n1 VPWR.n0 0.533915
R19 VPWR.n6 VPWR.n0 0.122949
R20 VPWR VPWR.n6 0.0617245
R21 VPB.t3 VPB.t5 495.43
R22 VPB VPB.t1 275.807
R23 VPB.t2 VPB.t4 263.038
R24 VPB.t0 VPB.t6 229.839
R25 VPB.t5 VPB.t0 229.839
R26 VPB.t4 VPB.t3 229.839
R27 VPB.t1 VPB.t2 229.839
R28 A2.n0 A2.t0 287.861
R29 A2.n0 A2.t1 191.194
R30 A2 A2.n0 156.96
R31 a_89_260.t2 a_89_260.n7 353.603
R32 a_89_260.n1 a_89_260.t4 242.388
R33 a_89_260.n0 a_89_260.t7 240.928
R34 a_89_260.n7 a_89_260.t3 205.619
R35 a_89_260.n1 a_89_260.t5 179.947
R36 a_89_260.n0 a_89_260.t6 179.947
R37 a_89_260.n3 a_89_260.n2 161.689
R38 a_89_260.n4 a_89_260.n3 92.5005
R39 a_89_260.n6 a_89_260.n5 92.5005
R40 a_89_260.n5 a_89_260.n4 87.5681
R41 a_89_260.n2 a_89_260.n1 30.396
R42 a_89_260.n2 a_89_260.n0 25.6895
R43 a_89_260.n5 a_89_260.t0 22.7032
R44 a_89_260.n4 a_89_260.t1 22.7032
R45 a_89_260.n6 a_89_260.n3 8.86204
R46 a_89_260.n7 a_89_260.n6 8.22543
R47 X.n2 X 589.85
R48 X.n2 X.n0 585
R49 X.n3 X.n2 585
R50 X X.n1 190.577
R51 X.n2 X.t0 26.3844
R52 X.n2 X.t1 26.3844
R53 X.n1 X.t2 22.7032
R54 X.n1 X.t3 22.7032
R55 X X.n3 12.9944
R56 X X.n0 11.249
R57 X X.n0 3.10353
R58 X.n3 X 1.35808
R59 C1.n0 C1.t0 308.135
R60 C1.n0 C1.t1 172.736
R61 C1 C1.n0 158.788
R62 a_515_392.n0 a_515_392.t2 1007.65
R63 a_515_392.n0 a_515_392.t1 29.5505
R64 a_515_392.t0 a_515_392.n0 29.5505
R65 B2.n0 B2.t0 298.572
R66 B2.n0 B2.t1 178.34
R67 B2 B2.n0 157.272
R68 B1.n0 B1.t1 242.349
R69 B1.n0 B1.t0 227.085
R70 B1 B1.n0 154.522
R71 VGND.n6 VGND.t2 239.703
R72 VGND.n2 VGND.n1 210.24
R73 VGND.n4 VGND.n3 199.873
R74 VGND.n3 VGND.t4 38.9194
R75 VGND.n3 VGND.t1 38.1086
R76 VGND.n1 VGND.t0 37.2978
R77 VGND.n1 VGND.t3 25.9464
R78 VGND.n5 VGND.n4 23.7181
R79 VGND.n6 VGND.n5 22.2123
R80 VGND.n7 VGND.n6 9.3005
R81 VGND.n5 VGND.n0 9.3005
R82 VGND.n4 VGND.n2 5.93461
R83 VGND.n2 VGND.n0 0.180378
R84 VGND.n7 VGND.n0 0.122949
R85 VGND VGND.n7 0.0617245
R86 VNB.t0 VNB.t2 2240.42
R87 VNB.t3 VNB.t6 1443.57
R88 VNB VNB.t4 1281.89
R89 VNB.t5 VNB.t1 1247.24
R90 VNB.t4 VNB.t3 993.177
R91 VNB.t2 VNB.t5 831.496
R92 VNB.t6 VNB.t0 831.496
R93 a_603_74.t0 a_603_74.t1 34.0546
R94 a_337_74.t0 a_337_74.t1 34.0546
C0 A2 B1 1.38e-19
C1 VPB B2 0.035659f
C2 X VGND 0.135312f
C3 A1 B1 0.067f
C4 VPB C1 0.045167f
C5 VPB VPWR 0.128188f
C6 VPB X 0.014005f
C7 A2 VPWR 0.027496f
C8 B1 B2 0.074214f
C9 A2 X 0.005275f
C10 A1 VPWR 0.021153f
C11 VPB VGND 0.00891f
C12 A2 VGND 0.015981f
C13 B2 C1 0.098293f
C14 B1 VPWR 0.007203f
C15 A1 X 5.43e-19
C16 A1 VGND 0.012258f
C17 B2 VPWR 0.00609f
C18 B1 X 7.83e-20
C19 C1 VPWR 0.010711f
C20 B1 VGND 0.011526f
C21 B2 X 2.52e-20
C22 VPB A2 0.043513f
C23 C1 X 1.65e-20
C24 B2 VGND 0.017524f
C25 VPB A1 0.047558f
C26 VPWR X 0.214506f
C27 C1 VGND 0.01458f
C28 VPB B1 0.057906f
C29 A2 A1 0.105155f
C30 VPWR VGND 0.070312f
C31 VGND VNB 0.558581f
C32 X VNB 0.065791f
C33 VPWR VNB 0.453487f
C34 C1 VNB 0.164843f
C35 B2 VNB 0.103842f
C36 B1 VNB 0.125726f
C37 A1 VNB 0.10954f
C38 A2 VNB 0.10898f
C39 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a221o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221o_1 VNB VPB VPWR VGND X C1 B2 A2 A1 B1
X0 VPWR.t2 A1.t0 a_310_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X1 a_310_392.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.199 ps=1.485 w=1 l=0.15
X2 a_148_260.t1 C1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.14295 ps=1.25 w=0.64 l=0.15
X3 VGND.t0 B2.t0 a_597_79.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.14295 pd=1.25 as=0.0672 ps=0.85 w=0.64 l=0.15
X4 a_509_392.t0 B2.t1 a_310_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X5 a_148_260.t2 C1.t1 a_509_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.165 ps=1.33 w=1 l=0.15
X6 a_310_392.t3 B1.t0 a_509_392.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X7 VGND.t2 a_148_260.t4 X.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.289475 pd=1.605 as=0.1961 ps=2.01 w=0.74 l=0.15
X8 VPWR.t1 a_148_260.t5 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.199 pd=1.485 as=0.308 ps=2.79 w=1.12 l=0.15
X9 a_417_79.t0 A2.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.289475 ps=1.605 w=0.64 l=0.15
X10 a_148_260.t0 A1.t1 a_417_79.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0672 ps=0.85 w=0.64 l=0.15
X11 a_597_79.t1 B1.t1 a_148_260.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1248 ps=1.03 w=0.64 l=0.15
R0 A1.n0 A1.t1 277.661
R1 A1.n0 A1.t0 237.47
R2 A1 A1.n0 154.133
R3 a_310_392.n1 a_310_392.n0 595.49
R4 a_310_392.n0 a_310_392.t2 29.5505
R5 a_310_392.n0 a_310_392.t3 29.5505
R6 a_310_392.n1 a_310_392.t1 29.5505
R7 a_310_392.t0 a_310_392.n1 29.5505
R8 VPWR.n1 VPWR.t2 350.983
R9 VPWR.n1 VPWR.n0 236.701
R10 VPWR.n0 VPWR.t0 42.3555
R11 VPWR.n0 VPWR.t1 27.4811
R12 VPWR VPWR.n1 0.629176
R13 VPB.t3 VPB.t5 495.43
R14 VPB VPB.t2 490.324
R15 VPB.t2 VPB.t0 263.038
R16 VPB.t4 VPB.t1 245.161
R17 VPB.t5 VPB.t4 229.839
R18 VPB.t0 VPB.t3 229.839
R19 A2.n0 A2.t1 311.986
R20 A2.n0 A2.t0 263.762
R21 A2 A2.n0 156.019
R22 C1.t0 C1.t1 460.31
R23 C1 C1.t0 327.349
R24 VGND.n5 VGND.n4 185
R25 VGND.n3 VGND.n0 185
R26 VGND.n2 VGND.n1 119.909
R27 VGND.n4 VGND.n3 109.689
R28 VGND.n1 VGND.t3 54.8797
R29 VGND.n1 VGND.t0 29.521
R30 VGND.n4 VGND.t1 26.2505
R31 VGND.n5 VGND.n2 24.6158
R32 VGND.n3 VGND.t2 20.4242
R33 VGND.n7 VGND.n6 9.3005
R34 VGND.n8 VGND.n0 7.43249
R35 VGND.n6 VGND.n0 6.50428
R36 VGND.n6 VGND.n5 1.59185
R37 VGND VGND.n8 0.276838
R38 VGND.n7 VGND.n2 0.217859
R39 VGND.n8 VGND.n7 0.153988
R40 a_148_260.n2 a_148_260.n1 360.49
R41 a_148_260.t2 a_148_260.n3 266.909
R42 a_148_260.n1 a_148_260.t5 264.298
R43 a_148_260.n3 a_148_260.t1 218.281
R44 a_148_260.n1 a_148_260.t4 204.048
R45 a_148_260.n2 a_148_260.n0 93.441
R46 a_148_260.n3 a_148_260.n2 86.8077
R47 a_148_260.n0 a_148_260.t3 36.563
R48 a_148_260.n0 a_148_260.t0 36.563
R49 VNB.t3 VNB.t1 2344.36
R50 VNB VNB.t3 2298.16
R51 VNB.t0 VNB.t4 1247.24
R52 VNB.t2 VNB.t5 1247.24
R53 VNB.t5 VNB.t0 831.496
R54 VNB.t1 VNB.t2 831.496
R55 B2.n0 B2.t0 260.281
R56 B2.n0 B2.t1 236.983
R57 B2 B2.n0 158.106
R58 a_597_79.t0 a_597_79.t1 39.3755
R59 a_509_392.n0 a_509_392.t2 604.808
R60 a_509_392.n0 a_509_392.t1 32.5055
R61 a_509_392.t0 a_509_392.n0 32.5055
R62 B1.n0 B1.t1 260.281
R63 B1.n0 B1.t0 236.983
R64 B1 B1.n0 162.438
R65 X.n1 X 587.066
R66 X.n1 X.n0 585
R67 X.n2 X.n1 585
R68 X X.t0 173.917
R69 X.n1 X.t1 26.3844
R70 X X.n2 5.5334
R71 X X.n0 4.79018
R72 X X.n0 1.32179
R73 X.n2 X 0.578565
R74 a_417_79.t0 a_417_79.t1 39.3755
C0 VPB X 0.041132f
C1 A1 B2 4.58e-20
C2 A2 C1 6.37e-20
C3 A2 X 0.005722f
C4 VPB VPWR 0.118262f
C5 B1 B2 0.107501f
C6 A1 C1 2.04e-20
C7 A2 VPWR 0.02725f
C8 A1 X 6.84e-19
C9 VPB VGND 0.00935f
C10 B1 X 9.88e-20
C11 A1 VPWR 0.022763f
C12 A2 VGND 0.025416f
C13 B2 C1 0.058699f
C14 A1 VGND 0.013318f
C15 B2 X 6.77e-20
C16 B1 VPWR 0.006573f
C17 B1 VGND 0.013251f
C18 B2 VPWR 0.007024f
C19 C1 X 1.72e-19
C20 VPB A2 0.049016f
C21 B2 VGND 0.01906f
C22 C1 VPWR 0.011153f
C23 VPB A1 0.061661f
C24 X VPWR 0.16714f
C25 C1 VGND 0.097711f
C26 A2 A1 0.121144f
C27 VPB B1 0.044548f
C28 X VGND 0.124238f
C29 VPB B2 0.040298f
C30 A2 B1 6.35e-19
C31 VPWR VGND 0.069626f
C32 A1 B1 0.079538f
C33 VPB C1 0.037109f
C34 A2 B2 1.18e-19
C35 VGND VNB 0.533566f
C36 VPWR VNB 0.420202f
C37 X VNB 0.137667f
C38 C1 VNB 0.208291f
C39 B2 VNB 0.111334f
C40 B1 VNB 0.10424f
C41 A1 VNB 0.120305f
C42 A2 VNB 0.161871f
C43 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a211oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a211oi_4 VNB VPB VPWR VGND Y C1 B1 A2 A1
X0 VGND.t4 A2.t0 a_92_74.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X2 Y.t0 A1.t0 a_92_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_901_368.t3 C1.t0 Y.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t7 C1.t1 a_901_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_77_368.t3 A1.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t2 A1.t2 a_77_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_92_74.t1 A1.t3 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_77_368.t1 A1.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VPWR.t0 A1.t5 a_77_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_92_74.t2 A1.t6 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_92_74.t6 A2.t1 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_901_368.t1 C1.t2 Y.t8 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 Y.t1 C1.t3 a_901_368.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_901_368.t7 B1.t0 a_77_368.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_92_74.t5 A2.t2 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 Y.t2 C1.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_77_368.t6 B1.t1 a_901_368.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X18 a_77_368.t5 B1.t2 a_901_368.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_901_368.t4 B1.t3 a_77_368.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_77_368.t11 A2.t3 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 Y.t5 A1.t7 a_92_74.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 Y.t9 B1.t4 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 VPWR.t6 A2.t4 a_77_368.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 VGND.t1 A2.t5 a_92_74.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 a_77_368.t9 A2.t6 VPWR.t5 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 VPWR.t4 A2.t7 a_77_368.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X27 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A2.n3 A2.t7 236.303
R1 A2.n0 A2.t3 226.809
R2 A2.n10 A2.t4 226.809
R3 A2.n2 A2.t6 226.809
R4 A2.n0 A2.t1 196.744
R5 A2.n3 A2.t0 196.013
R6 A2.n1 A2.t2 196.013
R7 A2.n11 A2.t5 196.013
R8 A2.n13 A2.n12 152
R9 A2.n9 A2.n8 152
R10 A2.n7 A2.n6 152
R11 A2.n5 A2.n4 152
R12 A2.n6 A2.n5 49.6611
R13 A2.n9 A2.n1 37.9763
R14 A2.n12 A2.n0 37.246
R15 A2.n12 A2.n11 24.8308
R16 A2.n10 A2.n9 21.1793
R17 A2.n8 A2.n7 10.1214
R18 A2.n4 A2 9.07957
R19 A2 A2.n13 7.29352
R20 A2.n13 A2 6.99585
R21 A2.n2 A2.n1 6.57323
R22 A2.n4 A2 5.2098
R23 A2.n6 A2.n2 5.11262
R24 A2.n11 A2.n10 3.65202
R25 A2.n8 A2 3.12608
R26 A2.n5 A2.n3 1.46111
R27 A2.n7 A2 1.04236
R28 a_92_74.n4 a_92_74.t1 321.276
R29 a_92_74.n1 a_92_74.t7 213.992
R30 a_92_74.n5 a_92_74.n4 185
R31 a_92_74.n1 a_92_74.n0 103.65
R32 a_92_74.n3 a_92_74.n2 86.3508
R33 a_92_74.n3 a_92_74.n1 80.4426
R34 a_92_74.n4 a_92_74.n3 53.841
R35 a_92_74.n2 a_92_74.t3 22.7032
R36 a_92_74.n2 a_92_74.t6 22.7032
R37 a_92_74.n0 a_92_74.t4 22.7032
R38 a_92_74.n0 a_92_74.t5 22.7032
R39 a_92_74.t0 a_92_74.n5 22.7032
R40 a_92_74.n5 a_92_74.t2 22.7032
R41 VGND.n7 VGND.t0 239.137
R42 VGND.n8 VGND.t5 231.946
R43 VGND.n22 VGND.n21 211.183
R44 VGND.n1 VGND.n0 211.183
R45 VGND.n10 VGND.n9 36.1417
R46 VGND.n10 VGND.n5 36.1417
R47 VGND.n14 VGND.n5 36.1417
R48 VGND.n15 VGND.n14 36.1417
R49 VGND.n16 VGND.n15 36.1417
R50 VGND.n16 VGND.n3 36.1417
R51 VGND.n20 VGND.n3 36.1417
R52 VGND.n24 VGND.n23 36.1417
R53 VGND.n21 VGND.t3 22.7032
R54 VGND.n21 VGND.t1 22.7032
R55 VGND.n0 VGND.t2 22.7032
R56 VGND.n0 VGND.t4 22.7032
R57 VGND.n9 VGND.n8 21.8358
R58 VGND.n26 VGND.n1 17.492
R59 VGND.n9 VGND.n6 9.3005
R60 VGND.n11 VGND.n10 9.3005
R61 VGND.n12 VGND.n5 9.3005
R62 VGND.n14 VGND.n13 9.3005
R63 VGND.n15 VGND.n4 9.3005
R64 VGND.n17 VGND.n16 9.3005
R65 VGND.n18 VGND.n3 9.3005
R66 VGND.n20 VGND.n19 9.3005
R67 VGND.n23 VGND.n2 9.3005
R68 VGND.n25 VGND.n24 9.3005
R69 VGND.n22 VGND.n20 9.03579
R70 VGND.n8 VGND.n7 6.68056
R71 VGND.n23 VGND.n22 2.25932
R72 VGND.n24 VGND.n1 1.50638
R73 VGND.n7 VGND.n6 0.662843
R74 VGND VGND.n26 0.163644
R75 VGND.n26 VGND.n25 0.144205
R76 VGND.n11 VGND.n6 0.122949
R77 VGND.n12 VGND.n11 0.122949
R78 VGND.n13 VGND.n12 0.122949
R79 VGND.n13 VGND.n4 0.122949
R80 VGND.n17 VGND.n4 0.122949
R81 VGND.n18 VGND.n17 0.122949
R82 VGND.n19 VGND.n18 0.122949
R83 VGND.n19 VGND.n2 0.122949
R84 VGND.n25 VGND.n2 0.122949
R85 VNB.t2 VNB.t9 5497.11
R86 VNB.t9 VNB.t1 1986.35
R87 VNB VNB.t8 1847.77
R88 VNB.t0 VNB.t2 993.177
R89 VNB.t3 VNB.t0 993.177
R90 VNB.t4 VNB.t3 993.177
R91 VNB.t7 VNB.t4 993.177
R92 VNB.t5 VNB.t7 993.177
R93 VNB.t6 VNB.t5 993.177
R94 VNB.t8 VNB.t6 993.177
R95 B1.n10 B1.t1 251.151
R96 B1.n2 B1.t0 242.835
R97 B1.n5 B1.t2 240.197
R98 B1.n0 B1.t3 240.197
R99 B1.n2 B1.t4 179.947
R100 B1.n4 B1.n1 179.947
R101 B1.n3 B1 152.934
R102 B1.n7 B1.n6 152
R103 B1.n9 B1.n8 152
R104 B1.n11 B1.n10 152
R105 B1.n10 B1.n9 49.6611
R106 B1.n6 B1.n0 44.549
R107 B1.n3 B1.n2 35.055
R108 B1.n4 B1.n3 27.752
R109 B1.n6 B1.n5 21.1793
R110 B1 B1.n11 12.1338
R111 B1.n8 B1 8.4005
R112 B1.n7 B1 8.13383
R113 B1.n9 B1.n0 5.11262
R114 B1 B1.n7 4.66717
R115 B1.n8 B1 4.4005
R116 B1.n5 B1.n4 0.730803
R117 B1.n11 B1 0.667167
R118 Y.n2 Y.n0 362.098
R119 Y.n2 Y.n1 304.724
R120 Y.n6 Y.n4 216.907
R121 Y.n6 Y.n5 185
R122 Y.n7 Y.n6 180.052
R123 Y.n7 Y.t9 154.728
R124 Y.n8 Y.t2 143.445
R125 Y.n8 Y.n7 57.029
R126 Y.n1 Y.t6 26.3844
R127 Y.n1 Y.t7 26.3844
R128 Y.n0 Y.t8 26.3844
R129 Y.n0 Y.t1 26.3844
R130 Y.n4 Y.t4 22.7032
R131 Y.n4 Y.t5 22.7032
R132 Y.n5 Y.t3 22.7032
R133 Y.n5 Y.t0 22.7032
R134 Y Y.n2 11.4354
R135 Y Y.n8 8.79086
R136 Y Y.n3 4.39568
R137 Y.n3 Y 3.00773
R138 Y.n3 Y 0.486576
R139 A1.n0 A1.t1 237.762
R140 A1.n2 A1.t2 226.809
R141 A1.n4 A1.t4 226.809
R142 A1.n6 A1.t5 226.809
R143 A1.n6 A1.t7 198.204
R144 A1.n5 A1.t6 196.013
R145 A1.n3 A1.t0 196.013
R146 A1.n0 A1.t3 196.013
R147 A1 A1.n1 157.209
R148 A1.n12 A1.n11 152
R149 A1.n10 A1.n9 152
R150 A1.n8 A1.n7 152
R151 A1.n11 A1.n10 49.6611
R152 A1.n7 A1.n5 40.8975
R153 A1.n2 A1.n1 37.246
R154 A1.n7 A1.n6 19.7187
R155 A1.n1 A1.n0 17.5278
R156 A1.n9 A1.n8 10.1214
R157 A1.n12 A1 9.37724
R158 A1.n3 A1.n2 8.03383
R159 A1.n5 A1.n4 5.11262
R160 A1 A1.n12 4.91213
R161 A1.n11 A1.n3 4.38232
R162 A1.n10 A1.n4 3.65202
R163 A1.n8 A1 3.42376
R164 A1.n9 A1 0.744686
R165 C1.n0 C1.t0 287.058
R166 C1.n0 C1.t1 226.809
R167 C1.n2 C1.t2 226.809
R168 C1.n4 C1.t3 226.809
R169 C1.n4 C1.n3 191.06
R170 C1.n7 C1.t4 186.374
R171 C1 C1.n1 153.042
R172 C1.n8 C1.n7 152
R173 C1.n6 C1.n5 152
R174 C1.n7 C1.n6 45.5227
R175 C1.n2 C1.n1 38.1588
R176 C1.n1 C1.n0 22.0922
R177 C1.n5 C1 9.37724
R178 C1 C1.n8 9.07957
R179 C1.n7 C1.n2 7.36439
R180 C1.n6 C1.n4 7.36439
R181 C1.n8 C1 5.2098
R182 C1.n5 C1 4.91213
R183 a_901_368.t3 a_901_368.n5 373.642
R184 a_901_368.n1 a_901_368.t6 372.606
R185 a_901_368.n5 a_901_368.n4 302.74
R186 a_901_368.n1 a_901_368.n0 302.719
R187 a_901_368.n3 a_901_368.n2 211.669
R188 a_901_368.n3 a_901_368.n1 46.6829
R189 a_901_368.n5 a_901_368.n3 42.9181
R190 a_901_368.n0 a_901_368.t5 26.3844
R191 a_901_368.n0 a_901_368.t4 26.3844
R192 a_901_368.n2 a_901_368.t0 26.3844
R193 a_901_368.n2 a_901_368.t7 26.3844
R194 a_901_368.n4 a_901_368.t2 26.3844
R195 a_901_368.n4 a_901_368.t1 26.3844
R196 VPB.t3 VPB.t10 495.43
R197 VPB VPB.t12 375.404
R198 VPB.t6 VPB.t7 229.839
R199 VPB.t5 VPB.t6 229.839
R200 VPB.t4 VPB.t5 229.839
R201 VPB.t11 VPB.t4 229.839
R202 VPB.t9 VPB.t11 229.839
R203 VPB.t8 VPB.t9 229.839
R204 VPB.t10 VPB.t8 229.839
R205 VPB.t2 VPB.t3 229.839
R206 VPB.t1 VPB.t2 229.839
R207 VPB.t0 VPB.t1 229.839
R208 VPB.t15 VPB.t0 229.839
R209 VPB.t14 VPB.t15 229.839
R210 VPB.t13 VPB.t14 229.839
R211 VPB.t12 VPB.t13 229.839
R212 VPWR.n13 VPWR.n1 331.5
R213 VPWR.n5 VPWR.n4 321.853
R214 VPWR.n3 VPWR.n2 316.353
R215 VPWR.n7 VPWR.n6 316.353
R216 VPWR.n12 VPWR.n11 36.1417
R217 VPWR.n8 VPWR.n7 32.7534
R218 VPWR.n1 VPWR.t5 26.3844
R219 VPWR.n1 VPWR.t4 26.3844
R220 VPWR.n2 VPWR.t7 26.3844
R221 VPWR.n2 VPWR.t6 26.3844
R222 VPWR.n6 VPWR.t1 26.3844
R223 VPWR.n6 VPWR.t0 26.3844
R224 VPWR.n4 VPWR.t3 26.3844
R225 VPWR.n4 VPWR.t2 26.3844
R226 VPWR.n14 VPWR.n13 25.7744
R227 VPWR.n13 VPWR.n12 18.0711
R228 VPWR.n8 VPWR.n3 10.1652
R229 VPWR.n9 VPWR.n8 9.3005
R230 VPWR.n11 VPWR.n10 9.3005
R231 VPWR.n12 VPWR.n0 9.3005
R232 VPWR.n7 VPWR.n5 6.08183
R233 VPWR.n11 VPWR.n3 1.12991
R234 VPWR.n9 VPWR.n5 0.593891
R235 VPWR VPWR.n14 0.163644
R236 VPWR.n14 VPWR.n0 0.144205
R237 VPWR.n10 VPWR.n9 0.122949
R238 VPWR.n10 VPWR.n0 0.122949
R239 a_77_368.n8 a_77_368.n7 360.557
R240 a_77_368.n8 a_77_368.n6 300.733
R241 a_77_368.n3 a_77_368.t8 272.759
R242 a_77_368.t3 a_77_368.n9 232.042
R243 a_77_368.n4 a_77_368.n1 208.423
R244 a_77_368.n5 a_77_368.n0 208.423
R245 a_77_368.n3 a_77_368.n2 206.078
R246 a_77_368.n5 a_77_368.n4 67.7652
R247 a_77_368.n9 a_77_368.n5 61.3652
R248 a_77_368.n4 a_77_368.n3 61.3652
R249 a_77_368.n9 a_77_368.n8 60.6123
R250 a_77_368.n6 a_77_368.t4 26.3844
R251 a_77_368.n6 a_77_368.t6 26.3844
R252 a_77_368.n7 a_77_368.t7 26.3844
R253 a_77_368.n7 a_77_368.t5 26.3844
R254 a_77_368.n1 a_77_368.t0 26.3844
R255 a_77_368.n1 a_77_368.t11 26.3844
R256 a_77_368.n0 a_77_368.t2 26.3844
R257 a_77_368.n0 a_77_368.t1 26.3844
R258 a_77_368.n2 a_77_368.t10 26.3844
R259 a_77_368.n2 a_77_368.t9 26.3844
C0 C1 Y 0.323955f
C1 B1 VGND 0.043432f
C2 VPWR Y 0.029212f
C3 C1 VGND 0.040552f
C4 VPB A2 0.146276f
C5 VPWR VGND 0.133564f
C6 VPB A1 0.138318f
C7 Y VGND 0.48246f
C8 VPB B1 0.139466f
C9 A2 A1 0.088805f
C10 A2 B1 6.1e-20
C11 VPB C1 0.137558f
C12 VPB VPWR 0.204113f
C13 A1 B1 0.035077f
C14 A2 VPWR 0.066567f
C15 VPB Y 0.014604f
C16 A2 Y 4.3e-20
C17 B1 C1 0.093802f
C18 VPB VGND 0.01215f
C19 A1 VPWR 0.08142f
C20 B1 VPWR 0.024444f
C21 A2 VGND 0.070588f
C22 A1 Y 0.130876f
C23 A1 VGND 0.027574f
C24 B1 Y 0.175551f
C25 C1 VPWR 0.02259f
C26 VGND VNB 1.01728f
C27 Y VNB 0.202227f
C28 VPWR VNB 0.791152f
C29 C1 VNB 0.351656f
C30 B1 VNB 0.348308f
C31 A1 VNB 0.406523f
C32 A2 VNB 0.449303f
C33 VPB VNB 2.01326f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a211oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a211oi_2 VNB VPB VPWR VGND Y C1 B1 A2 A1
X0 VGND.t2 C1.t0 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2664 ps=1.46 w=0.74 l=0.15
X1 VPWR.t1 A2.t0 a_114_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2 VGND.t3 A2.t1 a_38_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_114_368.t0 A2.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t0 B1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2664 pd=1.46 as=0.1961 ps=2.01 w=0.74 l=0.15
X5 VPWR.t3 A1.t0 a_114_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_38_74.t2 A1.t1 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 Y.t5 A1.t2 a_38_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X8 a_38_74.t0 A2.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2183 pd=2.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X9 a_114_368.t3 A1.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X10 a_497_368.t3 C1.t1 Y.t2 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t3 C1.t2 a_497_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_497_368.t1 B1.t1 a_114_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_114_368.t5 B1.t2 a_497_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
R0 C1.n1 C1.t1 272.574
R1 C1.n0 C1.t2 261.62
R2 C1.n0 C1.t0 160.814
R3 C1.n2 C1.n1 152
R4 C1.n1 C1.n0 54.7732
R5 C1.n2 C1 11.9356
R6 C1 C1.n2 4.67077
R7 Y.n3 Y.n1 339.291
R8 Y Y.n0 300.911
R9 Y.n3 Y.n2 70.8935
R10 Y.n2 Y.t4 57.7404
R11 Y.n2 Y.t0 44.7306
R12 Y.n0 Y.t2 26.3844
R13 Y.n0 Y.t3 26.3844
R14 Y.n1 Y.t1 22.7032
R15 Y.n1 Y.t5 22.7032
R16 Y Y.n3 1.94833
R17 VGND.n4 VGND.t0 292.372
R18 VGND.n1 VGND.n0 209.155
R19 VGND.n3 VGND.t2 160.541
R20 VGND.n6 VGND.n5 36.1417
R21 VGND.n8 VGND.n1 32.1234
R22 VGND.n0 VGND.t1 25.9464
R23 VGND.n0 VGND.t3 25.9464
R24 VGND.n5 VGND.n4 22.5887
R25 VGND.n6 VGND.n1 11.6711
R26 VGND.n7 VGND.n6 9.3005
R27 VGND.n5 VGND.n2 9.3005
R28 VGND.n4 VGND.n3 7.10562
R29 VGND VGND.n8 0.282382
R30 VGND.n3 VGND.n2 0.254824
R31 VGND.n8 VGND.n7 0.148529
R32 VGND.n7 VGND.n2 0.122949
R33 VNB.t2 VNB.t0 2263.52
R34 VNB.t0 VNB.t3 2009.45
R35 VNB VNB.t5 1224.15
R36 VNB.t4 VNB.t2 1085.56
R37 VNB.t1 VNB.t4 993.177
R38 VNB.t5 VNB.t1 993.177
R39 A2.n0 A2.t0 226.809
R40 A2.n1 A2.t2 226.809
R41 A2.n0 A2.t3 198.204
R42 A2.n1 A2.t1 196.744
R43 A2.n5 A2.n4 152
R44 A2.n3 A2.n2 152
R45 A2.n4 A2.n3 52.5823
R46 A2 A2.n5 11.1548
R47 A2.n4 A2.n0 10.955
R48 A2.n2 A2 10.7891
R49 A2.n2 A2 6.76621
R50 A2.n5 A2 6.4005
R51 A2.n3 A2.n1 2.19141
R52 a_114_368.n2 a_114_368.n0 376.808
R53 a_114_368.n2 a_114_368.n1 264.51
R54 a_114_368.n3 a_114_368.n2 204.838
R55 a_114_368.n1 a_114_368.t4 26.3844
R56 a_114_368.n1 a_114_368.t3 26.3844
R57 a_114_368.n0 a_114_368.t2 26.3844
R58 a_114_368.n0 a_114_368.t5 26.3844
R59 a_114_368.n3 a_114_368.t1 26.3844
R60 a_114_368.t0 a_114_368.n3 26.3844
R61 VPWR.n1 VPWR.t1 347.149
R62 VPWR.n3 VPWR.n2 316.683
R63 VPWR.n5 VPWR.t2 259.171
R64 VPWR.n5 VPWR.n4 27.4829
R65 VPWR.n2 VPWR.t0 26.3844
R66 VPWR.n2 VPWR.t3 26.3844
R67 VPWR.n4 VPWR.n3 21.4593
R68 VPWR.n4 VPWR.n0 9.3005
R69 VPWR.n6 VPWR.n5 9.3005
R70 VPWR.n3 VPWR.n1 6.76052
R71 VPWR.n1 VPWR.n0 0.611706
R72 VPWR.n6 VPWR.n0 0.122949
R73 VPWR VPWR.n6 0.0617245
R74 VPB.t1 VPB.t5 515.861
R75 VPB VPB.t3 252.823
R76 VPB.t6 VPB.t7 229.839
R77 VPB.t2 VPB.t6 229.839
R78 VPB.t5 VPB.t2 229.839
R79 VPB.t0 VPB.t1 229.839
R80 VPB.t4 VPB.t0 229.839
R81 VPB.t3 VPB.t4 229.839
R82 a_38_74.n0 a_38_74.t3 204.137
R83 a_38_74.n0 a_38_74.t0 182.638
R84 a_38_74.n1 a_38_74.n0 88.3446
R85 a_38_74.t1 a_38_74.n1 22.7032
R86 a_38_74.n1 a_38_74.t2 22.7032
R87 B1.n1 B1.t1 268.192
R88 B1.n0 B1.t2 261.62
R89 B1.n0 B1.t0 156.431
R90 B1.n2 B1.n1 152
R91 B1.n1 B1.n0 59.155
R92 B1.n2 B1 8.82212
R93 B1 B1.n2 7.78428
R94 A1.n0 A1.t0 261.62
R95 A1.n2 A1.t3 261.62
R96 A1 A1.n2 183.141
R97 A1.n0 A1.t1 156.431
R98 A1.n1 A1.t2 154.24
R99 A1.n1 A1.n0 60.6157
R100 A1.n2 A1.n1 5.11262
R101 a_497_368.n0 a_497_368.t0 383.885
R102 a_497_368.n1 a_497_368.n0 309.978
R103 a_497_368.n0 a_497_368.t3 303.128
R104 a_497_368.n1 a_497_368.t2 26.3844
R105 a_497_368.t1 a_497_368.n1 26.3844
C0 A2 VGND 0.02897f
C1 C1 VPWR 0.013204f
C2 B1 Y 0.195206f
C3 B1 VGND 0.022384f
C4 C1 Y 0.060967f
C5 C1 VGND 0.053306f
C6 VPWR Y 0.016265f
C7 VPB A1 0.070152f
C8 VPWR VGND 0.077005f
C9 VPB A2 0.072784f
C10 Y VGND 0.221242f
C11 VPB B1 0.062986f
C12 A1 A2 0.075608f
C13 VPB C1 0.064339f
C14 VPB VPWR 0.135539f
C15 A2 B1 0.020383f
C16 A1 VPWR 0.059019f
C17 VPB Y 0.013089f
C18 VPB VGND 0.009021f
C19 B1 C1 0.091943f
C20 A2 VPWR 0.041022f
C21 A1 Y 0.037817f
C22 A2 Y 0.146894f
C23 B1 VPWR 0.01192f
C24 A1 VGND 0.015019f
C25 VGND VNB 0.627008f
C26 Y VNB 0.055267f
C27 VPWR VNB 0.505818f
C28 C1 VNB 0.227404f
C29 B1 VNB 0.182038f
C30 A2 VNB 0.218441f
C31 A1 VNB 0.263661f
C32 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a211oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a211oi_1 VNB VPB VPWR VGND C1 Y B1 A2 A1
X0 a_71_368.t2 A1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2184 ps=1.51 w=1.12 l=0.15
X1 Y.t3 A1.t1 a_159_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X2 a_159_74.t0 A2.t0 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1961 ps=2.01 w=0.74 l=0.15
X3 VGND.t0 B1.t0 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X4 Y.t1 C1.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X5 VPWR.t0 A2.t1 a_71_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.308 ps=2.79 w=1.12 l=0.15
X6 a_354_368.t0 B1.t1 a_71_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t2 C1.t1 a_354_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1848 ps=1.45 w=1.12 l=0.15
R0 A1.n0 A1.t0 250.909
R1 A1.n0 A1.t1 220.113
R2 A1 A1.n0 154.522
R3 VPWR VPWR.n0 323.974
R4 VPWR.n0 VPWR.t1 38.6969
R5 VPWR.n0 VPWR.t0 29.9023
R6 a_71_368.t0 a_71_368.n0 483.243
R7 a_71_368.n0 a_71_368.t1 26.3844
R8 a_71_368.n0 a_71_368.t2 26.3844
R9 VPB VPB.t0 360.082
R10 VPB.t0 VPB.t3 275.807
R11 VPB.t1 VPB.t2 245.161
R12 VPB.t3 VPB.t1 229.839
R13 a_159_74.t0 a_159_74.t1 34.0546
R14 Y.n1 Y.n0 610.134
R15 Y.n2 Y.t2 279.219
R16 Y.n3 Y 195.024
R17 Y.n4 Y.n3 185
R18 Y.n0 Y.t1 143.78
R19 Y.n3 Y.t0 37.2978
R20 Y Y.n0 34.1338
R21 Y.n3 Y.t3 25.9464
R22 Y.n1 Y 16.1735
R23 Y Y.n4 4.21229
R24 Y.n4 Y 3.85592
R25 Y.n2 Y.n1 2.76807
R26 Y Y.n2 1.9032
R27 VNB VNB.t0 1662.99
R28 VNB.t1 VNB.t2 1247.24
R29 VNB.t3 VNB.t1 1247.24
R30 VNB.t0 VNB.t3 831.496
R31 A2.n0 A2.t1 250.909
R32 A2.n0 A2.t0 220.113
R33 A2 A2.n0 154.25
R34 VGND.n1 VGND.n0 208.904
R35 VGND.n1 VGND.t2 174.308
R36 VGND.n0 VGND.t1 37.2978
R37 VGND.n0 VGND.t0 25.9464
R38 VGND VGND.n1 0.264003
R39 B1.n0 B1.t1 250.909
R40 B1.n0 B1.t0 220.113
R41 B1 B1.n0 155.423
R42 C1.n0 C1.t1 261.62
R43 C1 C1.n0 222.325
R44 C1.n0 C1.t0 156.431
R45 a_354_368.t0 a_354_368.t1 58.0451
C0 Y VPB 0.02222f
C1 VPWR VGND 0.04779f
C2 VGND VPB 0.010661f
C3 Y VGND 0.224772f
C4 A2 A1 0.101689f
C5 A1 B1 0.087781f
C6 A2 VPWR 0.014286f
C7 A2 VPB 0.039218f
C8 B1 C1 0.05502f
C9 A2 Y 0.004962f
C10 A1 VPWR 0.015694f
C11 B1 VPWR 0.011024f
C12 A1 Y 0.035296f
C13 A2 VGND 0.037256f
C14 A1 VPB 0.032663f
C15 B1 VPB 0.032316f
C16 C1 VPWR 0.007265f
C17 B1 Y 0.089148f
C18 A1 VGND 0.013563f
C19 C1 VPB 0.05303f
C20 C1 Y 0.099823f
C21 B1 VGND 0.013345f
C22 VPWR VPB 0.084582f
C23 VPWR Y 0.062215f
C24 C1 VGND 0.016228f
C25 VGND VNB 0.433536f
C26 Y VNB 0.106495f
C27 VPWR VNB 0.318578f
C28 C1 VNB 0.192006f
C29 B1 VNB 0.104112f
C30 A1 VNB 0.100703f
C31 A2 VNB 0.14637f
C32 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a211o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a211o_4 VNB VPB VPWR VGND X C1 B1 A2 A1
X0 VGND.t5 a_105_280.t8 X.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.12205 pd=1.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_517_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.3275 ps=1.655 w=1 l=0.15
X2 VGND.t4 a_105_280.t9 X.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_105_280.t0 A1.t0 a_1064_123.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 a_105_280.t6 B1.t0 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.12205 ps=1.08 w=0.64 l=0.15
X5 a_517_392# B1.t1 a_602_392.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1525 pd=1.305 as=0.1625 ps=1.325 w=1 l=0.15
X6 X.t1 a_105_280.t10 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 VPWR.t4 a_105_280.t11 X.t7 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_602_392.t0 C1.t0 a_105_280.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1625 pd=1.325 as=0.15 ps=1.3 w=1 l=0.15
X9 VPWR.t0 A2.t0 a_517_392# VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.3275 pd=1.655 as=0.1525 ps=1.305 w=1 l=0.15
X10 X.t0 a_105_280.t12 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X11 VGND.t7 C1.t1 a_105_280.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.114925 pd=1.05 as=0.0896 ps=0.92 w=0.64 l=0.15
X12 X.t6 a_105_280.t13 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 VGND.t0 A2.t1 a_1064_123.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X14 VPWR.t2 a_105_280.t14 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_105_280.t3 C1.t2 a_602_392.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.175 ps=1.35 w=1 l=0.15
X16 a_105_280.t4 C1.t3 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.11055 pd=1.04 as=0.114925 ps=1.05 w=0.64 l=0.15
X17 a_1064_123.t2 A1.t1 a_105_280.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X18 a_602_392.t1 B1.t2 a_517_392# VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.275 ps=2.55 w=1 l=0.15
X19 a_517_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X20 X.t4 a_105_280.t15 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X21 VPWR.t5 A1.t2 a_517_392# VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X22 a_1064_123.t1 A2.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.2304 ps=1.36 w=0.64 l=0.15
X23 VGND.t9 B1.t3 a_105_280.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.2304 pd=1.36 as=0.11055 ps=1.04 w=0.64 l=0.15
R0 a_105_280.n13 a_105_280.n12 708.482
R1 a_105_280.n5 a_105_280.t15 397.382
R2 a_105_280.n3 a_105_280.n1 315.185
R3 a_105_280.n7 a_105_280.t13 272.954
R4 a_105_280.n5 a_105_280.t14 261.62
R5 a_105_280.n9 a_105_280.t11 261.62
R6 a_105_280.n11 a_105_280.t8 241
R7 a_105_280.n6 a_105_280.t12 212.081
R8 a_105_280.n3 a_105_280.n2 187.696
R9 a_105_280.n12 a_105_280.n11 164.19
R10 a_105_280.n8 a_105_280.t9 154.24
R11 a_105_280.n10 a_105_280.t10 154.24
R12 a_105_280.n4 a_105_280.n0 96.6897
R13 a_105_280.n7 a_105_280.n6 73.7211
R14 a_105_280.n4 a_105_280.n3 51.4797
R15 a_105_280.n9 a_105_280.n8 48.9308
R16 a_105_280.n12 a_105_280.n4 48.1787
R17 a_105_280.n6 a_105_280.n5 43.3805
R18 a_105_280.n2 a_105_280.t4 30.1551
R19 a_105_280.t2 a_105_280.n13 29.5505
R20 a_105_280.n13 a_105_280.t3 29.5505
R21 a_105_280.n2 a_105_280.t7 29.0932
R22 a_105_280.n0 a_105_280.t5 26.2505
R23 a_105_280.n0 a_105_280.t6 26.2505
R24 a_105_280.n1 a_105_280.t1 26.2505
R25 a_105_280.n1 a_105_280.t0 26.2505
R26 a_105_280.n10 a_105_280.n9 13.8763
R27 a_105_280.n11 a_105_280.n10 10.2247
R28 a_105_280.n8 a_105_280.n7 9.45779
R29 X.n2 X.n0 259.644
R30 X.n4 X.n3 222.746
R31 X.n2 X.n1 215.636
R32 X.n5 X 207.083
R33 X.n6 X.n5 185
R34 X X.n2 58.2362
R35 X.n1 X.t5 26.3844
R36 X.n1 X.t4 26.3844
R37 X.n0 X.t7 26.3844
R38 X.n0 X.t6 26.3844
R39 X.n3 X.t3 22.7032
R40 X.n3 X.t1 22.7032
R41 X.n5 X.t2 22.7032
R42 X.n5 X.t0 22.7032
R43 X X.n6 6.74459
R44 X.n6 X.n4 2.47792
R45 X X.n4 0.963941
R46 VGND.n6 VGND.n5 214.673
R47 VGND.n11 VGND.n10 208.856
R48 VGND.n18 VGND.n17 205.364
R49 VGND.n7 VGND.t0 172.37
R50 VGND.n0 VGND.t2 167.655
R51 VGND.n3 VGND.n2 115.659
R52 VGND.n5 VGND.t1 108.751
R53 VGND.n2 VGND.t8 37.5005
R54 VGND.n10 VGND.t6 37.3727
R55 VGND.n19 VGND.n18 36.1417
R56 VGND.n16 VGND.n3 28.6123
R57 VGND.n5 VGND.t9 26.2505
R58 VGND.n9 VGND.n6 25.977
R59 VGND.n12 VGND.n11 25.6005
R60 VGND.n10 VGND.t7 24.1459
R61 VGND.n17 VGND.t3 22.7032
R62 VGND.n17 VGND.t4 22.7032
R63 VGND.n2 VGND.t5 22.1988
R64 VGND.n11 VGND.n9 21.8358
R65 VGND.n12 VGND.n3 18.824
R66 VGND.n21 VGND.n0 15.2332
R67 VGND.n18 VGND.n16 11.2946
R68 VGND.n20 VGND.n19 9.3005
R69 VGND.n18 VGND.n1 9.3005
R70 VGND.n16 VGND.n15 9.3005
R71 VGND.n14 VGND.n3 9.3005
R72 VGND.n13 VGND.n12 9.3005
R73 VGND.n11 VGND.n4 9.3005
R74 VGND.n9 VGND.n8 9.3005
R75 VGND.n7 VGND.n6 7.01674
R76 VGND.n19 VGND.n0 3.76521
R77 VGND.n8 VGND.n7 0.164582
R78 VGND VGND.n21 0.163644
R79 VGND.n21 VGND.n20 0.144205
R80 VGND.n8 VGND.n4 0.122949
R81 VGND.n13 VGND.n4 0.122949
R82 VGND.n14 VGND.n13 0.122949
R83 VGND.n15 VGND.n14 0.122949
R84 VGND.n15 VGND.n1 0.122949
R85 VGND.n20 VGND.n1 0.122949
R86 VNB VNB.t4 2771.65
R87 VNB.t11 VNB.t1 2009.45
R88 VNB.t9 VNB.t8 1131.76
R89 VNB.t7 VNB.t10 1131.76
R90 VNB.t8 VNB.t11 1097.11
R91 VNB.t3 VNB.t0 993.177
R92 VNB.t2 VNB.t3 993.177
R93 VNB.t1 VNB.t2 993.177
R94 VNB.t10 VNB.t9 993.177
R95 VNB.t5 VNB.t7 993.177
R96 VNB.t6 VNB.t5 993.177
R97 VNB.t4 VNB.t6 993.177
R98 A1.n2 A1.n1 220.917
R99 A1.n0 A1.t2 212.883
R100 A1.n0 A1.t1 170.6
R101 A1.n2 A1.t0 165.488
R102 A1.n4 A1.n3 152
R103 A1.n3 A1.n0 54.7732
R104 A1.n4 A1 10.0853
R105 A1 A1.n4 8.53383
R106 A1.n3 A1.n2 2.92171
R107 VPWR.n6 VPWR.t5 352.123
R108 VPWR.n20 VPWR.n2 326.231
R109 VPWR.n14 VPWR.t4 270.3
R110 VPWR.n22 VPWR.t1 259.171
R111 VPWR.n7 VPWR.t0 203.18
R112 VPWR.n8 VPWR.n5 36.1417
R113 VPWR.n12 VPWR.n5 36.1417
R114 VPWR.n13 VPWR.n12 36.1417
R115 VPWR.n15 VPWR.n13 36.1417
R116 VPWR.n19 VPWR.n3 36.1417
R117 VPWR.n15 VPWR.n14 33.8829
R118 VPWR.n21 VPWR.n20 30.4946
R119 VPWR.n2 VPWR.t3 26.3844
R120 VPWR.n2 VPWR.t2 26.3844
R121 VPWR.n8 VPWR.n7 24.0946
R122 VPWR.n20 VPWR.n19 22.9652
R123 VPWR.n22 VPWR.n21 18.4476
R124 VPWR.n9 VPWR.n8 9.3005
R125 VPWR.n10 VPWR.n5 9.3005
R126 VPWR.n12 VPWR.n11 9.3005
R127 VPWR.n13 VPWR.n4 9.3005
R128 VPWR.n16 VPWR.n15 9.3005
R129 VPWR.n17 VPWR.n3 9.3005
R130 VPWR.n19 VPWR.n18 9.3005
R131 VPWR.n20 VPWR.n1 9.3005
R132 VPWR.n21 VPWR.n0 9.3005
R133 VPWR.n23 VPWR.n22 9.3005
R134 VPWR.n7 VPWR.n6 3.80607
R135 VPWR.n14 VPWR.n3 2.25932
R136 VPWR.n9 VPWR.n6 0.520877
R137 VPWR.n10 VPWR.n9 0.122949
R138 VPWR.n11 VPWR.n10 0.122949
R139 VPWR.n11 VPWR.n4 0.122949
R140 VPWR.n16 VPWR.n4 0.122949
R141 VPWR.n17 VPWR.n16 0.122949
R142 VPWR.n18 VPWR.n17 0.122949
R143 VPWR.n18 VPWR.n1 0.122949
R144 VPWR.n1 VPWR.n0 0.122949
R145 VPWR.n23 VPWR.n0 0.122949
R146 VPWR VPWR.n23 0.0617245
R147 VPB.t0 VPB.t7 640.995
R148 VPB.t5 VPB.t9 495.43
R149 VPB VPB.t2 314.113
R150 VPB.t9 VPB.t6 255.376
R151 VPB.t1 VPB.t8 242.608
R152 VPB.t8 VPB.t0 232.393
R153 VPB.t6 VPB.t1 229.839
R154 VPB.t4 VPB.t5 229.839
R155 VPB.t3 VPB.t4 229.839
R156 VPB.t2 VPB.t3 229.839
R157 a_1064_123.n1 a_1064_123.n0 346.986
R158 a_1064_123.n0 a_1064_123.t3 26.2505
R159 a_1064_123.n0 a_1064_123.t1 26.2505
R160 a_1064_123.n1 a_1064_123.t0 26.2505
R161 a_1064_123.t2 a_1064_123.n1 26.2505
R162 B1.n1 B1.t0 242.607
R163 B1.n0 B1.t1 231.629
R164 B1.n1 B1.t2 231.629
R165 B1 B1.n1 224.468
R166 B1.n0 B1.t3 196.013
R167 B1.n2 B1.n0 159.772
R168 B1 B1.n2 4.92358
R169 B1.n2 B1 3.04812
R170 a_602_392.n1 a_602_392.n0 1216.59
R171 a_602_392.n0 a_602_392.t1 39.4005
R172 a_602_392.t2 a_602_392.n1 32.5055
R173 a_602_392.n1 a_602_392.t0 31.5205
R174 a_602_392.n0 a_602_392.t3 29.5505
R175 C1.n0 C1.t0 255.728
R176 C1.n1 C1.t2 255.728
R177 C1.n1 C1.t1 164.319
R178 C1 C1.n2 161.504
R179 C1.n0 C1.t3 140.364
R180 C1.n2 C1.n0 39.4369
R181 C1.n2 C1.n1 26.2914
R182 A2.n1 A2.t1 622.948
R183 A2.t2 A2.t0 549.481
R184 A2.t1 A2.n0 463.257
R185 A2.n1 A2.t2 162.274
R186 A2.n2 A2.n1 158.656
R187 A2 A2.n2 5.4308
R188 A2.n2 A2 3.5845
C0 VPB VPWR 0.213727f
C1 C1 A2 0.002855f
C2 B1 A1 0.015045f
C3 C1 A1 6.41e-19
C4 VPB X 0.013305f
C5 B1 VPWR 0.023699f
C6 a_517_392# VPB 0.029643f
C7 C1 VPWR 0.012169f
C8 B1 X 7.19e-19
C9 A2 A1 0.140468f
C10 VPB VGND 0.017317f
C11 a_517_392# B1 0.07291f
C12 B1 VGND 0.032383f
C13 C1 X 1.66e-20
C14 A2 VPWR 0.037305f
C15 a_517_392# C1 0.017077f
C16 A1 VPWR 0.03785f
C17 C1 VGND 0.028416f
C18 a_517_392# A2 0.04361f
C19 A2 VGND 0.158317f
C20 a_517_392# A1 0.122085f
C21 VPWR X 0.423633f
C22 A1 VGND 0.011781f
C23 VPB B1 0.100984f
C24 a_517_392# VPWR 0.492972f
C25 VPWR VGND 0.126843f
C26 VPB C1 0.07142f
C27 X VGND 0.251844f
C28 a_517_392# VGND 0.019429f
C29 B1 C1 0.196714f
C30 VPB A2 0.088545f
C31 B1 A2 0.058509f
C32 VPB A1 0.084952f
C33 VGND VNB 0.959908f
C34 X VNB 0.051131f
C35 VPWR VNB 0.729428f
C36 A1 VNB 0.174068f
C37 A2 VNB 0.444184f
C38 C1 VNB 0.203139f
C39 B1 VNB 0.211085f
C40 VPB VNB 1.69186f
C41 a_517_392# VNB 0.040366f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a211o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a211o_2 VNB VPB VPWR VGND C1 B1 A2 A1 X
X0 a_85_270.t1 C1.t0 a_600_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t1 A2.t0 a_317_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.275 ps=2.55 w=1 l=0.15
X2 X.t3 a_85_270.t4 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X3 a_85_270.t0 A1.t0 a_399_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X4 a_600_392.t1 B1.t0 a_317_392.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X5 a_317_392.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X6 a_399_74.t0 A2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.2442 ps=1.4 w=0.74 l=0.15
X7 X.t0 a_85_270.t5 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X8 VGND.t2 B1.t1 a_85_270.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X9 a_85_270.t2 C1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X10 VPWR.t3 a_85_270.t6 X.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VGND.t3 a_85_270.t7 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2442 pd=1.4 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 C1.n0 C1.t1 245.821
R1 C1.n0 C1.t0 230.966
R2 C1 C1.n0 154.133
R3 a_600_392.t0 a_600_392.t1 53.1905
R4 a_85_270.t1 a_85_270.n5 424.026
R5 a_85_270.n2 a_85_270.t4 319.192
R6 a_85_270.n4 a_85_270.t6 244.097
R7 a_85_270.n1 a_85_270.t2 210.512
R8 a_85_270.n3 a_85_270.t7 203.873
R9 a_85_270.n2 a_85_270.t5 196.013
R10 a_85_270.n5 a_85_270.n4 152
R11 a_85_270.n5 a_85_270.n1 107.294
R12 a_85_270.n1 a_85_270.n0 98.6841
R13 a_85_270.n3 a_85_270.n2 62.6605
R14 a_85_270.n0 a_85_270.t3 37.2978
R15 a_85_270.n0 a_85_270.t0 25.9464
R16 a_85_270.n4 a_85_270.n3 9.43093
R17 VPB.t3 VPB.t2 495.43
R18 VPB.t2 VPB.t0 275.807
R19 VPB VPB.t4 263.038
R20 VPB.t0 VPB.t5 229.839
R21 VPB.t4 VPB.t3 229.839
R22 VPB.t5 VPB.t1 214.517
R23 A2.n0 A2.t0 288.933
R24 A2.n0 A2.t1 184.768
R25 A2 A2.n0 158.012
R26 a_317_392.n0 a_317_392.t1 677.351
R27 a_317_392.n0 a_317_392.t2 29.5505
R28 a_317_392.t0 a_317_392.n0 29.5505
R29 VPWR.n2 VPWR.n1 613.919
R30 VPWR.n3 VPWR.t3 342.31
R31 VPWR.n5 VPWR.t2 259.171
R32 VPWR.n1 VPWR.t0 43.3405
R33 VPWR.n1 VPWR.t1 33.4905
R34 VPWR.n5 VPWR.n4 25.977
R35 VPWR.n4 VPWR.n3 22.9652
R36 VPWR.n4 VPWR.n0 9.3005
R37 VPWR.n6 VPWR.n5 9.3005
R38 VPWR.n3 VPWR.n2 6.85679
R39 VPWR.n2 VPWR.n0 0.474531
R40 VPWR.n6 VPWR.n0 0.122949
R41 VPWR VPWR.n6 0.0617245
R42 X.n2 X 591.154
R43 X.n2 X.n0 585
R44 X.n3 X.n2 585
R45 X X.n1 119.433
R46 X.n2 X.t2 26.3844
R47 X.n2 X.t3 26.3844
R48 X.n1 X.t1 22.7032
R49 X.n1 X.t0 22.7032
R50 X X.n3 16.4928
R51 X X.n0 14.2774
R52 X X.n0 3.93896
R53 X.n3 X 1.72358
R54 A1.n0 A1.t1 295.36
R55 A1.n0 A1.t0 191.194
R56 A1 A1.n0 159.262
R57 a_399_74.t0 a_399_74.t1 34.0546
R58 VNB.t2 VNB.t0 1870.87
R59 VNB VNB.t3 1570.6
R60 VNB.t4 VNB.t1 1247.24
R61 VNB.t5 VNB.t4 1247.24
R62 VNB.t3 VNB.t2 993.177
R63 VNB.t0 VNB.t5 831.496
R64 B1.n0 B1.t0 287.861
R65 B1.n0 B1.t1 191.194
R66 B1 B1.n0 156.049
R67 VGND.n8 VGND.t4 273.74
R68 VGND.n4 VGND.n3 223.183
R69 VGND.n2 VGND.n1 104.704
R70 VGND.n1 VGND.t0 50.0805
R71 VGND.n1 VGND.t3 48.392
R72 VGND.n4 VGND.n2 40.2962
R73 VGND.n7 VGND.n6 36.1417
R74 VGND.n3 VGND.t1 31.6221
R75 VGND.n3 VGND.t2 31.6221
R76 VGND.n9 VGND.n8 13.8181
R77 VGND.n6 VGND.n5 9.3005
R78 VGND.n7 VGND.n0 9.3005
R79 VGND.n8 VGND.n7 6.77697
R80 VGND.n6 VGND.n2 3.38874
R81 VGND.n5 VGND.n4 0.256617
R82 VGND.n5 VGND.n0 0.122949
R83 VGND.n9 VGND.n0 0.122949
R84 VGND VGND.n9 0.0617245
C0 C1 X 6.15e-20
C1 B1 VGND 0.017634f
C2 C1 VGND 0.015788f
C3 VPWR X 0.180391f
C4 VPB A2 0.055287f
C5 VPWR VGND 0.071353f
C6 VPB A1 0.041999f
C7 X VGND 0.108456f
C8 A2 A1 0.117241f
C9 VPB B1 0.037961f
C10 VPB C1 0.051998f
C11 A1 B1 0.102606f
C12 VPB VPWR 0.123977f
C13 A2 VPWR 0.015603f
C14 VPB X 0.006341f
C15 B1 C1 0.101315f
C16 A1 VPWR 0.014785f
C17 A2 X 7.61e-19
C18 VPB VGND 0.009663f
C19 B1 VPWR 0.011221f
C20 A1 X 2.98e-19
C21 A2 VGND 0.017796f
C22 C1 VPWR 0.010983f
C23 A1 VGND 0.012111f
C24 B1 X 9.62e-20
C25 VGND VNB 0.518965f
C26 X VNB 0.04416f
C27 VPWR VNB 0.431871f
C28 C1 VNB 0.161345f
C29 B1 VNB 0.114238f
C30 A1 VNB 0.106733f
C31 A2 VNB 0.121913f
C32 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a211o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a211o_1 VNB VPB VPWR VGND X C1 B1 A2 A1
X0 a_366_136.t1 A2.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.156425 ps=1.35 w=0.64 l=0.15
X1 VGND.t0 B1.t0 a_81_264.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 a_81_264.t1 C1.t0 a_550_392.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.12 ps=1.24 w=1 l=0.15
X3 VGND.t2 a_81_264.t4 X.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.156425 pd=1.35 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 VPWR.t2 a_81_264.t5 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X5 a_550_392.t1 B1.t1 a_279_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.15 ps=1.3 w=1 l=0.15
X6 a_279_392.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR.t1 A2.t1 a_279_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.275 ps=2.55 w=1 l=0.15
X8 a_81_264.t3 C1.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.112 ps=0.99 w=0.64 l=0.15
X9 a_81_264.t0 A1.t1 a_366_136.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.104 ps=0.965 w=0.64 l=0.15
R0 A2.n0 A2.t1 236.983
R1 A2.n0 A2.t0 168.701
R2 A2 A2.n0 154.91
R3 VGND.n2 VGND.n1 255.684
R4 VGND.n2 VGND.n0 105.8
R5 VGND.n0 VGND.t1 43.4035
R6 VGND.n1 VGND.t0 39.3755
R7 VGND.n0 VGND.t2 37.6988
R8 VGND.n1 VGND.t3 26.2505
R9 VGND VGND.n2 0.41417
R10 a_366_136.t0 a_366_136.t1 60.938
R11 VNB VNB.t3 2783.2
R12 VNB.t3 VNB.t2 1270.34
R13 VNB.t1 VNB.t4 1154.86
R14 VNB.t2 VNB.t0 1097.11
R15 VNB.t0 VNB.t1 993.177
R16 B1.t0 B1.t1 442.904
R17 B1.n0 B1.t0 336.623
R18 B1 B1.n0 5.56572
R19 B1.n0 B1 3.45447
R20 a_81_264.n0 a_81_264.t5 282.373
R21 a_81_264.n3 a_81_264.t3 262.291
R22 a_81_264.t1 a_81_264.n3 259.06
R23 a_81_264.n0 a_81_264.t4 228.119
R24 a_81_264.n2 a_81_264.n1 185
R25 a_81_264.n2 a_81_264.n0 163.087
R26 a_81_264.n3 a_81_264.n2 37.7605
R27 a_81_264.n1 a_81_264.t2 26.2505
R28 a_81_264.n1 a_81_264.t0 26.2505
R29 C1.t1 C1.t0 430.546
R30 C1 C1.t1 349.659
R31 a_550_392.t0 a_550_392.t1 47.2805
R32 VPB.t3 VPB.t1 638.442
R33 VPB VPB.t3 252.823
R34 VPB.t1 VPB.t0 245.161
R35 VPB.t0 VPB.t4 229.839
R36 VPB.t4 VPB.t2 199.195
R37 X.n1 X 589.572
R38 X.n1 X.n0 585
R39 X.n2 X.n1 585
R40 X X.t0 215.255
R41 X.n1 X.t1 26.3844
R42 X X.n2 12.2519
R43 X X.n0 10.6062
R44 X X.n0 2.92621
R45 X.n2 X 1.2805
R46 VPWR.n1 VPWR.n0 339.714
R47 VPWR.n1 VPWR.t2 265.082
R48 VPWR.n0 VPWR.t0 32.5055
R49 VPWR.n0 VPWR.t1 32.5055
R50 VPWR VPWR.n1 0.304779
R51 a_279_392.n0 a_279_392.t1 485.7
R52 a_279_392.n0 a_279_392.t2 29.5505
R53 a_279_392.t0 a_279_392.n0 29.5505
R54 A1.n0 A1.t0 236.983
R55 A1.n0 A1.t1 168.701
R56 A1.n1 A1.n0 152
R57 A1 A1.n1 13.3823
R58 A1.n1 A1 5.23686
C0 X VGND 0.141537f
C1 X A2 0.003602f
C2 X A1 1.13e-19
C3 VPWR VPB 0.133752f
C4 X B1 3.16e-19
C5 VPWR VGND 0.061649f
C6 VGND VPB 0.012763f
C7 VPWR A2 0.015927f
C8 VPB A2 0.04998f
C9 X C1 1.3e-20
C10 VGND A2 0.01286f
C11 VPWR A1 0.017941f
C12 VPB A1 0.041018f
C13 VPWR B1 0.007499f
C14 VGND A1 0.007403f
C15 A2 A1 0.077525f
C16 VPB B1 0.028646f
C17 VGND B1 0.164824f
C18 VPWR C1 0.009963f
C19 VPB C1 0.045258f
C20 A2 B1 0.001048f
C21 VGND C1 0.099637f
C22 A1 B1 0.079133f
C23 A1 C1 0.00235f
C24 B1 C1 0.0846f
C25 X VPWR 0.130021f
C26 X VPB 0.016321f
C27 VGND VNB 0.500601f
C28 VPWR VNB 0.397225f
C29 X VNB 0.142495f
C30 C1 VNB 0.219773f
C31 B1 VNB 0.135276f
C32 A1 VNB 0.089858f
C33 A2 VNB 0.095192f
C34 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a221oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221oi_2 VNB VPB VPWR VGND Y B2 B1 A2 A1 C1
X0 a_675_74.t1 A2.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1 a_29_368.t5 B1.t0 a_294_368.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_294_368.t1 B2.t0 a_29_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VGND.t5 C1.t0 Y.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 a_293_74.t3 B1.t1 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_294_368.t6 B1.t2 a_29_368.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_29_368.t1 B2.t1 a_294_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1848 ps=1.45 w=1.12 l=0.15
X7 a_29_368.t3 C1.t1 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 Y.t5 B1.t3 a_293_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VGND.t2 A2.t1 a_675_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2479 ps=1.41 w=0.74 l=0.15
X10 a_294_368.t5 A2.t2 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t0 A1.t0 a_294_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VPWR.t2 A2.t3 a_294_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 Y.t0 C1.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.111 ps=1.04 w=0.74 l=0.15
X14 a_294_368.t3 A1.t1 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X15 VGND.t1 B2.t2 a_293_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1184 ps=1.06 w=0.74 l=0.15
X16 a_293_74.t0 B2.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1443 ps=1.13 w=0.74 l=0.15
X17 Y.t2 C1.t3 a_29_368.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X18 a_675_74.t3 A1.t2 Y.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2479 pd=1.41 as=0.1184 ps=1.06 w=0.74 l=0.15
X19 Y.t6 A1.t3 a_675_74.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A2.n0 A2.t2 230.459
R1 A2.n1 A2.t3 226.809
R2 A2.n1 A2.t1 206.969
R3 A2.n0 A2.t0 196.013
R4 A2.n3 A2.n2 152
R5 A2.n2 A2.n0 59.8853
R6 A2 A2.n3 9.69193
R7 A2.n3 A2 7.86336
R8 A2.n2 A2.n1 2.19141
R9 VGND.n4 VGND.n3 210.917
R10 VGND.n9 VGND.n8 209.686
R11 VGND.n2 VGND.n1 203.636
R12 VGND.n7 VGND.n6 36.1417
R13 VGND.n1 VGND.t4 34.8654
R14 VGND.n3 VGND.t3 29.1897
R15 VGND.n1 VGND.t1 28.3789
R16 VGND.n3 VGND.t2 27.5681
R17 VGND.n8 VGND.t0 24.3248
R18 VGND.n8 VGND.t5 24.3248
R19 VGND.n9 VGND.n7 21.8358
R20 VGND.n6 VGND.n2 19.577
R21 VGND.n6 VGND.n5 9.3005
R22 VGND.n7 VGND.n0 9.3005
R23 VGND.n4 VGND.n2 7.30931
R24 VGND.n10 VGND.n9 7.25439
R25 VGND.n5 VGND.n4 0.158565
R26 VGND VGND.n10 0.157727
R27 VGND.n10 VGND.n0 0.150046
R28 VGND.n5 VGND.n0 0.122949
R29 a_675_74.n1 a_675_74.n0 185.53
R30 a_675_74.n0 a_675_74.t3 47.5771
R31 a_675_74.n0 a_675_74.t0 45.4926
R32 a_675_74.n1 a_675_74.t2 22.7032
R33 a_675_74.t1 a_675_74.n1 22.7032
R34 VNB.t9 VNB.t2 1893.96
R35 VNB.t1 VNB.t4 1247.24
R36 VNB VNB.t7 1177.95
R37 VNB.t2 VNB.t3 1154.86
R38 VNB.t6 VNB.t9 1085.56
R39 VNB.t5 VNB.t1 1085.56
R40 VNB.t7 VNB.t0 1039.37
R41 VNB.t3 VNB.t8 993.177
R42 VNB.t4 VNB.t6 993.177
R43 VNB.t0 VNB.t5 993.177
R44 B1 B1.n1 255.462
R45 B1.n1 B1.t2 250.909
R46 B1.n0 B1.t0 250.909
R47 B1.n1 B1.t1 220.113
R48 B1.n0 B1.t3 220.113
R49 B1.n2 B1.n0 153.358
R50 B1.n2 B1 6.62506
R51 B1 B1.n2 4.15489
R52 a_294_368.n2 a_294_368.n0 645.519
R53 a_294_368.n2 a_294_368.n1 585
R54 a_294_368.n5 a_294_368.n4 340.063
R55 a_294_368.n4 a_294_368.n3 297.147
R56 a_294_368.n4 a_294_368.n2 94.4946
R57 a_294_368.n0 a_294_368.t2 29.0228
R58 a_294_368.n0 a_294_368.t6 29.0228
R59 a_294_368.n1 a_294_368.t7 26.3844
R60 a_294_368.n1 a_294_368.t1 26.3844
R61 a_294_368.n3 a_294_368.t4 26.3844
R62 a_294_368.n3 a_294_368.t3 26.3844
R63 a_294_368.t0 a_294_368.n5 26.3844
R64 a_294_368.n5 a_294_368.t5 26.3844
R65 a_29_368.n1 a_29_368.t5 906.754
R66 a_29_368.n1 a_29_368.n0 585
R67 a_29_368.n2 a_29_368.t2 393.745
R68 a_29_368.n3 a_29_368.n2 217.744
R69 a_29_368.n2 a_29_368.n1 66.069
R70 a_29_368.n0 a_29_368.t0 26.3844
R71 a_29_368.n0 a_29_368.t1 26.3844
R72 a_29_368.t4 a_29_368.n3 26.3844
R73 a_29_368.n3 a_29_368.t3 26.3844
R74 VPB.t9 VPB.t3 495.43
R75 VPB VPB.t6 252.823
R76 VPB.t8 VPB.t2 245.161
R77 VPB.t5 VPB.t0 229.839
R78 VPB.t4 VPB.t5 229.839
R79 VPB.t3 VPB.t4 229.839
R80 VPB.t1 VPB.t9 229.839
R81 VPB.t2 VPB.t1 229.839
R82 VPB.t7 VPB.t8 229.839
R83 VPB.t6 VPB.t7 229.839
R84 B2.n0 B2.t0 226.809
R85 B2.n1 B2.t1 226.809
R86 B2.n0 B2.t3 210.138
R87 B2.n1 B2.t2 198.204
R88 B2 B2.n2 154.522
R89 B2.n2 B2.n1 34.3247
R90 B2.n2 B2.n0 31.4035
R91 C1.n1 C1.t3 229
R92 C1.n0 C1.t1 226.809
R93 C1.n0 C1.t2 198.204
R94 C1.n1 C1.t0 196.013
R95 C1 C1.n2 155.423
R96 C1.n2 C1.n1 35.055
R97 C1.n2 C1.n0 28.4823
R98 Y Y.n0 334.772
R99 Y.n2 Y.t6 310.322
R100 Y.n5 Y.t1 155.404
R101 Y.n4 Y.n2 133.272
R102 Y.n2 Y.n1 110.052
R103 Y.n4 Y.n3 110.049
R104 Y.n5 Y.n4 53.4593
R105 Y.n1 Y.t7 29.1897
R106 Y.n0 Y.t3 26.3844
R107 Y.n0 Y.t2 26.3844
R108 Y.n3 Y.t4 22.7032
R109 Y.n3 Y.t0 22.7032
R110 Y.n1 Y.t5 22.7032
R111 Y Y.n5 5.77305
R112 a_293_74.n1 a_293_74.n0 242.569
R113 a_293_74.t1 a_293_74.n1 29.1897
R114 a_293_74.n0 a_293_74.t2 22.7032
R115 a_293_74.n0 a_293_74.t0 22.7032
R116 a_293_74.n1 a_293_74.t3 22.7032
R117 VPWR.n5 VPWR.t1 902.008
R118 VPWR.n3 VPWR.n1 618.13
R119 VPWR.n2 VPWR.t0 264.808
R120 VPWR.n5 VPWR.n4 35.7652
R121 VPWR.n1 VPWR.t3 26.3844
R122 VPWR.n1 VPWR.t2 26.3844
R123 VPWR.n4 VPWR.n3 25.6005
R124 VPWR.n3 VPWR.n2 17.6203
R125 VPWR.n4 VPWR.n0 9.3005
R126 VPWR.n6 VPWR.n5 6.77534
R127 VPWR VPWR.n6 0.882589
R128 VPWR.n2 VPWR.n0 0.696784
R129 VPWR.n6 VPWR.n0 0.163268
R130 A1.n1 A1.n0 278.712
R131 A1.n0 A1.t1 252.369
R132 A1.n2 A1.t0 250.909
R133 A1.n0 A1.t2 235.451
R134 A1.n2 A1.t3 220.113
R135 A1.n3 A1.n2 152
R136 A1 A1.n3 10.7891
R137 A1.n3 A1.n1 5.85193
R138 A1.n1 A1 0.914786
C0 VPB C1 0.063358f
C1 A1 VGND 0.025364f
C2 A2 VPWR 0.024693f
C3 VPB B1 0.076837f
C4 A2 VGND 0.023568f
C5 Y VPWR 0.017143f
C6 VPB B2 0.062107f
C7 C1 B1 0.083603f
C8 Y VGND 0.262952f
C9 C1 B2 5.81e-19
C10 VPB A1 0.098924f
C11 VPWR VGND 0.090508f
C12 VPB A2 0.063144f
C13 C1 A1 1.47e-19
C14 B1 B2 0.212969f
C15 VPB Y 0.010874f
C16 B1 A1 0.106825f
C17 C1 A2 7.9e-20
C18 VPB VPWR 0.155468f
C19 C1 Y 0.162209f
C20 C1 VPWR 0.012058f
C21 B1 Y 0.133669f
C22 VPB VGND 0.009576f
C23 C1 VGND 0.035711f
C24 B1 VPWR 0.018363f
C25 B2 Y 0.054732f
C26 A1 A2 0.238017f
C27 B2 VPWR 0.011311f
C28 A1 Y 0.127982f
C29 B1 VGND 0.02379f
C30 A1 VPWR 0.091205f
C31 A2 Y 0.081066f
C32 B2 VGND 0.026828f
C33 VGND VNB 0.691627f
C34 VPWR VNB 0.583876f
C35 Y VNB 0.174685f
C36 A2 VNB 0.200166f
C37 A1 VNB 0.292136f
C38 B2 VNB 0.195649f
C39 B1 VNB 0.206883f
C40 C1 VNB 0.219981f
C41 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a222o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a222o_1 VNB VPB VPWR VGND C2 X C1 B2 A2 A1 B1
X0 a_337_390.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.345 ps=2.69 w=1 l=0.15
X1 a_32_74.t4 B1.t0 a_386_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2512 pd=1.425 as=0.0768 ps=0.88 w=0.64 l=0.15
X2 a_119_74.t1 C1.t0 a_32_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X3 a_27_390.t3 B1.t1 a_337_390.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.22 ps=1.44 w=1 l=0.15
X4 X.t1 a_32_74.t5 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1997 ps=1.325 w=0.74 l=0.15
X5 VGND.t0 C2.t0 a_119_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2544 pd=1.435 as=0.0768 ps=0.88 w=0.64 l=0.15
X6 a_337_390.t2 B2.t0 a_27_390.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X7 a_32_74.t2 C1.t1 a_27_390.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2275 pd=1.455 as=0.295 ps=2.59 w=1 l=0.15
X8 VGND.t2 A2.t0 a_651_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1997 pd=1.325 as=0.0768 ps=0.88 w=0.64 l=0.15
X9 a_651_74.t0 A1.t1 a_32_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2512 ps=1.425 w=0.64 l=0.15
X10 a_386_74.t1 B2.t1 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2544 ps=1.435 w=0.64 l=0.15
X11 a_27_390.t1 C2.t1 a_32_74.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.2275 ps=1.455 w=1 l=0.15
X12 X.t0 a_32_74.t6 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2352 ps=1.555 w=1.12 l=0.15
X13 VPWR.t1 A2.t1 a_337_390.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.555 as=0.15 ps=1.3 w=1 l=0.15
R0 A1.n0 A1.t0 315.498
R1 A1.n0 A1.t1 162.274
R2 A1 A1.n0 154.91
R3 VPWR.n1 VPWR.t0 362.728
R4 VPWR.n1 VPWR.n0 228.732
R5 VPWR.n0 VPWR.t1 46.2955
R6 VPWR.n0 VPWR.t2 34.3111
R7 VPWR VPWR.n1 1.04253
R8 a_337_390.n1 a_337_390.n0 597.667
R9 a_337_390.n0 a_337_390.t1 47.2805
R10 a_337_390.n0 a_337_390.t2 39.4005
R11 a_337_390.n1 a_337_390.t3 29.5505
R12 a_337_390.t0 a_337_390.n1 29.5505
R13 VPB.t2 VPB.t0 541.399
R14 VPB.t1 VPB.t3 309.005
R15 VPB.t4 VPB.t2 301.344
R16 VPB.t5 VPB.t6 298.791
R17 VPB VPB.t1 257.93
R18 VPB.t3 VPB.t4 255.376
R19 VPB.t0 VPB.t5 229.839
R20 B1.n0 B1.t1 338.248
R21 B1.n0 B1.t0 157.571
R22 B1.n1 B1.n0 152
R23 B1.n1 B1 7.05844
R24 B1 B1.n1 1.79489
R25 a_386_74.t0 a_386_74.t1 45.0005
R26 a_32_74.n6 a_32_74.n5 377.224
R27 a_32_74.n0 a_32_74.t6 263.25
R28 a_32_74.n1 a_32_74.n0 260.745
R29 a_32_74.n0 a_32_74.t5 203
R30 a_32_74.n5 a_32_74.t0 157.055
R31 a_32_74.n5 a_32_74.n4 115.596
R32 a_32_74.n3 a_32_74.n2 94.688
R33 a_32_74.n4 a_32_74.n3 92.5005
R34 a_32_74.n2 a_32_74.n1 92.5005
R35 a_32_74.t2 a_32_74.n6 60.0855
R36 a_32_74.n6 a_32_74.t3 29.5505
R37 a_32_74.n2 a_32_74.t1 26.2505
R38 a_32_74.n3 a_32_74.t4 26.2505
R39 a_32_74.n4 a_32_74.n1 10.4263
R40 VNB.t0 VNB.t6 2182.68
R41 VNB.t5 VNB.t2 2159.58
R42 VNB.t4 VNB.t3 1697.64
R43 VNB VNB.t1 1201.05
R44 VNB.t2 VNB.t4 900.788
R45 VNB.t6 VNB.t5 900.788
R46 VNB.t1 VNB.t0 900.788
R47 C1.n0 C1.t1 319.781
R48 C1.n0 C1.t0 159.381
R49 C1.n1 C1.n0 152
R50 C1.n1 C1 8.88521
R51 C1 C1.n1 2.25932
R52 a_119_74.t0 a_119_74.t1 45.0005
R53 a_27_390.n1 a_27_390.t3 385.947
R54 a_27_390.t0 a_27_390.n1 297.257
R55 a_27_390.n1 a_27_390.n0 209.663
R56 a_27_390.n0 a_27_390.t1 39.4005
R57 a_27_390.n0 a_27_390.t2 29.5505
R58 VGND.n2 VGND.n1 191.651
R59 VGND.n5 VGND.n4 185
R60 VGND.n3 VGND.n0 185
R61 VGND.n4 VGND.n3 96.563
R62 VGND.n1 VGND.t1 58.2861
R63 VGND.n1 VGND.t2 47.813
R64 VGND.n8 VGND.n0 28.8576
R65 VGND.n4 VGND.t3 26.2505
R66 VGND.n3 VGND.t0 26.2505
R67 VGND.n7 VGND.n6 9.3005
R68 VGND.n6 VGND.n5 8.2224
R69 VGND.n5 VGND.n2 8.14073
R70 VGND.n6 VGND.n0 1.40196
R71 VGND VGND.n8 0.163644
R72 VGND.n7 VGND.n2 0.157634
R73 VGND.n8 VGND.n7 0.144205
R74 X.n1 X 589.508
R75 X.n1 X.n0 585
R76 X.n2 X.n1 585
R77 X X.t1 206.401
R78 X.n1 X.t0 26.3844
R79 X X.n2 12.0794
R80 X X.n0 10.4568
R81 X X.n0 2.88501
R82 X.n2 X 1.26247
R83 C2.n0 C2.t1 320.067
R84 C2.n0 C2.t0 185.244
R85 C2 C2.n0 154.201
R86 B2.n0 B2.t0 307.514
R87 B2.n0 B2.t1 181.554
R88 B2 B2.n0 155.752
R89 A2.n0 A2.t1 313.3
R90 A2.n0 A2.t0 162.274
R91 A2 A2.n0 156.368
R92 a_651_74.t0 a_651_74.t1 45.0005
C0 B1 VPWR 0.007614f
C1 B2 X 4.53e-20
C2 C2 VGND 0.019015f
C3 A1 A2 0.096463f
C4 VPB C1 0.04706f
C5 B2 VGND 0.01709f
C6 A1 VPWR 0.018103f
C7 B1 X 0.002198f
C8 VPB C2 0.045477f
C9 B1 VGND 0.012295f
C10 A1 X 7.36e-19
C11 A2 VPWR 0.023331f
C12 C1 C2 0.055985f
C13 VPB B2 0.044378f
C14 A1 VGND 0.009917f
C15 A2 X 0.002146f
C16 VPB B1 0.053903f
C17 A2 VGND 0.014302f
C18 VPWR X 0.130601f
C19 VPB A1 0.045639f
C20 C2 B2 0.105326f
C21 VPWR VGND 0.076653f
C22 C2 B1 0.001733f
C23 VPB A2 0.037569f
C24 X VGND 0.063974f
C25 VPB VPWR 0.127057f
C26 B2 B1 0.106466f
C27 C1 VPWR 0.006703f
C28 VPB X 0.017126f
C29 B1 A1 0.068334f
C30 VPB VGND 0.010465f
C31 C2 VPWR 0.006563f
C32 C2 X 2.88e-20
C33 C1 VGND 0.01313f
C34 B2 VPWR 0.006276f
C35 B1 A2 0.001383f
C36 VGND VNB 0.586542f
C37 X VNB 0.111955f
C38 VPWR VNB 0.464313f
C39 A2 VNB 0.119879f
C40 A1 VNB 0.127371f
C41 B1 VNB 0.139059f
C42 B2 VNB 0.121485f
C43 C2 VNB 0.143635f
C44 C1 VNB 0.18534f
C45 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a222o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a222o_2 VNB VPB VPWR VGND X C1 B2 B1 A2 C2 A1
X0 X.t3 a_27_82.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2077 ps=1.35 w=0.74 l=0.15
X1 a_116_392.t3 C1.t0 a_27_82.t1 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X2 VPWR.t2 a_27_82.t6 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2665 pd=1.65 as=0.168 ps=1.42 w=1.12 l=0.15
X3 a_114_82.t1 C1.t1 a_27_82.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X4 X.t0 a_27_82.t7 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.34065 ps=3.12 w=1.12 l=0.15
X5 a_639_368.t3 A1.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.28175 pd=1.685 as=0.2665 ps=1.65 w=1 l=0.15
X6 VGND.t3 C2.t0 a_114_82.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.2077 pd=1.35 as=0.0768 ps=0.88 w=0.64 l=0.15
X7 a_775_74.t1 B1.t0 a_27_82.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1504 ps=1.11 w=0.64 l=0.15
X8 a_639_368.t2 B2.t0 a_116_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X9 a_27_82.t4 A1.t1 a_557_74.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1504 pd=1.11 as=0.1971 ps=1.92 w=0.64 l=0.15
X10 a_116_392.t0 B1.t1 a_639_368.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.28175 ps=1.685 w=1 l=0.15
X11 a_27_82.t3 C2.t1 a_116_392.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X12 VGND.t1 a_27_82.t8 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2586 pd=2.67 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_557_74.t1 A2.t0 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1344 ps=1.06 w=0.64 l=0.15
X14 VPWR.t0 A2.t1 a_639_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.2 ps=1.4 w=1 l=0.15
X15 VGND.t0 B2.t1 a_775_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1344 pd=1.06 as=0.0768 ps=0.88 w=0.64 l=0.15
R0 a_27_82.n6 a_27_82.t3 815.39
R1 a_27_82.t1 a_27_82.n6 279.334
R2 a_27_82.n1 a_27_82.t5 268.606
R3 a_27_82.n3 a_27_82.t6 264.053
R4 a_27_82.n1 a_27_82.t7 250.909
R5 a_27_82.n4 a_27_82.n0 244.482
R6 a_27_82.n5 a_27_82.t2 219.734
R7 a_27_82.n4 a_27_82.n3 164.8
R8 a_27_82.n2 a_27_82.t8 154.24
R9 a_27_82.n5 a_27_82.n4 101.556
R10 a_27_82.n6 a_27_82.n5 78.0654
R11 a_27_82.n0 a_27_82.t4 46.8755
R12 a_27_82.n3 a_27_82.n2 46.7399
R13 a_27_82.n0 a_27_82.t0 41.2505
R14 a_27_82.n2 a_27_82.n1 3.65202
R15 VGND.n3 VGND.t1 300.387
R16 VGND.n5 VGND.n4 215.641
R17 VGND.n1 VGND.n0 214.185
R18 VGND.n0 VGND.t2 84.5361
R19 VGND.n4 VGND.t4 48.7505
R20 VGND.n8 VGND.n7 36.1417
R21 VGND.n9 VGND.n8 36.1417
R22 VGND.n4 VGND.t0 30.0005
R23 VGND.n0 VGND.t3 26.2505
R24 VGND.n11 VGND.n1 23.892
R25 VGND.n5 VGND.n3 19.8102
R26 VGND.n7 VGND.n6 9.3005
R27 VGND.n8 VGND.n2 9.3005
R28 VGND.n10 VGND.n9 9.3005
R29 VGND.n7 VGND.n3 7.6554
R30 VGND.n9 VGND.n1 1.12991
R31 VGND VGND.n11 0.163644
R32 VGND.n6 VGND.n5 0.162238
R33 VGND.n11 VGND.n10 0.144205
R34 VGND.n6 VGND.n2 0.122949
R35 VGND.n10 VGND.n2 0.122949
R36 X X.n0 591.737
R37 X X.n1 223.855
R38 X.n0 X.t1 26.3844
R39 X.n0 X.t0 26.3844
R40 X.n1 X.t2 22.7032
R41 X.n1 X.t3 22.7032
R42 VNB.t1 VNB.t6 2552.23
R43 VNB.t3 VNB.t2 1755.38
R44 VNB.t6 VNB.t4 1432.02
R45 VNB.t0 VNB.t7 1316.54
R46 VNB VNB.t5 1143.31
R47 VNB.t2 VNB.t1 993.177
R48 VNB.t4 VNB.t0 900.788
R49 VNB.t5 VNB.t3 900.788
R50 C1.n0 C1.t0 280.604
R51 C1.n0 C1.t1 200.263
R52 C1 C1.n0 155.067
R53 a_116_392.n1 a_116_392.n0 814.213
R54 a_116_392.n0 a_116_392.t2 29.5505
R55 a_116_392.n0 a_116_392.t3 29.5505
R56 a_116_392.n1 a_116_392.t1 29.5505
R57 a_116_392.t0 a_116_392.n1 29.5505
R58 VPB.t5 VPB.t1 559.274
R59 VPB.t6 VPB.t3 334.543
R60 VPB.t2 VPB.t6 316.668
R61 VPB.t4 VPB.t0 280.914
R62 VPB VPB.t7 257.93
R63 VPB.t3 VPB.t4 229.839
R64 VPB.t1 VPB.t2 229.839
R65 VPB.t7 VPB.t5 229.839
R66 VPWR.n7 VPWR.t1 778.611
R67 VPWR.n2 VPWR.n1 620.793
R68 VPWR.n3 VPWR.t0 426.325
R69 VPWR.n1 VPWR.t3 55.1605
R70 VPWR.n6 VPWR.n5 36.1417
R71 VPWR.n1 VPWR.t2 32.1543
R72 VPWR.n7 VPWR.n6 19.2005
R73 VPWR.n3 VPWR.n2 18.5562
R74 VPWR.n5 VPWR.n4 9.3005
R75 VPWR.n6 VPWR.n0 9.3005
R76 VPWR.n8 VPWR.n7 7.36287
R77 VPWR VPWR.n8 0.400061
R78 VPWR.n5 VPWR.n2 0.376971
R79 VPWR.n4 VPWR.n3 0.161319
R80 VPWR.n8 VPWR.n0 0.153815
R81 VPWR.n4 VPWR.n0 0.122949
R82 a_114_82.t0 a_114_82.t1 45.0005
R83 A1.n0 A1.t1 236.18
R84 A1.n0 A1.t0 231.629
R85 A1 A1.n0 154.522
R86 a_639_368.n1 a_639_368.n0 878.63
R87 a_639_368.n0 a_639_368.t1 50.2355
R88 a_639_368.n0 a_639_368.t3 49.2505
R89 a_639_368.t0 a_639_368.n1 39.4005
R90 a_639_368.n1 a_639_368.t2 39.4005
R91 C2.n0 C2.t1 287.861
R92 C2.n0 C2.t0 194.407
R93 C2 C2.n0 160.369
R94 B1.n0 B1.t0 231.478
R95 B1.n0 B1.t1 226.925
R96 B1 B1.n0 155.423
R97 a_775_74.t0 a_775_74.t1 45.0005
R98 B2.n0 B2.t1 236.18
R99 B2.n0 B2.t0 231.629
R100 B2 B2.n0 160.484
R101 a_557_74.n0 a_557_74.t1 500.353
R102 a_557_74.n0 a_557_74.t0 20.6255
R103 A2.n0 A2.t0 236.18
R104 A2.n0 A2.t1 231.629
R105 A2 A2.n0 155.126
C0 X A1 0.019498f
C1 VPWR B1 0.005747f
C2 VPB VGND 0.010528f
C3 C1 VGND 0.013503f
C4 X B1 5.8e-20
C5 VPWR B2 0.006215f
C6 A1 B1 0.084108f
C7 C2 VGND 0.016684f
C8 VPWR A2 0.052578f
C9 VPB C1 0.051164f
C10 VPWR VGND 0.084736f
C11 A1 B2 3.67e-19
C12 VPB C2 0.049109f
C13 X VGND 0.010627f
C14 A1 A2 1.73e-19
C15 B1 B2 0.10843f
C16 VPB VPWR 0.151437f
C17 C1 C2 0.118646f
C18 A1 VGND 0.007715f
C19 C1 VPWR 0.011068f
C20 VPB X 0.006646f
C21 B1 VGND 0.008301f
C22 B2 A2 0.080938f
C23 C2 VPWR 0.011224f
C24 VPB A1 0.042867f
C25 B2 VGND 0.017515f
C26 C2 X 0.002058f
C27 VPB B1 0.038723f
C28 A2 VGND 0.015929f
C29 VPB B2 0.034286f
C30 VPWR X 0.024741f
C31 C2 A1 8.21e-19
C32 VPB A2 0.039056f
C33 VPWR A1 0.016223f
C34 VGND VNB 0.655878f
C35 A2 VNB 0.163687f
C36 B2 VNB 0.109924f
C37 B1 VNB 0.115921f
C38 A1 VNB 0.128115f
C39 X VNB 0.00653f
C40 VPWR VNB 0.543587f
C41 C2 VNB 0.12315f
C42 C1 VNB 0.174183f
C43 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a222oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a222oi_1 VNB VPB VPWR VGND C2 C1 B1 A2 A1 Y B2
X0 a_369_392.t2 A2.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.225 ps=1.45 w=1 l=0.15
X1 a_697_74.t0 A1.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.2048 ps=1.28 w=0.64 l=0.15
X2 a_116_392.t3 C1.t0 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X3 a_369_392.t3 B1.t0 a_116_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X4 a_119_74.t1 C1.t1 Y.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.1824 ps=1.85 w=0.64 l=0.15
X5 Y.t1 B1.t1 a_461_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2048 pd=1.28 as=0.0768 ps=0.88 w=0.64 l=0.15
X6 a_461_74.t1 B2.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.3744 ps=1.81 w=0.64 l=0.15
X7 VGND.t0 C2.t0 a_119_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3744 pd=1.81 as=0.0768 ps=0.88 w=0.64 l=0.15
X8 Y.t2 C2.t1 a_116_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.175 ps=1.35 w=1 l=0.15
X9 a_116_392.t0 B2.t1 a_369_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.295 ps=2.59 w=1 l=0.15
X10 VGND.t1 A2.t1 a_697_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0768 ps=0.88 w=0.64 l=0.15
X11 VPWR.t0 A1.t1 a_369_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.45 as=0.175 ps=1.35 w=1 l=0.15
R0 A2.n0 A2.t0 301.414
R1 A2.n0 A2.t1 173.685
R2 A2.n1 A2.n0 152
R3 A2 A2.n1 9.11565
R4 A2.n1 A2 5.23686
R5 VPWR VPWR.n0 322.404
R6 VPWR.n0 VPWR.t1 49.2505
R7 VPWR.n0 VPWR.t0 39.4005
R8 a_369_392.t0 a_369_392.n1 379.853
R9 a_369_392.n1 a_369_392.t2 289.146
R10 a_369_392.n1 a_369_392.n0 205.383
R11 a_369_392.n0 a_369_392.t3 39.4005
R12 a_369_392.n0 a_369_392.t1 29.5505
R13 VPB.t1 VPB.t0 618.011
R14 VPB.t2 VPB.t3 306.452
R15 VPB VPB.t5 257.93
R16 VPB.t4 VPB.t2 255.376
R17 VPB.t0 VPB.t4 255.376
R18 VPB.t5 VPB.t1 255.376
R19 A1.n0 A1.t1 232.298
R20 A1.n1 A1.t0 160.266
R21 A1 A1.n0 153.03
R22 A1.n2 A1.n1 152
R23 A1.n1 A1.n0 45.5227
R24 A1 A1.n2 6.74336
R25 A1.n2 A1 1.71479
R26 Y.n1 Y.t2 336.411
R27 Y.n1 Y.t4 285.382
R28 Y.n2 Y.t3 208.256
R29 Y.n2 Y.n0 96.9278
R30 Y.n0 Y.t0 52.2017
R31 Y.n0 Y.t1 50.2717
R32 Y Y.n1 23.8263
R33 Y.n2 Y 14.2457
R34 Y Y.n2 1.03276
R35 a_697_74.t0 a_697_74.t1 45.0005
R36 VNB.t2 VNB.t3 3048.82
R37 VNB.t1 VNB.t0 1824.67
R38 VNB VNB.t5 1201.05
R39 VNB.t0 VNB.t4 900.788
R40 VNB.t3 VNB.t1 900.788
R41 VNB.t5 VNB.t2 900.788
R42 C1.n0 C1.t0 325.351
R43 C1.n0 C1.t1 162.274
R44 C1 C1.n0 157.255
R45 a_116_392.n1 a_116_392.n0 709.193
R46 a_116_392.n0 a_116_392.t3 39.4005
R47 a_116_392.t0 a_116_392.n1 39.4005
R48 a_116_392.n0 a_116_392.t1 29.5505
R49 a_116_392.n1 a_116_392.t2 29.5505
R50 B1.n0 B1.t0 234.306
R51 B1.n1 B1.t1 162.274
R52 B1 B1.n0 153.647
R53 B1.n2 B1.n1 152
R54 B1.n1 B1.n0 49.6611
R55 B1 B1.n2 10.7891
R56 B1.n2 B1 2.74336
R57 a_119_74.t0 a_119_74.t1 45.0005
R58 a_461_74.t0 a_461_74.t1 45.0005
R59 B2.n0 B2.t1 234.306
R60 B2.n1 B2.t0 162.274
R61 B2 B2.n0 153.745
R62 B2.n2 B2.n1 152
R63 B2.n1 B2.n0 49.6611
R64 B2 B2.n2 11.4429
R65 B2.n2 B2 2.90959
R66 VGND.n5 VGND.n4 185
R67 VGND.n8 VGND.n7 185
R68 VGND.n6 VGND.n0 185
R69 VGND.n3 VGND.t1 158.793
R70 VGND.n7 VGND.n5 83.438
R71 VGND.n7 VGND.n6 83.438
R72 VGND.n11 VGND.n0 28.8576
R73 VGND.n5 VGND.t2 26.2505
R74 VGND.n6 VGND.t0 26.2505
R75 VGND.n4 VGND.n3 10.3113
R76 VGND.n10 VGND.n9 9.3005
R77 VGND.n2 VGND.n1 9.3005
R78 VGND.n9 VGND.n8 6.91437
R79 VGND.n4 VGND.n2 6.26035
R80 VGND.n8 VGND.n2 2.05597
R81 VGND.n9 VGND.n0 1.40196
R82 VGND VGND.n11 0.163644
R83 VGND.n3 VGND.n1 0.162785
R84 VGND.n11 VGND.n10 0.144205
R85 VGND.n10 VGND.n1 0.122949
R86 C2.n0 C2.t1 226.774
R87 C2.n1 C2.t0 154.743
R88 C2 C2.n0 153.745
R89 C2.n2 C2.n1 152
R90 C2.n1 C2.n0 34.1422
R91 C2 C2.n2 11.4429
R92 C2.n2 C2 2.90959
C0 C1 VPWR 0.010786f
C1 VPB VGND 0.010661f
C2 B1 A1 0.10468f
C3 C2 Y 0.152496f
C4 B2 Y 0.098789f
C5 C1 VGND 0.012891f
C6 C2 VPWR 0.007113f
C7 A1 A2 0.131692f
C8 B1 Y 0.043576f
C9 C2 VGND 0.0195f
C10 B2 VPWR 0.005954f
C11 VPB C1 0.044063f
C12 B2 VGND 0.015665f
C13 A1 Y 0.026926f
C14 B1 VPWR 0.008489f
C15 VPB C2 0.057708f
C16 A1 VPWR 0.018692f
C17 A2 Y 0.003132f
C18 B1 VGND 0.006441f
C19 C1 C2 0.111646f
C20 VPB B2 0.048566f
C21 A2 VPWR 0.018736f
C22 A1 VGND 0.024619f
C23 VPB B1 0.041227f
C24 Y VPWR 0.057516f
C25 A2 VGND 0.047067f
C26 VPB A1 0.045695f
C27 C2 B2 0.024094f
C28 Y VGND 0.340545f
C29 VPB A2 0.051348f
C30 VPWR VGND 0.068034f
C31 VPB Y 0.040412f
C32 B2 B1 0.122586f
C33 C1 Y 0.110577f
C34 VPB VPWR 0.105152f
C35 VGND VNB 0.562632f
C36 VPWR VNB 0.423604f
C37 Y VNB 0.116221f
C38 A2 VNB 0.188728f
C39 A1 VNB 0.125742f
C40 B1 VNB 0.115962f
C41 B2 VNB 0.125737f
C42 C2 VNB 0.144367f
C43 C1 VNB 0.178671f
C44 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a222oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a222oi_2 VNB VPB VPWR VGND C1 B2 A2 A1 Y C2 B1
X0 a_116_392.t7 B2.t0 a_515_392.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.15 ps=1.3 w=1 l=0.15
X1 a_981_74.t2 A2.t0 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0928 ps=0.93 w=0.64 l=0.15
X2 a_116_392.t1 C2.t0 Y.t8 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X3 a_515_392.t6 B2.t1 a_116_392.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X4 VPWR.t1 A1.t0 a_515_392.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X5 a_515_392.t1 A1.t1 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.15
X6 a_116_392.t0 B1.t0 a_515_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.15
X7 a_515_392.t2 B1.t1 a_116_392.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X8 VPWR.t3 A2.t1 a_515_392.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X9 a_137_74.t1 C1.t0 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X10 a_515_392.t5 A2.t2 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.165 ps=1.33 w=1 l=0.15
X11 a_137_74.t3 C2.t1 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.264125 ps=2.13 w=0.64 l=0.15
X12 a_981_74.t0 A1.t2 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.112 pd=0.99 as=0.0896 ps=0.92 w=0.64 l=0.15
X13 a_593_74.t1 B1.t2 Y.t5 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X14 Y.t6 B1.t3 a_593_74.t0 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X15 VGND.t4 B2.t2 a_593_74.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.19325 pd=1.33 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 Y.t7 C2.t2 a_116_392.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.345 pd=2.69 as=0.15 ps=1.3 w=1 l=0.15
X17 Y.t3 C1.t1 a_116_392.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X18 a_116_392.t2 C1.t2 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.165 ps=1.33 w=1 l=0.15
X19 VGND.t0 C2.t3 a_137_74.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X20 a_593_74.t2 B2.t3 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.19325 ps=1.33 w=0.64 l=0.15
X21 VGND.t1 A2.t3 a_981_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0928 pd=0.93 as=0.112 ps=0.99 w=0.64 l=0.15
X22 Y.t0 C1.t3 a_137_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 B2.n0 B2.t0 263.762
R1 B2.n1 B2.t1 263.762
R2 B2.n1 B2.t2 194.115
R3 B2.n0 B2.t3 164.959
R4 B2 B2.n2 158.012
R5 B2.n2 B2.n0 40.1672
R6 B2.n2 B2.n1 25.5611
R7 a_515_392.n5 a_515_392.n4 585
R8 a_515_392.t0 a_515_392.n5 394.803
R9 a_515_392.n1 a_515_392.n0 298.363
R10 a_515_392.n1 a_515_392.t1 270.767
R11 a_515_392.n3 a_515_392.n2 197.494
R12 a_515_392.n5 a_515_392.n3 107.174
R13 a_515_392.n3 a_515_392.n1 46.5988
R14 a_515_392.n4 a_515_392.t7 29.5505
R15 a_515_392.n4 a_515_392.t6 29.5505
R16 a_515_392.n0 a_515_392.t4 29.5505
R17 a_515_392.n0 a_515_392.t5 29.5505
R18 a_515_392.n2 a_515_392.t3 29.5505
R19 a_515_392.n2 a_515_392.t2 29.5505
R20 a_116_392.n4 a_116_392.n0 620.001
R21 a_116_392.n5 a_116_392.n4 585
R22 a_116_392.n3 a_116_392.n1 347.565
R23 a_116_392.n3 a_116_392.n2 302.389
R24 a_116_392.n4 a_116_392.n3 93.5936
R25 a_116_392.n0 a_116_392.t4 38.4155
R26 a_116_392.n0 a_116_392.t7 38.4155
R27 a_116_392.n1 a_116_392.t3 29.5505
R28 a_116_392.n1 a_116_392.t1 29.5505
R29 a_116_392.n2 a_116_392.t5 29.5505
R30 a_116_392.n2 a_116_392.t2 29.5505
R31 a_116_392.t6 a_116_392.n5 29.5505
R32 a_116_392.n5 a_116_392.t0 29.5505
R33 VPB.t9 VPB.t0 541.399
R34 VPB.t11 VPB.t5 275.807
R35 VPB VPB.t1 257.93
R36 VPB.t6 VPB.t8 245.161
R37 VPB.t4 VPB.t2 245.161
R38 VPB.t7 VPB.t3 229.839
R39 VPB.t8 VPB.t7 229.839
R40 VPB.t5 VPB.t6 229.839
R41 VPB.t10 VPB.t11 229.839
R42 VPB.t0 VPB.t10 229.839
R43 VPB.t2 VPB.t9 229.839
R44 VPB.t1 VPB.t4 229.839
R45 A2.n0 A2.t0 244.945
R46 A2.n1 A2.t3 244.214
R47 A2.n1 A2.t2 215.075
R48 A2.n0 A2.t1 212.883
R49 A2 A2.n2 153.358
R50 A2.n2 A2.n0 43.0884
R51 A2.n2 A2.n1 20.449
R52 VGND.n18 VGND.t3 247.185
R53 VGND.n7 VGND.n4 211.06
R54 VGND.n6 VGND.n5 200.429
R55 VGND.n12 VGND.t0 151.525
R56 VGND.n5 VGND.t5 46.8755
R57 VGND.n5 VGND.t4 46.8755
R58 VGND.n11 VGND.n10 36.1417
R59 VGND.n16 VGND.n1 36.1417
R60 VGND.n17 VGND.n16 36.1417
R61 VGND.n7 VGND.n6 30.7154
R62 VGND.n10 VGND.n3 28.7263
R63 VGND.n4 VGND.t2 27.188
R64 VGND.n4 VGND.t1 27.188
R65 VGND.n12 VGND.n11 27.1064
R66 VGND.n12 VGND.n1 20.3299
R67 VGND.n18 VGND.n17 18.0711
R68 VGND.n19 VGND.n18 9.3005
R69 VGND.n17 VGND.n0 9.3005
R70 VGND.n16 VGND.n15 9.3005
R71 VGND.n14 VGND.n1 9.3005
R72 VGND.n13 VGND.n12 9.3005
R73 VGND.n8 VGND.n3 9.3005
R74 VGND.n10 VGND.n9 9.3005
R75 VGND.n11 VGND.n2 9.3005
R76 VGND.n6 VGND.n3 1.16414
R77 VGND.n8 VGND.n7 0.197101
R78 VGND.n9 VGND.n8 0.122949
R79 VGND.n9 VGND.n2 0.122949
R80 VGND.n13 VGND.n2 0.122949
R81 VGND.n14 VGND.n13 0.122949
R82 VGND.n15 VGND.n14 0.122949
R83 VGND.n15 VGND.n0 0.122949
R84 VGND.n19 VGND.n0 0.122949
R85 VGND VGND.n19 0.0617245
R86 a_981_74.n0 a_981_74.t2 283.264
R87 a_981_74.t1 a_981_74.n0 38.438
R88 a_981_74.n0 a_981_74.t0 27.188
R89 VNB.t1 VNB.t4 2286.61
R90 VNB.t10 VNB.t9 1501.31
R91 VNB VNB.t8 1408.92
R92 VNB.t2 VNB.t5 1154.86
R93 VNB.t5 VNB.t6 1016.27
R94 VNB.t7 VNB.t2 993.177
R95 VNB.t9 VNB.t7 993.177
R96 VNB.t4 VNB.t10 993.177
R97 VNB.t3 VNB.t1 993.177
R98 VNB.t0 VNB.t3 993.177
R99 VNB.t8 VNB.t0 993.177
R100 C2.n1 C2.t0 312.591
R101 C2.n0 C2.t2 252.206
R102 C2.n0 C2.t3 187.85
R103 C2.n1 C2.t1 176.025
R104 C2.n2 C2.n0 164.53
R105 C2.n2 C2.n1 152
R106 C2 C2.n2 3.74684
R107 Y Y.n0 590.715
R108 Y.n9 Y.n0 585
R109 Y.n8 Y.n0 585
R110 Y.n3 Y.t7 336.777
R111 Y Y.n6 335.113
R112 Y.n5 Y.n4 298.291
R113 Y.n2 Y.n1 224.53
R114 Y.n2 Y.t5 138.082
R115 Y.n3 Y.n2 73.3314
R116 Y.n7 Y.n5 52.7064
R117 Y.n5 Y.n3 50.4476
R118 Y.n4 Y.t1 32.5055
R119 Y.n4 Y.t3 32.5055
R120 Y.n0 Y.t8 29.5505
R121 Y.n1 Y.t2 26.2505
R122 Y.n1 Y.t6 26.2505
R123 Y.n6 Y.t4 26.2505
R124 Y.n6 Y.t0 26.2505
R125 Y Y.n9 10.5148
R126 Y Y.n8 9.82907
R127 Y.n9 Y 6.4005
R128 Y.n7 Y 6.4005
R129 Y.n8 Y.n7 0.686214
R130 A1.n2 A1.n1 268.313
R131 A1.n0 A1.t2 268.313
R132 A1.n3 A1.n0 255.358
R133 A1.n2 A1.t1 236.983
R134 A1.n0 A1.t0 236.983
R135 A1.n3 A1.n2 164.412
R136 A1 A1.n3 2.13383
R137 VPWR.n2 VPWR.n1 612.605
R138 VPWR.n2 VPWR.n0 610.403
R139 VPWR.n0 VPWR.t2 32.5055
R140 VPWR.n0 VPWR.t1 32.5055
R141 VPWR.n1 VPWR.t0 29.5505
R142 VPWR.n1 VPWR.t3 29.5505
R143 VPWR VPWR.n2 1.6565
R144 B1.n1 B1.t2 272.733
R145 B1.n0 B1.t3 268.313
R146 B1 B1.n0 264.57
R147 B1.n0 B1.t1 236.983
R148 B1.n1 B1.t0 229.619
R149 B1 B1.n1 159.565
R150 C1.n1 C1.t1 290.808
R151 C1.n0 C1.t2 289.2
R152 C1.n0 C1.t0 157.745
R153 C1 C1.n2 156.655
R154 C1.n1 C1.t3 152.633
R155 C1.n2 C1.n0 38.7066
R156 C1.n2 C1.n1 18.9884
R157 a_137_74.n1 a_137_74.n0 418.065
R158 a_137_74.n0 a_137_74.t0 26.2505
R159 a_137_74.n0 a_137_74.t3 26.2505
R160 a_137_74.n1 a_137_74.t2 26.2505
R161 a_137_74.t1 a_137_74.n1 26.2505
R162 a_593_74.n1 a_593_74.n0 437.031
R163 a_593_74.n0 a_593_74.t0 26.2505
R164 a_593_74.n0 a_593_74.t2 26.2505
R165 a_593_74.n1 a_593_74.t3 26.2505
R166 a_593_74.t1 a_593_74.n1 26.2505
C0 VPB C1 0.071938f
C1 A1 VPWR 0.042213f
C2 A2 Y 0.052788f
C3 B2 VGND 0.022441f
C4 C2 C1 0.246106f
C5 VPB B1 0.099554f
C6 A2 VPWR 0.029672f
C7 A1 VGND 0.02285f
C8 C2 B1 0.027444f
C9 VPB B2 0.078191f
C10 Y VPWR 0.065264f
C11 A2 VGND 0.027276f
C12 VPB A1 0.094867f
C13 Y VGND 0.241837f
C14 VPB A2 0.071094f
C15 VPWR VGND 0.102653f
C16 B1 B2 0.243778f
C17 VPB Y 0.039062f
C18 C2 Y 0.336411f
C19 VPB VPWR 0.151177f
C20 B1 A1 0.105958f
C21 VPB VGND 0.011093f
C22 B2 A1 3.73e-19
C23 C2 VPWR 0.018157f
C24 C1 Y 0.073192f
C25 C1 VPWR 0.010728f
C26 B1 Y 0.143794f
C27 C2 VGND 0.054484f
C28 B2 A2 2.6e-19
C29 B2 Y 0.064246f
C30 B1 VPWR 0.019475f
C31 C1 VGND 0.015045f
C32 A1 A2 0.243797f
C33 VPB C2 0.095468f
C34 B1 VGND 0.022503f
C35 B2 VPWR 0.012196f
C36 A1 Y 0.135595f
C37 VGND VNB 0.817789f
C38 VPWR VNB 0.623655f
C39 Y VNB 0.207885f
C40 A2 VNB 0.199156f
C41 A1 VNB 0.270158f
C42 B2 VNB 0.230462f
C43 B1 VNB 0.229402f
C44 C1 VNB 0.201337f
C45 C2 VNB 0.286267f
C46 VPB VNB 1.58472f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a311o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311o_1 VNB VPB VPWR VGND X C1 B1 A3 A2 A1
X0 a_258_392.t0 A3.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2809 ps=1.65 w=1 l=0.15
X1 a_546_392.t1 B1.t0 a_258_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.15 ps=1.3 w=1 l=0.15
X2 VGND.t2 B1.t1 a_89_270.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.136 pd=1.065 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 VPWR.t1 a_89_270.t4 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2809 pd=1.65 as=0.308 ps=2.79 w=1.12 l=0.15
X4 a_258_392.t2 A1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X5 a_359_123.t1 A2.t0 a_264_120.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1053 ps=0.98 w=0.64 l=0.15
X6 a_264_120.t0 A3.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1053 pd=0.98 as=0.12845 ps=1.1 w=0.64 l=0.15
X7 a_89_270.t2 C1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.136 ps=1.065 w=0.64 l=0.15
X8 a_89_270.t0 C1.t1 a_546_392.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.12 ps=1.24 w=1 l=0.15
X9 a_89_270.t3 A1.t1 a_359_123.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1024 ps=0.96 w=0.64 l=0.15
X10 VGND.t1 a_89_270.t5 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.12845 pd=1.1 as=0.1961 ps=2.01 w=0.74 l=0.15
X11 VPWR.t3 A2.t1 a_258_392.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.15 ps=1.3 w=1 l=0.15
R0 A3.n0 A3.t0 236.983
R1 A3.n0 A3.t1 194.407
R2 A3 A3.n0 155.298
R3 VPWR.n2 VPWR.n0 326.384
R4 VPWR.n2 VPWR.n1 219.381
R5 VPWR.n1 VPWR.t0 52.2055
R6 VPWR.n1 VPWR.t1 50.3459
R7 VPWR.n0 VPWR.t2 43.3405
R8 VPWR.n0 VPWR.t3 33.4905
R9 VPWR VPWR.n2 0.442502
R10 a_258_392.n1 a_258_392.n0 460.384
R11 a_258_392.n0 a_258_392.t1 29.5505
R12 a_258_392.n0 a_258_392.t2 29.5505
R13 a_258_392.n1 a_258_392.t3 29.5505
R14 a_258_392.t0 a_258_392.n1 29.5505
R15 VPB.t3 VPB.t0 347.312
R16 VPB.t5 VPB.t4 275.807
R17 VPB VPB.t3 273.253
R18 VPB.t4 VPB.t1 229.839
R19 VPB.t0 VPB.t5 229.839
R20 VPB.t1 VPB.t2 199.195
R21 B1.t1 B1.t0 456.293
R22 B1 B1.t1 319.029
R23 a_546_392.t0 a_546_392.t1 47.2805
R24 a_89_270.n3 a_89_270.t2 278.466
R25 a_89_270.n2 a_89_270.n0 269.517
R26 a_89_270.t0 a_89_270.n3 250.238
R27 a_89_270.n0 a_89_270.t4 248.597
R28 a_89_270.n2 a_89_270.n1 192.37
R29 a_89_270.n0 a_89_270.t5 176.03
R30 a_89_270.n3 a_89_270.n2 63.818
R31 a_89_270.n1 a_89_270.t1 26.2505
R32 a_89_270.n1 a_89_270.t3 26.2505
R33 VGND.n2 VGND.n1 251.036
R34 VGND.n2 VGND.n0 221.659
R35 VGND.n1 VGND.t2 41.2505
R36 VGND.n0 VGND.t0 41.2505
R37 VGND.n1 VGND.t3 38.438
R38 VGND.n0 VGND.t1 22.1988
R39 VGND VGND.n2 0.247415
R40 VNB VNB.t1 1697.64
R41 VNB.t2 VNB.t4 1328.08
R42 VNB.t1 VNB.t0 1177.95
R43 VNB.t0 VNB.t3 1097.11
R44 VNB.t3 VNB.t5 1085.56
R45 VNB.t5 VNB.t2 993.177
R46 X X.n0 589.572
R47 X.n2 X.n0 585
R48 X.n1 X.n0 585
R49 X X.t0 206.875
R50 X.n0 X.t1 26.3844
R51 X X.n1 11.1548
R52 X X.n2 10.0576
R53 X.n2 X 3.47479
R54 X.n1 X 2.37764
R55 A1.t1 A1.t0 460.31
R56 A1 A1.t1 319.317
R57 A2.n0 A2.t1 236.983
R58 A2.n0 A2.t0 189.588
R59 A2 A2.n0 157.625
R60 a_264_120.t0 a_264_120.t1 55.6399
R61 a_359_123.t0 a_359_123.t1 60.0005
R62 C1.t0 C1.t1 468.344
R63 C1 C1.t0 347.067
C0 A3 A2 0.082396f
C1 VPB A1 0.031432f
C2 X VGND 0.067156f
C3 VPB B1 0.029507f
C4 A3 A1 0.002049f
C5 VPWR VGND 0.063042f
C6 A2 A1 0.065362f
C7 VPB C1 0.045968f
C8 VPB X 0.01822f
C9 A2 B1 6.2e-19
C10 A2 C1 3.3e-19
C11 A3 X 0.004026f
C12 VPB VPWR 0.108075f
C13 A1 B1 0.112692f
C14 A2 X 3.06e-19
C15 A3 VPWR 0.023016f
C16 VPB VGND 0.010031f
C17 B1 C1 0.08453f
C18 A2 VPWR 0.014565f
C19 A3 VGND 0.011934f
C20 A1 X 1.5e-19
C21 A2 VGND 0.006014f
C22 B1 X 8.85e-20
C23 A1 VPWR 0.014391f
C24 B1 VPWR 0.006803f
C25 A1 VGND 0.093681f
C26 C1 X 6.52e-20
C27 VPB A3 0.044834f
C28 B1 VGND 0.091718f
C29 C1 VPWR 0.01048f
C30 VPB A2 0.041117f
C31 C1 VGND 0.107792f
C32 X VPWR 0.126095f
C33 VGND VNB 0.513889f
C34 VPWR VNB 0.392712f
C35 X VNB 0.11389f
C36 C1 VNB 0.227274f
C37 B1 VNB 0.121332f
C38 A1 VNB 0.137377f
C39 A2 VNB 0.093023f
C40 A3 VNB 0.099073f
C41 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a311o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311o_2 VNB VPB VPWR VGND C1 B1 A3 A2 A1 X
X0 a_21_270.t0 C1.t0 a_660_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t1 a_21_270.t4 X.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2015 pd=1.49 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_330_392.t0 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.27 ps=1.54 w=1 l=0.15
X3 a_660_392.t1 B1.t0 a_330_392.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X4 a_351_74.t0 A3.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1554 ps=1.16 w=0.74 l=0.15
X5 X.t1 a_21_270.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X6 a_21_270.t2 A1.t1 a_423_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X7 a_423_74.t1 A2.t0 a_351_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X8 VPWR.t4 A2.t1 a_330_392.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.27 pd=1.54 as=0.165 ps=1.33 w=1 l=0.15
X9 a_330_392.t1 A3.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.2015 ps=1.49 w=1 l=0.15
X10 X.t3 a_21_270.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X11 VGND.t4 B1.t1 a_21_270.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X12 a_21_270.t1 C1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X13 VGND.t1 a_21_270.t7 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 C1.n0 C1.t1 224.934
R1 C1.n0 C1.t0 216.972
R2 C1 C1.n0 211.035
R3 a_660_392.t0 a_660_392.t1 53.1905
R4 a_21_270.t0 a_21_270.n5 419.885
R5 a_21_270.n5 a_21_270.n2 301.608
R6 a_21_270.n0 a_21_270.t4 291.44
R7 a_21_270.n2 a_21_270.t5 226.809
R8 a_21_270.n0 a_21_270.t7 212.446
R9 a_21_270.n4 a_21_270.t1 198.948
R10 a_21_270.n1 a_21_270.t6 196.013
R11 a_21_270.n5 a_21_270.n4 168.66
R12 a_21_270.n4 a_21_270.n3 98.6841
R13 a_21_270.n1 a_21_270.n0 78.435
R14 a_21_270.n3 a_21_270.t3 37.2978
R15 a_21_270.n3 a_21_270.t2 25.9464
R16 a_21_270.n2 a_21_270.n1 10.955
R17 VPB.t5 VPB.t3 352.42
R18 VPB VPB.t1 309.005
R19 VPB.t2 VPB.t4 265.591
R20 VPB.t3 VPB.t6 245.161
R21 VPB.t4 VPB.t5 245.161
R22 VPB.t1 VPB.t2 229.839
R23 VPB.t6 VPB.t0 214.517
R24 X X.n0 597.965
R25 X X.n1 125.797
R26 X.n0 X.t2 26.3844
R27 X.n0 X.t1 26.3844
R28 X.n1 X.t0 22.7032
R29 X.n1 X.t3 22.7032
R30 VPWR.n6 VPWR.t0 848.062
R31 VPWR.n4 VPWR.n1 608.08
R32 VPWR.n3 VPWR.n2 591.077
R33 VPWR.n2 VPWR.t2 53.1905
R34 VPWR.n2 VPWR.t4 53.1905
R35 VPWR.n1 VPWR.t3 43.3405
R36 VPWR.n5 VPWR.n4 29.7417
R37 VPWR.n1 VPWR.t1 27.4811
R38 VPWR.n6 VPWR.n5 13.177
R39 VPWR.n5 VPWR.n0 9.3005
R40 VPWR.n7 VPWR.n6 9.3005
R41 VPWR.n4 VPWR.n3 6.55142
R42 VPWR.n3 VPWR.n0 0.380013
R43 VPWR.n7 VPWR.n0 0.122949
R44 VPWR VPWR.n7 0.0617245
R45 A1.n0 A1.t1 252.248
R46 A1.n0 A1.t0 236.983
R47 A1 A1.n0 156.462
R48 a_330_392.n1 a_330_392.n0 633.021
R49 a_330_392.n0 a_330_392.t2 35.4605
R50 a_330_392.t0 a_330_392.n1 35.4605
R51 a_330_392.n0 a_330_392.t1 29.5505
R52 a_330_392.n1 a_330_392.t3 29.5505
R53 B1.n0 B1.t0 287.861
R54 B1.n0 B1.t1 191.194
R55 B1.n1 B1.n0 152
R56 B1.n1 B1 7.50819
R57 B1 B1.n1 4.30819
R58 A3.n0 A3.t1 287.861
R59 A3.n0 A3.t0 191.194
R60 A3 A3.n0 158.841
R61 VGND.n4 VGND.n3 211.472
R62 VGND.n2 VGND.n1 203.72
R63 VGND.n8 VGND.t2 175.351
R64 VGND.n1 VGND.t1 39.7302
R65 VGND.n3 VGND.t0 37.2978
R66 VGND.n7 VGND.n6 36.1417
R67 VGND.n1 VGND.t3 28.3789
R68 VGND.n3 VGND.t4 25.9464
R69 VGND.n9 VGND.n8 13.8181
R70 VGND.n8 VGND.n7 12.8005
R71 VGND.n4 VGND.n2 11.3903
R72 VGND.n6 VGND.n5 9.3005
R73 VGND.n7 VGND.n0 9.3005
R74 VGND.n6 VGND.n2 2.25932
R75 VGND.n5 VGND.n4 0.174321
R76 VGND.n5 VGND.n0 0.122949
R77 VGND.n9 VGND.n0 0.122949
R78 VGND VGND.n9 0.0617245
R79 a_351_74.t0 a_351_74.t1 34.0546
R80 VNB VNB.t2 1570.6
R81 VNB.t1 VNB.t3 1316.54
R82 VNB.t5 VNB.t0 1247.24
R83 VNB.t4 VNB.t5 1247.24
R84 VNB.t6 VNB.t4 1247.24
R85 VNB.t2 VNB.t1 993.177
R86 VNB.t3 VNB.t6 831.496
R87 a_423_74.t0 a_423_74.t1 63.2437
R88 A2.n0 A2.t0 252.248
R89 A2.n0 A2.t1 236.983
R90 A2 A2.n0 154.133
C0 VPB A3 0.042261f
C1 B1 VGND 0.016319f
C2 VPB A2 0.042895f
C3 VPWR X 0.016412f
C4 C1 VGND 0.015946f
C5 A3 A2 0.101726f
C6 VPB A1 0.042895f
C7 VPWR VGND 0.070423f
C8 A3 A1 5.58e-19
C9 VPB B1 0.038899f
C10 X VGND 0.138164f
C11 A3 B1 0.003589f
C12 VPB C1 0.066956f
C13 A2 A1 0.077836f
C14 VPB VPWR 0.122375f
C15 A2 B1 4.13e-19
C16 A1 B1 0.084774f
C17 VPB X 0.00219f
C18 A3 VPWR 0.014915f
C19 VPB VGND 0.009638f
C20 A3 X 0.001131f
C21 A2 VPWR 0.013214f
C22 A1 VPWR 0.012705f
C23 B1 C1 0.112357f
C24 A2 X 3.26e-19
C25 A3 VGND 0.014529f
C26 B1 VPWR 0.010753f
C27 A1 X 1.35e-19
C28 A2 VGND 0.012056f
C29 A1 VGND 0.008593f
C30 C1 VPWR 0.010995f
C31 VGND VNB 0.587347f
C32 X VNB 0.014757f
C33 VPWR VNB 0.441746f
C34 C1 VNB 0.178959f
C35 B1 VNB 0.119329f
C36 A1 VNB 0.104414f
C37 A2 VNB 0.099914f
C38 A3 VNB 0.107004f
C39 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a311o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311o_4 VNB VPB VPWR X VGND C1 B1 A3 A2 A1
X0 a_888_105.t3 A2.t0 a_1081_39.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1088 ps=0.98 w=0.64 l=0.15
X1 VGND.t9 a_154_392.t8 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.12205 pd=1.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_154_392.t1 B1.t0 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 a_69_392.t1 B1.t1 a_334_392.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X4 a_154_392.t3 C1.t0 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X5 VGND.t5 A3.t0 a_888_105.t1 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X6 X.t2 a_154_392.t9 VGND.t8 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1165 ps=1.065 w=0.74 l=0.15
X7 VGND.t2 B1.t2 a_154_392.t2 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1165 pd=1.065 as=0.0896 ps=0.92 w=0.64 l=0.15
X8 a_1081_39.t1 A2.t1 a_888_105.t2 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X9 X.t1 a_154_392.t10 VGND.t7 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12155 ps=1.08 w=0.74 l=0.15
X10 VGND.t4 C1.t1 a_154_392.t4 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X11 VGND.t6 a_154_392.t11 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.12155 pd=1.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 VPWR.t7 a_154_392.t12 X.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.199 pd=1.485 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_154_392.t0 A1.t0 a_1081_39.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.3055 ps=2.71 w=0.64 l=0.15
X14 X.t6 a_154_392.t13 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_334_392.t2 B1.t3 a_69_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X16 VPWR.t5 a_154_392.t14 X.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 X.t4 a_154_392.t15 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X18 a_69_392.t2 C1.t2 a_154_392.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X19 a_154_392.t7 C1.t3 a_69_392.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X20 VPWR.t0 A1.t1 a_334_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X21 a_334_392.t4 A3.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.199 ps=1.485 w=1 l=0.15
X22 a_334_392.t5 A2.t2 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.165 ps=1.33 w=1 l=0.15
X23 a_1081_39.t3 A1.t2 a_154_392.t5 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1088 pd=0.98 as=0.0896 ps=0.92 w=0.64 l=0.15
X24 VPWR.t1 A3.t2 a_334_392.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X25 a_888_105.t0 A3.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.12205 ps=1.08 w=0.64 l=0.15
R0 A2.n1 A2.t2 214.793
R1 A2.n3 A2.n0 212.883
R2 A2 A2.n3 190.649
R3 A2.n1 A2.t0 175.127
R4 A2.n2 A2.t1 175.127
R5 A2.n2 A2.n1 62.8066
R6 A2.n3 A2.n2 0.730803
R7 a_1081_39.t0 a_1081_39.n1 580.169
R8 a_1081_39.n1 a_1081_39.n0 237.599
R9 a_1081_39.n1 a_1081_39.t1 128.471
R10 a_1081_39.n0 a_1081_39.t2 37.5005
R11 a_1081_39.n0 a_1081_39.t3 26.2505
R12 a_888_105.n1 a_888_105.n0 540.571
R13 a_888_105.n0 a_888_105.t1 26.2505
R14 a_888_105.n0 a_888_105.t0 26.2505
R15 a_888_105.t2 a_888_105.n1 26.2505
R16 a_888_105.n1 a_888_105.t3 26.2505
R17 VNB.t10 VNB.t5 2332.81
R18 VNB VNB.t8 1790.03
R19 VNB.t13 VNB.t12 1131.76
R20 VNB.t1 VNB.t0 1131.76
R21 VNB.t4 VNB.t3 1097.11
R22 VNB.t7 VNB.t2 1097.11
R23 VNB.t12 VNB.t11 993.177
R24 VNB.t5 VNB.t13 993.177
R25 VNB.t0 VNB.t10 993.177
R26 VNB.t3 VNB.t1 993.177
R27 VNB.t2 VNB.t4 993.177
R28 VNB.t6 VNB.t7 993.177
R29 VNB.t9 VNB.t6 993.177
R30 VNB.t8 VNB.t9 993.177
R31 a_154_392.n19 a_154_392.n18 651.26
R32 a_154_392.n7 a_154_392.n2 410.575
R33 a_154_392.n3 a_154_392.t12 327.187
R34 a_154_392.n3 a_154_392.t13 208.064
R35 a_154_392.n5 a_154_392.t14 208.064
R36 a_154_392.n11 a_154_392.t15 208.064
R37 a_154_392.n13 a_154_392.t9 193.697
R38 a_154_392.n12 a_154_392.t11 173.52
R39 a_154_392.n1 a_154_392.t10 168.701
R40 a_154_392.n4 a_154_392.t8 168.701
R41 a_154_392.n14 a_154_392.n13 152
R42 a_154_392.n10 a_154_392.n0 152
R43 a_154_392.n9 a_154_392.n8 152
R44 a_154_392.n7 a_154_392.n6 152
R45 a_154_392.n18 a_154_392.n17 120.731
R46 a_154_392.n16 a_154_392.n15 120.376
R47 a_154_392.n18 a_154_392.n16 50.824
R48 a_154_392.n16 a_154_392.n14 38.6881
R49 a_154_392.n10 a_154_392.n9 38.1121
R50 a_154_392.n6 a_154_392.n5 30.8261
R51 a_154_392.t6 a_154_392.n19 29.5505
R52 a_154_392.n19 a_154_392.t7 29.5505
R53 a_154_392.n13 a_154_392.n12 28.0238
R54 a_154_392.n2 a_154_392.t5 26.2505
R55 a_154_392.n2 a_154_392.t0 26.2505
R56 a_154_392.n15 a_154_392.t2 26.2505
R57 a_154_392.n15 a_154_392.t1 26.2505
R58 a_154_392.n17 a_154_392.t4 26.2505
R59 a_154_392.n17 a_154_392.t3 26.2505
R60 a_154_392.n6 a_154_392.n4 15.1331
R61 a_154_392.n8 a_154_392.n7 13.1884
R62 a_154_392.n8 a_154_392.n0 13.1884
R63 a_154_392.n14 a_154_392.n0 13.1884
R64 a_154_392.n9 a_154_392.n1 5.04469
R65 a_154_392.n11 a_154_392.n10 5.04469
R66 a_154_392.n12 a_154_392.n11 5.04469
R67 a_154_392.n4 a_154_392.n3 4.48422
R68 a_154_392.n5 a_154_392.n1 2.24236
R69 X.n5 X.n3 619.909
R70 X.n5 X.n4 585
R71 X.n6 X.n5 333.692
R72 X.n2 X.n0 148.536
R73 X.n2 X.n1 94.9818
R74 X.n4 X.t5 26.3844
R75 X.n4 X.t4 26.3844
R76 X.n3 X.t7 26.3844
R77 X.n3 X.t6 26.3844
R78 X.n1 X.t0 22.7032
R79 X.n1 X.t2 22.7032
R80 X.n0 X.t3 22.7032
R81 X.n0 X.t1 22.7032
R82 X.n6 X.n2 12.3667
R83 X X.n6 0.0466957
R84 VGND.n4 VGND.t5 319.861
R85 VGND.n16 VGND.t3 285.774
R86 VGND.n2 VGND.n1 225.704
R87 VGND.n7 VGND.n6 221.019
R88 VGND.n14 VGND.n13 116.436
R89 VGND.n4 VGND.n3 87.4775
R90 VGND.n5 VGND.n4 44.9924
R91 VGND.n3 VGND.t0 37.5005
R92 VGND.n16 VGND.n15 35.7652
R93 VGND.n8 VGND.n7 34.6358
R94 VGND.n12 VGND.n2 32.7534
R95 VGND.n1 VGND.t8 31.0986
R96 VGND.n1 VGND.t2 26.2505
R97 VGND.n13 VGND.t1 26.2505
R98 VGND.n13 VGND.t4 26.2505
R99 VGND.n6 VGND.t7 25.0707
R100 VGND.n6 VGND.t6 24.2431
R101 VGND.n3 VGND.t9 22.1988
R102 VGND.n8 VGND.n2 20.7064
R103 VGND.n15 VGND.n0 9.3005
R104 VGND.n12 VGND.n11 9.3005
R105 VGND.n10 VGND.n2 9.3005
R106 VGND.n9 VGND.n8 9.3005
R107 VGND.n14 VGND.n12 7.15344
R108 VGND.n7 VGND.n5 6.58549
R109 VGND.n17 VGND.n16 6.41781
R110 VGND.n15 VGND.n14 4.14168
R111 VGND.n9 VGND.n5 0.568226
R112 VGND.n17 VGND.n0 0.160917
R113 VGND VGND.n17 0.146712
R114 VGND.n10 VGND.n9 0.122949
R115 VGND.n11 VGND.n10 0.122949
R116 VGND.n11 VGND.n0 0.122949
R117 B1.n0 B1.t2 240.583
R118 B1.n1 B1.t0 237.787
R119 B1.n1 B1.t3 213.37
R120 B1.n0 B1.t1 207.529
R121 B1 B1.n2 156.073
R122 B1.n2 B1.n0 50.3914
R123 B1.n2 B1.n1 9.49444
R124 a_334_392.n2 a_334_392.n0 822.178
R125 a_334_392.n3 a_334_392.t5 316.817
R126 a_334_392.n2 a_334_392.n1 297.889
R127 a_334_392.t0 a_334_392.n3 224.733
R128 a_334_392.n3 a_334_392.n2 60.7765
R129 a_334_392.n1 a_334_392.t3 29.5505
R130 a_334_392.n1 a_334_392.t4 29.5505
R131 a_334_392.n0 a_334_392.t1 29.5505
R132 a_334_392.n0 a_334_392.t2 29.5505
R133 a_69_392.t1 a_69_392.n1 870.932
R134 a_69_392.n1 a_69_392.t3 867.797
R135 a_69_392.n1 a_69_392.n0 585
R136 a_69_392.n0 a_69_392.t0 29.5505
R137 a_69_392.n0 a_69_392.t2 29.5505
R138 VPB.t2 VPB.t8 495.43
R139 VPB.t3 VPB.t0 459.678
R140 VPB VPB.t7 354.974
R141 VPB.t11 VPB.t4 263.038
R142 VPB.t0 VPB.t5 245.161
R143 VPB.t4 VPB.t3 229.839
R144 VPB.t10 VPB.t11 229.839
R145 VPB.t9 VPB.t10 229.839
R146 VPB.t8 VPB.t9 229.839
R147 VPB.t1 VPB.t2 229.839
R148 VPB.t6 VPB.t1 229.839
R149 VPB.t7 VPB.t6 229.839
R150 C1.n0 C1.t1 238.935
R151 C1.n1 C1.t0 228.148
R152 C1.n0 C1.t2 207.529
R153 C1.n2 C1.t3 207.529
R154 C1 C1.n2 158.82
R155 C1.n1 C1.n0 49.5394
R156 C1.n2 C1.n1 10.7116
R157 A3.n0 A3.t3 252.644
R158 A3.n2 A3.t2 250.13
R159 A3.n1 A3.t1 220.917
R160 A3 A3.n2 158.222
R161 A3.n0 A3.t0 134.091
R162 A3.n2 A3.n1 36.5157
R163 A3.n1 A3.n0 23.7831
R164 VPWR.n15 VPWR.t4 878.553
R165 VPWR.n7 VPWR.t1 838.431
R166 VPWR.n13 VPWR.n2 606.333
R167 VPWR.n4 VPWR.n3 606.333
R168 VPWR.n6 VPWR.n5 319.423
R169 VPWR.n3 VPWR.t2 42.3555
R170 VPWR.n5 VPWR.t3 32.5055
R171 VPWR.n5 VPWR.t0 32.5055
R172 VPWR.n8 VPWR.n7 32.377
R173 VPWR.n14 VPWR.n13 30.4946
R174 VPWR.n3 VPWR.t7 27.4811
R175 VPWR.n2 VPWR.t6 26.3844
R176 VPWR.n2 VPWR.t5 26.3844
R177 VPWR.n12 VPWR.n4 25.977
R178 VPWR.n8 VPWR.n4 21.4593
R179 VPWR.n13 VPWR.n12 16.9417
R180 VPWR.n15 VPWR.n14 12.424
R181 VPWR.n9 VPWR.n8 9.3005
R182 VPWR.n10 VPWR.n4 9.3005
R183 VPWR.n12 VPWR.n11 9.3005
R184 VPWR.n13 VPWR.n1 9.3005
R185 VPWR.n14 VPWR.n0 9.3005
R186 VPWR.n16 VPWR.n15 7.61468
R187 VPWR.n7 VPWR.n6 6.53239
R188 VPWR VPWR.n16 0.649974
R189 VPWR.n9 VPWR.n6 0.588889
R190 VPWR.n16 VPWR.n0 0.15003
R191 VPWR.n10 VPWR.n9 0.122949
R192 VPWR.n11 VPWR.n10 0.122949
R193 VPWR.n11 VPWR.n1 0.122949
R194 VPWR.n1 VPWR.n0 0.122949
R195 A1.n1 A1.n0 216.536
R196 A1.n2 A1.t1 212.883
R197 A1.n1 A1.t0 175.127
R198 A1.n3 A1.t2 175.127
R199 A1.n4 A1.n3 153.462
R200 A1.n2 A1.n1 62.0763
R201 A1.n4 A1 12.8005
R202 A1 A1.n4 5.81868
R203 A1.n3 A1.n2 0.730803
C0 VPB A2 0.095552f
C1 B1 A3 7.18e-19
C2 VPB VPWR 0.206777f
C3 VPB X 0.038716f
C4 C1 VPWR 0.009878f
C5 A3 A1 0.04319f
C6 C1 X 0.081609f
C7 VPB VGND 0.008779f
C8 B1 VPWR 0.010681f
C9 B1 X 0.071646f
C10 C1 VGND 0.03287f
C11 A1 A2 0.106014f
C12 A3 VPWR 0.027589f
C13 A1 VPWR 0.037893f
C14 A3 X 0.002085f
C15 B1 VGND 0.026101f
C16 A1 X 2.44e-19
C17 A3 VGND 0.061798f
C18 A2 VPWR 0.073872f
C19 VPB C1 0.086538f
C20 A1 VGND 0.011946f
C21 A2 X 9.44e-20
C22 VPB B1 0.080427f
C23 VPWR X 0.112474f
C24 A2 VGND 0.010736f
C25 C1 B1 0.069668f
C26 VPB A3 0.087304f
C27 VPWR VGND 0.082808f
C28 VPB A1 0.079153f
C29 X VGND 0.479539f
C30 VGND VNB 0.929253f
C31 X VNB 0.112886f
C32 VPWR VNB 0.732388f
C33 A2 VNB 0.24791f
C34 A1 VNB 0.193714f
C35 A3 VNB 0.236914f
C36 B1 VNB 0.198615f
C37 C1 VNB 0.242646f
C38 VPB VNB 1.79899f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a311oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311oi_1 VNB VPB VPWR VGND C1 B1 A3 A2 A1 Y
X0 a_462_368.t1 B1.t0 a_156_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X1 Y.t3 C1.t0 a_462_368.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1848 ps=1.45 w=1.12 l=0.15
X2 a_156_368.t2 A1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2688 ps=1.6 w=1.12 l=0.15
X3 a_231_74.t1 A2.t0 a_159_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X4 a_159_74.t1 A3.t0 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1961 ps=2.01 w=0.74 l=0.15
X5 Y.t0 A1.t1 a_231_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X6 VGND.t0 B1.t1 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X7 Y.t2 C1.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X8 VPWR.t1 A2.t1 a_156_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2688 pd=1.6 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_156_368.t0 A3.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
R0 B1.n0 B1.t0 250.909
R1 B1.n0 B1.t1 220.113
R2 B1.n1 B1.n0 152
R3 B1 B1.n1 9.07957
R4 B1.n1 B1 5.2098
R5 a_156_368.n1 a_156_368.n0 651.938
R6 a_156_368.n0 a_156_368.t3 26.3844
R7 a_156_368.n0 a_156_368.t2 26.3844
R8 a_156_368.n1 a_156_368.t1 26.3844
R9 a_156_368.t0 a_156_368.n1 26.3844
R10 a_462_368.t0 a_462_368.t1 58.0451
R11 VPB VPB.t0 360.082
R12 VPB.t1 VPB.t2 321.774
R13 VPB.t4 VPB.t3 245.161
R14 VPB.t2 VPB.t4 229.839
R15 VPB.t0 VPB.t1 229.839
R16 C1.n0 C1.t0 226.809
R17 C1 C1.n0 209.294
R18 C1.n0 C1.t1 198.204
R19 Y Y.t3 468.005
R20 Y.n1 Y.t2 209.034
R21 Y.n1 Y.n0 92.5005
R22 Y.n0 Y.t1 37.2978
R23 Y.n0 Y.t0 25.9464
R24 Y Y.n1 4.01014
R25 A1.n0 A1.t0 250.909
R26 A1.n0 A1.t1 220.113
R27 A1 A1.n0 155.423
R28 VPWR.n1 VPWR.n0 607.636
R29 VPWR.n1 VPWR.t0 357.899
R30 VPWR.n0 VPWR.t2 42.2148
R31 VPWR.n0 VPWR.t1 42.2148
R32 VPWR VPWR.n1 0.395215
R33 A2.n0 A2.t1 250.909
R34 A2.n0 A2.t0 220.113
R35 A2 A2.n0 154.522
R36 a_159_74.t0 a_159_74.t1 34.0546
R37 a_231_74.t0 a_231_74.t1 63.2437
R38 VNB VNB.t4 1662.99
R39 VNB.t2 VNB.t3 1247.24
R40 VNB.t0 VNB.t2 1247.24
R41 VNB.t1 VNB.t0 1247.24
R42 VNB.t4 VNB.t1 831.496
R43 A3.n0 A3.t1 261.62
R44 A3.n1 A3.n0 206.774
R45 A3.n0 A3.t0 156.431
R46 A3 A3.n1 6.74645
R47 A3.n1 A3 6.05455
R48 VGND.n1 VGND.t1 240.637
R49 VGND.n1 VGND.n0 214.656
R50 VGND.n0 VGND.t2 37.2978
R51 VGND.n0 VGND.t0 25.9464
R52 VGND VGND.n1 0.165254
C0 VPB A3 0.052667f
C1 B1 VGND 0.016377f
C2 C1 Y 0.074876f
C3 VPB A2 0.033736f
C4 VPWR Y 0.073688f
C5 C1 VGND 0.017428f
C6 A3 A2 0.069458f
C7 VPB A1 0.033736f
C8 VPWR VGND 0.058743f
C9 VPB B1 0.033003f
C10 Y VGND 0.306929f
C11 A2 A1 0.081986f
C12 VPB C1 0.055165f
C13 VPB VPWR 0.104006f
C14 A3 VPWR 0.026143f
C15 A1 B1 0.092283f
C16 VPB Y 0.025373f
C17 VPB VGND 0.009494f
C18 A3 Y 0.080452f
C19 A2 VPWR 0.012285f
C20 A3 VGND 0.034515f
C21 A1 VPWR 0.013287f
C22 A2 Y 0.117252f
C23 B1 C1 0.104414f
C24 B1 VPWR 0.009654f
C25 A2 VGND 0.010125f
C26 A1 Y 0.079948f
C27 B1 Y 0.146793f
C28 A1 VGND 0.005271f
C29 C1 VPWR 0.011387f
C30 VGND VNB 0.467164f
C31 Y VNB 0.126538f
C32 VPWR VNB 0.377463f
C33 C1 VNB 0.181538f
C34 B1 VNB 0.106551f
C35 A1 VNB 0.104112f
C36 A2 VNB 0.100569f
C37 A3 VNB 0.192133f
C38 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a221oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221oi_4 VNB VPB VPWR VGND Y C1 B2 B1 A2 A1
X0 VPWR.t3 A1.t0 a_531_368.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t2 A1.t1 a_531_368.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2968 pd=1.65 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_534_74.t2 A1.t2 Y.t9 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_531_368.t7 A2.t0 VPWR.t4 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_531_368.t3 A1.t3 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 VPWR.t5 A2.t1 a_531_368.t8 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_531_368.t9 A2.t2 VPWR.t6 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t6 C1.t0 a_114_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t7 A2.t3 a_531_368.t10 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X9 a_114_368.t2 C1.t1 Y.t10 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_534_74.t3 A2.t4 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 Y.t11 B1.t0 a_1326_74.t0 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X12 Y.t0 C1.t2 a_114_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_531_368.t0 B2.t0 a_114_368.t11 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_534_74.t4 A2.t5 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_114_368.t10 B2.t1 a_531_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VGND.t9 B2.t2 a_1326_74.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t5 A2.t6 a_534_74.t5 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 VGND.t8 B2.t3 a_1326_74.t2 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 VGND.t0 C1.t3 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VGND.t4 A2.t7 a_534_74.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X21 VGND.t1 C1.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X22 Y.t12 B1.t1 a_1326_74.t1 VNB.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X23 a_114_368.t0 C1.t5 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X24 a_531_368.t6 B2.t4 a_114_368.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 Y.t8 A1.t4 a_534_74.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 a_114_368.t8 B2.t5 a_531_368.t11 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 Y.t4 C1.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 a_531_368.t12 B1.t2 a_114_368.t4 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 a_114_368.t5 B1.t3 a_531_368.t13 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_531_368.t14 B1.t4 a_114_368.t6 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X31 Y.t5 C1.t7 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X32 a_114_368.t7 B1.t5 a_531_368.t15 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X33 Y.t7 A1.t5 a_534_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X34 a_531_368.t2 A1.t6 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2968 ps=1.65 w=1.12 l=0.15
R0 A1.n1 A1.t6 263.885
R1 A1.n10 A1.t3 226.809
R2 A1.n5 A1.t0 226.809
R3 A1.n3 A1.t1 218.774
R4 A1.n5 A1.t5 196.416
R5 A1.n9 A1.t2 186.374
R6 A1.n1 A1.n0 186.374
R7 A1.n4 A1.t4 184.332
R8 A1 A1.n2 153.28
R9 A1.n12 A1.n11 152
R10 A1.n9 A1.n8 152
R11 A1.n7 A1.n6 152
R12 A1.n9 A1.n6 45.5227
R13 A1.n11 A1.n10 32.8033
R14 A1.n3 A1.n2 30.28
R15 A1 A1.n12 15.1776
R16 A1.n4 A1.n3 14.1622
R17 A1.n10 A1.n9 12.7199
R18 A1.n7 A1 12.6176
R19 A1.n11 A1.n4 11.7677
R20 A1.n8 A1 10.0576
R21 A1.n2 A1.n1 8.65178
R22 A1.n8 A1 7.49764
R23 A1 A1.n7 4.93764
R24 A1.n12 A1 2.37764
R25 A1.n6 A1.n5 2.00883
R26 a_531_368.n1 a_531_368.t10 366.743
R27 a_531_368.n9 a_531_368.n8 307.164
R28 a_531_368.n11 a_531_368.n10 307.164
R29 a_531_368.n13 a_531_368.n12 307.164
R30 a_531_368.n1 a_531_368.n0 297.44
R31 a_531_368.n3 a_531_368.n2 297.44
R32 a_531_368.n5 a_531_368.n4 297.44
R33 a_531_368.t0 a_531_368.n13 294.469
R34 a_531_368.n7 a_531_368.n6 288.443
R35 a_531_368.n7 a_531_368.n5 72.0079
R36 a_531_368.n9 a_531_368.n7 66.5625
R37 a_531_368.n11 a_531_368.n9 50.4476
R38 a_531_368.n13 a_531_368.n11 50.4476
R39 a_531_368.n3 a_531_368.n1 42.9181
R40 a_531_368.n5 a_531_368.n3 42.9181
R41 a_531_368.n6 a_531_368.t15 26.3844
R42 a_531_368.n6 a_531_368.t2 26.3844
R43 a_531_368.n0 a_531_368.t8 26.3844
R44 a_531_368.n0 a_531_368.t9 26.3844
R45 a_531_368.n2 a_531_368.t5 26.3844
R46 a_531_368.n2 a_531_368.t7 26.3844
R47 a_531_368.n4 a_531_368.t4 26.3844
R48 a_531_368.n4 a_531_368.t3 26.3844
R49 a_531_368.n8 a_531_368.t13 26.3844
R50 a_531_368.n8 a_531_368.t14 26.3844
R51 a_531_368.n10 a_531_368.t11 26.3844
R52 a_531_368.n10 a_531_368.t12 26.3844
R53 a_531_368.n12 a_531_368.t1 26.3844
R54 a_531_368.n12 a_531_368.t6 26.3844
R55 VPWR.n1 VPWR.n0 618.13
R56 VPWR.n10 VPWR.n3 618.13
R57 VPWR.n5 VPWR.n4 618.13
R58 VPWR.n7 VPWR.n6 604.931
R59 VPWR.n6 VPWR.t0 46.6121
R60 VPWR.n6 VPWR.t2 46.6121
R61 VPWR.n12 VPWR.n11 36.1417
R62 VPWR.n9 VPWR.n5 35.3887
R63 VPWR.n10 VPWR.n9 32.377
R64 VPWR.n12 VPWR.n1 27.8593
R65 VPWR.n0 VPWR.t6 26.3844
R66 VPWR.n0 VPWR.t7 26.3844
R67 VPWR.n3 VPWR.t4 26.3844
R68 VPWR.n3 VPWR.t5 26.3844
R69 VPWR.n4 VPWR.t1 26.3844
R70 VPWR.n4 VPWR.t3 26.3844
R71 VPWR.n14 VPWR.n1 15.9328
R72 VPWR.n9 VPWR.n8 9.3005
R73 VPWR.n11 VPWR.n2 9.3005
R74 VPWR.n13 VPWR.n12 9.3005
R75 VPWR.n7 VPWR.n5 8.09752
R76 VPWR.n11 VPWR.n10 3.76521
R77 VPWR VPWR.n14 0.773575
R78 VPWR.n8 VPWR.n7 0.435731
R79 VPWR.n14 VPWR.n13 0.14947
R80 VPWR.n8 VPWR.n2 0.122949
R81 VPWR.n13 VPWR.n2 0.122949
R82 VPB.t4 VPB.t14 592.473
R83 VPB.t7 VPB.t5 347.312
R84 VPB VPB.t3 252.823
R85 VPB.t1 VPB.t0 229.839
R86 VPB.t10 VPB.t1 229.839
R87 VPB.t15 VPB.t10 229.839
R88 VPB.t16 VPB.t15 229.839
R89 VPB.t17 VPB.t16 229.839
R90 VPB.t18 VPB.t17 229.839
R91 VPB.t19 VPB.t18 229.839
R92 VPB.t5 VPB.t19 229.839
R93 VPB.t6 VPB.t7 229.839
R94 VPB.t8 VPB.t6 229.839
R95 VPB.t11 VPB.t8 229.839
R96 VPB.t12 VPB.t11 229.839
R97 VPB.t13 VPB.t12 229.839
R98 VPB.t14 VPB.t13 229.839
R99 VPB.t9 VPB.t4 229.839
R100 VPB.t2 VPB.t9 229.839
R101 VPB.t3 VPB.t2 229.839
R102 Y.n11 Y.n10 585
R103 Y.n12 Y.n11 585
R104 Y.n11 Y.n9 585
R105 Y.n8 Y.t6 372.466
R106 Y.n1 Y.t12 308.358
R107 Y.n8 Y.n7 303.164
R108 Y.t2 Y.n14 286.887
R109 Y.n15 Y.t2 286.887
R110 Y.n1 Y.t11 275
R111 Y.n2 Y.t8 232.63
R112 Y.n4 Y.n3 209.927
R113 Y.n5 Y.n4 196.472
R114 Y.n5 Y.t4 155.638
R115 Y.n6 Y.n0 103.65
R116 Y.n2 Y.n1 65.3492
R117 Y.n6 Y.n5 58.3534
R118 Y.n13 Y.n6 58.3534
R119 Y.n9 Y.n8 57.9017
R120 Y.n4 Y.n2 50.4476
R121 Y.n11 Y.t3 26.3844
R122 Y.n7 Y.t10 26.3844
R123 Y.n7 Y.t0 26.3844
R124 Y.n3 Y.t9 22.7032
R125 Y.n3 Y.t7 22.7032
R126 Y.n0 Y.t1 22.7032
R127 Y.n0 Y.t5 22.7032
R128 Y.n12 Y 17.1525
R129 Y.n10 Y 14.8485
R130 Y.n15 Y 10.6672
R131 Y Y.n9 6.4005
R132 Y.n13 Y 4.32624
R133 Y.n14 Y.n13 4.26717
R134 Y.n14 Y 4.10306
R135 Y.n10 Y 4.0965
R136 Y Y.n12 1.7925
R137 Y Y.n15 1.47742
R138 a_534_74.n1 a_534_74.t6 276.296
R139 a_534_74.n1 a_534_74.n0 193.66
R140 a_534_74.n4 a_534_74.n3 153.802
R141 a_534_74.n3 a_534_74.n2 88.3446
R142 a_534_74.n3 a_534_74.n1 66.6668
R143 a_534_74.n2 a_534_74.t0 22.7032
R144 a_534_74.n2 a_534_74.t3 22.7032
R145 a_534_74.n0 a_534_74.t5 22.7032
R146 a_534_74.n0 a_534_74.t4 22.7032
R147 a_534_74.n4 a_534_74.t1 22.7032
R148 a_534_74.t2 a_534_74.n4 22.7032
R149 VNB.t6 VNB.t13 3187.4
R150 VNB.t3 VNB.t11 2529.13
R151 VNB.t12 VNB.t0 1986.35
R152 VNB.t14 VNB.t12 1986.35
R153 VNB.t13 VNB.t14 1986.35
R154 VNB VNB.t2 1443.57
R155 VNB.t7 VNB.t6 993.177
R156 VNB.t5 VNB.t7 993.177
R157 VNB.t8 VNB.t5 993.177
R158 VNB.t10 VNB.t8 993.177
R159 VNB.t9 VNB.t10 993.177
R160 VNB.t11 VNB.t9 993.177
R161 VNB.t1 VNB.t3 993.177
R162 VNB.t4 VNB.t1 993.177
R163 VNB.t2 VNB.t4 993.177
R164 A2.n0 A2.t0 234.72
R165 A2.n4 A2.t3 227.538
R166 A2.n2 A2.t1 226.809
R167 A2.n10 A2.t2 226.809
R168 A2.n4 A2.t7 196.013
R169 A2.n9 A2.t5 196.013
R170 A2.n3 A2.t6 196.013
R171 A2.n0 A2.t4 196.013
R172 A2 A2.n1 155.84
R173 A2.n12 A2.n11 152
R174 A2.n8 A2.n7 152
R175 A2.n6 A2.n5 152
R176 A2.n8 A2.n5 49.6611
R177 A2.n11 A2.n10 44.549
R178 A2.n1 A2.n0 29.2126
R179 A2.n2 A2.n1 28.4823
R180 A2.n11 A2.n3 16.0672
R181 A2.n7 A2.n6 12.4348
R182 A2.n5 A2.n4 10.2247
R183 A2.n12 A2 8.9605
R184 A2 A2.n12 8.59479
R185 A2.n3 A2.n2 5.11262
R186 A2.n7 A2 3.47479
R187 A2.n9 A2.n8 2.92171
R188 A2.n10 A2.n9 2.19141
R189 A2.n6 A2 1.64621
R190 B2.n4 B2.t5 234.841
R191 B2.n2 B2.t0 228.877
R192 B2.n12 B2.t1 226.809
R193 B2.n9 B2.t4 226.809
R194 B2.n2 B2.n1 196.744
R195 B2.n4 B2.t3 196.013
R196 B2.n10 B2.n3 196.013
R197 B2.n13 B2.t2 196.013
R198 B2.n15 B2.n14 152
R199 B2.n11 B2.n0 152
R200 B2.n8 B2.n7 152
R201 B2.n6 B2.n5 152
R202 B2.n8 B2.n5 49.6611
R203 B2.n11 B2.n10 39.4369
R204 B2.n14 B2.n2 35.7853
R205 B2.n14 B2.n13 26.2914
R206 B2.n12 B2.n11 21.1793
R207 B2.n6 B2 11.7586
R208 B2.n15 B2.n0 10.1214
R209 B2.n7 B2 7.5912
R210 B2.n7 B2 6.69817
R211 B2.n10 B2.n9 5.11262
R212 B2.n9 B2.n8 5.11262
R213 B2 B2.n0 3.42376
R214 B2.n5 B2.n4 2.92171
R215 B2 B2.n6 2.53073
R216 B2.n13 B2.n12 2.19141
R217 B2 B2.n15 0.744686
R218 VGND.n10 VGND.t9 239.326
R219 VGND.n11 VGND.t8 233.886
R220 VGND.n35 VGND.n2 211.183
R221 VGND.n38 VGND.n37 211.183
R222 VGND.n5 VGND.n4 204.201
R223 VGND.n30 VGND.n29 204.201
R224 VGND.n12 VGND.n9 36.1417
R225 VGND.n16 VGND.n9 36.1417
R226 VGND.n17 VGND.n16 36.1417
R227 VGND.n18 VGND.n17 36.1417
R228 VGND.n18 VGND.n7 36.1417
R229 VGND.n22 VGND.n7 36.1417
R230 VGND.n23 VGND.n22 36.1417
R231 VGND.n24 VGND.n23 36.1417
R232 VGND.n31 VGND.n1 36.1417
R233 VGND.n31 VGND.n30 31.624
R234 VGND.n12 VGND.n11 25.6005
R235 VGND.n36 VGND.n35 25.224
R236 VGND.n28 VGND.n5 24.0946
R237 VGND.n24 VGND.n5 23.3417
R238 VGND.n4 VGND.t7 22.7032
R239 VGND.n4 VGND.t5 22.7032
R240 VGND.n29 VGND.t6 22.7032
R241 VGND.n29 VGND.t4 22.7032
R242 VGND.n2 VGND.t2 22.7032
R243 VGND.n2 VGND.t0 22.7032
R244 VGND.n37 VGND.t3 22.7032
R245 VGND.n37 VGND.t1 22.7032
R246 VGND.n35 VGND.n1 22.2123
R247 VGND.n30 VGND.n28 15.8123
R248 VGND.n38 VGND.n36 14.6829
R249 VGND.n13 VGND.n12 9.3005
R250 VGND.n14 VGND.n9 9.3005
R251 VGND.n16 VGND.n15 9.3005
R252 VGND.n17 VGND.n8 9.3005
R253 VGND.n19 VGND.n18 9.3005
R254 VGND.n20 VGND.n7 9.3005
R255 VGND.n22 VGND.n21 9.3005
R256 VGND.n23 VGND.n6 9.3005
R257 VGND.n25 VGND.n24 9.3005
R258 VGND.n26 VGND.n5 9.3005
R259 VGND.n28 VGND.n27 9.3005
R260 VGND.n30 VGND.n3 9.3005
R261 VGND.n32 VGND.n31 9.3005
R262 VGND.n33 VGND.n1 9.3005
R263 VGND.n35 VGND.n34 9.3005
R264 VGND.n36 VGND.n0 9.3005
R265 VGND.n39 VGND.n38 7.59866
R266 VGND.n11 VGND.n10 6.50541
R267 VGND.n13 VGND.n10 0.648193
R268 VGND VGND.n39 0.162259
R269 VGND.n39 VGND.n0 0.145572
R270 VGND.n14 VGND.n13 0.122949
R271 VGND.n15 VGND.n14 0.122949
R272 VGND.n15 VGND.n8 0.122949
R273 VGND.n19 VGND.n8 0.122949
R274 VGND.n20 VGND.n19 0.122949
R275 VGND.n21 VGND.n20 0.122949
R276 VGND.n21 VGND.n6 0.122949
R277 VGND.n25 VGND.n6 0.122949
R278 VGND.n26 VGND.n25 0.122949
R279 VGND.n27 VGND.n26 0.122949
R280 VGND.n27 VGND.n3 0.122949
R281 VGND.n32 VGND.n3 0.122949
R282 VGND.n33 VGND.n32 0.122949
R283 VGND.n34 VGND.n33 0.122949
R284 VGND.n34 VGND.n0 0.122949
R285 a_1326_74.n0 a_1326_74.t0 326.824
R286 a_1326_74.n0 a_1326_74.t1 281.43
R287 a_1326_74.t3 a_1326_74.n1 233.337
R288 a_1326_74.n1 a_1326_74.t2 134.165
R289 a_1326_74.n1 a_1326_74.n0 55.5209
R290 C1.n5 C1.t5 244.214
R291 C1.n0 C1.t0 226.809
R292 C1.n3 C1.t1 226.809
R293 C1.n4 C1.t2 226.809
R294 C1.n0 C1.t6 198.228
R295 C1.n5 C1.t4 186.374
R296 C1.n10 C1.t7 186.374
R297 C1.n2 C1.t3 186.374
R298 C1 C1.n1 155.423
R299 C1.n12 C1.n11 152
R300 C1.n9 C1.n8 152
R301 C1.n7 C1.n6 152
R302 C1.n11 C1.n10 42.1755
R303 C1.n6 C1.n4 34.1422
R304 C1.n2 C1.n1 30.1255
R305 C1.n1 C1.n0 18.0755
R306 C1.n3 C1.n2 12.0505
R307 C1.n9 C1.n4 11.3811
R308 C1.n8 C1.n7 10.1214
R309 C1.n6 C1.n5 8.70328
R310 C1.n12 C1 7.5912
R311 C1 C1.n12 6.69817
R312 C1.n11 C1.n3 3.34772
R313 C1.n10 C1.n9 3.34772
R314 C1.n8 C1 2.53073
R315 C1.n7 C1 1.63771
R316 a_114_368.n8 a_114_368.n6 388.519
R317 a_114_368.n8 a_114_368.n7 348.938
R318 a_114_368.n2 a_114_368.n0 340.983
R319 a_114_368.n9 a_114_368.n8 299.76
R320 a_114_368.n2 a_114_368.n1 298.065
R321 a_114_368.n4 a_114_368.n3 298.065
R322 a_114_368.n6 a_114_368.n5 298.065
R323 a_114_368.n4 a_114_368.n2 42.9181
R324 a_114_368.n6 a_114_368.n4 42.9181
R325 a_114_368.n7 a_114_368.t1 26.3844
R326 a_114_368.n7 a_114_368.t0 26.3844
R327 a_114_368.n0 a_114_368.t11 26.3844
R328 a_114_368.n0 a_114_368.t10 26.3844
R329 a_114_368.n1 a_114_368.t9 26.3844
R330 a_114_368.n1 a_114_368.t8 26.3844
R331 a_114_368.n3 a_114_368.t4 26.3844
R332 a_114_368.n3 a_114_368.t5 26.3844
R333 a_114_368.n5 a_114_368.t6 26.3844
R334 a_114_368.n5 a_114_368.t7 26.3844
R335 a_114_368.t3 a_114_368.n9 26.3844
R336 a_114_368.n9 a_114_368.t2 26.3844
R337 B1.n7 B1.t5 237.762
R338 B1.n1 B1.t2 226.809
R339 B1.n4 B1.t3 226.809
R340 B1.n11 B1.t4 226.809
R341 B1.n1 B1.n0 210.138
R342 B1.n6 B1.t0 196.013
R343 B1.n12 B1.n5 196.013
R344 B1.n3 B1.t1 196.013
R345 B1 B1.n2 154.828
R346 B1.n14 B1.n13 152
R347 B1.n10 B1.n9 152
R348 B1.n8 B1.n7 152
R349 B1.n10 B1.n6 40.8975
R350 B1.n2 B1.n1 37.246
R351 B1.n13 B1.n12 27.752
R352 B1.n13 B1.n4 21.1793
R353 B1.n12 B1.n11 16.7975
R354 B1.n3 B1.n2 14.6066
R355 B1.n4 B1.n3 13.8763
R356 B1.n9 B1.n8 10.1214
R357 B1.n7 B1.n6 8.76414
R358 B1 B1.n14 7.29352
R359 B1.n14 B1 6.99585
R360 B1.n11 B1.n10 5.11262
R361 B1.n9 B1 3.12608
R362 B1.n8 B1 1.04236
C0 A1 Y 0.217819f
C1 C1 VGND 0.072097f
C2 B1 B2 0.102714f
C3 A2 VPWR 0.053887f
C4 B1 Y 0.185897f
C5 A1 VPWR 0.058903f
C6 A2 VGND 0.058234f
C7 B2 Y 1.12e-19
C8 B1 VPWR 0.024575f
C9 A1 VGND 0.028481f
C10 VPB C1 0.144f
C11 B2 VPWR 0.025067f
C12 B1 VGND 0.02633f
C13 VPB A2 0.143157f
C14 B2 VGND 0.073256f
C15 Y VPWR 0.264462f
C16 C1 A2 0.052155f
C17 VPB A1 0.15287f
C18 Y VGND 0.393532f
C19 VPB B1 0.135495f
C20 C1 A1 1.95e-19
C21 VPWR VGND 0.163412f
C22 VPB B2 0.138198f
C23 C1 B1 4.15e-19
C24 A2 A1 0.092164f
C25 VPB Y 0.034612f
C26 A2 B1 2.3e-19
C27 VPB VPWR 0.238845f
C28 C1 Y 0.289729f
C29 A1 B1 0.081012f
C30 C1 VPWR 0.024819f
C31 A2 Y 0.230511f
C32 VPB VGND 0.012054f
C33 VGND VNB 1.19689f
C34 VPWR VNB 0.935787f
C35 Y VNB 0.1993f
C36 B2 VNB 0.435091f
C37 B1 VNB 0.402438f
C38 A1 VNB 0.423908f
C39 A2 VNB 0.409297f
C40 C1 VNB 0.439158f
C41 VPB VNB 2.44181f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a311oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311oi_2 VNB VPB VGND VPWR Y C1 B1 A3 A2 A1
X0 VGND.t1 A3.t0 a_45_74.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X1 VPWR.t4 A1.t0 a_127_368.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_127_368.t5 A1.t1 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1848 ps=1.45 w=1.12 l=0.15
X3 VPWR.t5 A2.t0 a_127_368.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_300_74.t1 A2.t1 a_45_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_127_368.t1 A2.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VGND.t3 B1.t0 Y.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=1.43 as=0.1036 ps=1.02 w=0.74 l=0.15
X7 Y.t2 C1.t0 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.2553 ps=1.43 w=0.74 l=0.15
X8 VPWR.t2 A3.t1 a_127_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_45_74.t0 A2.t3 a_300_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_300_74.t2 A1.t2 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X11 Y.t0 C1.t1 a_692_368.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_692_368.t3 B1.t1 a_127_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X13 a_692_368.t0 C1.t2 Y.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_45_74.t2 A3.t2 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 a_127_368.t4 B1.t2 a_692_368.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X16 Y.t3 A1.t3 a_300_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_127_368.t2 A3.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
R0 A3.n1 A3.t3 262.349
R1 A3.n0 A3.t1 261.62
R2 A3.n3 A3.n2 157.786
R3 A3.n0 A3.t2 154.24
R4 A3.n1 A3.t0 154.24
R5 A3.n2 A3.n0 52.5823
R6 A3.n3 A3 27.2005
R7 A3.n2 A3.n1 10.2247
R8 A3 A3.n3 0.351185
R9 a_45_74.t0 a_45_74.n1 252.312
R10 a_45_74.n1 a_45_74.t3 196.292
R11 a_45_74.n1 a_45_74.n0 97.4026
R12 a_45_74.n0 a_45_74.t1 22.7032
R13 a_45_74.n0 a_45_74.t2 22.7032
R14 VGND.n2 VGND.n0 212.127
R15 VGND.n2 VGND.n1 97.9919
R16 VGND.n1 VGND.t2 50.8833
R17 VGND.n1 VGND.t3 50.8833
R18 VGND.n0 VGND.t0 22.7032
R19 VGND.n0 VGND.t1 22.7032
R20 VGND VGND.n2 0.198128
R21 VNB.t0 VNB.t4 2494.49
R22 VNB.t7 VNB.t5 1940.16
R23 VNB VNB.t3 1304.99
R24 VNB.t6 VNB.t7 993.177
R25 VNB.t4 VNB.t6 993.177
R26 VNB.t1 VNB.t0 993.177
R27 VNB.t2 VNB.t1 993.177
R28 VNB.t3 VNB.t2 993.177
R29 A1.n0 A1.t3 273.134
R30 A1.n3 A1.t1 236.321
R31 A1.n2 A1.t0 226.809
R32 A1 A1.n3 182.833
R33 A1.n1 A1.t2 179.947
R34 A1 A1.n0 152
R35 A1.n3 A1.n2 47.5663
R36 A1.n1 A1.n0 13.1652
R37 A1.n2 A1.n1 12.0505
R38 a_127_368.n5 a_127_368.n4 403.668
R39 a_127_368.n2 a_127_368.n0 253.62
R40 a_127_368.n2 a_127_368.n1 210.702
R41 a_127_368.n4 a_127_368.n3 207.35
R42 a_127_368.n4 a_127_368.n2 62.1181
R43 a_127_368.n3 a_127_368.t6 26.3844
R44 a_127_368.n3 a_127_368.t5 26.3844
R45 a_127_368.n0 a_127_368.t3 26.3844
R46 a_127_368.n0 a_127_368.t2 26.3844
R47 a_127_368.n1 a_127_368.t7 26.3844
R48 a_127_368.n1 a_127_368.t1 26.3844
R49 a_127_368.t0 a_127_368.n5 26.3844
R50 a_127_368.n5 a_127_368.t4 26.3844
R51 VPWR.n3 VPWR.t4 348.277
R52 VPWR.n2 VPWR.n1 335.577
R53 VPWR.n5 VPWR.n4 322.635
R54 VPWR.n11 VPWR.t1 259.171
R55 VPWR.n10 VPWR.n9 36.1417
R56 VPWR.n6 VPWR.n2 33.5064
R57 VPWR.n4 VPWR.t3 29.0228
R58 VPWR.n4 VPWR.t5 29.0228
R59 VPWR.n6 VPWR.n5 27.8593
R60 VPWR.n1 VPWR.t0 26.3844
R61 VPWR.n1 VPWR.t2 26.3844
R62 VPWR.n11 VPWR.n10 22.5887
R63 VPWR.n7 VPWR.n6 9.3005
R64 VPWR.n9 VPWR.n8 9.3005
R65 VPWR.n10 VPWR.n0 9.3005
R66 VPWR.n12 VPWR.n11 9.3005
R67 VPWR.n5 VPWR.n3 6.64362
R68 VPWR.n9 VPWR.n2 2.63579
R69 VPWR.n7 VPWR.n3 0.601517
R70 VPWR.n8 VPWR.n7 0.122949
R71 VPWR.n8 VPWR.n0 0.122949
R72 VPWR.n12 VPWR.n0 0.122949
R73 VPWR VPWR.n12 0.0617245
R74 VPB.t7 VPB.t5 495.43
R75 VPB VPB.t2 286.022
R76 VPB.t8 VPB.t6 245.161
R77 VPB.t4 VPB.t9 229.839
R78 VPB.t0 VPB.t4 229.839
R79 VPB.t5 VPB.t0 229.839
R80 VPB.t6 VPB.t7 229.839
R81 VPB.t1 VPB.t8 229.839
R82 VPB.t3 VPB.t1 229.839
R83 VPB.t2 VPB.t3 229.839
R84 A2.n0 A2.t0 261.62
R85 A2.n2 A2.t2 261.62
R86 A2.n4 A2.n0 169.319
R87 A2.n2 A2.t1 159.4
R88 A2.n1 A2.t3 154.24
R89 A2.n4 A2.n3 152
R90 A2.n3 A2.n1 46.7399
R91 A2.n5 A2 27.2005
R92 A2.n5 A2.n4 12.9944
R93 A2.n3 A2.n2 10.955
R94 A2.n1 A2.n0 8.03383
R95 A2 A2.n5 3.29747
R96 a_300_74.n1 a_300_74.n0 445.264
R97 a_300_74.n0 a_300_74.t3 22.7032
R98 a_300_74.n0 a_300_74.t2 22.7032
R99 a_300_74.n1 a_300_74.t0 22.7032
R100 a_300_74.t1 a_300_74.n1 22.7032
R101 B1.n3 B1.t1 237.762
R102 B1.n0 B1.t2 226.809
R103 B1.n0 B1.t0 198.204
R104 B1.n4 B1.n3 152
R105 B1.n2 B1.n1 152
R106 B1.n3 B1.n2 49.6611
R107 B1.n1 B1 9.82376
R108 B1 B1.n4 8.63306
R109 B1.n4 B1 5.65631
R110 B1.n2 B1.n0 5.11262
R111 B1.n1 B1 4.46562
R112 Y Y.n0 361.442
R113 Y.n2 Y.t4 314.192
R114 Y.n3 Y.t2 143.445
R115 Y.n2 Y.n1 96.2135
R116 Y.n3 Y.n2 78.9774
R117 Y.n0 Y.t5 26.3844
R118 Y.n0 Y.t0 26.3844
R119 Y.n1 Y.t1 22.7032
R120 Y.n1 Y.t3 22.7032
R121 Y Y.n3 9.02219
R122 C1.n1 C1.t2 248.718
R123 C1.n0 C1.t1 226.809
R124 C1.n0 C1.t0 206.969
R125 C1 C1.n1 154.522
R126 C1.n1 C1.n0 43.8187
R127 a_692_368.n0 a_692_368.t2 372.601
R128 a_692_368.n0 a_692_368.t0 372.325
R129 a_692_368.n1 a_692_368.n0 209.542
R130 a_692_368.t1 a_692_368.n1 26.3844
R131 a_692_368.n1 a_692_368.t3 26.3844
C0 A3 Y 2.07e-19
C1 A2 VPWR 0.037573f
C2 VPB VGND 0.009754f
C3 B1 C1 0.098458f
C4 A2 Y 0.002219f
C5 A3 VGND 0.031641f
C6 A1 VPWR 0.045783f
C7 A2 VGND 0.017797f
C8 B1 VPWR 0.013159f
C9 A1 Y 0.087031f
C10 B1 Y 0.117708f
C11 A1 VGND 0.01865f
C12 C1 VPWR 0.0111f
C13 VPB A3 0.06054f
C14 B1 VGND 0.023154f
C15 C1 Y 0.14008f
C16 VPB A2 0.06095f
C17 C1 VGND 0.016422f
C18 VPWR Y 0.015896f
C19 VPB A1 0.088467f
C20 A3 A2 0.087653f
C21 VPWR VGND 0.093284f
C22 VPB B1 0.069462f
C23 A3 A1 2.39e-19
C24 Y VGND 0.299853f
C25 A2 A1 0.063059f
C26 VPB C1 0.066678f
C27 A2 B1 1.24e-19
C28 VPB VPWR 0.163127f
C29 A2 C1 5.99e-20
C30 A1 B1 0.07502f
C31 A3 VPWR 0.037845f
C32 VPB Y 0.012064f
C33 VGND VNB 0.687576f
C34 Y VNB 0.135727f
C35 VPWR VNB 0.586594f
C36 C1 VNB 0.191885f
C37 B1 VNB 0.166463f
C38 A1 VNB 0.252564f
C39 A2 VNB 0.215551f
C40 A3 VNB 0.234176f
C41 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a311oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311oi_4 VNB VPB VPWR VGND Y C1 B1 A3 A2 A1
X0 VPWR.t5 A2.t0 a_114_368.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_1213_368.t4 B1.t0 a_114_368.t15 VPB.t18 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_114_368.t8 B1.t1 a_1213_368.t3 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X3 a_114_368.t4 A2.t1 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_465_74.t3 A2.t2 a_34_74.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VPWR.t3 A2.t3 a_114_368.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_114_368.t2 A2.t4 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 Y.t3 A1.t0 a_465_74.t4 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 VPWR.t6 A3.t0 a_114_368.t6 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VGND.t6 A3.t1 a_34_74.t7 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_114_368.t0 A3.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t1 A3.t3 a_114_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_34_74.t0 A3.t4 VGND.t5 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_465_74.t5 A1.t1 Y.t2 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_1213_368.t7 C1.t0 Y.t9 VPB.t19 sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_34_74.t5 A3.t5 VGND.t4 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_465_74.t6 A1.t2 Y.t1 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X17 VGND.t3 A3.t6 a_34_74.t6 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_114_368.t9 A1.t3 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 VPWR.t9 A1.t4 a_114_368.t10 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 VPWR.t10 A1.t5 a_114_368.t11 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X22 a_114_368.t7 A3.t7 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X23 a_34_74.t3 A2.t5 a_465_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 Y.t4 C1.t1 a_1213_368.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X25 a_34_74.t2 A2.t6 a_465_74.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 VGND.t2 B1.t2 Y.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.4181 pd=1.87 as=0.1036 ps=1.02 w=0.74 l=0.15
X27 a_1213_368.t5 C1.t2 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X28 Y.t0 C1.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X29 Y.t8 C1.t4 a_1213_368.t6 VPB.t17 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X30 a_1213_368.t2 B1.t3 a_114_368.t13 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X31 Y.t5 B1.t4 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.4181 ps=1.87 w=0.74 l=0.15
X32 a_114_368.t14 B1.t5 a_1213_368.t1 VPB.t16 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X33 a_465_74.t0 A2.t7 a_34_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X34 a_114_368.t12 A1.t6 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A2.n1 A2.t0 242.144
R1 A2.n11 A2.t1 226.809
R2 A2.n8 A2.t3 226.809
R3 A2.n3 A2.t4 226.809
R4 A2.n3 A2.t2 203.762
R5 A2.n2 A2.t6 196.013
R6 A2.n10 A2.t7 196.013
R7 A2.n1 A2.t5 196.013
R8 A2.n13 A2.n12 152
R9 A2.n9 A2.n0 152
R10 A2.n7 A2.n6 152
R11 A2.n5 A2.n4 152
R12 A2.n4 A2.n2 45.2793
R13 A2.n9 A2.n8 44.549
R14 A2.n12 A2.n11 28.4823
R15 A2.n12 A2.n1 21.9096
R16 A2.n11 A2.n10 12.4157
R17 A2.n4 A2.n3 10.955
R18 A2.n13 A2.n0 10.1214
R19 A2.n6 A2 9.67492
R20 A2.n5 A2 8.7819
R21 A2.n10 A2.n9 8.76414
R22 A2 A2.n5 5.50748
R23 A2.n8 A2.n7 5.11262
R24 A2.n6 A2 4.61445
R25 A2.n7 A2.n2 4.38232
R26 A2 A2.n13 3.72143
R27 A2 A2.n0 0.447012
R28 a_114_368.n5 a_114_368.n4 333.139
R29 a_114_368.n5 a_114_368.n3 298.229
R30 a_114_368.n12 a_114_368.n11 270.142
R31 a_114_368.n10 a_114_368.n0 208.897
R32 a_114_368.n9 a_114_368.n1 208.897
R33 a_114_368.n13 a_114_368.n12 208.897
R34 a_114_368.n7 a_114_368.n6 208.776
R35 a_114_368.n8 a_114_368.n2 207.35
R36 a_114_368.n7 a_114_368.n5 94.4946
R37 a_114_368.n9 a_114_368.n8 67.7652
R38 a_114_368.n10 a_114_368.n9 67.7652
R39 a_114_368.n12 a_114_368.n10 67.7652
R40 a_114_368.n8 a_114_368.n7 55.3417
R41 a_114_368.n0 a_114_368.t3 26.3844
R42 a_114_368.n0 a_114_368.t2 26.3844
R43 a_114_368.n1 a_114_368.t5 26.3844
R44 a_114_368.n1 a_114_368.t4 26.3844
R45 a_114_368.n2 a_114_368.t10 26.3844
R46 a_114_368.n2 a_114_368.t12 26.3844
R47 a_114_368.n11 a_114_368.t1 26.3844
R48 a_114_368.n11 a_114_368.t7 26.3844
R49 a_114_368.n3 a_114_368.t15 26.3844
R50 a_114_368.n3 a_114_368.t8 26.3844
R51 a_114_368.n4 a_114_368.t13 26.3844
R52 a_114_368.n4 a_114_368.t14 26.3844
R53 a_114_368.n6 a_114_368.t11 26.3844
R54 a_114_368.n6 a_114_368.t9 26.3844
R55 a_114_368.n13 a_114_368.t6 26.3844
R56 a_114_368.t0 a_114_368.n13 26.3844
R57 VPWR.n11 VPWR.t10 346.786
R58 VPWR.n12 VPWR.n10 323.406
R59 VPWR.n24 VPWR.n2 315.928
R60 VPWR.n4 VPWR.n3 315.928
R61 VPWR.n18 VPWR.n6 315.928
R62 VPWR.n8 VPWR.n7 315.928
R63 VPWR.n26 VPWR.t7 259.171
R64 VPWR.n14 VPWR.n13 36.1417
R65 VPWR.n18 VPWR.n17 35.0123
R66 VPWR.n19 VPWR.n4 30.4946
R67 VPWR.n26 VPWR.n25 27.4829
R68 VPWR.n2 VPWR.t0 26.3844
R69 VPWR.n2 VPWR.t1 26.3844
R70 VPWR.n3 VPWR.t2 26.3844
R71 VPWR.n3 VPWR.t6 26.3844
R72 VPWR.n6 VPWR.t4 26.3844
R73 VPWR.n6 VPWR.t3 26.3844
R74 VPWR.n7 VPWR.t11 26.3844
R75 VPWR.n7 VPWR.t5 26.3844
R76 VPWR.n10 VPWR.t8 26.3844
R77 VPWR.n10 VPWR.t9 26.3844
R78 VPWR.n24 VPWR.n23 25.977
R79 VPWR.n25 VPWR.n24 21.4593
R80 VPWR.n12 VPWR.n11 20.3395
R81 VPWR.n23 VPWR.n4 16.9417
R82 VPWR.n19 VPWR.n18 12.424
R83 VPWR.n13 VPWR.n9 9.3005
R84 VPWR.n15 VPWR.n14 9.3005
R85 VPWR.n17 VPWR.n16 9.3005
R86 VPWR.n18 VPWR.n5 9.3005
R87 VPWR.n20 VPWR.n19 9.3005
R88 VPWR.n21 VPWR.n4 9.3005
R89 VPWR.n23 VPWR.n22 9.3005
R90 VPWR.n24 VPWR.n1 9.3005
R91 VPWR.n25 VPWR.n0 9.3005
R92 VPWR.n27 VPWR.n26 9.3005
R93 VPWR.n17 VPWR.n8 7.90638
R94 VPWR.n13 VPWR.n12 3.38874
R95 VPWR.n14 VPWR.n8 3.38874
R96 VPWR.n11 VPWR.n9 1.31197
R97 VPWR.n15 VPWR.n9 0.122949
R98 VPWR.n16 VPWR.n15 0.122949
R99 VPWR.n16 VPWR.n5 0.122949
R100 VPWR.n20 VPWR.n5 0.122949
R101 VPWR.n21 VPWR.n20 0.122949
R102 VPWR.n22 VPWR.n21 0.122949
R103 VPWR.n22 VPWR.n1 0.122949
R104 VPWR.n1 VPWR.n0 0.122949
R105 VPWR.n27 VPWR.n0 0.122949
R106 VPWR VPWR.n27 0.0617245
R107 VPB.t13 VPB.t10 495.43
R108 VPB VPB.t9 252.823
R109 VPB.t2 VPB.t19 229.839
R110 VPB.t7 VPB.t2 229.839
R111 VPB.t17 VPB.t7 229.839
R112 VPB.t15 VPB.t17 229.839
R113 VPB.t16 VPB.t15 229.839
R114 VPB.t18 VPB.t16 229.839
R115 VPB.t10 VPB.t18 229.839
R116 VPB.t11 VPB.t13 229.839
R117 VPB.t12 VPB.t11 229.839
R118 VPB.t14 VPB.t12 229.839
R119 VPB.t6 VPB.t14 229.839
R120 VPB.t5 VPB.t6 229.839
R121 VPB.t4 VPB.t5 229.839
R122 VPB.t3 VPB.t4 229.839
R123 VPB.t8 VPB.t3 229.839
R124 VPB.t0 VPB.t8 229.839
R125 VPB.t1 VPB.t0 229.839
R126 VPB.t9 VPB.t1 229.839
R127 B1.n1 B1.t3 242.375
R128 B1.n5 B1.t1 237.032
R129 B1.n3 B1.t5 234.841
R130 B1.n6 B1.t0 234.841
R131 B1.n5 B1.t2 186.374
R132 B1.n1 B1.t4 186.374
R133 B1.n2 B1 159.969
R134 B1.n4 B1.n0 152
R135 B1.n8 B1.n7 152
R136 B1.n6 B1.n5 63.5369
R137 B1.n7 B1.n4 49.6611
R138 B1.n3 B1.n2 44.549
R139 B1.n2 B1.n1 13.146
R140 B1.n7 B1.n6 10.955
R141 B1.n8 B1.n0 9.26007
R142 B1.n4 B1.n3 5.11262
R143 B1 B1.n0 2.04305
R144 B1 B1.n8 1.77071
R145 a_1213_368.n4 a_1213_368.t3 372.512
R146 a_1213_368.n1 a_1213_368.n0 304.901
R147 a_1213_368.n5 a_1213_368.n4 303.212
R148 a_1213_368.n1 a_1213_368.t7 279.81
R149 a_1213_368.n3 a_1213_368.n2 210.508
R150 a_1213_368.n3 a_1213_368.n1 42.9181
R151 a_1213_368.n4 a_1213_368.n3 42.9181
R152 a_1213_368.n0 a_1213_368.t0 26.3844
R153 a_1213_368.n0 a_1213_368.t5 26.3844
R154 a_1213_368.n2 a_1213_368.t6 26.3844
R155 a_1213_368.n2 a_1213_368.t2 26.3844
R156 a_1213_368.n5 a_1213_368.t1 26.3844
R157 a_1213_368.t4 a_1213_368.n5 26.3844
R158 a_34_74.n1 a_34_74.t3 323.49
R159 a_34_74.n3 a_34_74.t6 197.988
R160 a_34_74.n1 a_34_74.n0 185
R161 a_34_74.n3 a_34_74.n2 104.579
R162 a_34_74.n5 a_34_74.n4 101.014
R163 a_34_74.n4 a_34_74.n3 57.2608
R164 a_34_74.n4 a_34_74.n1 48.5468
R165 a_34_74.n2 a_34_74.t7 22.7032
R166 a_34_74.n2 a_34_74.t5 22.7032
R167 a_34_74.n0 a_34_74.t1 22.7032
R168 a_34_74.n0 a_34_74.t2 22.7032
R169 a_34_74.n5 a_34_74.t4 22.7032
R170 a_34_74.t0 a_34_74.n5 22.7032
R171 a_465_74.n1 a_465_74.t5 323.413
R172 a_465_74.n4 a_465_74.n3 227.853
R173 a_465_74.n1 a_465_74.n0 185
R174 a_465_74.n3 a_465_74.n2 185
R175 a_465_74.n3 a_465_74.n1 81.9205
R176 a_465_74.n2 a_465_74.t2 22.7032
R177 a_465_74.n2 a_465_74.t0 22.7032
R178 a_465_74.n0 a_465_74.t4 22.7032
R179 a_465_74.n0 a_465_74.t6 22.7032
R180 a_465_74.n4 a_465_74.t1 22.7032
R181 a_465_74.t3 a_465_74.n4 22.7032
R182 VNB.t7 VNB.t6 2956.43
R183 VNB.t4 VNB.t12 2702.36
R184 VNB.t6 VNB.t0 1986.35
R185 VNB.t9 VNB.t7 1986.35
R186 VNB VNB.t11 1224.15
R187 VNB.t8 VNB.t9 993.177
R188 VNB.t12 VNB.t8 993.177
R189 VNB.t2 VNB.t4 993.177
R190 VNB.t3 VNB.t2 993.177
R191 VNB.t5 VNB.t3 993.177
R192 VNB.t1 VNB.t5 993.177
R193 VNB.t13 VNB.t1 993.177
R194 VNB.t10 VNB.t13 993.177
R195 VNB.t11 VNB.t10 993.177
R196 A1.n4 A1.t6 352.111
R197 A1.n9 A1.t5 226.809
R198 A1.n3 A1.t3 226.809
R199 A1.n11 A1.n1 209.16
R200 A1.n4 A1.t4 204.048
R201 A1.n10 A1.t1 196.013
R202 A1.n5 A1.t2 196.013
R203 A1.n2 A1.t0 196.013
R204 A1.n7 A1.n6 163.907
R205 A1.n12 A1.n11 152
R206 A1.n10 A1.n0 152
R207 A1.n8 A1.n7 152
R208 A1.n11 A1.n10 49.6611
R209 A1.n9 A1.n8 35.7853
R210 A1.n5 A1.n4 29.4146
R211 A1.n6 A1.n3 28.4823
R212 A1.n3 A1.n2 21.1793
R213 A1.n10 A1.n9 18.2581
R214 A1.n6 A1.n5 13.146
R215 A1.n12 A1.n0 10.1214
R216 A1.n8 A1.n2 8.76414
R217 A1.n7 A1 6.99585
R218 A1 A1.n0 4.0191
R219 A1 A1.n12 0.149337
R220 Y.n2 Y.n1 378.031
R221 Y.n4 Y.t1 317.733
R222 Y.n2 Y.n0 310.265
R223 Y.n4 Y.n3 185
R224 Y.n5 Y.t6 145.266
R225 Y.n6 Y.t5 137.635
R226 Y.n7 Y.t0 135.529
R227 Y.n6 Y.n5 104.963
R228 Y.n7 Y.n6 53.6019
R229 Y.n8 Y.n2 53.4593
R230 Y.n5 Y.n4 37.6933
R231 Y.n0 Y.t9 26.3844
R232 Y.n0 Y.t4 26.3844
R233 Y.n1 Y.t7 26.3844
R234 Y.n1 Y.t8 26.3844
R235 Y.n3 Y.t2 22.7032
R236 Y.n3 Y.t3 22.7032
R237 Y.n9 Y 13.2005
R238 Y Y.n9 6.0005
R239 Y.n9 Y.n8 1.64898
R240 Y.n8 Y 1.26111
R241 Y Y.n7 0.194439
R242 A3.n6 A3.t7 231.921
R243 A3.n0 A3.t0 230.459
R244 A3.n2 A3.t2 226.809
R245 A3.n5 A3.t3 226.809
R246 A3.n6 A3.t6 196.013
R247 A3.n4 A3.t5 196.013
R248 A3.n3 A3.t1 196.013
R249 A3.n0 A3.t4 196.013
R250 A3 A3.n1 155.423
R251 A3.n12 A3.n11 152
R252 A3.n10 A3.n9 152
R253 A3.n8 A3.n7 152
R254 A3.n11 A3.n10 49.6611
R255 A3.n2 A3.n1 46.0096
R256 A3.n7 A3.n5 37.246
R257 A3.n7 A3.n6 23.3702
R258 A3.n1 A3.n0 16.0672
R259 A3.n10 A3.n4 10.2247
R260 A3.n9 A3.n8 10.1214
R261 A3.n12 A3 7.5912
R262 A3 A3.n12 6.69817
R263 A3.n11 A3.n3 2.92171
R264 A3.n9 A3 2.53073
R265 A3.n5 A3.n4 2.19141
R266 A3.n8 A3 1.63771
R267 A3.n3 A3.n2 0.730803
R268 VGND.n10 VGND.t0 293.336
R269 VGND.n35 VGND.n34 219.56
R270 VGND.n32 VGND.n2 211.183
R271 VGND.n15 VGND.n14 185
R272 VGND.n13 VGND.n12 185
R273 VGND.n11 VGND.n9 185
R274 VGND.n13 VGND.n9 57.5681
R275 VGND.n14 VGND.n13 57.5681
R276 VGND.n16 VGND.n6 36.1417
R277 VGND.n20 VGND.n6 36.1417
R278 VGND.n21 VGND.n20 36.1417
R279 VGND.n22 VGND.n21 36.1417
R280 VGND.n22 VGND.n4 36.1417
R281 VGND.n26 VGND.n4 36.1417
R282 VGND.n27 VGND.n26 36.1417
R283 VGND.n28 VGND.n27 36.1417
R284 VGND.n28 VGND.n1 36.1417
R285 VGND.n9 VGND.t1 34.0546
R286 VGND.n14 VGND.t2 34.0546
R287 VGND.n32 VGND.n1 29.3652
R288 VGND.n35 VGND.n33 27.8593
R289 VGND.n2 VGND.t5 22.7032
R290 VGND.n2 VGND.t6 22.7032
R291 VGND.n34 VGND.t4 22.7032
R292 VGND.n34 VGND.t3 22.7032
R293 VGND.n33 VGND.n32 18.0711
R294 VGND.n8 VGND.n7 9.3005
R295 VGND.n17 VGND.n16 9.3005
R296 VGND.n18 VGND.n6 9.3005
R297 VGND.n20 VGND.n19 9.3005
R298 VGND.n21 VGND.n5 9.3005
R299 VGND.n23 VGND.n22 9.3005
R300 VGND.n24 VGND.n4 9.3005
R301 VGND.n26 VGND.n25 9.3005
R302 VGND.n27 VGND.n3 9.3005
R303 VGND.n29 VGND.n28 9.3005
R304 VGND.n30 VGND.n1 9.3005
R305 VGND.n32 VGND.n31 9.3005
R306 VGND.n33 VGND.n0 9.3005
R307 VGND.n16 VGND.n15 8.06844
R308 VGND.n36 VGND.n35 7.32393
R309 VGND.n11 VGND.n10 7.15613
R310 VGND.n12 VGND.n11 6.01904
R311 VGND.n15 VGND.n8 4.15414
R312 VGND.n12 VGND.n8 1.8654
R313 VGND.n10 VGND.n7 0.547153
R314 VGND VGND.n36 0.158642
R315 VGND.n36 VGND.n0 0.149142
R316 VGND.n17 VGND.n7 0.122949
R317 VGND.n18 VGND.n17 0.122949
R318 VGND.n19 VGND.n18 0.122949
R319 VGND.n19 VGND.n5 0.122949
R320 VGND.n23 VGND.n5 0.122949
R321 VGND.n24 VGND.n23 0.122949
R322 VGND.n25 VGND.n24 0.122949
R323 VGND.n25 VGND.n3 0.122949
R324 VGND.n29 VGND.n3 0.122949
R325 VGND.n30 VGND.n29 0.122949
R326 VGND.n31 VGND.n30 0.122949
R327 VGND.n31 VGND.n0 0.122949
R328 C1.n1 C1.t0 365.596
R329 C1.n1 C1.t1 261.62
R330 C1.n3 C1.t2 261.62
R331 C1.n6 C1.t4 261.62
R332 C1.n6 C1.n5 165.196
R333 C1.n2 C1 155.978
R334 C1 C1.n7 155.172
R335 C1.n4 C1.t3 154.24
R336 C1.n4 C1.n0 152
R337 C1.n7 C1.n4 49.6611
R338 C1.n3 C1.n2 35.7853
R339 C1.n2 C1.n1 29.9429
R340 C1.n4 C1.n3 13.8763
R341 C1 C1.n0 8.82212
R342 C1 C1.n0 7.78428
R343 C1.n7 C1.n6 2.19141
C0 A1 Y 0.155651f
C1 B1 VPWR 0.023159f
C2 A2 VGND 0.027852f
C3 B1 Y 0.121637f
C4 C1 VPWR 0.022955f
C5 A1 VGND 0.027907f
C6 VPB A3 0.13699f
C7 C1 Y 0.283657f
C8 B1 VGND 0.041805f
C9 VPB A2 0.134854f
C10 C1 VGND 0.040168f
C11 VPWR Y 0.021696f
C12 A3 A2 0.096361f
C13 VPB A1 0.167912f
C14 VPWR VGND 0.160884f
C15 VPB B1 0.134176f
C16 Y VGND 0.48984f
C17 A2 A1 0.048092f
C18 A3 B1 5.78e-20
C19 VPB C1 0.127835f
C20 VPB VPWR 0.250219f
C21 A2 B1 1.22e-19
C22 A1 B1 0.067111f
C23 A3 VPWR 0.082012f
C24 VPB Y 0.012008f
C25 A1 C1 1.42e-19
C26 VPB VGND 0.011868f
C27 A3 Y 8.22e-21
C28 A2 VPWR 0.075479f
C29 A2 Y 1.59e-19
C30 A1 VPWR 0.068472f
C31 A3 VGND 0.069271f
C32 B1 C1 0.078556f
C33 VGND VNB 1.14484f
C34 Y VNB 0.133251f
C35 VPWR VNB 0.950616f
C36 C1 VNB 0.378133f
C37 B1 VNB 0.343123f
C38 A1 VNB 0.444244f
C39 A2 VNB 0.407172f
C40 A3 VNB 0.43464f
C41 VPB VNB 2.33467f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2111o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111o_1 VNB VPB VPWR VGND X C1 B1 A2 A1 D1
X0 a_85_136.t1 D1.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1504 ps=1.11 w=0.64 l=0.15
X1 VGND.t4 C1.t0 a_85_136.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1504 pd=1.11 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 a_85_136.t2 D1.t1 a_431_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.12 ps=1.24 w=1 l=0.15
X3 X.t1 a_85_136.t5 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X4 VPWR.t0 A1.t0 a_80_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.17 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X5 a_431_392.t0 C1.t1 a_353_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.12 ps=1.24 w=1 l=0.15
X6 X.t0 a_85_136.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X7 VGND.t1 A2.t0 a_168_136.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0672 ps=0.85 w=0.64 l=0.15
X8 a_353_392.t1 B1.t0 a_80_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.15 ps=1.3 w=1 l=0.15
X9 a_80_392.t2 A2.t1 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.17 ps=1.34 w=1 l=0.15
X10 a_85_136.t0 B1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1248 ps=1.03 w=0.64 l=0.15
X11 a_168_136.t1 A1.t1 a_85_136.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1696 ps=1.81 w=0.64 l=0.15
R0 D1.n0 D1.t1 226.925
R1 D1.n0 D1.t0 170.424
R2 D1 D1.n0 154.347
R3 VGND.n4 VGND.n3 236.417
R4 VGND.n1 VGND.n0 234.695
R5 VGND.n5 VGND.t2 182.305
R6 VGND.n3 VGND.t4 61.8755
R7 VGND.n0 VGND.t0 46.8755
R8 VGND.n11 VGND.n1 42.3391
R9 VGND.n8 VGND.n7 36.1417
R10 VGND.n9 VGND.n8 36.1417
R11 VGND.n7 VGND.n4 32.377
R12 VGND.n3 VGND.t3 26.2505
R13 VGND.n0 VGND.t1 26.2505
R14 VGND.n5 VGND.n4 11.0959
R15 VGND.n10 VGND.n9 9.3005
R16 VGND.n8 VGND.n2 9.3005
R17 VGND.n7 VGND.n6 9.3005
R18 VGND.n9 VGND.n1 1.50638
R19 VGND.n6 VGND.n5 0.453235
R20 VGND VGND.n11 0.163644
R21 VGND.n11 VGND.n10 0.144205
R22 VGND.n6 VGND.n2 0.122949
R23 VGND.n10 VGND.n2 0.122949
R24 a_85_136.n2 a_85_136.t3 295.079
R25 a_85_136.t2 a_85_136.n4 284.149
R26 a_85_136.n0 a_85_136.t5 249.847
R27 a_85_136.n0 a_85_136.t6 194.952
R28 a_85_136.n2 a_85_136.n1 185
R29 a_85_136.n4 a_85_136.n0 167.904
R30 a_85_136.n3 a_85_136.t1 130.895
R31 a_85_136.n3 a_85_136.n2 84.7453
R32 a_85_136.n4 a_85_136.n3 47.8619
R33 a_85_136.n1 a_85_136.t4 26.2505
R34 a_85_136.n1 a_85_136.t0 26.2505
R35 VNB.t3 VNB.t2 2540.68
R36 VNB VNB.t4 1766.93
R37 VNB.t5 VNB.t3 1432.02
R38 VNB.t1 VNB.t0 1247.24
R39 VNB.t0 VNB.t5 993.177
R40 VNB.t4 VNB.t1 831.496
R41 C1.t0 C1.t1 442.904
R42 C1 C1.t0 328.45
R43 a_431_392.t0 a_431_392.t1 47.2805
R44 VPB.t3 VPB.t2 679.302
R45 VPB VPB.t0 383.065
R46 VPB.t0 VPB.t5 250.269
R47 VPB.t5 VPB.t4 229.839
R48 VPB.t1 VPB.t3 199.195
R49 VPB.t4 VPB.t1 199.195
R50 VPWR.n1 VPWR.n0 337.661
R51 VPWR.n1 VPWR.t1 265.808
R52 VPWR.n0 VPWR.t2 33.4905
R53 VPWR.n0 VPWR.t0 33.4905
R54 VPWR VPWR.n1 0.262473
R55 X.n3 X 589.777
R56 X.n3 X.n0 585
R57 X.n4 X.n3 585
R58 X.n2 X.t0 286.887
R59 X.t0 X.n1 286.887
R60 X.n3 X.t1 26.3844
R61 X X.n4 12.8005
R62 X.n1 X 11.6542
R63 X X.n0 11.0811
R64 X X.n2 8.59751
R65 X.n2 X 5.5408
R66 X X.n0 3.05722
R67 X.n1 X 2.48408
R68 X.n4 X 1.33781
R69 A1.t1 A1.t0 442.904
R70 A1 A1.t1 315.507
R71 a_80_392.t0 a_80_392.n0 485.187
R72 a_80_392.n0 a_80_392.t1 29.5505
R73 a_80_392.n0 a_80_392.t2 29.5505
R74 a_353_392.t0 a_353_392.t1 47.2805
R75 A2.n0 A2.t1 231.629
R76 A2.n0 A2.t0 175.127
R77 A2.n1 A2.n0 152
R78 A2 A2.n1 16.2138
R79 A2.n1 A2 4.26717
R80 a_168_136.t0 a_168_136.t1 39.3755
R81 B1.t1 B1.t0 440.791
R82 B1 B1.t1 329.077
C0 A2 C1 0.015736f
C1 VPB VPWR 0.148498f
C2 A1 VPWR 0.015963f
C3 A2 D1 0.026683f
C4 VPB X 0.015347f
C5 B1 C1 0.116253f
C6 A2 VPWR 0.026627f
C7 VPB VGND 0.014696f
C8 B1 VPWR 0.00631f
C9 A1 VGND 0.102081f
C10 C1 D1 0.054981f
C11 A2 VGND 0.015583f
C12 C1 VPWR 0.008571f
C13 C1 X 1.44e-19
C14 D1 VPWR 0.013449f
C15 B1 VGND 0.08338f
C16 VPB A1 0.041473f
C17 C1 VGND 0.082657f
C18 D1 X 3.47e-19
C19 VPB A2 0.046994f
C20 D1 VGND 0.013772f
C21 VPWR X 0.127488f
C22 VPB B1 0.029039f
C23 A1 A2 0.063336f
C24 VPWR VGND 0.071551f
C25 VPB C1 0.027658f
C26 A1 B1 0.008253f
C27 X VGND 0.101079f
C28 A2 B1 0.068222f
C29 VPB D1 0.053175f
C30 VGND VNB 0.586517f
C31 X VNB 0.109409f
C32 VPWR VNB 0.444943f
C33 D1 VNB 0.106021f
C34 C1 VNB 0.132217f
C35 B1 VNB 0.126767f
C36 A2 VNB 0.099958f
C37 A1 VNB 0.183089f
C38 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2111o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111o_2 VNB VPB VPWR VGND D1 C1 B1 A2 A1 X
X0 VPWR.t3 a_91_244.t5 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_630_368.t2 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.2184 ps=1.51 w=1.12 l=0.15
X2 X.t1 a_91_244.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X3 X.t2 a_91_244.t7 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X4 a_522_368.t1 C1.t0 a_444_368.t0 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1344 ps=1.36 w=1.12 l=0.15
X5 a_91_244.t3 C1.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1184 ps=1.06 w=0.74 l=0.15
X6 VGND.t0 D1.t0 a_91_244.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1961 ps=2.01 w=0.74 l=0.15
X7 a_771_74.t1 A2.t0 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.2109 ps=1.31 w=0.74 l=0.15
X8 a_91_244.t0 A1.t1 a_771_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.0777 ps=0.95 w=0.74 l=0.15
X9 VGND.t1 a_91_244.t8 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 VGND.t3 B1.t0 a_91_244.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=1.31 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_630_368.t0 B1.t1 a_522_368.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.2184 ps=1.51 w=1.12 l=0.15
X12 a_444_368.t1 D1.t1 a_91_244.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.36 as=0.308 ps=2.79 w=1.12 l=0.15
X13 VPWR.t1 A2.t1 a_630_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.2184 ps=1.51 w=1.12 l=0.15
R0 a_91_244.t4 a_91_244.n5 304.531
R1 a_91_244.n4 a_91_244.t7 263.81
R2 a_91_244.n0 a_91_244.t5 261.62
R3 a_91_244.n2 a_91_244.t0 241.57
R4 a_91_244.n5 a_91_244.n0 181.213
R5 a_91_244.n3 a_91_244.t1 155.638
R6 a_91_244.n4 a_91_244.t6 154.24
R7 a_91_244.n0 a_91_244.t8 154.24
R8 a_91_244.n2 a_91_244.n1 104.579
R9 a_91_244.n0 a_91_244.n4 63.5369
R10 a_91_244.n3 a_91_244.n2 54.9652
R11 a_91_244.n5 a_91_244.n3 47.4358
R12 a_91_244.n1 a_91_244.t2 22.7032
R13 a_91_244.n1 a_91_244.t3 22.7032
R14 X.n2 X 591.274
R15 X.n2 X.n0 585
R16 X.n3 X.n2 585
R17 X X.n1 145.815
R18 X.n2 X.t3 26.3844
R19 X.n2 X.t2 26.3844
R20 X.n1 X.t0 22.7032
R21 X.n1 X.t1 22.7032
R22 X X.n3 16.8162
R23 X X.n0 14.5574
R24 X X.n0 4.01619
R25 X.n3 X 1.75736
R26 VPWR.n3 VPWR.t3 342.31
R27 VPWR.n2 VPWR.n1 319.822
R28 VPWR.n5 VPWR.t2 259.171
R29 VPWR.n1 VPWR.t0 38.6969
R30 VPWR.n1 VPWR.t1 29.9023
R31 VPWR.n4 VPWR.n3 25.224
R32 VPWR.n5 VPWR.n4 23.7181
R33 VPWR.n4 VPWR.n0 9.3005
R34 VPWR.n6 VPWR.n5 9.3005
R35 VPWR.n3 VPWR.n2 7.06472
R36 VPWR.n2 VPWR.n0 0.159562
R37 VPWR.n6 VPWR.n0 0.122949
R38 VPWR VPWR.n6 0.0617245
R39 VPB.t4 VPB.t6 587.366
R40 VPB VPB.t3 278.361
R41 VPB.t2 VPB.t0 275.807
R42 VPB.t1 VPB.t2 275.807
R43 VPB.t5 VPB.t1 275.807
R44 VPB.t3 VPB.t4 229.839
R45 VPB.t6 VPB.t5 199.195
R46 A1.n0 A1.t0 226.809
R47 A1 A1.n0 209.294
R48 A1.n0 A1.t1 198.204
R49 a_630_368.n0 a_630_368.t2 489.699
R50 a_630_368.n0 a_630_368.t1 38.6969
R51 a_630_368.t0 a_630_368.n0 29.9023
R52 VGND.n10 VGND.t1 233.886
R53 VGND.n5 VGND.n4 208.351
R54 VGND.n3 VGND.n2 204.825
R55 VGND.n12 VGND.t2 167.655
R56 VGND.n2 VGND.t3 50.2708
R57 VGND.n2 VGND.t5 42.1627
R58 VGND.n6 VGND.n1 36.1417
R59 VGND.n4 VGND.t4 25.9464
R60 VGND.n4 VGND.t0 25.9464
R61 VGND.n11 VGND.n10 24.0946
R62 VGND.n10 VGND.n1 23.3417
R63 VGND.n12 VGND.n11 15.8123
R64 VGND.n5 VGND.n3 11.4978
R65 VGND.n13 VGND.n12 9.3005
R66 VGND.n7 VGND.n6 9.3005
R67 VGND.n8 VGND.n1 9.3005
R68 VGND.n10 VGND.n9 9.3005
R69 VGND.n11 VGND.n0 9.3005
R70 VGND.n6 VGND.n5 3.76521
R71 VGND.n7 VGND.n3 0.741596
R72 VGND.n8 VGND.n7 0.122949
R73 VGND.n9 VGND.n8 0.122949
R74 VGND.n9 VGND.n0 0.122949
R75 VGND.n13 VGND.n0 0.122949
R76 VGND VGND.n13 0.0617245
R77 VNB.t2 VNB.t0 2702.36
R78 VNB.t4 VNB.t6 1662.99
R79 VNB VNB.t3 1293.44
R80 VNB.t0 VNB.t5 1085.56
R81 VNB.t5 VNB.t4 993.177
R82 VNB.t3 VNB.t2 993.177
R83 VNB.t6 VNB.t1 831.496
R84 C1.n0 C1.t0 250.909
R85 C1.n0 C1.t1 220.113
R86 C1 C1.n0 154.522
R87 a_444_368.t0 a_444_368.t1 42.2148
R88 a_522_368.t0 a_522_368.t1 68.5987
R89 D1.n0 D1.t1 250.909
R90 D1.n0 D1.t0 220.113
R91 D1.n1 D1.n0 152
R92 D1.n1 D1 14.14
R93 D1 D1.n1 0.149337
R94 A2.n0 A2.t1 250.909
R95 A2.n0 A2.t0 220.113
R96 A2.n1 A2.n0 152
R97 A2 A2.n1 9.07957
R98 A2.n1 A2 5.2098
R99 a_771_74.t0 a_771_74.t1 34.0546
R100 B1.n0 B1.t1 250.909
R101 B1.n0 B1.t0 220.113
R102 B1 B1.n0 155.423
C0 VPB C1 0.036328f
C1 VPWR X 0.176697f
C2 A1 VGND 0.014766f
C3 VPB B1 0.034193f
C4 D1 C1 0.106901f
C5 VPWR VGND 0.090555f
C6 VPB A2 0.035131f
C7 X VGND 0.127985f
C8 VPB A1 0.056f
C9 C1 B1 0.097635f
C10 C1 A2 4.54e-19
C11 VPB VPWR 0.15666f
C12 VPB X 0.006402f
C13 C1 A1 2.05e-19
C14 D1 VPWR 0.011639f
C15 B1 A2 0.083884f
C16 VPB VGND 0.012641f
C17 C1 VPWR 0.034889f
C18 B1 VPWR 0.010649f
C19 D1 VGND 0.01593f
C20 A2 A1 0.115269f
C21 C1 VGND 0.015427f
C22 A2 VPWR 0.018741f
C23 A1 VPWR 0.018878f
C24 B1 VGND 0.014699f
C25 VPB D1 0.039616f
C26 A2 VGND 0.019848f
C27 VGND VNB 0.642125f
C28 X VNB 0.031749f
C29 VPWR VNB 0.52171f
C30 A1 VNB 0.177995f
C31 A2 VNB 0.105463f
C32 B1 VNB 0.104546f
C33 C1 VNB 0.10327f
C34 D1 VNB 0.11912f
C35 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21boi_2 VNB VPB VPWR VGND B1_N Y A2 A1
X0 VGND.t4 A2.t0 a_436_74.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_241_368.t5 A2.t1 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1792 ps=1.44 w=1.12 l=0.15
X2 Y.t3 a_62_94.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12205 ps=1.08 w=0.74 l=0.15
X3 a_436_74.t1 A2.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t2 a_62_94.t3 Y.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_436_74.t0 A1.t0 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 VPWR.t3 A2.t3 a_241_368.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_241_368.t3 A1.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VPWR.t0 A1.t2 a_241_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 a_62_94.t1 B1_N.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X10 a_241_368.t1 a_62_94.t4 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t0 a_62_94.t5 a_241_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X12 Y.t5 A1.t3 a_436_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X13 VGND.t0 B1_N.t1 a_62_94.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12205 pd=1.08 as=0.1696 ps=1.81 w=0.64 l=0.15
R0 A2.n1 A2.t3 265.271
R1 A2.n0 A2.t1 263.81
R2 A2.n3 A2.n2 156.694
R3 A2.n1 A2.t0 154.24
R4 A2.n0 A2.t2 154.24
R5 A2.n2 A2.n0 55.5035
R6 A2.n3 A2 27.2005
R7 A2.n2 A2.n1 7.30353
R8 A2 A2.n3 0.284944
R9 a_436_74.n0 a_436_74.t3 339.534
R10 a_436_74.n0 a_436_74.t1 216.023
R11 a_436_74.n1 a_436_74.n0 88.1937
R12 a_436_74.n1 a_436_74.t2 22.7032
R13 a_436_74.t0 a_436_74.n1 22.7032
R14 VGND.n4 VGND.t2 232.721
R15 VGND.n3 VGND.n2 212.613
R16 VGND.n1 VGND.n0 115.66
R17 VGND.n0 VGND.t0 37.5005
R18 VGND.n5 VGND.n4 31.624
R19 VGND.n2 VGND.t3 22.7032
R20 VGND.n2 VGND.t4 22.7032
R21 VGND.n0 VGND.t1 21.9089
R22 VGND.n7 VGND.n1 10.7156
R23 VGND.n6 VGND.n5 9.3005
R24 VGND.n5 VGND.n1 8.28285
R25 VGND.n4 VGND.n3 6.61607
R26 VGND.n6 VGND.n3 0.180314
R27 VGND VGND.n7 0.163644
R28 VGND.n7 VGND.n6 0.144205
R29 VNB.t3 VNB.t6 2194.23
R30 VNB VNB.t0 1501.31
R31 VNB.t0 VNB.t2 1131.76
R32 VNB.t5 VNB.t4 993.177
R33 VNB.t1 VNB.t5 993.177
R34 VNB.t6 VNB.t1 993.177
R35 VNB.t2 VNB.t3 993.177
R36 VPWR.n5 VPWR.n4 316.683
R37 VPWR.n12 VPWR.t1 260.599
R38 VPWR.n3 VPWR.n2 225.782
R39 VPWR.n6 VPWR.n1 36.1417
R40 VPWR.n10 VPWR.n1 36.1417
R41 VPWR.n11 VPWR.n10 36.1417
R42 VPWR.n2 VPWR.t4 28.1434
R43 VPWR.n2 VPWR.t3 28.1434
R44 VPWR.n6 VPWR.n5 26.7299
R45 VPWR.n4 VPWR.t2 26.3844
R46 VPWR.n4 VPWR.t0 26.3844
R47 VPWR.n12 VPWR.n11 20.7064
R48 VPWR.n7 VPWR.n6 9.3005
R49 VPWR.n8 VPWR.n1 9.3005
R50 VPWR.n10 VPWR.n9 9.3005
R51 VPWR.n11 VPWR.n0 9.3005
R52 VPWR.n13 VPWR.n12 9.3005
R53 VPWR.n5 VPWR.n3 6.50429
R54 VPWR.n7 VPWR.n3 0.595518
R55 VPWR.n8 VPWR.n7 0.122949
R56 VPWR.n9 VPWR.n8 0.122949
R57 VPWR.n9 VPWR.n0 0.122949
R58 VPWR.n13 VPWR.n0 0.122949
R59 VPWR VPWR.n13 0.0617245
R60 a_241_368.n1 a_241_368.t2 330.072
R61 a_241_368.n2 a_241_368.t5 309.408
R62 a_241_368.n3 a_241_368.n2 207.35
R63 a_241_368.n1 a_241_368.n0 184.756
R64 a_241_368.n2 a_241_368.n1 84.8443
R65 a_241_368.n0 a_241_368.t0 26.3844
R66 a_241_368.n0 a_241_368.t1 26.3844
R67 a_241_368.t4 a_241_368.n3 26.3844
R68 a_241_368.n3 a_241_368.t3 26.3844
R69 VPB.t3 VPB.t2 495.43
R70 VPB VPB.t3 298.791
R71 VPB.t5 VPB.t6 240.054
R72 VPB.t4 VPB.t5 229.839
R73 VPB.t0 VPB.t4 229.839
R74 VPB.t1 VPB.t0 229.839
R75 VPB.t2 VPB.t1 229.839
R76 a_62_94.n0 a_62_94.t4 319.728
R77 a_62_94.t1 a_62_94.n3 260.272
R78 a_62_94.n1 a_62_94.t3 230.558
R79 a_62_94.n0 a_62_94.t5 224.131
R80 a_62_94.n2 a_62_94.t2 199.519
R81 a_62_94.n3 a_62_94.t0 179.103
R82 a_62_94.n3 a_62_94.n2 165.189
R83 a_62_94.n1 a_62_94.n0 54.8949
R84 a_62_94.n2 a_62_94.n1 34.3247
R85 Y.n3 Y.n1 223.788
R86 Y Y.n0 218.724
R87 Y.n3 Y.n2 125.879
R88 Y.n1 Y.t1 26.3844
R89 Y.n1 Y.t0 26.3844
R90 Y.n2 Y.t2 22.7032
R91 Y.n2 Y.t3 22.7032
R92 Y.n0 Y.t4 22.7032
R93 Y.n0 Y.t5 22.7032
R94 Y Y.n3 8.7819
R95 A1.n1 A1.t2 244.335
R96 A1.n0 A1.t1 234.841
R97 A1.n0 A1.t0 193.963
R98 A1.n1 A1.t3 186.374
R99 A1 A1.n2 154.643
R100 A1.n2 A1.n0 37.246
R101 A1.n2 A1.n1 18.9884
R102 B1_N.n0 B1_N.t1 221.575
R103 B1_N.n0 B1_N.t0 212.883
R104 B1_N B1_N.n0 198.179
C0 Y VGND 0.161879f
C1 VPB B1_N 0.070382f
C2 VPB A1 0.061635f
C3 VPB A2 0.061322f
C4 VPB VPWR 0.128386f
C5 VPB Y 0.004332f
C6 A1 A2 0.073361f
C7 B1_N VPWR 0.044379f
C8 VPB VGND 0.008746f
C9 A1 VPWR 0.041199f
C10 B1_N Y 6.75e-19
C11 A1 Y 0.077221f
C12 B1_N VGND 0.018035f
C13 A2 VPWR 0.046047f
C14 A1 VGND 0.016716f
C15 A2 Y 0.003917f
C16 VPWR Y 0.012015f
C17 A2 VGND 0.031984f
C18 VPWR VGND 0.070105f
C19 VGND VNB 0.554337f
C20 Y VNB 0.033721f
C21 VPWR VNB 0.463372f
C22 A2 VNB 0.238957f
C23 A1 VNB 0.206309f
C24 B1_N VNB 0.177885f
C25 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2bb2oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2oi_2 VNB VPB VPWR VGND A2_N Y B2 B1 A1_N
X0 VGND.t2 A2_N.t0 a_212_102.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.12205 pd=1.08 as=0.104 ps=0.965 w=0.64 l=0.15
X1 Y.t5 a_212_102.t3 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12205 ps=1.08 w=0.74 l=0.15
X2 a_212_102.t1 A2_N.t1 a_209_392.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.12 ps=1.24 w=1 l=0.15
X3 a_424_368.t3 B1.t0 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VPWR.t3 B1.t1 a_424_368.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5 a_424_368.t0 B2.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t2 B2.t1 a_424_368.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_212_102.t2 A1_N.t0 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.1696 ps=1.81 w=0.64 l=0.15
X8 a_209_392.t0 A1_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.275 ps=2.55 w=1 l=0.15
X9 a_424_368.t5 a_212_102.t4 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t2 a_212_102.t5 a_424_368.t4 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X11 VGND.t1 B1.t2 a_615_74.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_615_74.t2 B1.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_615_74.t1 B2.t2 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 VGND.t5 a_212_102.t6 Y.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 Y.t1 B2.t3 a_615_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
R0 A2_N.n0 A2_N.t1 236.983
R1 A2_N.n0 A2_N.t0 223.327
R2 A2_N A2_N.n0 164.412
R3 a_212_102.n1 a_212_102.t4 345.142
R4 a_212_102.t1 a_212_102.n4 260.998
R5 a_212_102.n1 a_212_102.t5 241.035
R6 a_212_102.n3 a_212_102.t3 186.666
R7 a_212_102.n2 a_212_102.t6 173.52
R8 a_212_102.n4 a_212_102.n3 152
R9 a_212_102.n4 a_212_102.n0 149.216
R10 a_212_102.n3 a_212_102.n2 49.6611
R11 a_212_102.n0 a_212_102.t0 30.938
R12 a_212_102.n0 a_212_102.t2 30.0005
R13 a_212_102.n2 a_212_102.n1 7.16051
R14 VGND.n4 VGND.t5 232.721
R15 VGND.n5 VGND.n3 221.792
R16 VGND.n8 VGND.n2 213.898
R17 VGND.n10 VGND.t3 169.169
R18 VGND.n2 VGND.t2 37.5005
R19 VGND.n9 VGND.n8 27.8593
R20 VGND.n10 VGND.n9 25.977
R21 VGND.n3 VGND.t0 22.7032
R22 VGND.n3 VGND.t1 22.7032
R23 VGND.n2 VGND.t4 21.9089
R24 VGND.n4 VGND.n1 20.3299
R25 VGND.n8 VGND.n1 19.577
R26 VGND.n6 VGND.n1 9.3005
R27 VGND.n8 VGND.n7 9.3005
R28 VGND.n9 VGND.n0 9.3005
R29 VGND.n11 VGND.n10 7.40447
R30 VGND.n5 VGND.n4 7.29988
R31 VGND.n6 VGND.n5 0.167964
R32 VGND VGND.n11 0.159703
R33 VGND.n11 VGND.n0 0.148095
R34 VGND.n7 VGND.n6 0.122949
R35 VGND.n7 VGND.n0 0.122949
R36 VNB.t6 VNB.t3 2390.55
R37 VNB VNB.t5 2275.07
R38 VNB.t4 VNB.t7 1131.76
R39 VNB.t5 VNB.t4 1097.11
R40 VNB.t2 VNB.t0 993.177
R41 VNB.t1 VNB.t2 993.177
R42 VNB.t3 VNB.t1 993.177
R43 VNB.t7 VNB.t6 993.177
R44 Y.n2 Y.n0 328.526
R45 Y Y.n1 213.829
R46 Y Y.n3 127.862
R47 Y.n0 Y.t3 26.3844
R48 Y.n0 Y.t2 26.3844
R49 Y.n3 Y.t4 22.7032
R50 Y.n3 Y.t5 22.7032
R51 Y.n1 Y.t0 22.7032
R52 Y.n1 Y.t1 22.7032
R53 Y.n2 Y 11.461
R54 Y Y.n2 2.82841
R55 a_209_392.t0 a_209_392.t1 47.2805
R56 VPB.t5 VPB.t6 566.936
R57 VPB VPB.t0 495.43
R58 VPB.t4 VPB.t3 229.839
R59 VPB.t1 VPB.t4 229.839
R60 VPB.t2 VPB.t1 229.839
R61 VPB.t7 VPB.t2 229.839
R62 VPB.t6 VPB.t7 229.839
R63 VPB.t0 VPB.t5 199.195
R64 B1.n0 B1.t0 229
R65 B1.n1 B1.t1 227.538
R66 B1.n1 B1.t2 196.013
R67 B1.n0 B1.t3 196.013
R68 B1.n3 B1.n2 152
R69 B1.n2 B1.n0 52.5823
R70 B1.n3 B1 10.4191
R71 B1.n2 B1.n1 10.2247
R72 B1 B1.n3 3.87027
R73 VPWR.n4 VPWR.n3 321.438
R74 VPWR.n6 VPWR.n5 315.928
R75 VPWR.n14 VPWR.t0 252.012
R76 VPWR.n8 VPWR.n7 36.1417
R77 VPWR.n8 VPWR.n1 36.1417
R78 VPWR.n12 VPWR.n1 36.1417
R79 VPWR.n13 VPWR.n12 36.1417
R80 VPWR.n5 VPWR.t1 26.3844
R81 VPWR.n5 VPWR.t2 26.3844
R82 VPWR.n3 VPWR.t4 26.3844
R83 VPWR.n3 VPWR.t3 26.3844
R84 VPWR.n7 VPWR.n6 23.3417
R85 VPWR.n14 VPWR.n13 21.8358
R86 VPWR.n7 VPWR.n2 9.3005
R87 VPWR.n9 VPWR.n8 9.3005
R88 VPWR.n10 VPWR.n1 9.3005
R89 VPWR.n12 VPWR.n11 9.3005
R90 VPWR.n13 VPWR.n0 9.3005
R91 VPWR.n15 VPWR.n14 7.32393
R92 VPWR.n6 VPWR.n4 6.67638
R93 VPWR.n4 VPWR.n2 0.607026
R94 VPWR VPWR.n15 0.158642
R95 VPWR.n15 VPWR.n0 0.149142
R96 VPWR.n9 VPWR.n2 0.122949
R97 VPWR.n10 VPWR.n9 0.122949
R98 VPWR.n11 VPWR.n10 0.122949
R99 VPWR.n11 VPWR.n0 0.122949
R100 a_424_368.n2 a_424_368.t4 319.356
R101 a_424_368.t3 a_424_368.n3 293.408
R102 a_424_368.n3 a_424_368.n0 208.897
R103 a_424_368.n2 a_424_368.n1 186.73
R104 a_424_368.n3 a_424_368.n2 80.2951
R105 a_424_368.n0 a_424_368.t2 26.3844
R106 a_424_368.n0 a_424_368.t0 26.3844
R107 a_424_368.n1 a_424_368.t1 26.3844
R108 a_424_368.n1 a_424_368.t5 26.3844
R109 B2.n1 B2.t1 241.415
R110 B2.n0 B2.t0 234.841
R111 B2.n0 B2.t2 190.276
R112 B2.n1 B2.t3 186.374
R113 B2 B2.n2 155.685
R114 B2.n2 B2.n0 36.5157
R115 B2.n2 B2.n1 22.6399
R116 A1_N.t0 A1_N.t1 488.428
R117 A1_N A1_N.t0 483.584
R118 a_615_74.n0 a_615_74.t0 343.711
R119 a_615_74.n0 a_615_74.t2 221.232
R120 a_615_74.n1 a_615_74.n0 86.1054
R121 a_615_74.n1 a_615_74.t3 22.7032
R122 a_615_74.t1 a_615_74.n1 22.7032
C0 VPWR Y 0.011115f
C1 B1 VGND 0.032085f
C2 VPB A1_N 0.047393f
C3 VPWR VGND 0.095449f
C4 VPB A2_N 0.051172f
C5 Y VGND 0.156903f
C6 VPB B2 0.060254f
C7 A1_N A2_N 0.07322f
C8 VPB B1 0.066046f
C9 VPB VPWR 0.170765f
C10 A1_N VPWR 0.029573f
C11 VPB Y 0.005868f
C12 A1_N Y 4.64e-20
C13 B2 B1 0.093706f
C14 VPB VGND 0.016659f
C15 A2_N VPWR 0.022612f
C16 B2 VPWR 0.041166f
C17 A2_N Y 5.22e-19
C18 A1_N VGND 0.104004f
C19 B2 Y 0.076097f
C20 A2_N VGND 0.016297f
C21 B1 VPWR 0.041733f
C22 B2 VGND 0.016632f
C23 B1 Y 4.9e-19
C24 VGND VNB 0.687029f
C25 Y VNB 0.037229f
C26 VPWR VNB 0.545448f
C27 B1 VNB 0.23568f
C28 B2 VNB 0.200759f
C29 A2_N VNB 0.114715f
C30 A1_N VNB 0.263553f
C31 VPB VNB 1.26331f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2bb2oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2oi_1 VNB VPB VPWR VGND Y A2_N A1_N B2 B1
X0 a_126_112.t0 A1_N.t0 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.14575 ps=1.63 w=0.55 l=0.15
X1 Y.t0 a_126_112.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.245175 ps=1.54 w=0.74 l=0.15
X2 a_117_392.t0 A1_N.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.275 ps=2.55 w=1 l=0.15
X3 VGND.t2 B1.t0 a_488_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1184 ps=1.06 w=0.74 l=0.15
X4 a_488_74.t1 B2.t0 Y.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_126_112.t2 A2_N.t0 a_117_392.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.12 ps=1.24 w=1 l=0.15
X6 a_399_368.t0 B1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1848 ps=1.45 w=1.12 l=0.15
X7 VPWR.t0 B2.t1 a_399_368.t2 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X8 a_399_368.t1 a_126_112.t4 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X9 VGND.t3 A2_N.t1 a_126_112.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.245175 pd=1.54 as=0.077 ps=0.83 w=0.55 l=0.15
R0 A1_N.n0 A1_N.t1 263.762
R1 A1_N A1_N.n0 193.067
R2 A1_N.n0 A1_N.t0 143.732
R3 VGND.n11 VGND.t1 257.274
R4 VGND.n3 VGND.n1 185
R5 VGND.n5 VGND.n4 185
R6 VGND.n2 VGND.t2 165.654
R7 VGND.n4 VGND.n3 98.1823
R8 VGND.n3 VGND.t3 45.8187
R9 VGND.n5 VGND.n2 30.5782
R10 VGND.n10 VGND.n9 30.5183
R11 VGND.n4 VGND.t0 22.7275
R12 VGND.n11 VGND.n10 22.2123
R13 VGND.n12 VGND.n11 9.3005
R14 VGND.n7 VGND.n6 9.3005
R15 VGND.n9 VGND.n8 9.3005
R16 VGND.n10 VGND.n0 9.3005
R17 VGND.n6 VGND.n1 6.60176
R18 VGND.n9 VGND.n1 1.12754
R19 VGND.n6 VGND.n5 0.644525
R20 VGND.n7 VGND.n2 0.562535
R21 VGND.n8 VGND.n7 0.122949
R22 VGND.n8 VGND.n0 0.122949
R23 VGND.n12 VGND.n0 0.122949
R24 VGND VGND.n12 0.0617245
R25 a_126_112.t2 a_126_112.n2 284.087
R26 a_126_112.n1 a_126_112.t4 261.62
R27 a_126_112.n2 a_126_112.n0 236.345
R28 a_126_112.n2 a_126_112.n1 206.774
R29 a_126_112.n1 a_126_112.t3 156.431
R30 a_126_112.n0 a_126_112.t1 30.546
R31 a_126_112.n0 a_126_112.t0 30.546
R32 VNB.t4 VNB.t1 2194.23
R33 VNB VNB.t0 1281.89
R34 VNB.t3 VNB.t2 1085.56
R35 VNB.t1 VNB.t3 993.177
R36 VNB.t0 VNB.t4 993.177
R37 Y.n1 Y.t1 229.721
R38 Y.n1 Y.n0 168.706
R39 Y.n0 Y.t2 22.7032
R40 Y.n0 Y.t0 22.7032
R41 Y Y.n1 7.68715
R42 VPWR.n1 VPWR.n0 622.747
R43 VPWR.n1 VPWR.t2 258.858
R44 VPWR.n0 VPWR.t1 29.0228
R45 VPWR.n0 VPWR.t0 29.0228
R46 VPWR VPWR.n1 0.103195
R47 a_117_392.t0 a_117_392.t1 47.2805
R48 VPB.t4 VPB.t3 520.968
R49 VPB VPB.t2 260.485
R50 VPB.t0 VPB.t1 245.161
R51 VPB.t3 VPB.t0 229.839
R52 VPB.t2 VPB.t4 199.195
R53 B1.n0 B1.t1 277.687
R54 B1.n0 B1.t0 170.308
R55 B1 B1.n0 158.788
R56 a_488_74.t0 a_488_74.t1 51.8924
R57 B2.n0 B2.t1 285.719
R58 B2.n0 B2.t0 178.34
R59 B2 B2.n0 164.427
R60 A2_N.n0 A2_N.t0 228.281
R61 A2_N.n0 A2_N.t1 220.625
R62 A2_N A2_N.n0 166.352
R63 a_399_368.t0 a_399_368.n0 880.322
R64 a_399_368.n0 a_399_368.t2 26.3844
R65 a_399_368.n0 a_399_368.t1 26.3844
C0 VPB Y 0.012507f
C1 A1_N VPWR 0.054879f
C2 A2_N VPWR 0.023257f
C3 B2 B1 0.098738f
C4 VPB VGND 0.008727f
C5 A1_N VGND 0.042143f
C6 B2 VPWR 0.022901f
C7 A2_N Y 0.001351f
C8 A2_N VGND 0.013759f
C9 B1 VPWR 0.014178f
C10 B2 Y 0.084383f
C11 B2 VGND 0.025329f
C12 B1 Y 0.004858f
C13 VPWR Y 0.039063f
C14 B1 VGND 0.051913f
C15 VPB A1_N 0.050868f
C16 VPWR VGND 0.05769f
C17 VPB A2_N 0.050843f
C18 Y VGND 0.105904f
C19 A1_N A2_N 0.106602f
C20 VPB B2 0.033629f
C21 VPB B1 0.040625f
C22 A2_N B2 7.76e-20
C23 VPB VPWR 0.110137f
C24 VGND VNB 0.515031f
C25 Y VNB 0.018801f
C26 VPWR VNB 0.385555f
C27 B1 VNB 0.168155f
C28 B2 VNB 0.115462f
C29 A2_N VNB 0.112893f
C30 A1_N VNB 0.180145f
C31 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2bb2o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2o_4 VNB VPB VPWR VGND X B2 B1 A2_N A1_N
X0 VGND.t3 a_162_48.t5 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.18285 pd=1.27 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_162_48.t0 B2.t0 a_1009_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X2 VGND.t8 A2_N.t0 a_586_94.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.33325 pd=1.74 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 a_586_94.t1 A2_N.t1 a_583_368.t0 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1344 ps=1.36 w=1.12 l=0.15
X4 a_1009_74.t2 B2.t1 a_162_48.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 VPWR.t3 a_162_48.t6 X.t7 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.168 ps=1.42 w=1.12 l=0.15
X6 VPWR.t5 B1.t0 a_820_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X7 a_820_392.t1 a_586_94.t3 a_162_48.t2 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X8 X.t5 a_162_48.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 X.t2 a_162_48.t8 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_1009_74.t0 B1.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1024 ps=0.96 w=0.64 l=0.15
X11 VPWR.t1 a_162_48.t9 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_583_368.t1 A1_N.t0 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.1344 pd=1.36 as=0.2184 ps=1.51 w=1.12 l=0.15
X13 a_162_48.t3 a_586_94.t4 a_820_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X14 VPWR.t6 B2.t2 a_820_392.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X15 X.t0 a_162_48.t10 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X16 X.t4 a_162_48.t11 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X17 a_586_94.t2 A1_N.t1 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.18285 ps=1.27 w=0.64 l=0.15
X18 VGND.t0 a_162_48.t12 X.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X19 a_162_48.t4 a_586_94.t5 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.33325 ps=1.74 w=0.74 l=0.15
X20 VGND.t5 B1.t2 a_1009_74.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 a_162_48.n16 a_162_48.n15 365.009
R1 a_162_48.n15 a_162_48.n12 270.774
R2 a_162_48.n11 a_162_48.t6 251.882
R3 a_162_48.n14 a_162_48.n13 240.675
R4 a_162_48.n8 a_162_48.t8 240.197
R5 a_162_48.n1 a_162_48.t9 240.197
R6 a_162_48.n3 a_162_48.t10 240.197
R7 a_162_48.n3 a_162_48.t11 189.441
R8 a_162_48.n2 a_162_48.t12 179.947
R9 a_162_48.n7 a_162_48.t7 179.947
R10 a_162_48.n10 a_162_48.t5 179.947
R11 a_162_48.n5 a_162_48.n4 165.189
R12 a_162_48.n6 a_162_48.n5 152
R13 a_162_48.n9 a_162_48.n0 152
R14 a_162_48.n12 a_162_48.n11 152
R15 a_162_48.n14 a_162_48.t4 139.429
R16 a_162_48.n10 a_162_48.n9 43.0884
R17 a_162_48.n4 a_162_48.n3 36.5157
R18 a_162_48.n7 a_162_48.n6 29.9429
R19 a_162_48.t2 a_162_48.n16 29.5505
R20 a_162_48.n16 a_162_48.t3 29.5505
R21 a_162_48.n13 a_162_48.t1 26.2505
R22 a_162_48.n13 a_162_48.t0 26.2505
R23 a_162_48.n6 a_162_48.n1 20.449
R24 a_162_48.n4 a_162_48.n2 16.7975
R25 a_162_48.n15 a_162_48.n14 15.6751
R26 a_162_48.n8 a_162_48.n7 15.3369
R27 a_162_48.n12 a_162_48.n0 13.1884
R28 a_162_48.n5 a_162_48.n0 13.1884
R29 a_162_48.n2 a_162_48.n1 12.4157
R30 a_162_48.n11 a_162_48.n10 6.57323
R31 a_162_48.n9 a_162_48.n8 4.38232
R32 X.n2 X.n0 250.518
R33 X.n2 X.n1 207.6
R34 X.n5 X.n3 147.95
R35 X.n5 X.n4 102.019
R36 X.n0 X.t7 26.3844
R37 X.n0 X.t2 26.3844
R38 X.n1 X.t1 26.3844
R39 X.n1 X.t0 26.3844
R40 X X.n2 24.6885
R41 X.n3 X.t6 22.7032
R42 X.n3 X.t5 22.7032
R43 X.n4 X.t3 22.7032
R44 X.n4 X.t4 22.7032
R45 X X.n5 10.5046
R46 VGND.n24 VGND.t1 239.703
R47 VGND.n5 VGND.n4 223.159
R48 VGND.n15 VGND.n14 219.56
R49 VGND.n22 VGND.n21 217
R50 VGND.n6 VGND.n3 185
R51 VGND.n8 VGND.n7 185
R52 VGND.n7 VGND.n6 81.563
R53 VGND.n6 VGND.t8 79.688
R54 VGND.n14 VGND.t6 73.1255
R55 VGND.n13 VGND.n12 36.1417
R56 VGND.n16 VGND.n13 36.1417
R57 VGND.n20 VGND.n1 36.1417
R58 VGND.n24 VGND.n23 33.5064
R59 VGND.n4 VGND.t4 30.0005
R60 VGND.n4 VGND.t5 30.0005
R61 VGND.n8 VGND.n5 23.1042
R62 VGND.n21 VGND.t2 22.7032
R63 VGND.n21 VGND.t0 22.7032
R64 VGND.n14 VGND.t3 22.1988
R65 VGND.n7 VGND.t7 21.9089
R66 VGND.n16 VGND.n15 12.424
R67 VGND.n23 VGND.n22 12.424
R68 VGND.n10 VGND.n9 9.3005
R69 VGND.n12 VGND.n11 9.3005
R70 VGND.n13 VGND.n2 9.3005
R71 VGND.n17 VGND.n16 9.3005
R72 VGND.n18 VGND.n1 9.3005
R73 VGND.n20 VGND.n19 9.3005
R74 VGND.n23 VGND.n0 9.3005
R75 VGND.n12 VGND.n3 8.70613
R76 VGND.n25 VGND.n24 7.03525
R77 VGND.n15 VGND.n1 4.89462
R78 VGND.n22 VGND.n20 4.89462
R79 VGND.n9 VGND.n3 4.08266
R80 VGND.n9 VGND.n8 1.9378
R81 VGND.n10 VGND.n5 0.155444
R82 VGND VGND.n25 0.154841
R83 VGND.n25 VGND.n0 0.152893
R84 VGND.n11 VGND.n10 0.122949
R85 VGND.n11 VGND.n2 0.122949
R86 VGND.n17 VGND.n2 0.122949
R87 VGND.n18 VGND.n17 0.122949
R88 VGND.n19 VGND.n18 0.122949
R89 VGND.n19 VGND.n0 0.122949
R90 VNB.t10 VNB.t9 2656.17
R91 VNB.t9 VNB.t6 2194.23
R92 VNB VNB.t1 2044.09
R93 VNB.t3 VNB.t8 1570.6
R94 VNB.t5 VNB.t4 1085.56
R95 VNB.t7 VNB.t5 993.177
R96 VNB.t6 VNB.t7 993.177
R97 VNB.t8 VNB.t10 993.177
R98 VNB.t2 VNB.t3 993.177
R99 VNB.t0 VNB.t2 993.177
R100 VNB.t1 VNB.t0 993.177
R101 B2.n2 B2.t2 268.873
R102 B2.n1 B2.n0 263.762
R103 B2.n1 B2.t1 185.351
R104 B2.n2 B2.t0 183.161
R105 B2.n4 B2.n3 152
R106 B2.n3 B2.n1 33.5944
R107 B2.n3 B2.n2 27.0217
R108 B2.n4 B2 8.49281
R109 B2 B2.n4 3.32358
R110 a_1009_74.n0 a_1009_74.t3 296.382
R111 a_1009_74.n0 a_1009_74.t0 201.989
R112 a_1009_74.n1 a_1009_74.n0 97.0647
R113 a_1009_74.n1 a_1009_74.t1 26.2505
R114 a_1009_74.t2 a_1009_74.n1 26.2505
R115 A2_N.n0 A2_N.t1 243.73
R116 A2_N.n0 A2_N.t0 196.869
R117 A2_N A2_N.n0 154.084
R118 a_586_94.n1 a_586_94.t3 314.372
R119 a_586_94.n1 a_586_94.t5 312.498
R120 a_586_94.n2 a_586_94.n0 280.964
R121 a_586_94.n2 a_586_94.n1 278.63
R122 a_586_94.t1 a_586_94.n2 231.871
R123 a_586_94.n1 a_586_94.t4 227.612
R124 a_586_94.n0 a_586_94.t0 26.2505
R125 a_586_94.n0 a_586_94.t2 26.2505
R126 a_583_368.t0 a_583_368.t1 42.2148
R127 VPB.t7 VPB.t0 623.119
R128 VPB VPB.t3 485.216
R129 VPB.t9 VPB.t2 459.678
R130 VPB.t6 VPB.t8 275.807
R131 VPB.t1 VPB.t9 229.839
R132 VPB.t0 VPB.t1 229.839
R133 VPB.t5 VPB.t6 229.839
R134 VPB.t4 VPB.t5 229.839
R135 VPB.t3 VPB.t4 229.839
R136 VPB.t8 VPB.t7 199.195
R137 B1.n1 B1.n0 263.762
R138 B1.n2 B1.t0 263.762
R139 B1.n1 B1.t1 185.351
R140 B1.n2 B1.t2 183.891
R141 B1.n4 B1.n3 152
R142 B1.n3 B1.n2 40.8975
R143 B1.n3 B1.n1 24.8308
R144 B1.n4 B1 8.49281
R145 B1 B1.n4 3.32358
R146 VPWR.n7 VPWR.t5 367.733
R147 VPWR.n8 VPWR.t6 352.957
R148 VPWR.n23 VPWR.t0 351.637
R149 VPWR.n21 VPWR.n1 334.173
R150 VPWR.n16 VPWR.n4 219.417
R151 VPWR.n4 VPWR.t3 38.6969
R152 VPWR.n20 VPWR.n2 36.1417
R153 VPWR.n10 VPWR.n9 36.1417
R154 VPWR.n10 VPWR.n5 36.1417
R155 VPWR.n14 VPWR.n5 36.1417
R156 VPWR.n15 VPWR.n14 36.1417
R157 VPWR.n22 VPWR.n21 32.0005
R158 VPWR.n4 VPWR.t4 29.9023
R159 VPWR.n23 VPWR.n22 29.3652
R160 VPWR.n9 VPWR.n8 27.8593
R161 VPWR.n1 VPWR.t2 26.3844
R162 VPWR.n1 VPWR.t1 26.3844
R163 VPWR.n16 VPWR.n15 25.6005
R164 VPWR.n16 VPWR.n2 18.824
R165 VPWR.n9 VPWR.n6 9.3005
R166 VPWR.n11 VPWR.n10 9.3005
R167 VPWR.n12 VPWR.n5 9.3005
R168 VPWR.n14 VPWR.n13 9.3005
R169 VPWR.n15 VPWR.n3 9.3005
R170 VPWR.n17 VPWR.n16 9.3005
R171 VPWR.n18 VPWR.n2 9.3005
R172 VPWR.n20 VPWR.n19 9.3005
R173 VPWR.n22 VPWR.n0 9.3005
R174 VPWR.n24 VPWR.n23 7.25439
R175 VPWR.n8 VPWR.n7 6.93617
R176 VPWR.n21 VPWR.n20 4.14168
R177 VPWR.n7 VPWR.n6 0.462773
R178 VPWR VPWR.n24 0.157727
R179 VPWR.n24 VPWR.n0 0.150046
R180 VPWR.n11 VPWR.n6 0.122949
R181 VPWR.n12 VPWR.n11 0.122949
R182 VPWR.n13 VPWR.n12 0.122949
R183 VPWR.n13 VPWR.n3 0.122949
R184 VPWR.n17 VPWR.n3 0.122949
R185 VPWR.n18 VPWR.n17 0.122949
R186 VPWR.n19 VPWR.n18 0.122949
R187 VPWR.n19 VPWR.n0 0.122949
R188 a_820_392.n0 a_820_392.t0 401.555
R189 a_820_392.n0 a_820_392.t2 305.462
R190 a_820_392.n1 a_820_392.n0 187.292
R191 a_820_392.n1 a_820_392.t3 29.5505
R192 a_820_392.t1 a_820_392.n1 29.5505
R193 A1_N.n0 A1_N.t0 250.909
R194 A1_N.n0 A1_N.t1 204.048
R195 A1_N A1_N.n0 158.251
C0 VPB B2 0.074352f
C1 A1_N A2_N 0.066429f
C2 VPB B1 0.08029f
C3 VPB VPWR 0.217649f
C4 A1_N VPWR 0.046056f
C5 VPB X 0.029488f
C6 A2_N VPWR 0.014451f
C7 B2 B1 0.112751f
C8 VPB VGND 0.015736f
C9 A1_N X 0.002961f
C10 A1_N VGND 0.00679f
C11 B2 VPWR 0.035665f
C12 B2 X 9.47e-20
C13 A2_N VGND 0.00829f
C14 B1 VPWR 0.031301f
C15 B2 VGND 0.017158f
C16 B1 VGND 0.034121f
C17 VPWR X 0.423696f
C18 VPB A1_N 0.033038f
C19 VPWR VGND 0.116902f
C20 VPB A2_N 0.042492f
C21 X VGND 0.292131f
C22 VGND VNB 0.875228f
C23 X VNB 0.0834f
C24 VPWR VNB 0.697916f
C25 B1 VNB 0.264618f
C26 B2 VNB 0.22173f
C27 A2_N VNB 0.127087f
C28 A1_N VNB 0.106876f
C29 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2bb2o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2o_2 VNB VPB VPWR VGND B2 B1 A2_N X A1_N
X0 a_293_333.t0 A2_N.t0 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.2575 ps=1.59 w=0.55 l=0.15
X1 a_221_74.t0 B2.t0 a_149_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X2 a_61_392.t1 B2.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X3 VPWR.t0 B1.t0 a_61_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X4 VPWR.t1 A1_N.t0 a_546_378.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1959 pd=1.48 as=0.12 ps=1.24 w=1 l=0.15
X5 a_149_74.t0 B1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.2109 ps=2.05 w=0.74 l=0.15
X6 VGND.t5 a_293_333.t3 a_221_74.t1 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2575 pd=1.59 as=0.1443 ps=1.13 w=0.74 l=0.15
X7 VPWR.t3 a_221_74.t3 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t0 a_221_74.t4 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1959 ps=1.48 w=1.12 l=0.15
X9 a_546_378.t1 A2_N.t1 a_293_333.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.275 ps=2.55 w=1 l=0.15
X10 VGND.t4 A1_N.t1 a_293_333.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.131 pd=1.13 as=0.077 ps=0.83 w=0.55 l=0.15
X11 X.t3 a_221_74.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.131 ps=1.13 w=0.74 l=0.15
X12 a_221_74.t2 a_293_333.t4 a_61_392.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X13 VGND.t2 a_221_74.t6 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A2_N.n0 A2_N.t1 298.572
R1 A2_N.n0 A2_N.t0 196.013
R2 A2_N A2_N.n0 156.671
R3 VGND.n5 VGND.n4 216.155
R4 VGND.n10 VGND.n9 185
R5 VGND.n8 VGND.n7 185
R6 VGND.n3 VGND.t2 181.968
R7 VGND.n17 VGND.t0 156.062
R8 VGND.n9 VGND.n8 117.819
R9 VGND.n4 VGND.t1 46.9117
R10 VGND.n16 VGND.n15 36.1417
R11 VGND.n15 VGND.n1 34.3915
R12 VGND.n4 VGND.t4 31.6369
R13 VGND.n6 VGND.n5 30.8711
R14 VGND.n9 VGND.t5 30.548
R15 VGND.n8 VGND.t3 30.546
R16 VGND.n18 VGND.n17 13.0652
R17 VGND.n7 VGND.n6 11.8331
R18 VGND.n16 VGND.n0 9.3005
R19 VGND.n15 VGND.n14 9.3005
R20 VGND.n13 VGND.n1 9.3005
R21 VGND.n12 VGND.n11 9.3005
R22 VGND.n6 VGND.n2 9.3005
R23 VGND.n17 VGND.n16 7.52991
R24 VGND.n5 VGND.n3 6.74296
R25 VGND.n11 VGND.n10 5.84951
R26 VGND.n11 VGND.n7 3.30646
R27 VGND.n10 VGND.n1 2.28924
R28 VGND.n3 VGND.n2 0.436958
R29 VGND.n12 VGND.n2 0.122949
R30 VGND.n13 VGND.n12 0.122949
R31 VGND.n14 VGND.n13 0.122949
R32 VGND.n14 VGND.n0 0.122949
R33 VGND.n18 VGND.n0 0.122949
R34 VGND VGND.n18 0.0617245
R35 a_293_333.t1 a_293_333.n2 364.12
R36 a_293_333.n1 a_293_333.t4 280.632
R37 a_293_333.n2 a_293_333.n0 267.24
R38 a_293_333.n2 a_293_333.n1 216.268
R39 a_293_333.n1 a_293_333.t3 154.24
R40 a_293_333.n0 a_293_333.t2 30.546
R41 a_293_333.n0 a_293_333.t0 30.546
R42 VNB.t4 VNB.t5 2309.71
R43 VNB VNB.t0 1547.51
R44 VNB.t6 VNB.t2 1247.24
R45 VNB.t1 VNB.t4 1247.24
R46 VNB.t2 VNB.t3 993.177
R47 VNB.t5 VNB.t6 993.177
R48 VNB.t0 VNB.t1 831.496
R49 B2.n0 B2.t1 298.572
R50 B2.n0 B2.t0 178.34
R51 B2 B2.n0 152.173
R52 a_149_74.t0 a_149_74.t1 34.0546
R53 a_221_74.n4 a_221_74.n3 419.296
R54 a_221_74.n1 a_221_74.t5 273.938
R55 a_221_74.n1 a_221_74.t4 246.892
R56 a_221_74.n3 a_221_74.t3 226.809
R57 a_221_74.t2 a_221_74.n4 219.07
R58 a_221_74.n2 a_221_74.t6 196.013
R59 a_221_74.n4 a_221_74.n0 189.648
R60 a_221_74.n2 a_221_74.n1 91.2884
R61 a_221_74.n0 a_221_74.t1 31.6221
R62 a_221_74.n0 a_221_74.t0 31.6221
R63 a_221_74.n3 a_221_74.n2 5.11262
R64 VPWR.n3 VPWR.t3 883.885
R65 VPWR.n5 VPWR.n4 604.201
R66 VPWR.n12 VPWR.n1 318.087
R67 VPWR.n6 VPWR.n2 36.1417
R68 VPWR.n10 VPWR.n2 36.1417
R69 VPWR.n11 VPWR.n10 36.1417
R70 VPWR.n4 VPWR.t1 35.4605
R71 VPWR.n6 VPWR.n5 35.0123
R72 VPWR.n4 VPWR.t4 32.13
R73 VPWR.n1 VPWR.t2 29.5505
R74 VPWR.n1 VPWR.t0 29.5505
R75 VPWR.n12 VPWR.n11 11.6711
R76 VPWR.n7 VPWR.n6 9.3005
R77 VPWR.n8 VPWR.n2 9.3005
R78 VPWR.n10 VPWR.n9 9.3005
R79 VPWR.n11 VPWR.n0 9.3005
R80 VPWR.n13 VPWR.n12 7.69275
R81 VPWR.n5 VPWR.n3 5.3337
R82 VPWR.n7 VPWR.n3 0.62172
R83 VPWR VPWR.n13 0.163498
R84 VPWR.n13 VPWR.n0 0.144349
R85 VPWR.n8 VPWR.n7 0.122949
R86 VPWR.n9 VPWR.n8 0.122949
R87 VPWR.n9 VPWR.n0 0.122949
R88 a_61_392.t0 a_61_392.n0 536.523
R89 a_61_392.n0 a_61_392.t2 29.5505
R90 a_61_392.n0 a_61_392.t1 29.5505
R91 VPB.t3 VPB.t4 561.828
R92 VPB VPB.t0 334.543
R93 VPB.t1 VPB.t5 260.485
R94 VPB.t5 VPB.t6 229.839
R95 VPB.t2 VPB.t3 229.839
R96 VPB.t0 VPB.t2 229.839
R97 VPB.t4 VPB.t1 199.195
R98 B1.n0 B1.t0 274.473
R99 B1 B1.n0 215.022
R100 B1.n0 B1.t1 156.431
R101 A1_N.n0 A1_N.t0 279.829
R102 A1_N.n0 A1_N.t1 208.868
R103 A1_N.n1 A1_N.n0 152
R104 A1_N A1_N.n1 7.56414
R105 A1_N.n1 A1_N 6.78838
R106 a_546_378.t0 a_546_378.t1 47.2805
R107 X X.n0 586.03
R108 X.n3 X.n2 185
R109 X.n2 X.n1 185
R110 X.n0 X.t1 26.3844
R111 X.n0 X.t0 26.3844
R112 X.n2 X.t2 22.7032
R113 X.n2 X.t3 22.7032
R114 X.n1 X 9.56372
R115 X X.n3 7.2097
R116 X.n3 X 3.67866
R117 X.n1 X 1.32464
C0 VPB VPWR 0.144625f
C1 B1 B2 0.121101f
C2 VPB A2_N 0.038952f
C3 B1 VPWR 0.022458f
C4 B2 VPWR 0.021003f
C5 VPB A1_N 0.0373f
C6 VPB X 0.002421f
C7 VPB VGND 0.013787f
C8 VPWR A2_N 0.0061f
C9 B1 VGND 0.040332f
C10 VPWR A1_N 0.018167f
C11 VPWR X 0.017781f
C12 B2 VGND 0.027838f
C13 A2_N A1_N 0.115932f
C14 A2_N X 4.01e-19
C15 VPWR VGND 0.0811f
C16 A2_N VGND 0.015392f
C17 A1_N X 0.069452f
C18 VPB B1 0.057916f
C19 A1_N VGND 0.037974f
C20 VPB B2 0.03554f
C21 X VGND 0.165553f
C22 VGND VNB 0.671875f
C23 X VNB 0.019176f
C24 A1_N VNB 0.124232f
C25 A2_N VNB 0.129077f
C26 VPWR VNB 0.486897f
C27 B2 VNB 0.106836f
C28 B1 VNB 0.185311f
C29 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2o_1 VNB VPB VPWR VGND B2 A1_N X B1 A2_N
X0 a_258_392.t1 A1_N.t0 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1.24 as=0.199 ps=1.485 w=1 l=0.15
X1 a_257_126.t2 A1_N.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.118675 ps=1.08 w=0.55 l=0.15
X2 a_530_392.t0 a_257_126.t3 a_93_264.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X3 a_93_264.t0 a_257_126.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.212 ps=1.37 w=0.64 l=0.15
X4 VGND.t3 A2_N.t0 a_257_126.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.212 pd=1.37 as=0.077 ps=0.83 w=0.55 l=0.15
X5 a_605_126.t0 B2.t0 a_93_264.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0896 ps=0.92 w=0.64 l=0.15
X6 VGND.t2 a_93_264.t3 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.118675 pd=1.08 as=0.1961 ps=2.01 w=0.74 l=0.15
X7 VGND.t1 B1.t0 a_605_126.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1248 ps=1.03 w=0.64 l=0.15
X8 VPWR.t2 a_93_264.t4 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.199 pd=1.485 as=0.308 ps=2.79 w=1.12 l=0.15
X9 a_257_126.t1 A2_N.t1 a_258_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.12 ps=1.24 w=1 l=0.15
X10 VPWR.t1 B2.t1 a_530_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X11 a_530_392.t1 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.165 ps=1.33 w=1 l=0.15
R0 A1_N.n0 A1_N.t0 279.829
R1 A1_N A1_N.n0 163.834
R2 A1_N.n0 A1_N.t1 147.814
R3 VPWR.n2 VPWR.n0 324.077
R4 VPWR.n2 VPWR.n1 319.969
R5 VPWR.n0 VPWR.t3 42.3555
R6 VPWR.n1 VPWR.t0 32.5055
R7 VPWR.n1 VPWR.t1 32.5055
R8 VPWR.n0 VPWR.t2 27.4811
R9 VPWR VPWR.n2 0.234694
R10 a_258_392.t0 a_258_392.t1 47.2805
R11 VPB.t4 VPB.t1 495.43
R12 VPB VPB.t3 357.527
R13 VPB.t3 VPB.t5 263.038
R14 VPB.t2 VPB.t0 245.161
R15 VPB.t1 VPB.t2 229.839
R16 VPB.t5 VPB.t4 199.195
R17 VGND.n6 VGND.t1 301.683
R18 VGND.n5 VGND.n4 168.659
R19 VGND.n1 VGND.n0 123.008
R20 VGND.n4 VGND.t3 82.5992
R21 VGND.n4 VGND.t0 56.9974
R22 VGND.n0 VGND.t4 44.7031
R23 VGND.n9 VGND.n3 36.1417
R24 VGND.n10 VGND.n9 36.1417
R25 VGND.n11 VGND.n10 36.1417
R26 VGND.n0 VGND.t2 22.147
R27 VGND.n6 VGND.n5 21.7759
R28 VGND.n5 VGND.n3 15.8123
R29 VGND.n13 VGND.n1 11.4685
R30 VGND.n12 VGND.n11 9.3005
R31 VGND.n10 VGND.n2 9.3005
R32 VGND.n9 VGND.n8 9.3005
R33 VGND.n7 VGND.n3 9.3005
R34 VGND.n11 VGND.n1 7.52991
R35 VGND.n7 VGND.n6 6.35487
R36 VGND VGND.n13 0.163644
R37 VGND.n13 VGND.n12 0.144205
R38 VGND.n8 VGND.n7 0.122949
R39 VGND.n8 VGND.n2 0.122949
R40 VGND.n12 VGND.n2 0.122949
R41 a_257_126.t1 a_257_126.n1 593.699
R42 a_257_126.t4 a_257_126.n0 559.153
R43 a_257_126.n1 a_257_126.t3 236.983
R44 a_257_126.n1 a_257_126.t4 184.768
R45 a_257_126.n0 a_257_126.t0 30.546
R46 a_257_126.n0 a_257_126.t2 30.546
R47 VNB.t3 VNB.t0 2032.55
R48 VNB VNB.t2 1662.99
R49 VNB.t5 VNB.t1 1247.24
R50 VNB.t2 VNB.t4 1131.76
R51 VNB.t0 VNB.t5 993.177
R52 VNB.t4 VNB.t3 993.177
R53 a_93_264.t1 a_93_264.n2 853.639
R54 a_93_264.n2 a_93_264.n0 325.8
R55 a_93_264.n1 a_93_264.t4 258.942
R56 a_93_264.n2 a_93_264.n1 214.518
R57 a_93_264.n1 a_93_264.t3 187.981
R58 a_93_264.n0 a_93_264.t2 26.2505
R59 a_93_264.n0 a_93_264.t0 26.2505
R60 a_530_392.n0 a_530_392.t1 510.469
R61 a_530_392.n0 a_530_392.t2 29.5505
R62 a_530_392.t0 a_530_392.n0 29.5505
R63 A2_N.n0 A2_N.t1 285.719
R64 A2_N A2_N.n0 162.282
R65 A2_N.n0 A2_N.t0 147.814
R66 B2.n0 B2.t1 236.983
R67 B2.n0 B2.t0 184.768
R68 B2 B2.n0 153.244
R69 a_605_126.t0 a_605_126.t1 73.1255
R70 X.n1 X 588.678
R71 X.n1 X.n0 585
R72 X.n2 X.n1 585
R73 X X.t0 198.847
R74 X.n1 X.t1 26.3844
R75 X X.n2 9.85797
R76 X X.n0 8.53383
R77 X X.n0 2.35452
R78 X.n2 X 1.03039
R79 B1.t0 B1.t1 456.293
R80 B1.n0 B1.t0 310.057
R81 B1.n0 B1 10.6415
R82 B1 B1.n0 4.16436
C0 B2 VGND 0.026971f
C1 B1 VPWR 0.020568f
C2 X VPWR 0.117214f
C3 B1 VGND 0.185369f
C4 VPB A1_N 0.038618f
C5 X VGND 0.095014f
C6 VPB A2_N 0.043201f
C7 VPWR VGND 0.070984f
C8 VPB B2 0.040875f
C9 A1_N A2_N 0.103911f
C10 VPB B1 0.043165f
C11 VPB X 0.023244f
C12 VPB VPWR 0.120321f
C13 A1_N X 0.005656f
C14 A1_N VPWR 0.016863f
C15 VPB VGND 0.01421f
C16 B2 B1 0.056593f
C17 A2_N X 1.9e-19
C18 A1_N VGND 0.020474f
C19 A2_N VPWR 0.005825f
C20 B2 VPWR 0.018384f
C21 A2_N VGND 0.014153f
C22 VGND VNB 0.586296f
C23 VPWR VNB 0.438396f
C24 X VNB 0.12094f
C25 B1 VNB 0.202358f
C26 B2 VNB 0.102708f
C27 A2_N VNB 0.110634f
C28 A1_N VNB 0.106259f
C29 VPB VNB 1.04904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21boi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21boi_1 VNB VPB VPWR VGND B1_N Y A2 A1
X0 VPWR.t1 B1_N.t0 a_29_424.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.231 pd=2.23 as=0.231 ps=2.23 w=0.84 l=0.15
X1 Y.t0 a_29_424.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.170925 ps=1.27 w=0.74 l=0.15
X2 VGND.t2 B1_N.t1 a_29_424.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.170925 pd=1.27 as=0.14575 ps=1.63 w=0.55 l=0.15
X3 VGND.t0 A2.t0 a_437_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X4 a_437_74.t1 A1.t0 Y.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VPWR.t0 A1.t1 a_348_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_348_368.t1 A2.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.1848 ps=1.45 w=1.12 l=0.15
X7 a_348_368.t2 a_29_424.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
R0 B1_N.n0 B1_N.t0 295.166
R1 B1_N.n1 B1_N.t1 255.46
R2 B1_N B1_N.n0 160.922
R3 B1_N.n4 B1_N.n3 152
R4 B1_N.n3 B1_N.n2 119.749
R5 B1_N.n1 B1_N.n0 19.9453
R6 B1_N.n3 B1_N.n1 17.7292
R7 B1_N.n4 B1_N 10.0853
R8 B1_N.n2 B1_N 7.92216
R9 B1_N.n2 B1_N 6.07479
R10 B1_N B1_N.n4 4.26717
R11 a_29_424.t1 a_29_424.n1 459.236
R12 a_29_424.n0 a_29_424.t3 278.541
R13 a_29_424.n1 a_29_424.t0 236.052
R14 a_29_424.n1 a_29_424.n0 175.468
R15 a_29_424.n0 a_29_424.t2 171.161
R16 VPWR.n1 VPWR.t1 427.476
R17 VPWR.n1 VPWR.n0 321.897
R18 VPWR.n0 VPWR.t2 29.0228
R19 VPWR.n0 VPWR.t0 29.0228
R20 VPWR VPWR.n1 0.227504
R21 VPB.t2 VPB.t1 597.582
R22 VPB VPB.t2 252.823
R23 VPB.t0 VPB.t3 245.161
R24 VPB.t1 VPB.t0 229.839
R25 VGND.n1 VGND.t0 162.512
R26 VGND.n1 VGND.n0 105.578
R27 VGND.n0 VGND.t2 64.131
R28 VGND.n0 VGND.t1 40.0184
R29 VGND VGND.n1 0.429336
R30 Y.n2 Y 588.636
R31 Y.n2 Y.n0 585
R32 Y.n3 Y.n2 585
R33 Y Y.n1 175.841
R34 Y.n2 Y.t1 26.3844
R35 Y.n1 Y.t2 22.7032
R36 Y.n1 Y.t0 22.7032
R37 Y Y.n3 9.74595
R38 Y Y.n0 8.43686
R39 Y Y.n0 2.32777
R40 Y.n3 Y 1.01868
R41 VNB VNB.t2 2309.71
R42 VNB.t2 VNB.t1 1570.6
R43 VNB.t3 VNB.t0 1085.56
R44 VNB.t1 VNB.t3 993.177
R45 A2.n0 A2.t1 285.719
R46 A2.n0 A2.t0 178.34
R47 A2.n1 A2.n0 152
R48 A2.n1 A2 12.6275
R49 A2 A2.n1 3.97888
R50 a_437_74.t0 a_437_74.t1 51.8924
R51 A1.n0 A1.t1 250.909
R52 A1.n0 A1.t0 220.113
R53 A1 A1.n0 155.328
R54 a_348_368.n0 a_348_368.t1 578.764
R55 a_348_368.t0 a_348_368.n0 26.3844
R56 a_348_368.n0 a_348_368.t2 26.3844
C0 VPWR VGND 0.054956f
C1 Y VGND 0.11245f
C2 VPB B1_N 0.086728f
C3 VPB A1 0.032907f
C4 VPB A2 0.040765f
C5 VPB VPWR 0.111596f
C6 B1_N VPWR 0.020247f
C7 A1 A2 0.075863f
C8 VPB Y 0.02406f
C9 A1 VPWR 0.01626f
C10 VPB VGND 0.011193f
C11 B1_N Y 0.00376f
C12 A1 Y 0.054124f
C13 A2 VPWR 0.019359f
C14 B1_N VGND 0.081368f
C15 A2 Y 0.009487f
C16 A1 VGND 0.015587f
C17 A2 VGND 0.058201f
C18 VPWR Y 0.120622f
C19 VGND VNB 0.474756f
C20 Y VNB 0.022657f
C21 VPWR VNB 0.354238f
C22 A2 VNB 0.161068f
C23 A1 VNB 0.107359f
C24 B1_N VNB 0.410245f
C25 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21bo_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21bo_4 VNB VPB VPWR VGND B1_N A2 A1 X
X0 a_864_123.t1 A1.t0 a_187_338.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 X.t7 a_187_338.t6 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.161225 ps=1.195 w=0.74 l=0.15
X2 VPWR.t3 a_187_338.t7 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VGND.t8 A2.t0 a_864_123.t3 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 VGND.t0 a_187_338.t8 X.t6 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 X.t2 a_187_338.t9 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_187_338.t3 a_29_392.t2 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.12335 ps=1.095 w=0.64 l=0.15
X7 a_864_123.t2 A2.t1 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1088 pd=0.98 as=0.2016 ps=1.27 w=0.64 l=0.15
X8 VPWR.t1 a_187_338.t10 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 X.t0 a_187_338.t11 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.199 ps=1.485 w=1.12 l=0.15
X10 a_596_392.t1 A1.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR.t7 B1_N.t0 a_29_392.t1 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.199 pd=1.485 as=0.275 ps=2.55 w=1 l=0.15
X12 VPWR.t6 A2.t2 a_596_392.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X13 VPWR.t4 A1.t2 a_596_392.t0 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X14 X.t5 a_187_338.t12 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X15 VGND.t2 a_187_338.t13 X.t4 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.12335 pd=1.095 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_596_392.t3 a_29_392.t3 a_187_338.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X17 VGND.t7 a_29_392.t4 a_187_338.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.2016 pd=1.27 as=0.0896 ps=0.92 w=0.64 l=0.15
X18 a_187_338.t2 a_29_392.t5 a_596_392.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X19 VGND.t4 B1_N.t1 a_29_392.t0 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.161225 pd=1.195 as=0.1696 ps=1.81 w=0.64 l=0.15
X20 a_187_338.t1 A1.t3 a_864_123.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1088 ps=0.98 w=0.64 l=0.15
R0 A1.n1 A1.t1 220.917
R1 A1.n0 A1.t2 212.883
R2 A1.n0 A1.t0 171.148
R3 A1.n1 A1.t3 165.488
R4 A1.n3 A1.n2 152
R5 A1.n2 A1.n0 54.7732
R6 A1.n3 A1 10.8611
R7 A1 A1.n3 7.75808
R8 A1.n2 A1.n1 2.92171
R9 a_187_338.n15 a_187_338.n14 345.315
R10 a_187_338.n1 a_187_338.t11 262.764
R11 a_187_338.n8 a_187_338.t7 226.809
R12 a_187_338.n5 a_187_338.t9 226.809
R13 a_187_338.n2 a_187_338.t10 226.809
R14 a_187_338.n14 a_187_338.n13 181.315
R15 a_187_338.n9 a_187_338.t13 170.308
R16 a_187_338.n4 a_187_338.n0 165.189
R17 a_187_338.n1 a_187_338.t6 154.24
R18 a_187_338.n3 a_187_338.t8 154.24
R19 a_187_338.n7 a_187_338.t12 154.24
R20 a_187_338.n6 a_187_338.n0 152
R21 a_187_338.n10 a_187_338.n9 152
R22 a_187_338.n12 a_187_338.n11 99.0723
R23 a_187_338.n12 a_187_338.n10 45.6333
R24 a_187_338.n8 a_187_338.n7 35.7853
R25 a_187_338.n3 a_187_338.n2 32.8641
R26 a_187_338.n2 a_187_338.n1 29.9429
R27 a_187_338.n15 a_187_338.t4 29.5505
R28 a_187_338.t2 a_187_338.n15 29.5505
R29 a_187_338.n6 a_187_338.n5 27.0217
R30 a_187_338.n13 a_187_338.t0 26.2505
R31 a_187_338.n13 a_187_338.t1 26.2505
R32 a_187_338.n11 a_187_338.t5 26.2505
R33 a_187_338.n11 a_187_338.t3 26.2505
R34 a_187_338.n5 a_187_338.n4 22.6399
R35 a_187_338.n10 a_187_338.n0 13.1884
R36 a_187_338.n9 a_187_338.n8 10.955
R37 a_187_338.n4 a_187_338.n3 10.2247
R38 a_187_338.n14 a_187_338.n12 4.14168
R39 a_187_338.n7 a_187_338.n6 2.92171
R40 a_864_123.n1 a_864_123.n0 374.995
R41 a_864_123.n0 a_864_123.t2 37.5005
R42 a_864_123.n0 a_864_123.t0 26.2505
R43 a_864_123.n1 a_864_123.t3 26.2505
R44 a_864_123.t1 a_864_123.n1 26.2505
R45 VNB.t9 VNB.t7 1801.57
R46 VNB VNB.t6 1535.96
R47 VNB.t6 VNB.t3 1362.73
R48 VNB.t7 VNB.t4 1131.76
R49 VNB.t0 VNB.t8 1131.76
R50 VNB.t5 VNB.t10 993.177
R51 VNB.t4 VNB.t5 993.177
R52 VNB.t8 VNB.t9 993.177
R53 VNB.t1 VNB.t0 993.177
R54 VNB.t2 VNB.t1 993.177
R55 VNB.t3 VNB.t2 993.177
R56 VGND.n8 VGND.n6 236.953
R57 VGND.n4 VGND.n3 224.68
R58 VGND.n16 VGND.n15 218.792
R59 VGND.n7 VGND.t8 183.272
R60 VGND.n1 VGND.n0 131.118
R61 VGND.n6 VGND.t5 91.8755
R62 VGND.n8 VGND.n7 37.7524
R63 VGND.n10 VGND.n9 36.1417
R64 VGND.n18 VGND.n17 36.1417
R65 VGND.n3 VGND.t6 35.0202
R66 VGND.n0 VGND.t4 33.3822
R67 VGND.n14 VGND.n4 32.7534
R68 VGND.n0 VGND.t1 31.6698
R69 VGND.n6 VGND.t7 26.2505
R70 VGND.n15 VGND.t3 22.7032
R71 VGND.n15 VGND.t0 22.7032
R72 VGND.n3 VGND.t2 22.4442
R73 VGND.n10 VGND.n4 20.7064
R74 VGND.n20 VGND.n1 13.3508
R75 VGND.n16 VGND.n14 13.177
R76 VGND.n18 VGND.n1 11.6711
R77 VGND.n9 VGND.n5 9.3005
R78 VGND.n11 VGND.n10 9.3005
R79 VGND.n12 VGND.n4 9.3005
R80 VGND.n14 VGND.n13 9.3005
R81 VGND.n17 VGND.n2 9.3005
R82 VGND.n19 VGND.n18 9.3005
R83 VGND.n9 VGND.n8 6.02403
R84 VGND.n17 VGND.n16 4.14168
R85 VGND.n7 VGND.n5 0.16513
R86 VGND VGND.n20 0.163644
R87 VGND.n20 VGND.n19 0.144205
R88 VGND.n11 VGND.n5 0.122949
R89 VGND.n12 VGND.n11 0.122949
R90 VGND.n13 VGND.n12 0.122949
R91 VGND.n13 VGND.n2 0.122949
R92 VGND.n19 VGND.n2 0.122949
R93 X.n4 X.n3 623.452
R94 X.n6 X.n5 585
R95 X.n2 X.n0 147.032
R96 X.n2 X.n1 99.5845
R97 X.n4 X.n2 28.4148
R98 X.n5 X.t1 26.3844
R99 X.n5 X.t0 26.3844
R100 X.n3 X.t3 26.3844
R101 X.n3 X.t2 26.3844
R102 X.n1 X.t6 22.7032
R103 X.n1 X.t7 22.7032
R104 X.n0 X.t4 22.7032
R105 X.n0 X.t5 22.7032
R106 X X.n6 13.0174
R107 X.n6 X.n4 2.16999
R108 VPWR.n4 VPWR.t3 875.164
R109 VPWR.n19 VPWR.n1 606.528
R110 VPWR.n17 VPWR.n3 606.528
R111 VPWR.n8 VPWR.t4 358.646
R112 VPWR.n7 VPWR.n6 323.406
R113 VPWR.n1 VPWR.t7 42.3555
R114 VPWR.n11 VPWR.n10 36.1417
R115 VPWR.n12 VPWR.n11 36.1417
R116 VPWR.n6 VPWR.t5 29.5505
R117 VPWR.n6 VPWR.t6 29.5505
R118 VPWR.n12 VPWR.n4 27.8593
R119 VPWR.n1 VPWR.t0 27.3314
R120 VPWR.n3 VPWR.t2 26.3844
R121 VPWR.n3 VPWR.t1 26.3844
R122 VPWR.n18 VPWR.n17 24.0946
R123 VPWR.n17 VPWR.n16 23.3417
R124 VPWR.n16 VPWR.n4 19.577
R125 VPWR.n19 VPWR.n18 18.824
R126 VPWR.n10 VPWR.n7 15.8123
R127 VPWR.n10 VPWR.n9 9.3005
R128 VPWR.n11 VPWR.n5 9.3005
R129 VPWR.n13 VPWR.n12 9.3005
R130 VPWR.n14 VPWR.n4 9.3005
R131 VPWR.n16 VPWR.n15 9.3005
R132 VPWR.n17 VPWR.n2 9.3005
R133 VPWR.n18 VPWR.n0 9.3005
R134 VPWR.n8 VPWR.n7 8.75696
R135 VPWR.n20 VPWR.n19 7.44972
R136 VPWR.n9 VPWR.n8 0.521381
R137 VPWR VPWR.n20 0.160299
R138 VPWR.n20 VPWR.n0 0.147507
R139 VPWR.n9 VPWR.n5 0.122949
R140 VPWR.n13 VPWR.n5 0.122949
R141 VPWR.n14 VPWR.n13 0.122949
R142 VPWR.n15 VPWR.n14 0.122949
R143 VPWR.n15 VPWR.n2 0.122949
R144 VPWR.n2 VPWR.n0 0.122949
R145 VPB.t3 VPB.t6 495.43
R146 VPB.t9 VPB.t0 263.038
R147 VPB VPB.t9 252.823
R148 VPB.t5 VPB.t4 229.839
R149 VPB.t7 VPB.t5 229.839
R150 VPB.t8 VPB.t7 229.839
R151 VPB.t6 VPB.t8 229.839
R152 VPB.t2 VPB.t3 229.839
R153 VPB.t1 VPB.t2 229.839
R154 VPB.t0 VPB.t1 229.839
R155 A2.n1 A2.t0 639.308
R156 A2.t0 A2.n0 460.31
R157 A2.t1 A2.t2 460.31
R158 A2.n1 A2.t1 158.831
R159 A2 A2.n1 157.042
R160 a_29_392.n3 a_29_392.n2 376.606
R161 a_29_392.n0 a_29_392.t3 352.527
R162 a_29_392.n3 a_29_392.t0 258.76
R163 a_29_392.t1 a_29_392.n3 225.696
R164 a_29_392.n1 a_29_392.t5 212.883
R165 a_29_392.n2 a_29_392.t2 178.632
R166 a_29_392.n0 a_29_392.t4 162.385
R167 a_29_392.n2 a_29_392.n1 29.9429
R168 a_29_392.n1 a_29_392.n0 26.4733
R169 a_596_392.n1 a_596_392.t2 420.572
R170 a_596_392.n2 a_596_392.n1 285.695
R171 a_596_392.n1 a_596_392.n0 183.911
R172 a_596_392.n0 a_596_392.t4 29.5505
R173 a_596_392.n0 a_596_392.t3 29.5505
R174 a_596_392.n2 a_596_392.t0 29.5505
R175 a_596_392.t1 a_596_392.n2 29.5505
R176 B1_N.t1 B1_N.t0 465.933
R177 B1_N.n0 B1_N.t1 331.38
R178 B1_N B1_N.n0 6.59444
R179 B1_N.n0 B1_N 4.3525
C0 B1_N VPWR 0.0149f
C1 A2 A1 0.143514f
C2 VPB X 0.00851f
C3 B1_N X 0.019033f
C4 A2 VPWR 0.035522f
C5 VPB VGND 0.013502f
C6 A1 VPWR 0.027469f
C7 B1_N VGND 0.10866f
C8 A2 VGND 0.139808f
C9 VPWR X 0.043815f
C10 A1 VGND 0.00834f
C11 VPWR VGND 0.103621f
C12 X VGND 0.276067f
C13 VPB B1_N 0.045764f
C14 VPB A2 0.070755f
C15 B1_N A2 9.77e-19
C16 VPB A1 0.075554f
C17 VPB VPWR 0.171401f
C18 VGND VNB 0.816828f
C19 X VNB 0.020094f
C20 VPWR VNB 0.589313f
C21 A1 VNB 0.169883f
C22 A2 VNB 0.42084f
C23 B1_N VNB 0.219101f
C24 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21bo_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21bo_2 VNB VPB VPWR VGND B1_N A2 A1 X
X0 VPWR.t2 a_187_244.t3 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X1 X.t2 a_187_244.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1918 ps=1.485 w=1.12 l=0.15
X2 VGND.t0 A2.t0 a_587_74.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1184 ps=1.06 w=0.74 l=0.15
X3 a_587_74.t1 A1.t0 a_187_244.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VPWR.t4 B1_N.t0 a_32_368.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1918 pd=1.485 as=0.231 ps=2.23 w=0.84 l=0.15
X5 VGND.t4 B1_N.t1 a_32_368.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.13295 pd=1.125 as=0.14575 ps=1.63 w=0.55 l=0.15
X6 a_504_392.t0 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X7 VPWR.t3 A1.t1 a_504_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X8 a_504_392.t1 a_32_368.t2 a_187_244.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X9 X.t1 a_187_244.t5 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.13295 ps=1.125 w=0.74 l=0.15
X10 VGND.t1 a_187_244.t6 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_187_244.t2 a_32_368.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.24605 ps=1.405 w=0.74 l=0.15
R0 a_187_244.t0 a_187_244.n4 474.76
R1 a_187_244.n1 a_187_244.t4 361.233
R2 a_187_244.n3 a_187_244.t3 285.719
R3 a_187_244.n4 a_187_244.n3 229.161
R4 a_187_244.n2 a_187_244.t6 165.196
R5 a_187_244.n1 a_187_244.t5 154.24
R6 a_187_244.n4 a_187_244.n0 109.445
R7 a_187_244.n2 a_187_244.n1 56.2338
R8 a_187_244.n0 a_187_244.t1 22.7032
R9 a_187_244.n0 a_187_244.t2 22.7032
R10 a_187_244.n3 a_187_244.n2 13.146
R11 X X.n1 649.716
R12 X X.n0 211.786
R13 X.n1 X.t3 26.3844
R14 X.n1 X.t2 26.3844
R15 X.n0 X.t0 22.7032
R16 X.n0 X.t1 22.7032
R17 VPWR.n4 VPWR.t2 854.837
R18 VPWR.n6 VPWR.n1 654.255
R19 VPWR.n3 VPWR.n2 623.016
R20 VPWR.n1 VPWR.t4 52.7684
R21 VPWR.n2 VPWR.t0 29.5505
R22 VPWR.n2 VPWR.t3 29.5505
R23 VPWR.n1 VPWR.t1 28.2153
R24 VPWR.n5 VPWR.n4 25.224
R25 VPWR.n6 VPWR.n5 17.6946
R26 VPWR.n5 VPWR.n0 9.3005
R27 VPWR.n7 VPWR.n6 7.49287
R28 VPWR.n4 VPWR.n3 6.99282
R29 VPWR.n3 VPWR.n0 0.230598
R30 VPWR VPWR.n7 0.160867
R31 VPWR.n7 VPWR.n0 0.146947
R32 VPB.t3 VPB.t1 495.43
R33 VPB.t5 VPB.t2 263.038
R34 VPB VPB.t5 260.485
R35 VPB.t4 VPB.t0 229.839
R36 VPB.t1 VPB.t4 229.839
R37 VPB.t2 VPB.t3 229.839
R38 A2.n0 A2.t0 244.715
R39 A2.n0 A2.t1 229.452
R40 A2 A2.n0 154.133
R41 a_587_74.t0 a_587_74.t1 51.8924
R42 VGND.n1 VGND.n0 234.014
R43 VGND.n4 VGND.t0 166.722
R44 VGND.n5 VGND.n3 92.1689
R45 VGND.n0 VGND.t4 52.3641
R46 VGND.n3 VGND.t3 49.4131
R47 VGND.n3 VGND.t1 49.4131
R48 VGND.n7 VGND.n6 36.1417
R49 VGND.n0 VGND.t2 22.3201
R50 VGND.n9 VGND.n1 14.1038
R51 VGND.n7 VGND.n1 10.9181
R52 VGND.n8 VGND.n7 9.3005
R53 VGND.n6 VGND.n2 9.3005
R54 VGND.n5 VGND.n4 7.11628
R55 VGND.n6 VGND.n5 4.14168
R56 VGND.n4 VGND.n2 0.245265
R57 VGND VGND.n9 0.163644
R58 VGND.n9 VGND.n8 0.144205
R59 VGND.n8 VGND.n2 0.122949
R60 VNB.t2 VNB.t4 1882.41
R61 VNB VNB.t5 1501.31
R62 VNB.t5 VNB.t3 1235.7
R63 VNB.t1 VNB.t0 1085.56
R64 VNB.t4 VNB.t1 993.177
R65 VNB.t3 VNB.t2 993.177
R66 A1.n0 A1.t1 287.861
R67 A1.n0 A1.t0 191.194
R68 A1 A1.n0 155.815
R69 B1_N.n0 B1_N.t0 231.226
R70 B1_N B1_N.n0 158.573
R71 B1_N.n0 B1_N.t1 138.306
R72 a_32_368.t1 a_32_368.n1 420.048
R73 a_32_368.n1 a_32_368.n0 331.183
R74 a_32_368.n1 a_32_368.t0 325.075
R75 a_32_368.n0 a_32_368.t2 271.26
R76 a_32_368.n0 a_32_368.t3 167.094
R77 a_504_392.t0 a_504_392.n0 588.841
R78 a_504_392.n0 a_504_392.t2 29.5505
R79 a_504_392.n0 a_504_392.t1 29.5505
C0 A2 VGND 0.041081f
C1 VPWR X 0.015538f
C2 VPWR VGND 0.063781f
C3 B1_N X 0.001359f
C4 B1_N VGND 0.013788f
C5 X VGND 0.114514f
C6 VPB A1 0.038685f
C7 VPB A2 0.05263f
C8 VPB VPWR 0.123042f
C9 A1 A2 0.102481f
C10 A1 VPWR 0.01942f
C11 VPB B1_N 0.047594f
C12 A2 VPWR 0.015295f
C13 VPB X 0.003082f
C14 VPB VGND 0.010063f
C15 VPWR B1_N 0.010409f
C16 A1 VGND 0.024331f
C17 VGND VNB 0.535546f
C18 X VNB 0.009833f
C19 B1_N VNB 0.179942f
C20 VPWR VNB 0.393362f
C21 A2 VNB 0.161755f
C22 A1 VNB 0.113023f
C23 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21bo_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21bo_1 VNB VPB VPWR VGND X B1_N A1 A2
X0 a_122_136.t0 A2.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1696 ps=1.81 w=0.64 l=0.15
X1 a_194_136.t1 a_272_110.t2 a_34_392.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X2 a_34_392.t0 A1.t0 VPWR.t3 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.165 ps=1.33 w=1 l=0.15
X3 X.t0 a_194_136.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.203 ps=1.505 w=1.12 l=0.15
X4 VPWR.t1 B1_N.t0 a_272_110.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.231 ps=2.23 w=0.84 l=0.15
X5 a_194_136.t0 A1.t1 a_122_136.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0672 ps=0.85 w=0.64 l=0.15
X6 VPWR.t0 A2.t1 a_34_392.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.275 ps=2.55 w=1 l=0.15
X7 VGND.t3 a_272_110.t3 a_194_136.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1248 ps=1.03 w=0.64 l=0.15
X8 X.t1 a_194_136.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.113125 ps=1.065 w=0.74 l=0.15
X9 VGND.t2 B1_N.t1 a_272_110.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.113125 pd=1.065 as=0.15675 ps=1.67 w=0.55 l=0.15
R0 A2.t0 A2.t1 442.904
R1 A2 A2.t0 332.426
R2 VGND.n1 VGND.t3 292.106
R3 VGND.n7 VGND.t1 282.611
R4 VGND.n3 VGND.n2 231.031
R5 VGND.n8 VGND.n7 43.1829
R6 VGND.n6 VGND.n5 36.1417
R7 VGND.n2 VGND.t2 34.9096
R8 VGND.n2 VGND.t0 29.4571
R9 VGND.n5 VGND.n1 21.4593
R10 VGND.n5 VGND.n4 9.3005
R11 VGND.n6 VGND.n0 9.3005
R12 VGND.n3 VGND.n1 7.18202
R13 VGND.n7 VGND.n6 2.25932
R14 VGND.n4 VGND.n3 0.233531
R15 VGND.n4 VGND.n0 0.122949
R16 VGND.n8 VGND.n0 0.122949
R17 VGND VGND.n8 0.0617245
R18 a_122_136.t0 a_122_136.t1 39.3755
R19 VNB.t4 VNB.t2 3083.46
R20 VNB.t3 VNB.t4 1247.24
R21 VNB VNB.t1 1235.7
R22 VNB.t2 VNB.t0 1097.11
R23 VNB.t1 VNB.t3 831.496
R24 a_272_110.t1 a_272_110.n1 817.283
R25 a_272_110.n0 a_272_110.t2 295.894
R26 a_272_110.n1 a_272_110.t0 249.103
R27 a_272_110.n1 a_272_110.n0 205.667
R28 a_272_110.n0 a_272_110.t3 147.011
R29 a_34_392.n0 a_34_392.t1 485.414
R30 a_34_392.n0 a_34_392.t2 29.5505
R31 a_34_392.t0 a_34_392.n0 29.5505
R32 a_194_136.n2 a_194_136.n0 314.149
R33 a_194_136.n0 a_194_136.t3 258.942
R34 a_194_136.t1 a_194_136.n2 227.877
R35 a_194_136.n0 a_194_136.t4 210.474
R36 a_194_136.n2 a_194_136.n1 193.179
R37 a_194_136.n1 a_194_136.t2 43.1255
R38 a_194_136.n1 a_194_136.t0 30.0005
R39 VPB.t4 VPB.t2 666.533
R40 VPB.t2 VPB.t3 273.253
R41 VPB VPB.t1 265.591
R42 VPB.t1 VPB.t0 245.161
R43 VPB.t0 VPB.t4 229.839
R44 A1.n0 A1.t0 236.983
R45 A1.n0 A1.t1 168.701
R46 A1 A1.n0 157.042
R47 VPWR.n2 VPWR.n0 657.49
R48 VPWR.n2 VPWR.n1 337.241
R49 VPWR.n0 VPWR.t1 55.1136
R50 VPWR.n1 VPWR.t3 32.5055
R51 VPWR.n1 VPWR.t0 32.5055
R52 VPWR.n0 VPWR.t2 29.6087
R53 VPWR VPWR.n2 0.195732
R54 X.n1 X 589.923
R55 X.n1 X.n0 585
R56 X.n2 X.n1 585
R57 X X.t1 208.173
R58 X.n1 X.t0 26.3844
R59 X X.n2 13.1943
R60 X X.n0 11.422
R61 X X.n0 3.15127
R62 X.n2 X 1.37896
R63 B1_N.n0 B1_N.t0 240.732
R64 B1_N.n0 B1_N.t1 208.868
R65 B1_N B1_N.n0 158.788
C0 VPB A1 0.042255f
C1 VPB VPWR 0.126114f
C2 A2 A1 0.065479f
C3 VPB B1_N 0.040009f
C4 A2 VPWR 0.017499f
C5 A1 VPWR 0.018233f
C6 A2 B1_N 9.98e-19
C7 VPB X 0.016937f
C8 VPB VGND 0.014198f
C9 A2 X 8.06e-20
C10 A2 VGND 0.137501f
C11 VPWR B1_N 0.009319f
C12 A1 VGND 0.023743f
C13 VPWR X 0.071044f
C14 VPWR VGND 0.063454f
C15 B1_N X 0.007072f
C16 B1_N VGND 0.019503f
C17 X VGND 0.096309f
C18 VPB A2 0.038346f
C19 VGND VNB 0.54678f
C20 X VNB 0.122637f
C21 B1_N VNB 0.137823f
C22 VPWR VNB 0.390883f
C23 A1 VNB 0.101369f
C24 A2 VNB 0.204818f
C25 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a2bb2oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2oi_4 VNB VPB VPWR VGND A2_N Y B2 B1 A1_N
X0 Y.t10 B2.t0 a_914_74# VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 Y.t1 a_114_392.t4 VGND.t5 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_29_392.t1 A1_N.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X3 a_539_368.t3 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 Y.t9 B2.t1 a_914_74# VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X5 VPWR.t1 A1_N.t1 a_29_392.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X6 a_29_392.t2 A2_N.t0 a_114_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X7 VPWR.t7 B1.t1 a_539_368.t2 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8 VGND.t0 A1_N.t2 a_114_392.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_539_368.t11 B2.t2 VPWR.t6 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 VPWR.t5 B2.t3 a_539_368.t10 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 VPWR.t4 B2.t4 a_539_368.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 VGND.t4 a_114_392.t5 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VGND.t6 B1.t2 a_914_74# VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X14 a_539_368.t7 a_114_392.t6 Y.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_539_368.t8 B2.t5 VPWR.t3 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 VGND.t3 a_114_392.t7 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 VGND.t7 B1.t3 a_914_74# VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 Y.t4 a_114_392.t8 a_539_368.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_539_368.t5 a_114_392.t9 Y.t5 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 a_914_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 Y.t6 a_114_392.t10 a_539_368.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X22 a_114_392.t2 A2_N.t1 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X23 a_914_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X24 a_114_392.t3 A2_N.t2 a_29_392.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X25 a_914_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X26 Y.t7 a_114_392.t11 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1184 ps=1.06 w=0.74 l=0.15
X27 a_914_74# B2.t6 Y.t8 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 a_539_368.t1 B1.t4 VPWR.t8 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X29 VPWR.t9 B1.t5 a_539_368.t0 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 B2.n5 B2.t3 236.303
R1 B2.n1 B2.t2 226.809
R2 B2.n4 B2.t4 226.809
R3 B2.n10 B2.t5 226.809
R4 B2.n1 B2.n0 196.744
R5 B2.n5 B2.t1 196.013
R6 B2.n11 B2.t6 196.013
R7 B2.n3 B2.t0 196.013
R8 B2 B2.n2 152.744
R9 B2.n13 B2.n12 152
R10 B2.n9 B2.n8 152
R11 B2.n7 B2.n6 152
R12 B2.n9 B2.n6 49.6611
R13 B2.n12 B2.n11 37.9763
R14 B2.n2 B2.n1 37.246
R15 B2.n3 B2.n2 24.8308
R16 B2.n12 B2.n4 21.1793
R17 B2.n7 B2 13.247
R18 B2 B2.n13 9.37724
R19 B2.n8 B2 9.07957
R20 B2.n11 B2.n10 6.57323
R21 B2.n8 B2 5.2098
R22 B2.n10 B2.n9 5.11262
R23 B2.n13 B2 4.91213
R24 B2.n4 B2.n3 3.65202
R25 B2.n6 B2.n5 1.46111
R26 B2 B2.n7 1.04236
R27 Y.n2 Y.n0 362.596
R28 Y.n2 Y.n1 314.017
R29 Y.n4 Y.t10 305.579
R30 Y.n4 Y.n3 185
R31 Y.n7 Y.n6 155.244
R32 Y.n7 Y.n5 97.4026
R33 Y Y.n7 51.577
R34 Y.n8 Y.n4 37.8672
R35 Y.n0 Y.t5 26.3844
R36 Y.n0 Y.t6 26.3844
R37 Y.n1 Y.t0 26.3844
R38 Y.n1 Y.t4 26.3844
R39 Y Y.n2 26.2626
R40 Y.n5 Y.t2 22.7032
R41 Y.n5 Y.t1 22.7032
R42 Y.n6 Y.t3 22.7032
R43 Y.n6 Y.t7 22.7032
R44 Y.n3 Y.t8 22.7032
R45 Y.n3 Y.t9 22.7032
R46 Y.n8 Y 4.32991
R47 Y Y.n8 3.53153
R48 VNB.t1 VNB.t7 3233.6
R49 VNB VNB.t5 3048.82
R50 VNB.t10 VNB.t9 1986.35
R51 VNB.t8 VNB.t10 1986.35
R52 VNB.t2 VNB.t4 1085.56
R53 VNB.t6 VNB.t8 993.177
R54 VNB.t7 VNB.t6 993.177
R55 VNB.t0 VNB.t1 993.177
R56 VNB.t3 VNB.t0 993.177
R57 VNB.t4 VNB.t3 993.177
R58 VNB.t5 VNB.t2 993.177
R59 a_114_392.n11 a_114_392.n10 392.844
R60 a_114_392.n1 a_114_392.t6 368.462
R61 a_114_392.n1 a_114_392.t8 281.702
R62 a_114_392.n7 a_114_392.t11 279.269
R63 a_114_392.n3 a_114_392.t9 261.62
R64 a_114_392.n6 a_114_392.t10 261.62
R65 a_114_392.n5 a_114_392.t4 154.24
R66 a_114_392.n7 a_114_392.t7 154.24
R67 a_114_392.n2 a_114_392.t5 154.24
R68 a_114_392.n9 a_114_392.n8 152
R69 a_114_392.n10 a_114_392.n0 112.686
R70 a_114_392.n2 a_114_392.n1 97.715
R71 a_114_392.n10 a_114_392.n9 83.3349
R72 a_114_392.n9 a_114_392.n4 78.1582
R73 a_114_392.n8 a_114_392.n6 44.549
R74 a_114_392.n4 a_114_392.n3 33.1053
R75 a_114_392.t1 a_114_392.n11 29.5505
R76 a_114_392.n11 a_114_392.t3 29.5505
R77 a_114_392.n0 a_114_392.t0 22.7032
R78 a_114_392.n0 a_114_392.t2 22.7032
R79 a_114_392.n5 a_114_392.n4 20.7371
R80 a_114_392.n8 a_114_392.n7 13.146
R81 a_114_392.n6 a_114_392.n5 5.11262
R82 a_114_392.n3 a_114_392.n2 2.19141
R83 VGND.n17 VGND.t4 295.89
R84 VGND.n7 VGND.t6 249.677
R85 VGND.n6 VGND.t7 242.263
R86 VGND.n26 VGND.n25 216.78
R87 VGND.n19 VGND.n18 205.364
R88 VGND.n28 VGND.t1 138.751
R89 VGND.n10 VGND.n5 36.1417
R90 VGND.n11 VGND.n10 36.1417
R91 VGND.n12 VGND.n11 36.1417
R92 VGND.n12 VGND.n3 36.1417
R93 VGND.n16 VGND.n3 36.1417
R94 VGND.n24 VGND.n1 36.1417
R95 VGND.n20 VGND.n17 33.1299
R96 VGND.n28 VGND.n27 30.8711
R97 VGND.n25 VGND.t2 25.9464
R98 VGND.n25 VGND.t0 25.9464
R99 VGND.n18 VGND.t5 22.7032
R100 VGND.n18 VGND.t3 22.7032
R101 VGND.n6 VGND.n5 15.0593
R102 VGND.n17 VGND.n16 14.3064
R103 VGND.n8 VGND.n5 9.3005
R104 VGND.n10 VGND.n9 9.3005
R105 VGND.n11 VGND.n4 9.3005
R106 VGND.n13 VGND.n12 9.3005
R107 VGND.n14 VGND.n3 9.3005
R108 VGND.n16 VGND.n15 9.3005
R109 VGND.n17 VGND.n2 9.3005
R110 VGND.n21 VGND.n20 9.3005
R111 VGND.n22 VGND.n1 9.3005
R112 VGND.n24 VGND.n23 9.3005
R113 VGND.n27 VGND.n0 9.3005
R114 VGND.n7 VGND.n6 9.04071
R115 VGND.n27 VGND.n26 9.03579
R116 VGND.n20 VGND.n19 6.77697
R117 VGND.n29 VGND.n28 6.69578
R118 VGND.n26 VGND.n24 5.27109
R119 VGND.n19 VGND.n1 4.51815
R120 VGND.n8 VGND.n7 0.990573
R121 VGND VGND.n29 0.267593
R122 VGND.n29 VGND.n0 0.163093
R123 VGND.n9 VGND.n8 0.122949
R124 VGND.n9 VGND.n4 0.122949
R125 VGND.n13 VGND.n4 0.122949
R126 VGND.n14 VGND.n13 0.122949
R127 VGND.n15 VGND.n14 0.122949
R128 VGND.n15 VGND.n2 0.122949
R129 VGND.n21 VGND.n2 0.122949
R130 VGND.n22 VGND.n21 0.122949
R131 VGND.n23 VGND.n22 0.122949
R132 VGND.n23 VGND.n0 0.122949
R133 A1_N.n0 A1_N.t1 266.171
R134 A1_N.n1 A1_N.t2 258.673
R135 A1_N.n0 A1_N.t0 218.482
R136 A1_N.n2 A1_N.n1 152
R137 A1_N.n1 A1_N.n0 13.146
R138 A1_N A1_N.n2 11.8308
R139 A1_N.n2 A1_N 6.78838
R140 VPWR.n10 VPWR.n9 343.06
R141 VPWR.n15 VPWR.n14 331.5
R142 VPWR.n13 VPWR.n6 323.406
R143 VPWR.n8 VPWR.n7 323.406
R144 VPWR.n28 VPWR.n1 323.156
R145 VPWR.n20 VPWR.n4 36.1417
R146 VPWR.n21 VPWR.n20 36.1417
R147 VPWR.n22 VPWR.n21 36.1417
R148 VPWR.n22 VPWR.n2 36.1417
R149 VPWR.n26 VPWR.n2 36.1417
R150 VPWR.n27 VPWR.n26 36.1417
R151 VPWR.n28 VPWR.n27 34.2593
R152 VPWR.n16 VPWR.n15 33.8829
R153 VPWR.n1 VPWR.t2 29.5505
R154 VPWR.n1 VPWR.t1 29.5505
R155 VPWR.n16 VPWR.n13 27.4829
R156 VPWR.n14 VPWR.t3 26.3844
R157 VPWR.n14 VPWR.t5 26.3844
R158 VPWR.n6 VPWR.t6 26.3844
R159 VPWR.n6 VPWR.t4 26.3844
R160 VPWR.n7 VPWR.t0 26.3844
R161 VPWR.n7 VPWR.t7 26.3844
R162 VPWR.n9 VPWR.t8 26.3844
R163 VPWR.n9 VPWR.t9 26.3844
R164 VPWR.n13 VPWR.n12 25.977
R165 VPWR.n12 VPWR.n8 16.9417
R166 VPWR.n12 VPWR.n11 9.3005
R167 VPWR.n13 VPWR.n5 9.3005
R168 VPWR.n17 VPWR.n16 9.3005
R169 VPWR.n18 VPWR.n4 9.3005
R170 VPWR.n20 VPWR.n19 9.3005
R171 VPWR.n21 VPWR.n3 9.3005
R172 VPWR.n23 VPWR.n22 9.3005
R173 VPWR.n24 VPWR.n2 9.3005
R174 VPWR.n26 VPWR.n25 9.3005
R175 VPWR.n27 VPWR.n0 9.3005
R176 VPWR.n10 VPWR.n8 7.44802
R177 VPWR.n29 VPWR.n28 6.88046
R178 VPWR.n15 VPWR.n4 2.25932
R179 VPWR.n11 VPWR.n10 0.72842
R180 VPWR VPWR.n29 0.392383
R181 VPWR.n29 VPWR.n0 0.161373
R182 VPWR.n11 VPWR.n5 0.122949
R183 VPWR.n17 VPWR.n5 0.122949
R184 VPWR.n18 VPWR.n17 0.122949
R185 VPWR.n19 VPWR.n18 0.122949
R186 VPWR.n19 VPWR.n3 0.122949
R187 VPWR.n23 VPWR.n3 0.122949
R188 VPWR.n24 VPWR.n23 0.122949
R189 VPWR.n25 VPWR.n24 0.122949
R190 VPWR.n25 VPWR.n0 0.122949
R191 a_29_392.n1 a_29_392.t3 325.712
R192 a_29_392.t1 a_29_392.n1 314.111
R193 a_29_392.n1 a_29_392.n0 184.216
R194 a_29_392.n0 a_29_392.t0 29.5505
R195 a_29_392.n0 a_29_392.t2 29.5505
R196 VPB.t2 VPB.t5 612.904
R197 VPB VPB.t4 252.823
R198 VPB.t15 VPB.t14 229.839
R199 VPB.t0 VPB.t15 229.839
R200 VPB.t13 VPB.t0 229.839
R201 VPB.t12 VPB.t13 229.839
R202 VPB.t10 VPB.t12 229.839
R203 VPB.t9 VPB.t10 229.839
R204 VPB.t11 VPB.t9 229.839
R205 VPB.t8 VPB.t11 229.839
R206 VPB.t7 VPB.t8 229.839
R207 VPB.t6 VPB.t7 229.839
R208 VPB.t5 VPB.t6 229.839
R209 VPB.t1 VPB.t2 229.839
R210 VPB.t3 VPB.t1 229.839
R211 VPB.t4 VPB.t3 229.839
R212 B1.n2 B1.t4 237.762
R213 B1.n12 B1.t5 226.809
R214 B1.n3 B1.t0 226.809
R215 B1.n6 B1.t1 226.809
R216 B1.n6 B1.t3 198.204
R217 B1.n2 B1.n1 196.013
R218 B1.n5 B1.n4 196.013
R219 B1.n11 B1.t2 196.013
R220 B1.n2 B1.n0 152
R221 B1.n14 B1.n13 152
R222 B1.n10 B1.n9 152
R223 B1.n8 B1.n7 152
R224 B1.n13 B1.n2 49.6611
R225 B1.n7 B1.n6 37.246
R226 B1.n11 B1.n10 36.5157
R227 B1.n7 B1.n5 23.3702
R228 B1.n10 B1.n3 21.1793
R229 B1.n0 B1 11.7586
R230 B1.n9 B1.n8 10.1214
R231 B1.n12 B1.n11 8.03383
R232 B1 B1.n14 7.5912
R233 B1.n14 B1 6.69817
R234 B1.n13 B1.n12 5.11262
R235 B1.n5 B1.n3 5.11262
R236 B1.n9 B1 3.42376
R237 B1 B1.n0 2.53073
R238 B1.n8 B1 0.744686
R239 a_539_368.n3 a_539_368.n2 304.901
R240 a_539_368.n3 a_539_368.t4 279.81
R241 a_539_368.n8 a_539_368.t1 274.788
R242 a_539_368.n7 a_539_368.n0 207.35
R243 a_539_368.n6 a_539_368.n5 205.487
R244 a_539_368.n9 a_539_368.n8 205.486
R245 a_539_368.n4 a_539_368.n1 189.115
R246 a_539_368.n4 a_539_368.n3 62.9747
R247 a_539_368.n6 a_539_368.n4 59.2902
R248 a_539_368.n8 a_539_368.n7 55.3417
R249 a_539_368.n7 a_539_368.n6 55.3417
R250 a_539_368.n0 a_539_368.t2 26.3844
R251 a_539_368.n0 a_539_368.t11 26.3844
R252 a_539_368.n1 a_539_368.t10 26.3844
R253 a_539_368.n1 a_539_368.t7 26.3844
R254 a_539_368.n2 a_539_368.t6 26.3844
R255 a_539_368.n2 a_539_368.t5 26.3844
R256 a_539_368.n5 a_539_368.t9 26.3844
R257 a_539_368.n5 a_539_368.t8 26.3844
R258 a_539_368.n9 a_539_368.t0 26.3844
R259 a_539_368.t3 a_539_368.n9 26.3844
R260 A2_N.n0 A2_N.t1 242.26
R261 A2_N.n0 A2_N.t0 215.561
R262 A2_N.n1 A2_N.t2 215.561
R263 A2_N.n4 A2_N.n3 190.113
R264 A2_N.n5 A2_N.n4 152
R265 A2_N A2_N.n2 81.7369
R266 A2_N.n1 A2_N.n0 45.188
R267 A2_N.n4 A2_N.n2 39.4232
R268 A2_N.n2 A2_N.n1 17.0332
R269 A2_N A2_N.n5 11.055
R270 A2_N.n3 A2_N 9.89141
R271 A2_N.n3 A2_N 4.46111
R272 A2_N.n5 A2_N 3.29747
C0 VPB Y 0.00845f
C1 A2_N VPWR 0.014337f
C2 VPB VGND 0.014046f
C3 B2 B1 0.075758f
C4 A2_N Y 0.001005f
C5 A1_N VPWR 0.03494f
C6 A2_N VGND 0.091121f
C7 A1_N Y 0.005013f
C8 B2 VPWR 0.068937f
C9 a_914_74# VPB 7.44e-19
C10 B1 VPWR 0.067994f
C11 A1_N VGND 0.018491f
C12 B2 Y 0.193541f
C13 a_914_74# A2_N 2.37e-19
C14 B1 Y 2.52e-19
C15 B2 VGND 0.029018f
C16 VPWR Y 0.020657f
C17 B1 VGND 0.063417f
C18 VPB A2_N 0.099244f
C19 a_914_74# B2 0.036729f
C20 VPWR VGND 0.136796f
C21 VPB A1_N 0.087303f
C22 a_914_74# B1 0.196999f
C23 Y VGND 0.29866f
C24 a_914_74# VPWR 0.004866f
C25 VPB B2 0.133818f
C26 A2_N A1_N 0.059593f
C27 a_914_74# Y 0.187872f
C28 VPB B1 0.143012f
C29 a_914_74# VGND 0.479182f
C30 VPB VPWR 0.21931f
C31 VGND VNB 1.03452f
C32 Y VNB 0.06263f
C33 VPWR VNB 0.796686f
C34 B1 VNB 0.446162f
C35 B2 VNB 0.404134f
C36 A1_N VNB 0.152609f
C37 A2_N VNB 0.44357f
C38 VPB VNB 2.01326f
C39 a_914_74# VNB 0.070067f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21o_4 VNB VPB VPWR VGND X B1 A2 A1
X0 VPWR.t5 a_91_48.t6 X.t3 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t1 A2.t0 a_503_392.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X2 X.t7 a_91_48.t7 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_503_392.t4 A1.t0 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X4 a_503_392.t1 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X5 a_700_74.t1 A2.t2 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X6 VPWR.t6 A1.t1 a_503_392.t3 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X7 VGND.t7 B1.t0 a_91_48.t3 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X8 a_503_392.t0 B1.t1 a_91_48.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X9 a_91_48.t5 B1.t2 a_503_392.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X10 VGND.t2 a_91_48.t8 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.12205 pd=1.08 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 X.t2 a_91_48.t9 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X12 VGND.t1 a_91_48.t10 X.t5 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 X.t4 a_91_48.t11 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X14 a_91_48.t2 B1.t3 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.12205 ps=1.08 w=0.64 l=0.15
X15 VGND.t5 A2.t3 a_700_74.t0 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X16 a_91_48.t4 A1.t2 a_700_74.t3 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X17 a_700_74.t2 A1.t3 a_91_48.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X18 VPWR.t3 a_91_48.t12 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X19 X.t0 a_91_48.t13 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 a_91_48.n16 a_91_48.n15 332.827
R1 a_91_48.n15 a_91_48.n0 259.498
R2 a_91_48.n11 a_91_48.t12 251.151
R3 a_91_48.n9 a_91_48.t13 240.197
R4 a_91_48.n2 a_91_48.t6 240.197
R5 a_91_48.n4 a_91_48.t9 240.197
R6 a_91_48.n4 a_91_48.t11 182.138
R7 a_91_48.n11 a_91_48.t8 179.947
R8 a_91_48.n3 a_91_48.t10 179.947
R9 a_91_48.n8 a_91_48.t7 179.947
R10 a_91_48.n6 a_91_48.n5 165.189
R11 a_91_48.n7 a_91_48.n6 152
R12 a_91_48.n10 a_91_48.n1 152
R13 a_91_48.n12 a_91_48.n11 152
R14 a_91_48.n14 a_91_48.n13 107.782
R15 a_91_48.n11 a_91_48.n10 49.6611
R16 a_91_48.n5 a_91_48.n4 37.246
R17 a_91_48.n8 a_91_48.n7 36.5157
R18 a_91_48.t1 a_91_48.n16 29.5505
R19 a_91_48.n16 a_91_48.t5 29.5505
R20 a_91_48.n13 a_91_48.t3 26.2505
R21 a_91_48.n13 a_91_48.t2 26.2505
R22 a_91_48.n0 a_91_48.t0 26.2505
R23 a_91_48.n0 a_91_48.t4 26.2505
R24 a_91_48.n15 a_91_48.n14 24.3
R25 a_91_48.n5 a_91_48.n3 23.3702
R26 a_91_48.n14 a_91_48.n12 21.6254
R27 a_91_48.n7 a_91_48.n2 21.1793
R28 a_91_48.n12 a_91_48.n1 13.1884
R29 a_91_48.n6 a_91_48.n1 13.1884
R30 a_91_48.n9 a_91_48.n8 8.03383
R31 a_91_48.n10 a_91_48.n9 5.11262
R32 a_91_48.n3 a_91_48.n2 5.11262
R33 X.n2 X.n1 262.94
R34 X.n2 X.n0 212.668
R35 X.n5 X.n4 154.35
R36 X.n5 X.n3 100.181
R37 X X.n2 48.2215
R38 X X.n5 38.5478
R39 X.n1 X.t1 26.3844
R40 X.n1 X.t0 26.3844
R41 X.n0 X.t3 26.3844
R42 X.n0 X.t2 26.3844
R43 X.n3 X.t5 22.7032
R44 X.n3 X.t4 22.7032
R45 X.n4 X.t6 22.7032
R46 X.n4 X.t7 22.7032
R47 VPWR.n19 VPWR.t4 420.425
R48 VPWR.n17 VPWR.n2 325.255
R49 VPWR.n6 VPWR.n5 323.406
R50 VPWR.n8 VPWR.n7 321.207
R51 VPWR.n3 VPWR.t3 257.433
R52 VPWR.n11 VPWR.n10 36.1417
R53 VPWR.n12 VPWR.n11 36.1417
R54 VPWR.n5 VPWR.t7 29.5505
R55 VPWR.n5 VPWR.t6 29.5505
R56 VPWR.n7 VPWR.t0 29.5505
R57 VPWR.n7 VPWR.t1 29.5505
R58 VPWR.n17 VPWR.n16 28.2358
R59 VPWR.n16 VPWR.n3 26.7299
R60 VPWR.n12 VPWR.n3 26.7299
R61 VPWR.n2 VPWR.t2 26.3844
R62 VPWR.n2 VPWR.t5 26.3844
R63 VPWR.n18 VPWR.n17 25.224
R64 VPWR.n19 VPWR.n18 17.6946
R65 VPWR.n10 VPWR.n6 16.9417
R66 VPWR.n10 VPWR.n9 9.3005
R67 VPWR.n11 VPWR.n4 9.3005
R68 VPWR.n13 VPWR.n12 9.3005
R69 VPWR.n14 VPWR.n3 9.3005
R70 VPWR.n16 VPWR.n15 9.3005
R71 VPWR.n17 VPWR.n1 9.3005
R72 VPWR.n18 VPWR.n0 9.3005
R73 VPWR.n20 VPWR.n19 9.3005
R74 VPWR.n8 VPWR.n6 7.54965
R75 VPWR.n9 VPWR.n8 0.585966
R76 VPWR.n9 VPWR.n4 0.122949
R77 VPWR.n13 VPWR.n4 0.122949
R78 VPWR.n14 VPWR.n13 0.122949
R79 VPWR.n15 VPWR.n14 0.122949
R80 VPWR.n15 VPWR.n1 0.122949
R81 VPWR.n1 VPWR.n0 0.122949
R82 VPWR.n20 VPWR.n0 0.122949
R83 VPWR VPWR.n20 0.0617245
R84 VPB.t4 VPB.t9 495.43
R85 VPB VPB.t5 278.361
R86 VPB.t2 VPB.t0 229.839
R87 VPB.t8 VPB.t2 229.839
R88 VPB.t7 VPB.t8 229.839
R89 VPB.t1 VPB.t7 229.839
R90 VPB.t9 VPB.t1 229.839
R91 VPB.t3 VPB.t4 229.839
R92 VPB.t6 VPB.t3 229.839
R93 VPB.t5 VPB.t6 229.839
R94 A2.n1 A2.t0 268.873
R95 A2.n0 A2.t1 263.762
R96 A2.n0 A2.t2 185.351
R97 A2.n1 A2.t3 183.161
R98 A2 A2.n2 158.524
R99 A2.n2 A2.n0 54.7732
R100 A2.n2 A2.n1 5.84292
R101 a_503_392.n1 a_503_392.t5 336.437
R102 a_503_392.n2 a_503_392.t1 292.913
R103 a_503_392.n3 a_503_392.n2 208.775
R104 a_503_392.n1 a_503_392.n0 183.911
R105 a_503_392.n2 a_503_392.n1 80.3282
R106 a_503_392.n0 a_503_392.t3 29.5505
R107 a_503_392.n0 a_503_392.t0 29.5505
R108 a_503_392.t2 a_503_392.n3 29.5505
R109 a_503_392.n3 a_503_392.t4 29.5505
R110 VGND.n6 VGND.t7 240.73
R111 VGND.n16 VGND.t0 231.946
R112 VGND.n9 VGND.n8 221.096
R113 VGND.n14 VGND.n2 217
R114 VGND.n5 VGND.n4 213.742
R115 VGND.n8 VGND.t6 37.5005
R116 VGND.n10 VGND.n7 36.1417
R117 VGND.n14 VGND.n1 31.624
R118 VGND.n4 VGND.t4 26.2505
R119 VGND.n4 VGND.t5 26.2505
R120 VGND.n2 VGND.t3 22.7032
R121 VGND.n2 VGND.t1 22.7032
R122 VGND.n8 VGND.t2 22.1988
R123 VGND.n15 VGND.n14 21.8358
R124 VGND.n16 VGND.n15 18.0711
R125 VGND.n9 VGND.n1 14.3064
R126 VGND.n7 VGND.n6 11.2946
R127 VGND.n17 VGND.n16 9.3005
R128 VGND.n15 VGND.n0 9.3005
R129 VGND.n14 VGND.n13 9.3005
R130 VGND.n12 VGND.n1 9.3005
R131 VGND.n7 VGND.n3 9.3005
R132 VGND.n11 VGND.n10 9.3005
R133 VGND.n6 VGND.n5 7.63801
R134 VGND.n10 VGND.n9 3.01226
R135 VGND.n5 VGND.n3 0.161883
R136 VGND.n11 VGND.n3 0.122949
R137 VGND.n12 VGND.n11 0.122949
R138 VGND.n13 VGND.n12 0.122949
R139 VGND.n13 VGND.n0 0.122949
R140 VGND.n17 VGND.n0 0.122949
R141 VGND VGND.n17 0.0617245
R142 VNB.t8 VNB.t9 2540.68
R143 VNB VNB.t1 1224.15
R144 VNB.t3 VNB.t7 1131.76
R145 VNB.t5 VNB.t6 993.177
R146 VNB.t0 VNB.t5 993.177
R147 VNB.t9 VNB.t0 993.177
R148 VNB.t7 VNB.t8 993.177
R149 VNB.t4 VNB.t3 993.177
R150 VNB.t2 VNB.t4 993.177
R151 VNB.t1 VNB.t2 993.177
R152 A1.n0 A1.t3 254.827
R153 A1.n1 A1.t2 244.214
R154 A1.n1 A1.t1 223.839
R155 A1.n0 A1.t0 212.883
R156 A1.n2 A1.n1 152
R157 A1.n1 A1.n0 54.7732
R158 A1.n2 A1 12.6066
R159 A1 A1.n2 6.01262
R160 a_700_74.t1 a_700_74.n1 218.421
R161 a_700_74.n1 a_700_74.t3 212.448
R162 a_700_74.n1 a_700_74.n0 86.3508
R163 a_700_74.n0 a_700_74.t0 26.2505
R164 a_700_74.n0 a_700_74.t2 26.2505
R165 B1.n0 B1.t1 282.627
R166 B1.n2 B1.t3 248.157
R167 B1.n0 B1.t2 216.9
R168 B1.n1 B1.t0 207.261
R169 B1 B1.n2 153.299
R170 B1.n2 B1.n1 21.9096
R171 B1.n1 B1.n0 18.2581
C0 VPWR VGND 0.095495f
C1 X VGND 0.284169f
C2 VPB B1 0.112009f
C3 VPB A1 0.074534f
C4 VPB A2 0.080982f
C5 B1 A1 0.047875f
C6 VPB VPWR 0.173747f
C7 B1 A2 2.59e-20
C8 A1 A2 0.101188f
C9 VPB X 0.016905f
C10 B1 VPWR 0.01708f
C11 A1 VPWR 0.035236f
C12 B1 X 0.003238f
C13 VPB VGND 0.01256f
C14 A2 VPWR 0.037033f
C15 A1 X 1.69e-19
C16 B1 VGND 0.031411f
C17 A1 VGND 0.012965f
C18 VPWR X 0.40715f
C19 A2 VGND 0.032388f
C20 VGND VNB 0.730138f
C21 X VNB 0.077649f
C22 VPWR VNB 0.579887f
C23 A2 VNB 0.256288f
C24 A1 VNB 0.216082f
C25 B1 VNB 0.249529f
C26 VPB VNB 1.37045f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21o_2 VNB VPB VPWR VGND B1 A2 A1 X
X0 VGND.t2 a_84_244.t3 X.t3 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2442 pd=1.4 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 a_401_392.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X2 VPWR.t3 A1.t0 a_401_392.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X3 a_401_392.t2 B1.t0 a_84_244.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X4 X.t1 a_84_244.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X5 a_484_74.t1 A1.t1 a_84_244.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X6 a_84_244.t0 B1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2442 ps=1.4 w=0.74 l=0.15
X7 VPWR.t1 a_84_244.t5 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t2 a_84_244.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X9 VGND.t3 A2.t1 a_484_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1184 ps=1.06 w=0.74 l=0.15
R0 a_84_244.n1 a_84_244.t4 285.719
R1 a_84_244.t2 a_84_244.n4 277.361
R2 a_84_244.n2 a_84_244.t5 261.62
R3 a_84_244.n4 a_84_244.n3 170.258
R4 a_84_244.n4 a_84_244.n0 168.119
R5 a_84_244.n1 a_84_244.t6 154.24
R6 a_84_244.n3 a_84_244.t3 154.24
R7 a_84_244.n2 a_84_244.n1 41.6278
R8 a_84_244.n0 a_84_244.t1 22.7032
R9 a_84_244.n0 a_84_244.t0 22.7032
R10 a_84_244.n3 a_84_244.n2 21.1793
R11 X.n2 X 590.715
R12 X.n2 X.n0 585
R13 X.n3 X.n2 585
R14 X X.n1 140.09
R15 X.n2 X.t0 26.3844
R16 X.n2 X.t1 26.3844
R17 X.n1 X.t3 22.7032
R18 X.n1 X.t2 22.7032
R19 X X.n3 15.3148
R20 X X.n0 13.2576
R21 X X.n0 3.65764
R22 X.n3 X 1.6005
R23 VGND.n3 VGND.n1 185
R24 VGND.n5 VGND.n4 185
R25 VGND.n11 VGND.t1 175.351
R26 VGND.n2 VGND.t3 166.083
R27 VGND.n4 VGND.n3 61.6221
R28 VGND.n5 VGND.n2 36.2871
R29 VGND.n10 VGND.n9 36.1417
R30 VGND.n4 VGND.t0 22.7032
R31 VGND.n3 VGND.t2 22.7032
R32 VGND.n12 VGND.n11 13.4417
R33 VGND.n11 VGND.n10 13.177
R34 VGND.n7 VGND.n6 9.3005
R35 VGND.n9 VGND.n8 9.3005
R36 VGND.n10 VGND.n0 9.3005
R37 VGND.n6 VGND.n1 6.10381
R38 VGND.n9 VGND.n1 3.49345
R39 VGND.n7 VGND.n2 0.581012
R40 VGND.n6 VGND.n5 0.339573
R41 VGND.n8 VGND.n7 0.122949
R42 VGND.n8 VGND.n0 0.122949
R43 VGND.n12 VGND.n0 0.122949
R44 VGND VGND.n12 0.0617245
R45 VNB.t2 VNB.t0 1870.87
R46 VNB VNB.t1 1559.06
R47 VNB.t3 VNB.t4 1085.56
R48 VNB.t0 VNB.t3 993.177
R49 VNB.t1 VNB.t2 993.177
R50 A2.n0 A2.t0 305.082
R51 A2.n0 A2.t1 169.684
R52 A2 A2.n0 158.788
R53 VPWR.n5 VPWR.t2 259.171
R54 VPWR.n3 VPWR.t1 248.62
R55 VPWR.n2 VPWR.n1 227.459
R56 VPWR.n1 VPWR.t0 29.5505
R57 VPWR.n1 VPWR.t3 29.5505
R58 VPWR.n5 VPWR.n4 26.3534
R59 VPWR.n4 VPWR.n3 22.5887
R60 VPWR.n4 VPWR.n0 9.3005
R61 VPWR.n6 VPWR.n5 9.3005
R62 VPWR.n3 VPWR.n2 7.1337
R63 VPWR.n2 VPWR.n0 0.22781
R64 VPWR.n6 VPWR.n0 0.122949
R65 VPWR VPWR.n6 0.0617245
R66 a_401_392.t0 a_401_392.n0 524.865
R67 a_401_392.n0 a_401_392.t1 29.5505
R68 a_401_392.n0 a_401_392.t2 29.5505
R69 VPB.t1 VPB.t4 495.43
R70 VPB VPB.t2 260.485
R71 VPB.t3 VPB.t0 229.839
R72 VPB.t4 VPB.t3 229.839
R73 VPB.t2 VPB.t1 229.839
R74 A1.n0 A1.t0 298.572
R75 A1.n0 A1.t1 178.34
R76 A1 A1.n0 158.573
R77 B1.n0 B1.t0 313.738
R78 B1.n0 B1.t1 178.34
R79 B1 B1.n0 160.293
R80 a_484_74.t0 a_484_74.t1 51.8924
C0 VPB VGND 0.008159f
C1 B1 X 5.73e-19
C2 A1 VPWR 0.022793f
C3 B1 VGND 0.016661f
C4 A2 VPWR 0.022786f
C5 A1 VGND 0.025271f
C6 VPWR X 0.204828f
C7 A2 VGND 0.050091f
C8 VPWR VGND 0.065443f
C9 X VGND 0.133076f
C10 VPB B1 0.045075f
C11 VPB A1 0.036099f
C12 B1 A1 0.094064f
C13 VPB A2 0.04919f
C14 VPB VPWR 0.116291f
C15 B1 VPWR 0.015573f
C16 A1 A2 0.10373f
C17 VPB X 0.006181f
C18 VGND VNB 0.507483f
C19 X VNB 0.028066f
C20 VPWR VNB 0.390997f
C21 A2 VNB 0.172759f
C22 A1 VNB 0.107158f
C23 B1 VNB 0.112274f
C24 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21o_1 VNB VPB VPWR VGND X A1 B1 A2
X0 a_81_264.t1 B1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.14225 ps=1.14 w=0.64 l=0.15
X1 VGND.t1 A2.t0 a_452_136.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.104 ps=0.965 w=0.64 l=0.15
X2 VGND.t0 a_81_264.t3 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.14225 pd=1.14 as=0.1961 ps=2.01 w=0.74 l=0.15
X3 a_452_136.t0 A1.t0 a_81_264.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.104 pd=0.965 as=0.0896 ps=0.92 w=0.64 l=0.15
X4 VPWR.t2 a_81_264.t4 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.308 ps=2.79 w=1.12 l=0.15
X5 VPWR.t0 A1.t1 a_364_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X6 a_364_392.t1 A2.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.165 ps=1.33 w=1 l=0.15
X7 a_364_392.t2 B1.t1 a_81_264.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
R0 B1.n0 B1.t1 236.983
R1 B1.n0 B1.t0 168.701
R2 B1 B1.n0 154.91
R3 VGND.n1 VGND.t1 309.113
R4 VGND.n1 VGND.n0 221.226
R5 VGND.n0 VGND.t2 48.7505
R6 VGND.n0 VGND.t0 21.3263
R7 VGND VGND.n1 0.715943
R8 a_81_264.n1 a_81_264.t3 311.693
R9 a_81_264.t2 a_81_264.n2 259.786
R10 a_81_264.n1 a_81_264.t4 248.718
R11 a_81_264.n2 a_81_264.n1 180.703
R12 a_81_264.n2 a_81_264.n0 136.4
R13 a_81_264.n0 a_81_264.t0 26.2505
R14 a_81_264.n0 a_81_264.t1 26.2505
R15 VNB VNB.t1 2783.2
R16 VNB.t1 VNB.t3 1270.34
R17 VNB.t0 VNB.t2 1097.11
R18 VNB.t3 VNB.t0 993.177
R19 A2.t0 A2.t1 442.904
R20 A2 A2.t0 319.709
R21 a_452_136.t0 a_452_136.t1 60.938
R22 X.n1 X 589.572
R23 X.n1 X.n0 585
R24 X.n2 X.n1 585
R25 X X.t0 321.438
R26 X.n1 X.t1 26.3844
R27 X X.n2 12.2519
R28 X X.n0 10.6062
R29 X X.n0 2.92621
R30 X.n2 X 1.2805
R31 A1.n0 A1.t1 236.983
R32 A1.n0 A1.t0 168.701
R33 A1 A1.n0 157.237
R34 VPWR.n1 VPWR.n0 340.399
R35 VPWR.n1 VPWR.t2 265.171
R36 VPWR.n0 VPWR.t1 32.5055
R37 VPWR.n0 VPWR.t0 32.5055
R38 VPWR VPWR.n1 0.216971
R39 VPB.t2 VPB.t3 638.442
R40 VPB VPB.t2 252.823
R41 VPB.t0 VPB.t1 245.161
R42 VPB.t3 VPB.t0 229.839
R43 a_364_392.n0 a_364_392.t1 485.416
R44 a_364_392.t0 a_364_392.n0 29.5505
R45 a_364_392.n0 a_364_392.t2 29.5505
C0 X VGND 0.064045f
C1 B1 X 6.09e-19
C2 VPB VPWR 0.11808f
C3 VPWR VGND 0.055006f
C4 B1 VPWR 0.012361f
C5 VPB VGND 0.014088f
C6 VPB B1 0.04869f
C7 B1 VGND 0.010718f
C8 A1 VPWR 0.014368f
C9 VPB A1 0.040522f
C10 A1 VGND 0.017921f
C11 A2 VPWR 0.015432f
C12 VPB A2 0.040677f
C13 B1 A1 0.081198f
C14 A2 VGND 0.154331f
C15 A1 A2 0.05628f
C16 X VPWR 0.129116f
C17 VPB X 0.015614f
C18 VGND VNB 0.510322f
C19 VPWR VNB 0.361074f
C20 X VNB 0.117307f
C21 A2 VNB 0.196652f
C22 A1 VNB 0.098376f
C23 B1 VNB 0.094899f
C24 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21boi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21boi_4 VNB VPB VPWR VGND B1_N Y A2 A1
X0 VPWR.t7 A1.t0 a_31_368.t10 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X1 a_31_368.t11 a_803_323.t2 Y.t3 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_31_368.t2 a_803_323.t3 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t7 a_803_323.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 VGND.t0 A2.t0 a_46_74.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 Y.t8 A1.t1 a_46_74.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X6 Y.t1 a_803_323.t5 a_31_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 VGND.t1 A2.t1 a_46_74.t2 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_31_368.t3 A2.t2 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X9 VPWR.t1 A2.t3 a_31_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X10 a_31_368.t5 A2.t4 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 Y.t11 A1.t2 a_46_74.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_46_74.t1 A2.t5 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t3 A2.t6 a_31_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_31_368.t9 A1.t3 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 VGND.t4 a_803_323.t6 Y.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VPWR.t5 A1.t4 a_31_368.t8 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 a_46_74.t5 A1.t5 Y.t10 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X18 a_31_368.t7 A1.t6 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 a_46_74.t4 A1.t7 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 VGND.t3 a_803_323.t7 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 Y.t4 a_803_323.t8 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X22 VPWR.t8 B1_N.t0 a_803_323.t0 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.231 pd=2.23 as=0.126 ps=1.14 w=0.84 l=0.15
X23 a_803_323.t1 B1_N.t1 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.231 ps=2.23 w=0.84 l=0.15
X24 a_46_74.t0 A2.t7 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 Y.t0 a_803_323.t9 a_31_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A1.n4 A1.t0 236.303
R1 A1.n0 A1.t3 226.809
R2 A1.n3 A1.t4 226.809
R3 A1.n9 A1.t6 226.809
R4 A1.n0 A1.t5 196.744
R5 A1.n4 A1.t1 196.013
R6 A1.n10 A1.t7 196.013
R7 A1.n2 A1.t2 196.013
R8 A1 A1.n1 152.184
R9 A1.n12 A1.n11 152
R10 A1.n8 A1.n7 152
R11 A1.n6 A1.n5 152
R12 A1.n8 A1.n5 49.6611
R13 A1.n11 A1.n10 37.9763
R14 A1.n1 A1.n0 37.246
R15 A1.n2 A1.n1 24.8308
R16 A1.n11 A1.n3 21.1793
R17 A1.n6 A1 15.5434
R18 A1 A1.n12 12.2519
R19 A1.n7 A1 10.4234
R20 A1.n7 A1 7.13193
R21 A1.n10 A1.n9 6.57323
R22 A1.n12 A1 5.30336
R23 A1.n9 A1.n8 5.11262
R24 A1.n3 A1.n2 3.65202
R25 A1 A1.n6 2.01193
R26 A1.n5 A1.n4 1.46111
R27 a_31_368.n1 a_31_368.n0 308.902
R28 a_31_368.n4 a_31_368.t10 296.526
R29 a_31_368.n1 a_31_368.t2 290.063
R30 a_31_368.n4 a_31_368.n3 208.897
R31 a_31_368.n5 a_31_368.n2 207.35
R32 a_31_368.n7 a_31_368.n6 205.487
R33 a_31_368.n9 a_31_368.n8 188.095
R34 a_31_368.n8 a_31_368.n1 74.0228
R35 a_31_368.n5 a_31_368.n4 67.7652
R36 a_31_368.n8 a_31_368.n7 62.1501
R37 a_31_368.n7 a_31_368.n5 55.3417
R38 a_31_368.n3 a_31_368.t8 26.3844
R39 a_31_368.n3 a_31_368.t7 26.3844
R40 a_31_368.n2 a_31_368.t6 26.3844
R41 a_31_368.n2 a_31_368.t9 26.3844
R42 a_31_368.n6 a_31_368.t4 26.3844
R43 a_31_368.n6 a_31_368.t5 26.3844
R44 a_31_368.n0 a_31_368.t1 26.3844
R45 a_31_368.n0 a_31_368.t11 26.3844
R46 a_31_368.t0 a_31_368.n9 26.3844
R47 a_31_368.n9 a_31_368.t3 26.3844
R48 VPWR.n12 VPWR.t8 431.106
R49 VPWR.n11 VPWR.t9 352.079
R50 VPWR.n22 VPWR.n7 331.5
R51 VPWR.n5 VPWR.n4 323.406
R52 VPWR.n28 VPWR.n3 315.928
R53 VPWR.n30 VPWR.n1 315.926
R54 VPWR.n15 VPWR.n10 36.1417
R55 VPWR.n16 VPWR.n15 36.1417
R56 VPWR.n17 VPWR.n16 36.1417
R57 VPWR.n17 VPWR.n8 36.1417
R58 VPWR.n21 VPWR.n8 36.1417
R59 VPWR.n24 VPWR.n23 36.1417
R60 VPWR.n28 VPWR.n27 27.4829
R61 VPWR.n1 VPWR.t4 26.3844
R62 VPWR.n1 VPWR.t7 26.3844
R63 VPWR.n3 VPWR.t6 26.3844
R64 VPWR.n3 VPWR.t5 26.3844
R65 VPWR.n4 VPWR.t2 26.3844
R66 VPWR.n4 VPWR.t3 26.3844
R67 VPWR.n7 VPWR.t0 26.3844
R68 VPWR.n7 VPWR.t1 26.3844
R69 VPWR.n23 VPWR.n22 23.3417
R70 VPWR.n30 VPWR.n29 22.9652
R71 VPWR.n29 VPWR.n28 19.9534
R72 VPWR.n27 VPWR.n5 15.4358
R73 VPWR.n12 VPWR.n11 15.2558
R74 VPWR.n22 VPWR.n21 12.8005
R75 VPWR.n13 VPWR.n10 9.3005
R76 VPWR.n15 VPWR.n14 9.3005
R77 VPWR.n16 VPWR.n9 9.3005
R78 VPWR.n18 VPWR.n17 9.3005
R79 VPWR.n19 VPWR.n8 9.3005
R80 VPWR.n21 VPWR.n20 9.3005
R81 VPWR.n23 VPWR.n6 9.3005
R82 VPWR.n25 VPWR.n24 9.3005
R83 VPWR.n27 VPWR.n26 9.3005
R84 VPWR.n28 VPWR.n2 9.3005
R85 VPWR.n29 VPWR.n0 9.3005
R86 VPWR.n31 VPWR.n30 7.27223
R87 VPWR.n11 VPWR.n10 2.63579
R88 VPWR.n24 VPWR.n5 1.88285
R89 VPWR.n13 VPWR.n12 1.17896
R90 VPWR VPWR.n31 0.157962
R91 VPWR.n31 VPWR.n0 0.149814
R92 VPWR.n14 VPWR.n13 0.122949
R93 VPWR.n14 VPWR.n9 0.122949
R94 VPWR.n18 VPWR.n9 0.122949
R95 VPWR.n19 VPWR.n18 0.122949
R96 VPWR.n20 VPWR.n19 0.122949
R97 VPWR.n20 VPWR.n6 0.122949
R98 VPWR.n25 VPWR.n6 0.122949
R99 VPWR.n26 VPWR.n25 0.122949
R100 VPWR.n26 VPWR.n2 0.122949
R101 VPWR.n2 VPWR.n0 0.122949
R102 VPB.t2 VPB.t12 495.43
R103 VPB VPB.t10 257.93
R104 VPB.t12 VPB.t11 229.839
R105 VPB.t1 VPB.t2 229.839
R106 VPB.t13 VPB.t1 229.839
R107 VPB.t0 VPB.t13 229.839
R108 VPB.t3 VPB.t0 229.839
R109 VPB.t4 VPB.t3 229.839
R110 VPB.t5 VPB.t4 229.839
R111 VPB.t6 VPB.t5 229.839
R112 VPB.t9 VPB.t6 229.839
R113 VPB.t8 VPB.t9 229.839
R114 VPB.t7 VPB.t8 229.839
R115 VPB.t10 VPB.t7 229.839
R116 a_803_323.n9 a_803_323.n8 378.517
R117 a_803_323.n0 a_803_323.t5 326
R118 a_803_323.n1 a_803_323.t4 266.808
R119 a_803_323.n6 a_803_323.t3 234.841
R120 a_803_323.n3 a_803_323.t9 234.841
R121 a_803_323.n0 a_803_323.t2 223.743
R122 a_803_323.n7 a_803_323.t6 199.519
R123 a_803_323.n5 a_803_323.t8 186.374
R124 a_803_323.n2 a_803_323.t7 186.374
R125 a_803_323.n8 a_803_323.n7 152
R126 a_803_323.n2 a_803_323.n1 97.715
R127 a_803_323.n8 a_803_323.n4 81.6328
R128 a_803_323.n7 a_803_323.n6 44.549
R129 a_803_323.t0 a_803_323.n9 35.1791
R130 a_803_323.n9 a_803_323.t1 35.1791
R131 a_803_323.n1 a_803_323.n0 34.7921
R132 a_803_323.n4 a_803_323.n3 33.3172
R133 a_803_323.n5 a_803_323.n4 20.5774
R134 a_803_323.n6 a_803_323.n5 5.11262
R135 a_803_323.n3 a_803_323.n2 2.19141
R136 Y.n10 Y.n8 235.083
R137 Y.n1 Y.n0 230.298
R138 Y.n7 Y.n2 204.282
R139 Y.n10 Y.n9 185
R140 Y Y.n10 167.126
R141 Y.n5 Y.n3 148.974
R142 Y.n5 Y.n4 106.118
R143 Y.n2 Y.t3 26.3844
R144 Y.n2 Y.t1 26.3844
R145 Y.n0 Y.t2 26.3844
R146 Y.n0 Y.t0 26.3844
R147 Y Y.n1 22.9652
R148 Y.n9 Y.t10 22.7032
R149 Y.n9 Y.t11 22.7032
R150 Y.n8 Y.t9 22.7032
R151 Y.n8 Y.t8 22.7032
R152 Y.n3 Y.t6 22.7032
R153 Y.n3 Y.t4 22.7032
R154 Y.n4 Y.t5 22.7032
R155 Y.n4 Y.t7 22.7032
R156 Y.n6 Y 16.9417
R157 Y.n7 Y.n1 12.4957
R158 Y.n6 Y 10.9181
R159 Y Y.n5 10.9181
R160 Y Y.n7 6.95702
R161 Y.n7 Y 1.94833
R162 Y Y.n6 1.85557
R163 VGND.n5 VGND.t5 244.311
R164 VGND.n4 VGND.n3 218.024
R165 VGND.n12 VGND.n11 204.201
R166 VGND.n15 VGND.n14 204.201
R167 VGND.n2 VGND.t4 143.445
R168 VGND.n6 VGND.n4 36.1417
R169 VGND.n10 VGND.n1 36.1417
R170 VGND.n15 VGND.n13 33.8829
R171 VGND.n3 VGND.t2 22.7032
R172 VGND.n3 VGND.t3 22.7032
R173 VGND.n11 VGND.t7 22.7032
R174 VGND.n11 VGND.t0 22.7032
R175 VGND.n14 VGND.t6 22.7032
R176 VGND.n14 VGND.t1 22.7032
R177 VGND.n6 VGND.n5 9.78874
R178 VGND.n13 VGND.n0 9.3005
R179 VGND.n10 VGND.n9 9.3005
R180 VGND.n8 VGND.n1 9.3005
R181 VGND.n7 VGND.n6 9.3005
R182 VGND.n5 VGND.n1 7.52991
R183 VGND.n16 VGND.n15 6.43412
R184 VGND.n4 VGND.n2 6.33642
R185 VGND.n13 VGND.n12 6.02403
R186 VGND.n12 VGND.n10 5.27109
R187 VGND VGND.n16 0.631067
R188 VGND.n7 VGND.n2 0.552852
R189 VGND.n16 VGND.n0 0.168639
R190 VGND.n8 VGND.n7 0.122949
R191 VGND.n9 VGND.n8 0.122949
R192 VGND.n9 VGND.n0 0.122949
R193 VNB.t7 VNB.t5 2263.52
R194 VNB VNB.t11 1316.54
R195 VNB.t2 VNB.t4 993.177
R196 VNB.t3 VNB.t2 993.177
R197 VNB.t5 VNB.t3 993.177
R198 VNB.t0 VNB.t7 993.177
R199 VNB.t6 VNB.t0 993.177
R200 VNB.t1 VNB.t6 993.177
R201 VNB.t9 VNB.t1 993.177
R202 VNB.t10 VNB.t9 993.177
R203 VNB.t8 VNB.t10 993.177
R204 VNB.t11 VNB.t8 993.177
R205 A2.n0 A2.t2 237.642
R206 A2.n9 A2.t3 226.809
R207 A2.n2 A2.t4 226.809
R208 A2.n4 A2.t6 226.809
R209 A2.n4 A2.t1 198.204
R210 A2.n3 A2.t5 196.013
R211 A2.n8 A2.t0 196.013
R212 A2.n0 A2.t7 196.013
R213 A2 A2.n1 153.28
R214 A2 A2.n5 152.915
R215 A2.n11 A2.n10 152
R216 A2.n7 A2.n6 152
R217 A2.n10 A2.n1 49.6611
R218 A2.n8 A2.n7 40.8975
R219 A2.n5 A2.n4 32.8641
R220 A2.n5 A2.n3 27.752
R221 A2.n7 A2.n2 16.7975
R222 A2.n6 A2 11.5205
R223 A2 A2.n11 11.1548
R224 A2.n9 A2.n8 8.03383
R225 A2.n11 A2 6.4005
R226 A2.n6 A2 6.03479
R227 A2.n3 A2.n2 5.11262
R228 A2.n1 A2.n0 4.38232
R229 A2.n10 A2.n9 0.730803
R230 a_46_74.n4 a_46_74.t0 271.688
R231 a_46_74.n5 a_46_74.n4 186.882
R232 a_46_74.n1 a_46_74.n0 185
R233 a_46_74.n3 a_46_74.n2 185
R234 a_46_74.n1 a_46_74.t7 184.815
R235 a_46_74.n4 a_46_74.n3 66.6358
R236 a_46_74.n3 a_46_74.n1 53.4443
R237 a_46_74.n2 a_46_74.t2 22.7032
R238 a_46_74.n2 a_46_74.t5 22.7032
R239 a_46_74.n0 a_46_74.t6 22.7032
R240 a_46_74.n0 a_46_74.t4 22.7032
R241 a_46_74.t3 a_46_74.n5 22.7032
R242 a_46_74.n5 a_46_74.t1 22.7032
R243 B1_N.n1 B1_N.n0 273.517
R244 B1_N.n2 B1_N.t0 269.702
R245 B1_N.n1 B1_N.t1 219.31
R246 B1_N.n3 B1_N.n2 152
R247 B1_N.n2 B1_N.n1 15.3369
R248 B1_N B1_N.n3 13.3823
R249 B1_N.n3 B1_N 5.23686
C0 A2 VGND 0.052494f
C1 B1_N Y 0.001429f
C2 VPWR Y 0.026553f
C3 B1_N VGND 0.037986f
C4 VPWR VGND 0.122944f
C5 Y VGND 0.325608f
C6 VPB A1 0.138558f
C7 VPB A2 0.131924f
C8 A1 A2 0.072725f
C9 VPB B1_N 0.133615f
C10 VPB VPWR 0.216394f
C11 A1 VPWR 0.084421f
C12 VPB Y 0.009522f
C13 A1 Y 0.112156f
C14 A2 VPWR 0.062083f
C15 VPB VGND 0.013049f
C16 B1_N VPWR 0.057698f
C17 A1 VGND 0.030526f
C18 A2 Y 0.188099f
C19 VGND VNB 0.920581f
C20 Y VNB 0.062153f
C21 VPWR VNB 0.744944f
C22 B1_N VNB 0.223783f
C23 A2 VNB 0.398842f
C24 A1 VNB 0.443059f
C25 VPB VNB 1.79899f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a22o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a22o_2 VNB VPB VPWR VGND X B2 B1 A2 A1
X0 a_81_48.t2 A1.t0 a_304_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VGND.t3 B2.t0 a_491_74.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0925 ps=0.99 w=0.74 l=0.15
X2 VGND.t1 a_81_48.t4 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 X.t2 a_81_48.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 a_388_368.t3 B2.t1 a_81_48.t1 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.185 pd=1.37 as=0.175 ps=1.35 w=1 l=0.15
X5 a_304_74.t1 A2.t0 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1443 ps=1.13 w=0.74 l=0.15
X6 a_491_74.t0 B1.t0 a_81_48.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.0925 pd=0.99 as=0.1295 ps=1.09 w=0.74 l=0.15
X7 VPWR.t1 a_81_48.t6 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2109 pd=1.51 as=0.168 ps=1.42 w=1.12 l=0.15
X8 X.t0 a_81_48.t7 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X9 a_81_48.t0 B1.t1 a_388_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.35 as=0.15 ps=1.3 w=1 l=0.15
X10 a_388_368.t2 A1.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2109 ps=1.51 w=1 l=0.15
X11 VPWR.t2 A2.t1 a_388_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.185 ps=1.37 w=1 l=0.15
R0 A1.n0 A1.t1 231.629
R1 A1.n0 A1.t0 220.113
R2 A1 A1.n0 157.805
R3 a_304_74.t0 a_304_74.t1 529.841
R4 a_81_48.n5 a_81_48.n4 423.531
R5 a_81_48.n3 a_81_48.t6 272.574
R6 a_81_48.n1 a_81_48.t7 261.62
R7 a_81_48.n4 a_81_48.n0 253.29
R8 a_81_48.n1 a_81_48.t5 211.935
R9 a_81_48.n2 a_81_48.t4 154.24
R10 a_81_48.n4 a_81_48.n3 152
R11 a_81_48.n3 a_81_48.n2 49.6611
R12 a_81_48.n5 a_81_48.t1 39.4005
R13 a_81_48.n0 a_81_48.t2 34.0546
R14 a_81_48.t0 a_81_48.n5 29.5505
R15 a_81_48.n0 a_81_48.t3 22.7032
R16 a_81_48.n2 a_81_48.n1 5.11262
R17 VNB.t1 VNB.t3 2240.42
R18 VNB.t2 VNB.t5 1247.24
R19 VNB.t3 VNB.t4 1154.86
R20 VNB VNB.t0 1108.66
R21 VNB.t0 VNB.t1 993.177
R22 VNB.t4 VNB.t2 923.885
R23 B2.n0 B2.t1 231.629
R24 B2.n0 B2.t0 220.113
R25 B2 B2.n0 156.912
R26 a_491_74.t0 a_491_74.t1 40.541
R27 VGND.n3 VGND.t1 242.263
R28 VGND.n2 VGND.n1 217.356
R29 VGND.n5 VGND.t0 175.351
R30 VGND.n1 VGND.t2 34.0546
R31 VGND.n1 VGND.t3 29.1897
R32 VGND.n5 VGND.n4 27.8593
R33 VGND.n4 VGND.n3 24.0946
R34 VGND.n6 VGND.n5 9.3005
R35 VGND.n4 VGND.n0 9.3005
R36 VGND.n3 VGND.n2 7.39693
R37 VGND.n2 VGND.n0 0.166031
R38 VGND.n6 VGND.n0 0.122949
R39 VGND VGND.n6 0.0617245
R40 X X.n0 352.735
R41 X.n3 X.n2 185
R42 X.n2 X.n1 185
R43 X.n0 X.t1 26.3844
R44 X.n0 X.t0 26.3844
R45 X.n2 X.t3 22.7032
R46 X.n2 X.t2 22.7032
R47 X.n1 X 12.6066
R48 X X.n3 9.50353
R49 X.n3 X 4.84898
R50 X.n1 X 1.74595
R51 a_388_368.n1 a_388_368.n0 564.942
R52 a_388_368.n0 a_388_368.t1 41.3705
R53 a_388_368.n0 a_388_368.t3 31.5205
R54 a_388_368.t0 a_388_368.n1 29.5505
R55 a_388_368.n1 a_388_368.t2 29.5505
R56 VPB VPB.t2 446.909
R57 VPB.t3 VPB.t4 275.807
R58 VPB.t5 VPB.t1 265.591
R59 VPB.t0 VPB.t5 255.376
R60 VPB.t4 VPB.t0 229.839
R61 VPB.t2 VPB.t3 229.839
R62 A2.n0 A2.t1 223.758
R63 A2.n0 A2.t0 212.244
R64 A2 A2.n0 154.522
R65 B1.n0 B1.t1 231.629
R66 B1.n0 B1.t0 220.113
R67 B1 B1.n0 159.591
R68 VPWR.n1 VPWR.t2 433.245
R69 VPWR.n5 VPWR.t0 428.991
R70 VPWR.n3 VPWR.n2 319.616
R71 VPWR.n2 VPWR.t3 47.2805
R72 VPWR.n5 VPWR.n4 35.0123
R73 VPWR.n2 VPWR.t1 27.6909
R74 VPWR.n4 VPWR.n3 13.9299
R75 VPWR.n4 VPWR.n0 9.3005
R76 VPWR.n3 VPWR.n1 7.55201
R77 VPWR.n6 VPWR.n5 6.94346
R78 VPWR.n1 VPWR.n0 0.163292
R79 VPWR.n6 VPWR.n0 0.154086
R80 VPWR VPWR.n6 0.153633
C0 B1 B2 0.09404f
C1 X VGND 0.147767f
C2 A1 VGND 0.006514f
C3 B2 A2 0.095448f
C4 B1 VGND 0.006593f
C5 VPB VPWR 0.134447f
C6 B2 VGND 0.018262f
C7 VPB X 0.010002f
C8 A2 VGND 0.017139f
C9 VPB A1 0.036034f
C10 VPWR X 0.190534f
C11 VPWR A1 0.016327f
C12 VPB B1 0.033158f
C13 X A1 0.00118f
C14 VPB B2 0.034614f
C15 VPWR B1 0.005693f
C16 VPWR B2 0.006475f
C17 VPB A2 0.045492f
C18 X B1 2.46e-19
C19 VPB VGND 0.014659f
C20 VPWR A2 0.053079f
C21 A1 B1 0.095845f
C22 VPWR VGND 0.068474f
C23 VGND VNB 0.527618f
C24 A2 VNB 0.166072f
C25 B2 VNB 0.10281f
C26 B1 VNB 0.101212f
C27 A1 VNB 0.106847f
C28 X VNB 0.038628f
C29 VPWR VNB 0.454427f
C30 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a22o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a22o_1 VNB VPB VPWR VGND X B2 B1 A2 A1
X0 a_222_392.t2 B1.t0 a_230_79.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_52_123.t1 A1.t0 a_222_392.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 a_222_392.t0 B2.t0 a_132_392.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X3 a_132_392.t0 B1.t1 a_222_392.t1 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X4 X.t0 a_222_392.t4 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.3065 ps=1.7 w=1.12 l=0.15
X5 VGND.t0 A2.t0 a_52_123.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.12325 pd=1.185 as=0.1696 ps=1.81 w=0.64 l=0.15
X6 X.t1 a_222_392.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X7 VPWR.t2 A1.t1 a_132_392.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.3065 pd=1.7 as=0.195 ps=1.39 w=1 l=0.15
X8 a_132_392.t1 A2.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X9 a_230_79.t1 B2.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.12325 ps=1.185 w=0.64 l=0.15
R0 B1.n0 B1.t0 252.136
R1 B1.n0 B1.t1 231.629
R2 B1 B1.n0 153.904
R3 a_230_79.t0 a_230_79.t1 39.3755
R4 a_222_392.n3 a_222_392.n2 411.288
R5 a_222_392.n2 a_222_392.n0 264.043
R6 a_222_392.n1 a_222_392.t4 261.692
R7 a_222_392.n1 a_222_392.t5 204.113
R8 a_222_392.n2 a_222_392.n1 152
R9 a_222_392.n3 a_222_392.t1 35.4605
R10 a_222_392.t0 a_222_392.n3 29.5505
R11 a_222_392.n0 a_222_392.t3 26.2505
R12 a_222_392.n0 a_222_392.t2 26.2505
R13 VNB.t4 VNB.t1 2332.81
R14 VNB VNB.t2 1385.83
R15 VNB.t2 VNB.t3 1097.11
R16 VNB.t0 VNB.t4 993.177
R17 VNB.t3 VNB.t0 831.496
R18 A1.n0 A1.t1 263.762
R19 A1.n0 A1.t0 236.18
R20 A1 A1.n0 154.522
R21 a_52_123.t0 a_52_123.t1 606.547
R22 B2.n0 B2.t1 266.707
R23 B2.n0 B2.t0 231.629
R24 B2 B2.n0 168.097
R25 a_132_392.n1 a_132_392.n0 566.874
R26 a_132_392.t0 a_132_392.n1 40.3855
R27 a_132_392.n1 a_132_392.t2 36.4455
R28 a_132_392.n0 a_132_392.t3 29.5505
R29 a_132_392.n0 a_132_392.t1 29.5505
R30 VPB.t3 VPB.t1 372.849
R31 VPB VPB.t2 298.791
R32 VPB.t0 VPB.t3 275.807
R33 VPB.t4 VPB.t0 245.161
R34 VPB.t2 VPB.t4 229.839
R35 VPWR.n1 VPWR.n0 298.887
R36 VPWR.n1 VPWR.t1 267.3
R37 VPWR.n0 VPWR.t2 56.2686
R38 VPWR.n0 VPWR.t0 53.3913
R39 VPWR VPWR.n1 0.104606
R40 X.n3 X 589.85
R41 X.n3 X.n0 585
R42 X.n4 X.n3 585
R43 X.n2 X.t1 286.887
R44 X.t1 X.n1 286.887
R45 X.n3 X.t0 26.3844
R46 X X.n4 12.9944
R47 X.n1 X 12.6066
R48 X X.n0 11.249
R49 X X.n2 9.50353
R50 X.n2 X 4.84898
R51 X X.n0 3.10353
R52 X.n1 X 1.74595
R53 X.n4 X 1.35808
R54 A2.t0 A2.t1 460.31
R55 A2.n0 A2.t0 328.053
R56 A2 A2.n0 6.59444
R57 A2.n0 A2 4.3525
R58 VGND.n1 VGND.t1 248.752
R59 VGND.n1 VGND.n0 237.529
R60 VGND.n0 VGND.t2 34.8666
R61 VGND.n0 VGND.t0 33.438
R62 VGND VGND.n1 0.21682
C0 A2 VGND 0.099952f
C1 B1 VPWR 0.006237f
C2 A1 VPWR 0.017267f
C3 B2 VGND 0.016985f
C4 B1 X 1.97e-19
C5 A1 X 0.001166f
C6 B1 VGND 0.007845f
C7 VPWR X 0.093961f
C8 A1 VGND 0.008848f
C9 VPB A2 0.037429f
C10 VPWR VGND 0.056326f
C11 VPB B2 0.046185f
C12 X VGND 0.079755f
C13 VPB B1 0.042584f
C14 A2 B2 0.079314f
C15 VPB A1 0.049896f
C16 A2 A1 1.74e-19
C17 VPB VPWR 0.099892f
C18 B2 B1 0.102924f
C19 VPB X 0.016636f
C20 A2 VPWR 0.016026f
C21 B2 A1 2.95e-19
C22 A2 X 1.01e-19
C23 VPB VGND 0.00764f
C24 B1 A1 0.095545f
C25 B2 VPWR 0.034445f
C26 VGND VNB 0.446769f
C27 X VNB 0.112111f
C28 VPWR VNB 0.381293f
C29 A1 VNB 0.137415f
C30 B1 VNB 0.108688f
C31 B2 VNB 0.128304f
C32 A2 VNB 0.207562f
C33 VPB VNB 0.834768f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21oi_4 VNB VPB VPWR VGND Y B1 A2 A1
X0 a_69_368.t10 A1.t0 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t6 A1.t1 a_69_368.t9 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_69_368.t8 A1.t2 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 Y.t8 A1.t3 a_84_74.t7 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 VGND.t1 B1.t0 Y.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X5 VPWR.t4 A1.t4 a_69_368.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6 a_69_368.t3 A2.t0 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7 a_84_74.t6 A1.t5 Y.t7 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 Y.t4 B1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_84_74.t5 A1.t6 Y.t6 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X10 a_84_74.t0 A2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 VPWR.t1 A2.t2 a_69_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X12 a_84_74.t1 A2.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 a_69_368.t5 A2.t4 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR.t3 A2.t5 a_69_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X15 VGND.t4 A2.t6 a_84_74.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 VGND.t5 A2.t7 a_84_74.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X17 a_69_368.t11 B1.t2 Y.t9 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 a_69_368.t2 B1.t3 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X19 Y.t0 B1.t4 a_69_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 Y.t1 B1.t5 a_69_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X21 Y.t5 A1.t7 a_84_74.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 A1.n0 A1.t0 237.762
R1 A1.n7 A1.t1 226.809
R2 A1.n4 A1.t2 226.809
R3 A1.n2 A1.t4 226.809
R4 A1.n2 A1.t3 198.204
R5 A1.n0 A1.t5 196.013
R6 A1.n3 A1.t6 196.013
R7 A1.n6 A1.t7 196.013
R8 A1 A1.n0 159.591
R9 A1.n9 A1.n8 152
R10 A1.n5 A1.n1 152
R11 A1.n3 A1.n2 60.6157
R12 A1.n8 A1.n0 49.6611
R13 A1.n6 A1.n5 36.5157
R14 A1.n5 A1.n4 21.1793
R15 A1.n9 A1.n1 10.1214
R16 A1.n7 A1.n6 8.03383
R17 A1.n8 A1.n7 5.11262
R18 A1.n4 A1.n3 5.11262
R19 A1 A1.n9 2.53073
R20 A1.n1 A1 1.63771
R21 VPWR.n5 VPWR.n4 625.544
R22 VPWR.n7 VPWR.n6 611.88
R23 VPWR.n3 VPWR.n2 331.5
R24 VPWR.n13 VPWR.n1 323.406
R25 VPWR.n12 VPWR.n11 36.1417
R26 VPWR.n8 VPWR.n7 29.7417
R27 VPWR.n1 VPWR.t2 26.3844
R28 VPWR.n1 VPWR.t3 26.3844
R29 VPWR.n2 VPWR.t0 26.3844
R30 VPWR.n2 VPWR.t1 26.3844
R31 VPWR.n6 VPWR.t5 26.3844
R32 VPWR.n6 VPWR.t4 26.3844
R33 VPWR.n4 VPWR.t7 26.3844
R34 VPWR.n4 VPWR.t6 26.3844
R35 VPWR.n8 VPWR.n3 25.6005
R36 VPWR.n13 VPWR.n12 14.6829
R37 VPWR.n11 VPWR.n3 10.5417
R38 VPWR.n14 VPWR.n13 10.3391
R39 VPWR.n9 VPWR.n8 9.3005
R40 VPWR.n11 VPWR.n10 9.3005
R41 VPWR.n12 VPWR.n0 9.3005
R42 VPWR.n7 VPWR.n5 6.85408
R43 VPWR.n9 VPWR.n5 0.451374
R44 VPWR VPWR.n14 0.163644
R45 VPWR.n14 VPWR.n0 0.144205
R46 VPWR.n10 VPWR.n9 0.122949
R47 VPWR.n10 VPWR.n0 0.122949
R48 a_69_368.n7 a_69_368.n6 305.901
R49 a_69_368.n7 a_69_368.t2 303.128
R50 a_69_368.n5 a_69_368.n4 299.053
R51 a_69_368.n9 a_69_368.n8 287.964
R52 a_69_368.n1 a_69_368.t6 280.985
R53 a_69_368.n1 a_69_368.n0 205.487
R54 a_69_368.n3 a_69_368.n2 196.025
R55 a_69_368.n8 a_69_368.n7 79.3988
R56 a_69_368.n8 a_69_368.n5 56.0877
R57 a_69_368.n3 a_69_368.n1 55.6691
R58 a_69_368.n5 a_69_368.n3 53.4028
R59 a_69_368.n2 a_69_368.t7 26.3844
R60 a_69_368.n2 a_69_368.t3 26.3844
R61 a_69_368.n0 a_69_368.t4 26.3844
R62 a_69_368.n0 a_69_368.t5 26.3844
R63 a_69_368.n4 a_69_368.t9 26.3844
R64 a_69_368.n4 a_69_368.t8 26.3844
R65 a_69_368.n6 a_69_368.t1 26.3844
R66 a_69_368.n6 a_69_368.t11 26.3844
R67 a_69_368.n9 a_69_368.t0 26.3844
R68 a_69_368.t10 a_69_368.n9 26.3844
R69 VPB VPB.t6 354.974
R70 VPB.t1 VPB.t2 229.839
R71 VPB.t11 VPB.t1 229.839
R72 VPB.t0 VPB.t11 229.839
R73 VPB.t10 VPB.t0 229.839
R74 VPB.t9 VPB.t10 229.839
R75 VPB.t8 VPB.t9 229.839
R76 VPB.t7 VPB.t8 229.839
R77 VPB.t3 VPB.t7 229.839
R78 VPB.t4 VPB.t3 229.839
R79 VPB.t5 VPB.t4 229.839
R80 VPB.t6 VPB.t5 229.839
R81 a_84_74.n1 a_84_74.t6 325.339
R82 a_84_74.n3 a_84_74.t3 213.992
R83 a_84_74.n1 a_84_74.n0 185
R84 a_84_74.n3 a_84_74.n2 103.65
R85 a_84_74.n5 a_84_74.n4 84.741
R86 a_84_74.n4 a_84_74.n3 83.6621
R87 a_84_74.n4 a_84_74.n1 79.2686
R88 a_84_74.n2 a_84_74.t2 22.7032
R89 a_84_74.n2 a_84_74.t1 22.7032
R90 a_84_74.n0 a_84_74.t4 22.7032
R91 a_84_74.n0 a_84_74.t5 22.7032
R92 a_84_74.n5 a_84_74.t7 22.7032
R93 a_84_74.t0 a_84_74.n5 22.7032
R94 Y.n2 Y.n0 342.868
R95 Y.n2 Y.n1 299.952
R96 Y.n3 Y.t4 212.042
R97 Y.n7 Y.n6 187.022
R98 Y.n5 Y.n4 185
R99 Y.n3 Y.t2 147.544
R100 Y Y.n2 145.792
R101 Y.n5 Y.n3 42.2654
R102 Y.n7 Y.n5 38.6138
R103 Y.n0 Y.t3 26.3844
R104 Y.n0 Y.t1 26.3844
R105 Y.n1 Y.t9 26.3844
R106 Y.n1 Y.t0 26.3844
R107 Y.n6 Y.t6 22.7032
R108 Y.n6 Y.t8 22.7032
R109 Y.n4 Y.t7 22.7032
R110 Y.n4 Y.t5 22.7032
R111 Y.n7 Y 4.26717
R112 Y Y.n8 3.62717
R113 Y.n8 Y 1.67007
R114 Y.n8 Y.n7 0.427167
R115 VNB.t8 VNB.t0 2332.81
R116 VNB VNB.t5 1755.38
R117 VNB.t0 VNB.t1 993.177
R118 VNB.t6 VNB.t8 993.177
R119 VNB.t7 VNB.t6 993.177
R120 VNB.t9 VNB.t7 993.177
R121 VNB.t2 VNB.t9 993.177
R122 VNB.t4 VNB.t2 993.177
R123 VNB.t3 VNB.t4 993.177
R124 VNB.t5 VNB.t3 993.177
R125 B1.n0 B1.t3 344.606
R126 B1.n5 B1.t4 242.023
R127 B1.n1 B1.t5 226.809
R128 B1.n4 B1.t2 226.809
R129 B1.n3 B1.t0 196.013
R130 B1.n0 B1.t1 196.013
R131 B1 B1.n2 155.721
R132 B1.n5 B1 154.233
R133 B1.n7 B1.n6 152
R134 B1.n6 B1.n5 49.6611
R135 B1.n3 B1.n2 43.8187
R136 B1.n2 B1.n1 16.7975
R137 B1.n7 B1 7.88887
R138 B1 B1.n7 6.4005
R139 B1.n4 B1.n3 5.11262
R140 B1.n1 B1.n0 2.19141
R141 B1.n6 B1.n4 0.730803
R142 VGND.n3 VGND.n2 214.655
R143 VGND.n5 VGND.n4 208.079
R144 VGND.n1 VGND.n0 208.079
R145 VGND.n6 VGND.n5 35.3887
R146 VGND.n2 VGND.t0 22.7032
R147 VGND.n2 VGND.t1 22.7032
R148 VGND.n4 VGND.t2 22.7032
R149 VGND.n4 VGND.t4 22.7032
R150 VGND.n0 VGND.t3 22.7032
R151 VGND.n0 VGND.t5 22.7032
R152 VGND.n8 VGND.n1 14.4803
R153 VGND.n7 VGND.n6 9.3005
R154 VGND.n5 VGND.n3 6.28589
R155 VGND.n6 VGND.n1 4.51815
R156 VGND.n7 VGND.n3 0.171081
R157 VGND VGND.n8 0.163644
R158 VGND.n8 VGND.n7 0.144205
R159 A2.n4 A2.t5 236.303
R160 A2.n1 A2.t0 226.809
R161 A2.n8 A2.t2 226.809
R162 A2.n3 A2.t4 226.809
R163 A2.n1 A2.t1 196.744
R164 A2.n4 A2.t7 196.013
R165 A2.n2 A2.t3 196.013
R166 A2.n9 A2.t6 196.013
R167 A2 A2.n5 156.912
R168 A2.n12 A2.n11 152
R169 A2.n10 A2.n0 152
R170 A2.n7 A2.n6 152
R171 A2.n11 A2.n10 49.6611
R172 A2.n8 A2.n7 44.549
R173 A2.n5 A2.n3 28.4823
R174 A2.n5 A2.n4 27.752
R175 A2.n7 A2.n2 14.6066
R176 A2.n11 A2.n1 10.955
R177 A2.n12 A2.n0 10.1214
R178 A2.n6 A2 9.07957
R179 A2.n3 A2.n2 6.57323
R180 A2.n6 A2 5.2098
R181 A2.n9 A2.n8 3.65202
R182 A2 A2.n12 3.12608
R183 A2.n10 A2.n9 1.46111
R184 A2 A2.n0 1.04236
C0 VPB A1 0.131161f
C1 A2 A1 0.061082f
C2 VPB B1 0.136443f
C3 VPB VPWR 0.157432f
C4 VPB Y 0.009275f
C5 A1 B1 0.065186f
C6 A2 VPWR 0.060375f
C7 VPB VGND 0.011179f
C8 A1 VPWR 0.05371f
C9 A2 Y 0.031349f
C10 A1 Y 0.307184f
C11 A2 VGND 0.063804f
C12 B1 VPWR 0.022536f
C13 A1 VGND 0.023104f
C14 B1 Y 0.266671f
C15 B1 VGND 0.041353f
C16 VPWR Y 0.04237f
C17 VPWR VGND 0.100446f
C18 Y VGND 0.208223f
C19 VPB A2 0.139515f
C20 VGND VNB 0.760639f
C21 Y VNB 0.089914f
C22 VPWR VNB 0.597005f
C23 B1 VNB 0.357612f
C24 A1 VNB 0.39542f
C25 A2 VNB 0.434889f
C26 VPB VNB 1.47758f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21oi_2 VNB VPB VPWR VGND Y B1 A2 A1
X0 a_131_368.t4 A1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X1 VPWR.t0 A2.t0 a_131_368.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.168 ps=1.42 w=1.12 l=0.15
X2 a_131_368.t1 B1.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3 VPWR.t1 A1.t1 a_131_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_131_368.t5 A2.t1 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2016 ps=1.48 w=1.12 l=0.15
X5 Y.t0 B1.t1 a_131_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X6 Y.t2 B1.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X7 Y.t4 A1.t2 a_280_107.t3 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_280_107.t2 A1.t3 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_280_107.t1 A2.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.19365 ps=1.405 w=0.74 l=0.15
X10 VGND.t1 A2.t3 a_280_107.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.19365 pd=1.405 as=0.25175 ps=2.22 w=0.74 l=0.15
R0 A1.n1 A1.t1 229
R1 A1.n0 A1.t0 227.538
R2 A1.n1 A1.t2 196.013
R3 A1.n0 A1.t3 196.013
R4 A1 A1.n2 156.465
R5 A1.n2 A1.n1 44.549
R6 A1.n2 A1.n0 18.2581
R7 VPWR.n2 VPWR.n1 626.035
R8 VPWR.n2 VPWR.n0 616.499
R9 VPWR.n0 VPWR.t3 36.0585
R10 VPWR.n0 VPWR.t0 27.2639
R11 VPWR.n1 VPWR.t2 26.3844
R12 VPWR.n1 VPWR.t1 26.3844
R13 VPWR VPWR.n2 0.87081
R14 a_131_368.t4 a_131_368.n3 368.354
R15 a_131_368.n1 a_131_368.t0 304.615
R16 a_131_368.n3 a_131_368.n2 299.053
R17 a_131_368.n1 a_131_368.n0 288.443
R18 a_131_368.n3 a_131_368.n1 59.2079
R19 a_131_368.n0 a_131_368.t2 26.3844
R20 a_131_368.n0 a_131_368.t1 26.3844
R21 a_131_368.n2 a_131_368.t3 26.3844
R22 a_131_368.n2 a_131_368.t5 26.3844
R23 VPB VPB.t0 513.307
R24 VPB.t2 VPB.t5 260.485
R25 VPB.t3 VPB.t4 229.839
R26 VPB.t5 VPB.t3 229.839
R27 VPB.t1 VPB.t2 229.839
R28 VPB.t0 VPB.t1 229.839
R29 A2.n0 A2.t1 226.809
R30 A2.n1 A2.t0 226.809
R31 A2.n0 A2.t2 201.125
R32 A2.n1 A2.t3 160.513
R33 A2.n3 A2.n2 152
R34 A2.n2 A2.n1 72.3005
R35 A2.n3 A2 6.93383
R36 A2 A2.n3 3.30717
R37 A2.n2 A2.n0 2.19141
R38 B1.n0 B1.t0 348.647
R39 B1.n1 B1.t2 223.327
R40 B1.n0 B1.t1 204.048
R41 B1 B1.n1 186.94
R42 B1.n1 B1.n0 155.555
R43 Y.n3 Y.n2 349.733
R44 Y.n1 Y.n0 214.007
R45 Y.n3 Y.t2 145.738
R46 Y Y.n3 34.0108
R47 Y.n0 Y.t1 26.3844
R48 Y.n0 Y.t0 26.3844
R49 Y.n2 Y.t3 22.7032
R50 Y.n2 Y.t4 22.7032
R51 Y Y.n1 15.6759
R52 Y.n1 Y 3.29747
R53 VGND.n1 VGND.n0 223.959
R54 VGND.n1 VGND.t2 174.686
R55 VGND.n0 VGND.t1 61.3164
R56 VGND.n0 VGND.t0 24.3603
R57 VGND VGND.n1 0.109886
R58 VNB.t2 VNB.t0 3048.82
R59 VNB.t0 VNB.t1 1501.31
R60 VNB VNB.t2 1108.66
R61 VNB.t4 VNB.t3 993.177
R62 VNB.t1 VNB.t4 993.177
R63 a_280_107.n0 a_280_107.t0 554.524
R64 a_280_107.n1 a_280_107.n0 231.381
R65 a_280_107.n0 a_280_107.t2 139.209
R66 a_280_107.n1 a_280_107.t3 22.7032
R67 a_280_107.t1 a_280_107.n1 22.7032
C0 VPB Y 0.00484f
C1 VPB VPWR 0.10856f
C2 A2 A1 0.101599f
C3 B1 Y 0.093964f
C4 VPB VGND 0.010914f
C5 A2 Y 0.071205f
C6 B1 VPWR 0.018861f
C7 A1 Y 0.029501f
C8 B1 VGND 0.046579f
C9 A2 VPWR 0.030822f
C10 A2 VGND 0.028668f
C11 A1 VPWR 0.025659f
C12 Y VPWR 0.014598f
C13 A1 VGND 0.013222f
C14 Y VGND 0.202842f
C15 VPWR VGND 0.063213f
C16 VPB B1 0.115545f
C17 VPB A2 0.071388f
C18 B1 A2 0.027042f
C19 VPB A1 0.063136f
C20 VGND VNB 0.533118f
C21 VPWR VNB 0.386446f
C22 Y VNB 0.068807f
C23 A1 VNB 0.217199f
C24 A2 VNB 0.229489f
C25 B1 VNB 0.259624f
C26 VPB VNB 0.941904f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a21oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21oi_1 VNB VPB VPWR VGND B1 Y A2 A1
X0 Y.t0 A1.t0 a_117_74.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X1 VGND.t1 B1.t0 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1443 ps=1.13 w=0.74 l=0.15
X2 a_117_74.t0 A2.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1961 ps=2.01 w=0.74 l=0.15
X3 Y.t2 B1.t1 a_29_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X4 a_29_368.t2 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1848 ps=1.45 w=1.12 l=0.15
X5 VPWR.t0 A2.t1 a_29_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.308 ps=2.79 w=1.12 l=0.15
R0 A1.n0 A1.t1 250.909
R1 A1.n0 A1.t0 220.113
R2 A1 A1.n0 161.674
R3 a_117_74.t0 a_117_74.t1 34.0546
R4 Y.n2 Y 591.4
R5 Y.n2 Y.n0 585
R6 Y.n3 Y.n2 585
R7 Y Y.n1 180.512
R8 Y.n1 Y.t1 37.2978
R9 Y.n2 Y.t2 26.3844
R10 Y.n1 Y.t0 25.9464
R11 Y Y.n3 17.1525
R12 Y Y.n0 14.8485
R13 Y Y.n0 4.0965
R14 Y.n3 Y 1.7925
R15 VNB.t1 VNB.t2 1247.24
R16 VNB VNB.t0 1177.95
R17 VNB.t0 VNB.t1 831.496
R18 B1.n0 B1.t1 278.188
R19 B1.n0 B1.t0 170.81
R20 B1 B1.n0 160.785
R21 VGND.n0 VGND.t0 165.871
R22 VGND.n0 VGND.t1 159.133
R23 VGND VGND.n0 0.184018
R24 A2.n0 A2.t1 278.188
R25 A2.n0 A2.t0 170.81
R26 A2 A2.n0 158.788
R27 a_29_368.t0 a_29_368.n0 567.265
R28 a_29_368.n0 a_29_368.t1 26.3844
R29 a_29_368.n0 a_29_368.t2 26.3844
R30 VPB VPB.t0 252.823
R31 VPB.t0 VPB.t2 245.161
R32 VPB.t2 VPB.t1 229.839
R33 VPWR VPWR.n0 321.096
R34 VPWR.n0 VPWR.t1 29.0228
R35 VPWR.n0 VPWR.t0 29.0228
C0 A1 VPB 0.033291f
C1 B1 VPB 0.038383f
C2 A2 VPB 0.039467f
C3 A1 B1 0.056293f
C4 A2 A1 0.091984f
C5 VPWR VPB 0.054807f
C6 A1 VPWR 0.020251f
C7 Y VPB 0.015287f
C8 B1 VPWR 0.011419f
C9 A1 Y 0.064526f
C10 A2 VPWR 0.01841f
C11 VGND VPB 0.004976f
C12 A1 VGND 0.021272f
C13 B1 Y 0.093655f
C14 A2 Y 0.009899f
C15 B1 VGND 0.039989f
C16 VPWR Y 0.035724f
C17 A2 VGND 0.051917f
C18 VPWR VGND 0.032164f
C19 Y VGND 0.121769f
C20 VGND VNB 0.344532f
C21 Y VNB 0.076144f
C22 VPWR VNB 0.224633f
C23 B1 VNB 0.166709f
C24 A1 VNB 0.109919f
C25 A2 VNB 0.165389f
C26 VPB VNB 0.51336f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a22o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a22o_4 VNB VPB VPWR VGND X B2 B1 A2 A1
X0 a_645_120.t3 B1.t0 a_95_306.t5 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1053 pd=0.98 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 X.t3 a_95_306.t8 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X2 a_95_306.t0 A1.t0 a_1064_123.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X3 X.t7 a_95_306.t9 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4 a_555_392.t3 B2.t0 a_95_306.t6 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X5 a_95_306.t3 B1.t1 a_555_392.t2 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X6 VPWR.t0 A2.t0 a_555_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2575 pd=1.515 as=0.165 ps=1.33 w=1 l=0.15
X7 VGND.t6 A2.t1 a_1064_123.t0 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X8 VGND.t2 a_95_306.t10 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.12685 pd=1.095 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 a_1064_123.t2 A1.t1 a_95_306.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X10 a_555_392.t1 B1.t2 a_95_306.t2 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X11 a_95_306.t7 B2.t1 a_555_392.t4 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X12 VPWR.t3 a_95_306.t11 X.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X13 X.t1 a_95_306.t12 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 X.t5 a_95_306.t13 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X15 VPWR.t1 a_95_306.t14 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X16 a_645_120.t0 B2.t2 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.12685 ps=1.095 w=0.64 l=0.15
X17 VPWR.t5 A1.t2 a_555_392.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND.t5 B2.t3 a_645_120.t1 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1952 pd=1.25 as=0.1053 ps=0.98 w=0.64 l=0.15
X19 VGND.t0 a_95_306.t15 X.t4 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X20 a_1064_123.t1 A2.t2 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1952 ps=1.25 w=0.64 l=0.15
X21 a_95_306.t4 B1.t3 a_645_120.t2 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 B1.n0 B1.t1 219.091
R1 B1.n1 B1.t2 217.631
R2 B1.n1 B1.t3 165.488
R3 B1.n0 B1.t0 165.488
R4 B1 B1.n2 157.625
R5 B1.n2 B1.n0 51.1217
R6 B1.n2 B1.n1 11.6853
R7 a_95_306.n13 a_95_306.n1 619.49
R8 a_95_306.n14 a_95_306.n13 585
R9 a_95_306.n5 a_95_306.t8 352.111
R10 a_95_306.n4 a_95_306.n2 333.988
R11 a_95_306.n7 a_95_306.t12 226.809
R12 a_95_306.n9 a_95_306.t11 226.809
R13 a_95_306.n6 a_95_306.t13 212.081
R14 a_95_306.n5 a_95_306.t14 204.048
R15 a_95_306.n4 a_95_306.n3 185
R16 a_95_306.n0 a_95_306.n10 168.874
R17 a_95_306.n12 a_95_306.t10 167.386
R18 a_95_306.n8 a_95_306.t15 154.24
R19 a_95_306.n11 a_95_306.t9 154.24
R20 a_95_306.n0 a_95_306.n12 152
R21 a_95_306.n13 a_95_306.n0 144.383
R22 a_95_306.n6 a_95_306.n5 98.7934
R23 a_95_306.n8 a_95_306.n7 89.6817
R24 a_95_306.n0 a_95_306.n4 87.4627
R25 a_95_306.n12 a_95_306.n11 49.6611
R26 a_95_306.n7 a_95_306.n6 35.3472
R27 a_95_306.n10 a_95_306.n9 29.9429
R28 a_95_306.n1 a_95_306.t6 29.5505
R29 a_95_306.n1 a_95_306.t3 29.5505
R30 a_95_306.t2 a_95_306.n14 29.5505
R31 a_95_306.n14 a_95_306.t7 29.5505
R32 a_95_306.n3 a_95_306.t5 26.2505
R33 a_95_306.n3 a_95_306.t4 26.2505
R34 a_95_306.n2 a_95_306.t1 26.2505
R35 a_95_306.n2 a_95_306.t0 26.2505
R36 a_95_306.n9 a_95_306.n8 18.9884
R37 a_95_306.n11 a_95_306.n10 13.8763
R38 a_645_120.n1 a_645_120.n0 415.057
R39 a_645_120.n0 a_645_120.t1 28.3002
R40 a_645_120.n0 a_645_120.t3 27.3402
R41 a_645_120.t2 a_645_120.n1 26.2505
R42 a_645_120.n1 a_645_120.t0 26.2505
R43 VNB VNB.t3 3129.66
R44 VNB.t7 VNB.t11 1755.38
R45 VNB.t4 VNB.t6 1166.4
R46 VNB.t9 VNB.t7 1097.11
R47 VNB.t1 VNB.t10 993.177
R48 VNB.t0 VNB.t1 993.177
R49 VNB.t11 VNB.t0 993.177
R50 VNB.t8 VNB.t9 993.177
R51 VNB.t6 VNB.t8 993.177
R52 VNB.t5 VNB.t4 993.177
R53 VNB.t2 VNB.t5 993.177
R54 VNB.t3 VNB.t2 993.177
R55 A1.n2 A1.n1 220.917
R56 A1.n0 A1.t2 212.883
R57 A1.n0 A1.t1 170.6
R58 A1.n2 A1.t0 165.488
R59 A1.n4 A1.n3 152
R60 A1.n3 A1.n0 54.7732
R61 A1.n4 A1 10.0853
R62 A1 A1.n4 8.53383
R63 A1.n3 A1.n2 2.92171
R64 VPWR.n7 VPWR.t0 356.594
R65 VPWR.n6 VPWR.t5 352.173
R66 VPWR.n3 VPWR.t3 258.772
R67 VPWR.n21 VPWR.t4 250.081
R68 VPWR.n19 VPWR.n2 232.787
R69 VPWR.n8 VPWR.n5 36.1417
R70 VPWR.n12 VPWR.n5 36.1417
R71 VPWR.n13 VPWR.n12 36.1417
R72 VPWR.n14 VPWR.n13 36.1417
R73 VPWR.n8 VPWR.n7 35.7652
R74 VPWR.n18 VPWR.n3 28.2358
R75 VPWR.n20 VPWR.n19 26.7299
R76 VPWR.n19 VPWR.n18 26.7299
R77 VPWR.n2 VPWR.t2 26.3844
R78 VPWR.n2 VPWR.t1 26.3844
R79 VPWR.n14 VPWR.n3 25.224
R80 VPWR.n21 VPWR.n20 16.1887
R81 VPWR.n9 VPWR.n8 9.3005
R82 VPWR.n10 VPWR.n5 9.3005
R83 VPWR.n12 VPWR.n11 9.3005
R84 VPWR.n13 VPWR.n4 9.3005
R85 VPWR.n15 VPWR.n14 9.3005
R86 VPWR.n16 VPWR.n3 9.3005
R87 VPWR.n18 VPWR.n17 9.3005
R88 VPWR.n19 VPWR.n1 9.3005
R89 VPWR.n20 VPWR.n0 9.3005
R90 VPWR.n22 VPWR.n21 9.3005
R91 VPWR.n7 VPWR.n6 4.08171
R92 VPWR.n9 VPWR.n6 0.48579
R93 VPWR.n10 VPWR.n9 0.122949
R94 VPWR.n11 VPWR.n10 0.122949
R95 VPWR.n11 VPWR.n4 0.122949
R96 VPWR.n15 VPWR.n4 0.122949
R97 VPWR.n16 VPWR.n15 0.122949
R98 VPWR.n17 VPWR.n16 0.122949
R99 VPWR.n17 VPWR.n1 0.122949
R100 VPWR.n1 VPWR.n0 0.122949
R101 VPWR.n22 VPWR.n0 0.122949
R102 VPWR VPWR.n22 0.0617245
R103 a_555_392.n3 a_555_392.n2 585
R104 a_555_392.n2 a_555_392.t4 395.348
R105 a_555_392.n1 a_555_392.t5 313.259
R106 a_555_392.n1 a_555_392.n0 194.833
R107 a_555_392.n2 a_555_392.n1 66.4813
R108 a_555_392.n0 a_555_392.t0 35.4605
R109 a_555_392.n0 a_555_392.t3 29.5505
R110 a_555_392.t2 a_555_392.n3 29.5505
R111 a_555_392.n3 a_555_392.t1 29.5505
R112 VPB.t3 VPB.t8 618.011
R113 VPB.t0 VPB.t9 569.49
R114 VPB VPB.t4 288.575
R115 VPB.t7 VPB.t0 245.161
R116 VPB.t6 VPB.t7 229.839
R117 VPB.t5 VPB.t6 229.839
R118 VPB.t8 VPB.t5 229.839
R119 VPB.t2 VPB.t3 229.839
R120 VPB.t1 VPB.t2 229.839
R121 VPB.t4 VPB.t1 229.839
R122 X.n6 X.n0 236.762
R123 X.n5 X.n1 223.968
R124 X.n4 X.n2 131.974
R125 X.n4 X.n3 97.4922
R126 X.n1 X.t2 26.3844
R127 X.n1 X.t1 26.3844
R128 X.n0 X.t0 26.3844
R129 X.n0 X.t3 26.3844
R130 X.n2 X.t6 22.7032
R131 X.n2 X.t7 22.7032
R132 X.n3 X.t4 22.7032
R133 X.n3 X.t5 22.7032
R134 X.n6 X.n5 15.4358
R135 X.n5 X.n4 8.53383
R136 X X.n7 3.31902
R137 X.n7 X.n6 2.13383
R138 X.n7 X 1.75736
R139 a_1064_123.n1 a_1064_123.n0 346.986
R140 a_1064_123.n0 a_1064_123.t3 26.2505
R141 a_1064_123.n0 a_1064_123.t1 26.2505
R142 a_1064_123.n1 a_1064_123.t0 26.2505
R143 a_1064_123.t2 a_1064_123.n1 26.2505
R144 VGND.n19 VGND.t1 248.919
R145 VGND.n4 VGND.n3 223.912
R146 VGND.n17 VGND.n16 218.792
R147 VGND.n10 VGND.n9 214.091
R148 VGND.n5 VGND.t6 172.368
R149 VGND.n3 VGND.t7 88.1255
R150 VGND.n9 VGND.t4 40.313
R151 VGND.n8 VGND.n7 36.1417
R152 VGND.n11 VGND.n8 36.1417
R153 VGND.n15 VGND.n1 36.1417
R154 VGND.n7 VGND.n4 34.2593
R155 VGND.n19 VGND.n18 34.2593
R156 VGND.n3 VGND.t5 26.2505
R157 VGND.n16 VGND.t3 22.7032
R158 VGND.n16 VGND.t0 22.7032
R159 VGND.n9 VGND.t2 22.1988
R160 VGND.n18 VGND.n17 11.6711
R161 VGND.n18 VGND.n0 9.3005
R162 VGND.n15 VGND.n14 9.3005
R163 VGND.n13 VGND.n1 9.3005
R164 VGND.n12 VGND.n11 9.3005
R165 VGND.n8 VGND.n2 9.3005
R166 VGND.n7 VGND.n6 9.3005
R167 VGND.n11 VGND.n10 7.15344
R168 VGND.n20 VGND.n19 6.88467
R169 VGND.n5 VGND.n4 6.87459
R170 VGND.n17 VGND.n15 5.64756
R171 VGND.n10 VGND.n1 4.14168
R172 VGND VGND.n20 0.270511
R173 VGND.n6 VGND.n5 0.167141
R174 VGND.n20 VGND.n0 0.160218
R175 VGND.n6 VGND.n2 0.122949
R176 VGND.n12 VGND.n2 0.122949
R177 VGND.n13 VGND.n12 0.122949
R178 VGND.n14 VGND.n13 0.122949
R179 VGND.n14 VGND.n0 0.122949
R180 B2.n1 B2.t1 241
R181 B2.n0 B2.t0 239.661
R182 B2.n1 B2.t2 189.588
R183 B2 B2.n1 188.213
R184 B2.n0 B2.t3 186.374
R185 B2 B2.n0 186.01
R186 A2.n1 A2.t1 622.948
R187 A2.t2 A2.t0 504.493
R188 A2.t1 A2.n0 460.31
R189 A2.n1 A2.t2 162.274
R190 A2.n2 A2.n1 157.888
R191 A2 A2.n2 6.59444
R192 A2.n2 A2 4.3525
C0 VPB A1 0.080045f
C1 B2 A2 0.056739f
C2 B2 A1 0.009748f
C3 VPB VPWR 0.21249f
C4 B1 A2 2.93e-19
C5 B1 A1 5.95e-21
C6 VPB X 0.015569f
C7 B2 VPWR 0.018255f
C8 A2 A1 0.133061f
C9 B2 X 5.92e-19
C10 B1 VPWR 0.009124f
C11 VPB VGND 0.017715f
C12 B2 VGND 0.025563f
C13 A2 VPWR 0.035665f
C14 B1 X 1.45e-20
C15 A1 VPWR 0.03404f
C16 A2 X 1.7e-21
C17 B1 VGND 0.010335f
C18 A2 VGND 0.152568f
C19 A1 X 2.28e-21
C20 A1 VGND 0.010417f
C21 VPWR X 0.460585f
C22 VPB B2 0.100007f
C23 VPWR VGND 0.118883f
C24 VPB B1 0.070183f
C25 X VGND 0.275806f
C26 VPB A2 0.082422f
C27 B2 B1 0.231798f
C28 VGND VNB 0.981682f
C29 X VNB 0.083031f
C30 VPWR VNB 0.716725f
C31 A1 VNB 0.17043f
C32 A2 VNB 0.431126f
C33 B1 VNB 0.172523f
C34 B2 VNB 0.197999f
C35 VPB VNB 1.69186f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a22oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a22oi_1 VNB VPB VPWR VGND B2 Y B1 A2 A1
X0 Y.t2 B1.t0 a_159_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X1 a_159_74.t1 B2.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1961 ps=2.01 w=0.74 l=0.15
X2 a_339_74.t1 A1.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1443 ps=1.13 w=0.74 l=0.15
X3 VGND.t0 A2.t0 a_339_74.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1443 ps=1.13 w=0.74 l=0.15
X4 VPWR.t0 A1.t1 a_71_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.2184 pd=1.51 as=0.1848 ps=1.45 w=1.12 l=0.15
X5 a_71_368.t1 B1.t1 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t3 B2.t1 a_71_368.t3 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X7 a_71_368.t2 A2.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.2184 ps=1.51 w=1.12 l=0.15
R0 B1.n0 B1.t1 250.909
R1 B1.n0 B1.t0 220.113
R2 B1 B1.n0 154.522
R3 a_159_74.t0 a_159_74.t1 34.0546
R4 Y Y.n0 333.207
R5 Y Y.n1 128.055
R6 Y.n1 Y.t0 31.6221
R7 Y.n1 Y.t2 31.6221
R8 Y.n0 Y.t1 26.3844
R9 Y.n0 Y.t3 26.3844
R10 VNB VNB.t3 1662.99
R11 VNB.t0 VNB.t1 1247.24
R12 VNB.t2 VNB.t0 1247.24
R13 VNB.t3 VNB.t2 831.496
R14 B2.n0 B2.t1 261.62
R15 B2.n1 B2.n0 215.536
R16 B2.n0 B2.t0 156.431
R17 B2 B2.n1 7.56414
R18 B2.n1 B2 6.78838
R19 VGND.n0 VGND.t1 240.635
R20 VGND.n0 VGND.t0 174.841
R21 VGND VGND.n0 0.167461
R22 A1.n0 A1.t1 250.909
R23 A1.n0 A1.t0 220.113
R24 A1 A1.n0 155.423
R25 a_339_74.t0 a_339_74.t1 63.2437
R26 A2.n0 A2.t1 250.909
R27 A2.n0 A2.t0 220.113
R28 A2.n1 A2.n0 152
R29 A2 A2.n1 9.07957
R30 A2.n1 A2 5.2098
R31 a_71_368.n0 a_71_368.t3 392.096
R32 a_71_368.n0 a_71_368.t2 300.195
R33 a_71_368.n1 a_71_368.n0 189.115
R34 a_71_368.t0 a_71_368.n1 31.6612
R35 a_71_368.n1 a_71_368.t1 26.3844
R36 VPWR VPWR.n0 321.101
R37 VPWR.n0 VPWR.t1 36.938
R38 VPWR.n0 VPWR.t0 31.6612
R39 VPB VPB.t3 360.082
R40 VPB.t0 VPB.t2 275.807
R41 VPB.t1 VPB.t0 245.161
R42 VPB.t3 VPB.t1 229.839
C0 VPB A1 0.033119f
C1 B2 B1 0.069458f
C2 VPB A2 0.044356f
C3 VPB Y 0.008552f
C4 B1 A1 0.086353f
C5 VPB VPWR 0.079242f
C6 B2 Y 0.087548f
C7 B1 Y 0.08992f
C8 A1 A2 0.088678f
C9 VPB VGND 0.009467f
C10 B2 VPWR 0.009807f
C11 A1 Y 0.012667f
C12 B2 VGND 0.030067f
C13 B1 VPWR 0.005972f
C14 B1 VGND 0.012396f
C15 A1 VPWR 0.017502f
C16 A2 Y 0.003428f
C17 A1 VGND 0.0169f
C18 A2 VPWR 0.018508f
C19 A2 VGND 0.0514f
C20 Y VPWR 0.009782f
C21 VPB B2 0.05525f
C22 Y VGND 0.116181f
C23 VPB B1 0.031827f
C24 VPWR VGND 0.046438f
C25 VGND VNB 0.457657f
C26 VPWR VNB 0.310602f
C27 Y VNB 0.051086f
C28 A2 VNB 0.159216f
C29 A1 VNB 0.10514f
C30 B1 VNB 0.100569f
C31 B2 VNB 0.198256f
C32 VPB VNB 0.727632f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a22oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a22oi_2 VNB VPB VPWR VGND B2 A2 A1 Y B1
X0 VPWR.t3 A1.t0 a_66_368.t4 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X1 VGND.t2 A2.t0 a_148_74.t3 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 a_558_74.t1 B2.t0 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 a_148_74.t1 A1.t1 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 Y.t2 B1.t0 a_558_74.t2 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VGND.t0 B2.t1 a_558_74.t0 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1443 ps=1.13 w=0.74 l=0.15
X6 a_558_74.t3 B1.t1 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.1998 ps=1.28 w=0.74 l=0.15
X7 Y.t4 A1.t2 a_148_74.t0 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=1.28 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_66_368.t7 B1.t2 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X9 Y.t6 B1.t3 a_66_368.t5 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.168 ps=1.42 w=1.12 l=0.15
X10 Y.t1 B2.t2 a_66_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X11 a_66_368.t0 B2.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1848 ps=1.45 w=1.12 l=0.15
X12 a_66_368.t3 A1.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3416 ps=1.73 w=1.12 l=0.15
X13 a_148_74.t2 A2.t1 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X14 VPWR.t0 A2.t2 a_66_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.3416 pd=1.73 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_66_368.t2 A2.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
R0 A1 A1.n0 272.515
R1 A1.n1 A1.t0 250.909
R2 A1.n0 A1.t3 241.268
R3 A1.n1 A1.t1 220.113
R4 A1.n0 A1.t2 210.474
R5 A1.n2 A1.n1 152
R6 A1.n2 A1 16.4576
R7 A1 A1.n2 1.09764
R8 a_66_368.n4 a_66_368.t7 372.702
R9 a_66_368.n5 a_66_368.n4 303.401
R10 a_66_368.n2 a_66_368.n1 296.705
R11 a_66_368.n2 a_66_368.t4 275.812
R12 a_66_368.n3 a_66_368.n0 192.103
R13 a_66_368.n3 a_66_368.n2 73.5533
R14 a_66_368.n4 a_66_368.n3 61.4576
R15 a_66_368.n0 a_66_368.t5 26.3844
R16 a_66_368.n0 a_66_368.t3 26.3844
R17 a_66_368.n1 a_66_368.t1 26.3844
R18 a_66_368.n1 a_66_368.t2 26.3844
R19 a_66_368.n5 a_66_368.t6 26.3844
R20 a_66_368.t0 a_66_368.n5 26.3844
R21 VPWR.n2 VPWR.n0 618.254
R22 VPWR.n2 VPWR.n1 590.885
R23 VPWR.n1 VPWR.t2 53.6478
R24 VPWR.n1 VPWR.t0 53.6478
R25 VPWR.n0 VPWR.t1 26.3844
R26 VPWR.n0 VPWR.t3 26.3844
R27 VPWR VPWR.n2 0.414099
R28 VPB.t1 VPB.t3 388.173
R29 VPB VPB.t4 347.312
R30 VPB.t5 VPB.t0 245.161
R31 VPB.t6 VPB.t7 229.839
R32 VPB.t0 VPB.t6 229.839
R33 VPB.t3 VPB.t5 229.839
R34 VPB.t2 VPB.t1 229.839
R35 VPB.t4 VPB.t2 229.839
R36 A2.n0 A2.t2 226.809
R37 A2.n1 A2.t3 226.809
R38 A2.n1 A2.t0 201.125
R39 A2.n0 A2.t1 198.204
R40 A2 A2.n2 155.657
R41 A2.n2 A2.n0 53.3126
R42 A2.n2 A2.n1 12.4157
R43 a_148_74.n1 a_148_74.n0 351.613
R44 a_148_74.n0 a_148_74.t3 22.7032
R45 a_148_74.n0 a_148_74.t1 22.7032
R46 a_148_74.t0 a_148_74.n1 22.7032
R47 a_148_74.n1 a_148_74.t2 22.7032
R48 VGND.n2 VGND.n0 210.345
R49 VGND.n2 VGND.n1 209.833
R50 VGND.n1 VGND.t1 34.0546
R51 VGND.n0 VGND.t3 22.7032
R52 VGND.n0 VGND.t0 22.7032
R53 VGND.n1 VGND.t2 22.7032
R54 VGND VGND.n2 0.326924
R55 VNB.t2 VNB.t1 1593.7
R56 VNB VNB.t3 1535.96
R57 VNB.t1 VNB.t4 1247.24
R58 VNB.t6 VNB.t5 1154.86
R59 VNB.t7 VNB.t0 993.177
R60 VNB.t4 VNB.t7 993.177
R61 VNB.t5 VNB.t2 993.177
R62 VNB.t3 VNB.t6 993.177
R63 B2.n0 B2.t2 231.921
R64 B2.n1 B2.t3 226.809
R65 B2.n1 B2.t1 198.204
R66 B2.n0 B2.t0 196.013
R67 B2 B2.n2 154.522
R68 B2.n2 B2.n1 43.8187
R69 B2.n2 B2.n0 16.7975
R70 a_558_74.n1 a_558_74.n0 243.847
R71 a_558_74.n0 a_558_74.t3 34.0546
R72 a_558_74.n0 a_558_74.t0 29.1897
R73 a_558_74.n1 a_558_74.t2 22.7032
R74 a_558_74.t1 a_558_74.n1 22.7032
R75 Y.n2 Y.n1 300.733
R76 Y.n3 Y.n0 300.021
R77 Y.n4 Y.t5 273.053
R78 Y.n2 Y.t2 263.959
R79 Y.n6 Y.n5 94.176
R80 Y.n4 Y.n3 84.8518
R81 Y.n3 Y.n2 63.0068
R82 Y.n5 Y.t3 47.8383
R83 Y.n5 Y.t4 39.7302
R84 Y.n0 Y.t0 29.0228
R85 Y.n0 Y.t6 29.0228
R86 Y.n1 Y.t7 26.3844
R87 Y.n1 Y.t1 26.3844
R88 Y.n6 Y.n4 6.78613
R89 Y Y.n6 1.59803
R90 B1.n1 B1.t3 285.719
R91 B1.n0 B1.t2 264.298
R92 B1 B1.n0 225.763
R93 B1.n0 B1.t0 204.048
R94 B1.n1 B1.t1 178.34
R95 B1 B1.n1 158.4
C0 B2 VPWR 0.01134f
C1 B1 Y 0.222852f
C2 B1 VPB 0.06503f
C3 B1 VGND 0.030013f
C4 B2 Y 0.078735f
C5 B2 VPB 0.060882f
C6 B1 A1 0.0506f
C7 B2 VGND 0.025392f
C8 VPWR Y 0.028182f
C9 VPWR VPB 0.118381f
C10 VPWR VGND 0.07527f
C11 VPWR A1 0.055555f
C12 Y VPB 0.020331f
C13 Y VGND 0.149574f
C14 VGND VPB 0.008506f
C15 VPWR A2 0.024323f
C16 Y A1 0.197068f
C17 VPB A1 0.094422f
C18 VGND A1 0.024541f
C19 Y A2 0.057077f
C20 VPB A2 0.063976f
C21 VGND A2 0.024585f
C22 A1 A2 0.213367f
C23 B1 B2 0.207684f
C24 B1 VPWR 0.013289f
C25 VGND VNB 0.588935f
C26 Y VNB 0.171054f
C27 VPWR VNB 0.461716f
C28 B2 VNB 0.186381f
C29 B1 VNB 0.253341f
C30 A2 VNB 0.190026f
C31 A1 VNB 0.284228f
C32 VPB VNB 1.15618f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a22oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a22oi_4 VNB VPB VPWR VGND Y B2 B1 A2 A1
X0 Y.t8 B2.t0 a_45_368.t11 VPB.t12 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1 a_45_368.t10 B2.t1 Y.t7 VPB.t11 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y.t2 B1.t0 a_48_74.t7 VNB.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3 Y.t0 A1.t0 a_840_74.t3 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X4 Y.t3 B1.t1 a_48_74.t6 VNB.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 a_45_368.t3 A2.t0 VPWR.t7 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X6 Y.t6 B2.t2 a_45_368.t9 VPB.t10 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.308 ps=2.79 w=1.12 l=0.15
X7 VGND.t5 B2.t3 a_48_74.t3 VNB.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8 a_840_74.t2 A1.t1 Y.t9 VNB.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X9 VGND.t4 B2.t4 a_48_74.t2 VNB.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1961 ps=2.01 w=0.74 l=0.15
X10 a_840_74.t5 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X11 a_48_74.t1 B2.t5 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X12 a_840_74.t4 A2.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 VPWR.t6 A2.t3 a_45_368.t1 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X14 a_45_368.t2 A2.t4 VPWR.t5 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X15 a_48_74.t0 B2.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X16 a_840_74.t1 A1.t2 Y.t10 VNB.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X17 a_45_368.t5 A1.t3 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X18 VPWR.t4 A2.t5 a_45_368.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X19 VPWR.t2 A1.t4 a_45_368.t6 VPB.t6 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 VPWR.t1 A1.t5 a_45_368.t7 VPB.t7 sky130_fd_pr__pfet_01v8 ad=0.2968 pd=1.65 as=0.168 ps=1.42 w=1.12 l=0.15
X21 a_45_368.t8 A1.t6 VPWR.t0 VPB.t8 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.2968 ps=1.65 w=1.12 l=0.15
X22 a_45_368.t4 B1.t2 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X23 Y.t11 B1.t3 a_45_368.t13 VPB.t13 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X24 a_48_74.t5 B1.t4 Y.t12 VNB.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.1961 pd=2.01 as=0.1036 ps=1.02 w=0.74 l=0.15
X25 a_45_368.t14 B1.t5 Y.t13 VPB.t14 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X26 Y.t14 B1.t6 a_45_368.t15 VPB.t15 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X27 a_48_74.t4 B1.t7 Y.t15 VNB.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X28 a_45_368.t12 B2.t7 Y.t5 VPB.t9 sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X29 Y.t4 A1.t7 a_840_74.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
R0 B2.n0 B2.t7 234.841
R1 B2.n5 B2.t2 228.877
R2 B2.n2 B2.t0 226.809
R3 B2.n3 B2.t1 226.809
R4 B2.n5 B2.t4 196.744
R5 B2.n4 B2.t6 196.013
R6 B2.n10 B2.t3 196.013
R7 B2.n0 B2.t5 196.013
R8 B2 B2.n1 157.805
R9 B2.n12 B2.n11 152
R10 B2.n9 B2.n8 152
R11 B2.n7 B2.n6 152
R12 B2.n10 B2.n9 48.2005
R13 B2.n2 B2.n1 46.0096
R14 B2.n6 B2.n4 35.055
R15 B2.n6 B2.n5 27.0217
R16 B2.n9 B2.n3 12.4157
R17 B2.n1 B2.n0 11.6853
R18 B2.n8 B2.n7 10.1214
R19 B2.n12 B2 9.97259
R20 B2 B2.n12 4.31678
R21 B2.n7 B2 4.0191
R22 B2.n11 B2.n2 3.65202
R23 B2.n4 B2.n3 2.19141
R24 B2.n11 B2.n10 1.46111
R25 B2.n8 B2 0.149337
R26 a_45_368.n3 a_45_368.n2 303.495
R27 a_45_368.n5 a_45_368.n4 303.495
R28 a_45_368.n7 a_45_368.n6 303.495
R29 a_45_368.n1 a_45_368.t3 293.408
R30 a_45_368.n3 a_45_368.t9 290.704
R31 a_45_368.n1 a_45_368.n0 208.897
R32 a_45_368.n13 a_45_368.n12 206.404
R33 a_45_368.n11 a_45_368.n10 205.589
R34 a_45_368.n9 a_45_368.n8 186.73
R35 a_45_368.n11 a_45_368.n9 73.8951
R36 a_45_368.n9 a_45_368.n7 71.569
R37 a_45_368.n12 a_45_368.n1 61.3652
R38 a_45_368.n12 a_45_368.n11 60.2358
R39 a_45_368.n5 a_45_368.n3 42.9181
R40 a_45_368.n7 a_45_368.n5 42.9181
R41 a_45_368.n8 a_45_368.t6 26.3844
R42 a_45_368.n8 a_45_368.t4 26.3844
R43 a_45_368.n2 a_45_368.t11 26.3844
R44 a_45_368.n2 a_45_368.t10 26.3844
R45 a_45_368.n4 a_45_368.t15 26.3844
R46 a_45_368.n4 a_45_368.t12 26.3844
R47 a_45_368.n6 a_45_368.t13 26.3844
R48 a_45_368.n6 a_45_368.t14 26.3844
R49 a_45_368.n10 a_45_368.t7 26.3844
R50 a_45_368.n10 a_45_368.t5 26.3844
R51 a_45_368.n0 a_45_368.t1 26.3844
R52 a_45_368.n0 a_45_368.t2 26.3844
R53 a_45_368.t0 a_45_368.n13 26.3844
R54 a_45_368.n13 a_45_368.t8 26.3844
R55 Y.n3 Y.n2 360.558
R56 Y.n6 Y.n5 304.724
R57 Y.n3 Y.n1 300.733
R58 Y.n4 Y.n0 300.733
R59 Y.n14 Y.n12 243.052
R60 Y.n9 Y.n7 222.638
R61 Y.n14 Y.n13 185
R62 Y.n9 Y.n8 185
R63 Y.n4 Y.n3 67.7652
R64 Y.n6 Y.n4 61.3652
R65 Y.n11 Y.n6 37.817
R66 Y.n10 Y.n9 37.7761
R67 Y.n5 Y.t1 26.3844
R68 Y.n5 Y.t11 26.3844
R69 Y.n1 Y.t5 26.3844
R70 Y.n1 Y.t8 26.3844
R71 Y.n0 Y.t13 26.3844
R72 Y.n0 Y.t14 26.3844
R73 Y.n2 Y.t7 26.3844
R74 Y.n2 Y.t6 26.3844
R75 Y.n13 Y.t12 22.7032
R76 Y.n13 Y.t2 22.7032
R77 Y.n12 Y.t15 22.7032
R78 Y.n12 Y.t3 22.7032
R79 Y.n8 Y.t9 22.7032
R80 Y.n8 Y.t0 22.7032
R81 Y.n7 Y.t10 22.7032
R82 Y.n7 Y.t4 22.7032
R83 Y.n11 Y.n10 7.85117
R84 Y Y.n14 3.38053
R85 Y.n10 Y 1.56148
R86 Y Y.n11 0.2565
R87 VPB.t7 VPB.t8 347.312
R88 VPB VPB.t10 293.683
R89 VPB.t1 VPB.t3 229.839
R90 VPB.t2 VPB.t1 229.839
R91 VPB.t0 VPB.t2 229.839
R92 VPB.t8 VPB.t0 229.839
R93 VPB.t5 VPB.t7 229.839
R94 VPB.t6 VPB.t5 229.839
R95 VPB.t4 VPB.t6 229.839
R96 VPB.t13 VPB.t4 229.839
R97 VPB.t14 VPB.t13 229.839
R98 VPB.t15 VPB.t14 229.839
R99 VPB.t9 VPB.t15 229.839
R100 VPB.t12 VPB.t9 229.839
R101 VPB.t11 VPB.t12 229.839
R102 VPB.t10 VPB.t11 229.839
R103 B1.n0 B1.t2 244.883
R104 B1.n1 B1.t3 226.809
R105 B1.n4 B1.t5 226.809
R106 B1.n5 B1.t6 226.809
R107 B1.n5 B1.t1 198.175
R108 B1.n7 B1.t7 186.374
R109 B1.n2 B1.t0 186.374
R110 B1.n0 B1.t4 186.374
R111 B1.n6 B1 155.721
R112 B1 B1.n3 154.233
R113 B1.n9 B1.n8 152
R114 B1.n1 B1.n0 42.1755
R115 B1.n7 B1.n6 40.1672
R116 B1.n4 B1.n3 38.1588
R117 B1.n2 B1.n1 15.3977
R118 B1 B1.n9 7.88887
R119 B1.n8 B1.n4 7.36439
R120 B1.n6 B1.n5 7.36439
R121 B1.n3 B1.n2 6.69494
R122 B1.n9 B1 6.4005
R123 B1.n8 B1.n7 5.35606
R124 a_48_74.n1 a_48_74.t5 318.795
R125 a_48_74.n3 a_48_74.t2 201.567
R126 a_48_74.n1 a_48_74.n0 185
R127 a_48_74.n3 a_48_74.n2 104.579
R128 a_48_74.n5 a_48_74.n4 84.741
R129 a_48_74.n4 a_48_74.n1 83.804
R130 a_48_74.n4 a_48_74.n3 77.2621
R131 a_48_74.n2 a_48_74.t3 22.7032
R132 a_48_74.n2 a_48_74.t0 22.7032
R133 a_48_74.n0 a_48_74.t7 22.7032
R134 a_48_74.n0 a_48_74.t4 22.7032
R135 a_48_74.t6 a_48_74.n5 22.7032
R136 a_48_74.n5 a_48_74.t1 22.7032
R137 VNB.t9 VNB.t0 2194.23
R138 VNB.t1 VNB.t2 1986.35
R139 VNB.t13 VNB.t1 1986.35
R140 VNB VNB.t6 1339.63
R141 VNB.t3 VNB.t13 993.177
R142 VNB.t12 VNB.t3 993.177
R143 VNB.t0 VNB.t12 993.177
R144 VNB.t11 VNB.t9 993.177
R145 VNB.t8 VNB.t11 993.177
R146 VNB.t10 VNB.t8 993.177
R147 VNB.t5 VNB.t10 993.177
R148 VNB.t7 VNB.t5 993.177
R149 VNB.t4 VNB.t7 993.177
R150 VNB.t6 VNB.t4 993.177
R151 A1.n2 A1.t4 374.949
R152 A1.n1 A1.t6 226.809
R153 A1.n8 A1.t5 226.809
R154 A1.n3 A1.t3 226.809
R155 A1.n2 A1.t0 208.358
R156 A1.n1 A1.t2 206.969
R157 A1.n6 A1.t1 196.013
R158 A1.n9 A1.t7 196.013
R159 A1.n11 A1.n10 152
R160 A1.n7 A1.n0 152
R161 A1.n5 A1.n4 152
R162 A1.n10 A1.n1 50.3914
R163 A1.n9 A1.n8 47.4702
R164 A1.n6 A1.n5 35.055
R165 A1.n5 A1.n3 15.3369
R166 A1.n7 A1.n6 14.6066
R167 A1.n11 A1.n0 10.1214
R168 A1.n3 A1.n2 8.90371
R169 A1.n4 A1 7.5912
R170 A1.n4 A1 6.69817
R171 A1 A1.n0 3.42376
R172 A1.n10 A1.n9 1.46111
R173 A1 A1.n11 0.744686
R174 A1.n8 A1.n7 0.730803
R175 a_840_74.t3 a_840_74.n3 328.872
R176 a_840_74.n0 a_840_74.t5 198.651
R177 a_840_74.n3 a_840_74.n2 185
R178 a_840_74.n0 a_840_74.t4 152.905
R179 a_840_74.n1 a_840_74.t1 134.165
R180 a_840_74.n1 a_840_74.n0 68.8201
R181 a_840_74.n3 a_840_74.n1 57.1345
R182 a_840_74.n2 a_840_74.t0 22.7032
R183 a_840_74.n2 a_840_74.t2 22.7032
R184 A2.n10 A2.t5 234.841
R185 A2.n2 A2.t0 227.538
R186 A2.n5 A2.t3 226.809
R187 A2.n8 A2.t4 226.809
R188 A2.n10 A2.n9 196.013
R189 A2.n7 A2.t2 196.013
R190 A2.n4 A2.n1 196.013
R191 A2.n2 A2.t1 196.013
R192 A2.n3 A2.n0 162.121
R193 A2.n6 A2.n0 152
R194 A2.n14 A2.n13 152
R195 A2.n12 A2.n11 152
R196 A2.n13 A2.n12 49.6611
R197 A2.n7 A2.n6 39.4369
R198 A2.n3 A2.n2 36.5157
R199 A2.n4 A2.n3 26.2914
R200 A2.n6 A2.n5 21.1793
R201 A2.n11 A2 10.8656
R202 A2 A2.n14 7.5912
R203 A2.n14 A2 6.69817
R204 A2.n8 A2.n7 5.11262
R205 A2.n13 A2.n8 5.11262
R206 A2.n11 A2 3.42376
R207 A2.n12 A2.n10 2.92171
R208 A2 A2.n0 2.53073
R209 A2.n5 A2.n4 2.19141
R210 VPWR.n7 VPWR.n6 322.065
R211 VPWR.n5 VPWR.n4 316.683
R212 VPWR.n12 VPWR.n1 316.682
R213 VPWR.n10 VPWR.n3 309.861
R214 VPWR.n3 VPWR.t0 46.6121
R215 VPWR.n3 VPWR.t1 46.6121
R216 VPWR.n12 VPWR.n11 35.7652
R217 VPWR.n10 VPWR.n9 26.7299
R218 VPWR.n1 VPWR.t3 26.3844
R219 VPWR.n1 VPWR.t2 26.3844
R220 VPWR.n4 VPWR.t5 26.3844
R221 VPWR.n4 VPWR.t4 26.3844
R222 VPWR.n6 VPWR.t7 26.3844
R223 VPWR.n6 VPWR.t6 26.3844
R224 VPWR.n9 VPWR.n5 19.9534
R225 VPWR.n11 VPWR.n10 10.9181
R226 VPWR.n9 VPWR.n8 9.3005
R227 VPWR.n10 VPWR.n2 9.3005
R228 VPWR.n11 VPWR.n0 9.3005
R229 VPWR.n7 VPWR.n5 6.81595
R230 VPWR.n13 VPWR.n12 6.24654
R231 VPWR VPWR.n13 1.12018
R232 VPWR.n8 VPWR.n7 0.622084
R233 VPWR.n13 VPWR.n0 0.171605
R234 VPWR.n8 VPWR.n2 0.122949
R235 VPWR.n2 VPWR.n0 0.122949
R236 VGND.n8 VGND.t1 283.863
R237 VGND.n7 VGND.t0 277.608
R238 VGND.n26 VGND.n25 219.56
R239 VGND.n23 VGND.n2 211.183
R240 VGND.n11 VGND.n6 36.1417
R241 VGND.n12 VGND.n11 36.1417
R242 VGND.n13 VGND.n12 36.1417
R243 VGND.n13 VGND.n4 36.1417
R244 VGND.n17 VGND.n4 36.1417
R245 VGND.n18 VGND.n17 36.1417
R246 VGND.n19 VGND.n18 36.1417
R247 VGND.n19 VGND.n1 36.1417
R248 VGND.n23 VGND.n1 25.6005
R249 VGND.n26 VGND.n24 24.0946
R250 VGND.n7 VGND.n6 23.3417
R251 VGND.n2 VGND.t3 22.7032
R252 VGND.n2 VGND.t5 22.7032
R253 VGND.n25 VGND.t2 22.7032
R254 VGND.n25 VGND.t4 22.7032
R255 VGND.n24 VGND.n23 21.8358
R256 VGND.n9 VGND.n6 9.3005
R257 VGND.n11 VGND.n10 9.3005
R258 VGND.n12 VGND.n5 9.3005
R259 VGND.n14 VGND.n13 9.3005
R260 VGND.n15 VGND.n4 9.3005
R261 VGND.n17 VGND.n16 9.3005
R262 VGND.n18 VGND.n3 9.3005
R263 VGND.n20 VGND.n19 9.3005
R264 VGND.n21 VGND.n1 9.3005
R265 VGND.n23 VGND.n22 9.3005
R266 VGND.n24 VGND.n0 9.3005
R267 VGND.n27 VGND.n26 7.47871
R268 VGND.n8 VGND.n7 6.903
R269 VGND.n9 VGND.n8 0.654684
R270 VGND VGND.n27 0.16068
R271 VGND.n27 VGND.n0 0.14713
R272 VGND.n10 VGND.n9 0.122949
R273 VGND.n10 VGND.n5 0.122949
R274 VGND.n14 VGND.n5 0.122949
R275 VGND.n15 VGND.n14 0.122949
R276 VGND.n16 VGND.n15 0.122949
R277 VGND.n16 VGND.n3 0.122949
R278 VGND.n20 VGND.n3 0.122949
R279 VGND.n21 VGND.n20 0.122949
R280 VGND.n22 VGND.n21 0.122949
R281 VGND.n22 VGND.n0 0.122949
C0 A1 VGND 0.027227f
C1 A2 VPWR 0.083089f
C2 A2 VGND 0.065144f
C3 Y VPWR 0.037213f
C4 VPB B2 0.137232f
C5 Y VGND 0.047974f
C6 VPB B1 0.133339f
C7 VPWR VGND 0.128886f
C8 VPB A1 0.15257f
C9 B2 B1 0.08559f
C10 VPB A2 0.139051f
C11 VPB Y 0.008343f
C12 B1 A1 0.038984f
C13 B2 Y 0.164672f
C14 VPB VPWR 0.187358f
C15 A1 A2 0.100123f
C16 VPB VGND 0.010634f
C17 B2 VPWR 0.024299f
C18 B1 Y 0.340412f
C19 A1 Y 0.156697f
C20 B2 VGND 0.068803f
C21 B1 VPWR 0.023352f
C22 A2 Y 2.98e-19
C23 A1 VPWR 0.075935f
C24 B1 VGND 0.022512f
C25 VGND VNB 0.94116f
C26 VPWR VNB 0.740959f
C27 Y VNB 0.046336f
C28 A2 VNB 0.435f
C29 A1 VNB 0.41862f
C30 B1 VNB 0.400385f
C31 B2 VNB 0.432665f
C32 VPB VNB 1.90613f
.ends

* NGSPICE file created from sky130_fd_sc_hs__a31o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31o_1 VNB VPB VPWR VGND X A3 A2 A1 B1
X0 VGND.t1 a_81_270.t3 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.20655 pd=1.33 as=0.1961 ps=2.01 w=0.74 l=0.15
X1 VGND.t2 B1.t0 a_81_270.t2 VNB.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.1408 ps=1.08 w=0.64 l=0.15
X2 a_337_120.t1 A2.t0 a_265_120.t1 VNB.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.125625 pd=1.045 as=0.0672 ps=0.85 w=0.64 l=0.15
X3 a_81_270.t1 A1.t0 a_337_120.t0 VNB.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.1408 pd=1.08 as=0.125625 ps=1.045 w=0.64 l=0.15
X4 a_265_120.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.20655 ps=1.33 w=0.64 l=0.15
X5 VPWR.t3 A2.t1 a_250_392.t3 VPB.t4 sky130_fd_pr__pfet_01v8 ad=0.24 pd=1.48 as=0.15 ps=1.3 w=1 l=0.15
X6 a_250_392.t1 A3.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.2809 ps=1.65 w=1 l=0.15
X7 VPWR.t2 a_81_270.t4 X.t0 VPB.t3 sky130_fd_pr__pfet_01v8 ad=0.2809 pd=1.65 as=0.308 ps=2.79 w=1.12 l=0.15
X8 a_81_270.t0 B1.t1 a_250_392.t0 VPB.t0 sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.15 ps=1.3 w=1 l=0.15
X9 a_250_392.t2 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.24 ps=1.48 w=1 l=0.15
R0 a_81_270.t0 a_81_270.n2 300.745
R1 a_81_270.n2 a_81_270.n0 278.156
R2 a_81_270.n0 a_81_270.t4 249.531
R3 a_81_270.n2 a_81_270.n1 185
R4 a_81_270.n0 a_81_270.t3 176.964
R5 a_81_270.n1 a_81_270.t2 41.2505
R6 a_81_270.n1 a_81_270.t1 41.2505
R7 X X.n0 589.572
R8 X.n2 X.n0 585
R9 X.n1 X.n0 585
R10 X X.t1 196.423
R11 X.n0 X.t0 26.3844
R12 X X.n1 11.1548
R13 X X.n2 10.0576
R14 X.n2 X 3.47479
R15 X.n1 X 2.37764
R16 VGND.n1 VGND.t2 284.83
R17 VGND.n1 VGND.n0 99.5809
R18 VGND.n0 VGND.t0 51.0775
R19 VGND.n0 VGND.t1 43.5421
R20 VGND VGND.n1 0.251227
R21 VNB.t2 VNB.t0 1709.19
R22 VNB.t3 VNB.t4 1362.73
R23 VNB.t1 VNB.t3 1247.24
R24 VNB VNB.t2 1177.95
R25 VNB.t0 VNB.t1 831.496
R26 B1.t0 B1.t1 461.918
R27 B1 B1.t0 317.433
R28 A2.n0 A2.t1 231.629
R29 A2.n0 A2.t0 200.833
R30 A2 A2.n0 156.335
R31 a_265_120.t0 a_265_120.t1 39.3755
R32 a_337_120.t0 a_337_120.t1 68.1199
R33 A1.n0 A1.t1 231.629
R34 A1.n0 A1.t0 196.013
R35 A1 A1.n0 158.814
R36 A3.n0 A3.t1 231.629
R37 A3.n0 A3.t0 200.833
R38 A3 A3.n0 154.133
R39 a_250_392.n1 a_250_392.n0 467.031
R40 a_250_392.n0 a_250_392.t3 29.5505
R41 a_250_392.n0 a_250_392.t1 29.5505
R42 a_250_392.t0 a_250_392.n1 29.5505
R43 a_250_392.n1 a_250_392.t2 29.5505
R44 VPWR.n2 VPWR.n0 316.704
R45 VPWR.n2 VPWR.n1 219.501
R46 VPWR.n1 VPWR.t0 52.2055
R47 VPWR.n1 VPWR.t2 50.3459
R48 VPWR.n0 VPWR.t1 47.2805
R49 VPWR.n0 VPWR.t3 47.2805
R50 VPWR VPWR.n2 0.40776
R51 VPB.t3 VPB.t1 347.312
R52 VPB.t4 VPB.t2 321.774
R53 VPB VPB.t3 252.823
R54 VPB.t2 VPB.t0 229.839
R55 VPB.t1 VPB.t4 229.839
C0 VPB A3 0.045835f
C1 X VGND 0.075136f
C2 VPB A2 0.041266f
C3 VPWR VGND 0.057696f
C4 VPB A1 0.041636f
C5 A3 A2 0.091127f
C6 VPB B1 0.037817f
C7 VPB X 0.017134f
C8 A3 B1 9.97e-19
C9 A2 A1 0.073487f
C10 VPB VPWR 0.095688f
C11 A2 B1 0.008162f
C12 A3 X 0.005148f
C13 A1 B1 0.067154f
C14 VPB VGND 0.009719f
C15 A2 X 5.46e-19
C16 A3 VPWR 0.028251f
C17 A2 VPWR 0.016065f
C18 A1 X 2.84e-19
C19 A3 VGND 0.014408f
C20 A2 VGND 0.007713f
C21 A1 VPWR 0.016324f
C22 B1 X 8.66e-20
C23 B1 VPWR 0.009583f
C24 A1 VGND 0.006012f
C25 X VPWR 0.124474f
C26 B1 VGND 0.214039f
C27 VGND VNB 0.479723f
C28 VPWR VNB 0.347822f
C29 X VNB 0.106474f
C30 B1 VNB 0.188346f
C31 A1 VNB 0.095155f
C32 A2 VNB 0.09198f
C33 A3 VNB 0.097393f
C34 VPB VNB 0.834768f
.ends

