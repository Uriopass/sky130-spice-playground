INV1 cell simulation
.include "prelude.spice"

.include "inv_hd_nopex.spice"
.include "inv_hs.spice"

.param cval={{cval}}
.param risefall=0.01666n

xcell  A Vgnd Vgnd Vdd Vdd Y {{celltype}}

Vgnd Vgnd 0 0
Vdd Vdd Vgnd 1.8

Va  A  Vgnd pulse(0 1.8 0 {risefall} {risefall} 15n 20n)

Ccout Y  Vgnd {cval}

.tran 3p 5n 0

* .measure tran t_start_fall when V(A)=0.9 cross=1
* .measure tran t_end_fall   when V(Y)=0.9 cross=1
* .measure tran diff_time_fall PARAM='t_end_fall - t_start_fall'
* .measure tran t_start_rise when V(A)=0.9 cross=2
* .measure tran t_end_rise   when V(Y)=0.9 cross=2
* .measure tran diff_time_rise PARAM='t_end_rise - t_start_rise'

.control

* let loops = 6
* let i = 0
* let fall_times = vector(loops)
* let rise_times = vector(loops)
* let cval_vec   = vector(loops)
* set cvals = ( 1.6818300000p )
*
* foreach cval_l $cvals
*     alterparam cval = $cval_l
*     reset
*     run
*     meas tran t_start_fall when V(A)=0.9 cross=1
*     meas tran t_end_fall   when V(Y)=0.9 cross=1
*
*     meas tran t_start_rise when V(A)=0.9 cross=2
*     meas tran t_end_rise   when V(Y)=0.9 cross=2
*     let fall_times[i] = t_end_fall - t_start_fall
*     let rise_times[i] = t_end_rise - t_start_rise
*     let cval_vec[i] = $cval_l
*     let i = i + 1
*
*     plot V(A) V(Y) V(A2) V(Y2)
*     print t_end_fall - t_start_fall
*     print t_end_rise - t_start_rise
* end

* print (fall_times[1] - fall_times[0]) / (cval_vec[1] - cval_vec[0])
* print (rise_times[1] - rise_times[0]) / (cval_vec[1] - cval_vec[0])

* plot fall_times vs cval_vec rise_times vs cval_vec
* plot V(A) V(Y) V(A2) V(Y2)

run

*meas tran t_start_fall when V(A)=0.9 cross=2
*meas tran t_end_fall   when V(Y)=0.9 cross=2

meas tran t_start_rise when V(A)=0.9 cross=1
meas tran t_end_rise   when V(Y)=0.9 cross=1

.endc
