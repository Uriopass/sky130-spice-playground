.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y.t1 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
R0 A.n0 A.t1 230.576
R1 A A.n0 158.667
R2 A.n0 A.t0 158.275
R3 VGND VGND.t0 166.951
R4 Y.n0 Y.t0 235.56
R5 Y Y.t1 152.889
R6 Y Y.n0 2.22659
R7 Y.n0 Y 1.55202
R8 VNB VNB.t0 1612.5
R9 VPWR VPWR.t0 264.904
R10 VPB VPB.t0 350.853
C0 VPWR A 0.037031f
C1 VGND A 0.040045f
C2 A VPB 0.045062f
C3 VGND VPWR 0.033816f
C4 VPWR VPB 0.054478f
C5 Y A 0.047605f
C6 VGND VPB 0.009478f
C7 Y VPWR 0.127579f
C8 VGND Y 0.099841f
C9 Y VPB 0.017744f
C10 VGND VNB 0.251126f
C11 Y VNB 0.096099f
C12 VPWR VNB 0.218922f
C13 A VNB 0.166643f
C14 VPB VNB 0.338976f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t0 A.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n0 A.t3 212.081
R1 A.n1 A.t0 212.081
R2 A A.n1 189.073
R3 A.n0 A.t1 139.78
R4 A.n1 A.t2 139.78
R5 A.n1 A.n0 61.346
R6 VPWR.n0 VPWR.t0 262.851
R7 VPWR.n0 VPWR.t1 259.721
R8 VPWR VPWR.n0 0.491471
R9 Y.n2 Y.n1 208.965
R10 Y Y.n0 96.8352
R11 Y.n1 Y.t0 26.5955
R12 Y.n1 Y.t1 26.5955
R13 Y.n0 Y.t3 24.9236
R14 Y.n0 Y.t2 24.9236
R15 Y.n3 Y 11.2645
R16 Y Y.n3 6.1445
R17 Y.n3 Y 4.65505
R18 Y Y.n2 2.0485
R19 Y.n2 Y 1.55202
R20 VPB.t1 VPB.t0 248.599
R21 VPB VPB.t1 198.287
R22 VGND.n0 VGND.t1 169.418
R23 VGND.n0 VGND.t0 166.787
R24 VGND VGND.n0 0.491471
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 954.045
C0 Y VGND 0.154601f
C1 VPB A 0.074183f
C2 VPB VPWR 0.052063f
C3 A VPWR 0.06305f
C4 VGND VPB 0.006491f
C5 VGND A 0.063754f
C6 VGND VPWR 0.042274f
C7 Y VPB 0.006097f
C8 Y A 0.089386f
C9 Y VPWR 0.209105f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR.t3 A.t0 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t3 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t1 A.t3 Y.t7 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t2 A.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t6 A.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND.t1 A.t6 Y.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t4 A.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n2 A.t1 212.081
R2 A.n7 A.t3 212.081
R3 A.n3 A.t5 212.081
R4 A.n4 A.n3 188.516
R5 A A.n1 154.304
R6 A.n9 A.n8 152
R7 A.n6 A.n5 152
R8 A.n0 A.t6 139.78
R9 A.n2 A.t7 139.78
R10 A.n7 A.t4 139.78
R11 A.n3 A.t2 139.78
R12 A.n1 A.n0 30.6732
R13 A.n2 A.n1 30.6732
R14 A.n8 A.n2 30.6732
R15 A.n8 A.n7 30.6732
R16 A.n7 A.n6 30.6732
R17 A.n6 A.n3 30.6732
R18 A A.n9 19.2005
R19 A.n5 A 17.1525
R20 A A.n4 17.1525
R21 A.n5 A 6.4005
R22 A.n4 A 6.4005
R23 A.n9 A 4.3525
R24 Y.n5 Y.n4 244.069
R25 Y.n2 Y.n0 236.589
R26 Y.n5 Y.n3 204.893
R27 Y.n2 Y.n1 200.321
R28 Y.n3 Y.t1 26.5955
R29 Y.n3 Y.t0 26.5955
R30 Y.n4 Y.t7 26.5955
R31 Y.n4 Y.t6 26.5955
R32 Y.n0 Y.t2 24.9236
R33 Y.n0 Y.t3 24.9236
R34 Y.n1 Y.t5 24.9236
R35 Y.n1 Y.t4 24.9236
R36 Y Y.n5 18.4569
R37 Y.n6 Y 14.008
R38 Y.n6 Y.n2 12.0894
R39 Y Y.n6 2.41559
R40 VPWR.n2 VPWR.t3 884.006
R41 VPWR.n3 VPWR.n1 320.976
R42 VPWR.n5 VPWR.t0 248.843
R43 VPWR.n4 VPWR.n3 34.6358
R44 VPWR.n1 VPWR.t2 26.5955
R45 VPWR.n1 VPWR.t1 26.5955
R46 VPWR.n5 VPWR.n4 22.2123
R47 VPWR.n4 VPWR.n0 9.3005
R48 VPWR.n6 VPWR.n5 9.3005
R49 VPWR.n3 VPWR.n2 7.2029
R50 VPWR.n2 VPWR.n0 0.531054
R51 VPWR.n6 VPWR.n0 0.120292
R52 VPWR VPWR.n6 0.0226354
R53 VPB.t2 VPB.t3 248.599
R54 VPB.t1 VPB.t2 248.599
R55 VPB.t0 VPB.t1 248.599
R56 VPB VPB.t0 221.964
R57 VGND.n2 VGND.t1 292.346
R58 VGND.n5 VGND.t3 286.433
R59 VGND.n3 VGND.n1 207.213
R60 VGND.n4 VGND.n3 34.6358
R61 VGND.n1 VGND.t0 24.9236
R62 VGND.n1 VGND.t2 24.9236
R63 VGND.n5 VGND.n4 22.2123
R64 VGND.n6 VGND.n5 9.3005
R65 VGND.n4 VGND.n0 9.3005
R66 VGND.n3 VGND.n2 7.2029
R67 VGND.n2 VGND.n0 0.531054
R68 VGND.n6 VGND.n0 0.120292
R69 VGND VGND.n6 0.0226354
R70 VNB.t0 VNB.t1 1196.12
R71 VNB.t2 VNB.t0 1196.12
R72 VNB.t3 VNB.t2 1196.12
R73 VNB VNB.t3 1067.96
C0 VPB VPWR 0.065385f
C1 VPWR VGND 0.050092f
C2 A VPB 0.141975f
C3 A VGND 0.081909f
C4 VPB Y 0.015896f
C5 A VPWR 0.098226f
C6 Y VGND 0.262586f
C7 VPWR Y 0.361779f
C8 A Y 0.359887f
C9 VPB VGND 0.006668f
C10 VGND VNB 0.326816f
C11 Y VNB 0.084947f
C12 VPWR VNB 0.296394f
C13 A VNB 0.451855f
C14 VPB VNB 0.516168f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
X0 VPWR.t7 A.t0 Y.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t9 A.t2 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t12 A.t3 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t5 A.t4 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t3 A.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y.t11 A.t6 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR.t3 A.t7 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t10 A.t8 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t7 A.t9 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t1 A.t10 Y.t6 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t3 A.t11 Y.t15 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t2 A.t12 Y.t14 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t1 A.t13 Y.t13 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t5 A.t14 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t0 A.t15 Y.t8 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n1 A.t7 212.081
R1 A.n18 A.t9 212.081
R2 A.n16 A.t10 212.081
R3 A.n2 A.t14 212.081
R4 A.n11 A.t0 212.081
R5 A.n3 A.t1 212.081
R6 A.n6 A.t4 212.081
R7 A.n4 A.t5 212.081
R8 A.n5 A 163.264
R9 A A.n19 152
R10 A.n17 A.n0 152
R11 A.n15 A.n14 152
R12 A.n13 A.n12 152
R13 A.n10 A.n9 152
R14 A.n8 A.n7 152
R15 A.n1 A.t15 139.78
R16 A.n18 A.t3 139.78
R17 A.n16 A.t13 139.78
R18 A.n2 A.t2 139.78
R19 A.n11 A.t12 139.78
R20 A.n3 A.t8 139.78
R21 A.n6 A.t11 139.78
R22 A.n4 A.t6 139.78
R23 A.n19 A.n1 30.6732
R24 A.n19 A.n18 30.6732
R25 A.n18 A.n17 30.6732
R26 A.n17 A.n16 30.6732
R27 A.n16 A.n15 30.6732
R28 A.n15 A.n2 30.6732
R29 A.n12 A.n2 30.6732
R30 A.n12 A.n11 30.6732
R31 A.n11 A.n10 30.6732
R32 A.n10 A.n3 30.6732
R33 A.n7 A.n3 30.6732
R34 A.n7 A.n6 30.6732
R35 A.n6 A.n5 30.6732
R36 A.n5 A.n4 30.6732
R37 A A.n0 21.5045
R38 A.n14 A 19.4565
R39 A A.n13 17.4085
R40 A.n9 A 15.3605
R41 A A.n8 13.3125
R42 A.n8 A 10.2405
R43 A.n9 A 8.1925
R44 A.n13 A 6.1445
R45 A.n14 A 4.0965
R46 A A.n0 2.0485
R47 Y.n1 Y.n0 205.28
R48 Y.n3 Y.n2 205.28
R49 Y.n5 Y.n4 205.28
R50 Y.n7 Y.n6 205.28
R51 Y.n9 Y.n8 99.1759
R52 Y.n11 Y.n10 99.1759
R53 Y.n13 Y.n12 99.1759
R54 Y.n15 Y.n14 99.1759
R55 Y.n3 Y.n1 38.4005
R56 Y.n5 Y.n3 38.4005
R57 Y.n7 Y.n5 38.4005
R58 Y Y.n1 36.4472
R59 Y Y.n7 34.4358
R60 Y.n11 Y.n9 34.3584
R61 Y.n13 Y.n11 34.3584
R62 Y.n15 Y.n13 34.3584
R63 Y Y.n15 27.7875
R64 Y.n0 Y.t4 26.5955
R65 Y.n0 Y.t3 26.5955
R66 Y.n2 Y.t1 26.5955
R67 Y.n2 Y.t0 26.5955
R68 Y.n4 Y.t6 26.5955
R69 Y.n4 Y.t5 26.5955
R70 Y.n6 Y.t2 26.5955
R71 Y.n6 Y.t7 26.5955
R72 Y.n9 Y 25.611
R73 Y.n8 Y.t8 24.9236
R74 Y.n8 Y.t12 24.9236
R75 Y.n10 Y.t13 24.9236
R76 Y.n10 Y.t9 24.9236
R77 Y.n12 Y.t14 24.9236
R78 Y.n12 Y.t10 24.9236
R79 Y.n14 Y.t15 24.9236
R80 Y.n14 Y.t11 24.9236
R81 VPWR.n7 VPWR.t3 345.505
R82 VPWR.n17 VPWR.t4 342.375
R83 VPWR.n2 VPWR.n1 320.976
R84 VPWR.n10 VPWR.n4 320.976
R85 VPWR.n6 VPWR.n5 320.976
R86 VPWR.n12 VPWR.n11 34.6358
R87 VPWR.n16 VPWR.n15 34.6358
R88 VPWR.n10 VPWR.n9 32.0005
R89 VPWR.n9 VPWR.n6 31.2476
R90 VPWR.n1 VPWR.t6 26.5955
R91 VPWR.n1 VPWR.t5 26.5955
R92 VPWR.n4 VPWR.t0 26.5955
R93 VPWR.n4 VPWR.t7 26.5955
R94 VPWR.n5 VPWR.t2 26.5955
R95 VPWR.n5 VPWR.t1 26.5955
R96 VPWR.n12 VPWR.n2 25.977
R97 VPWR.n17 VPWR.n16 13.5534
R98 VPWR.n18 VPWR.n17 11.1829
R99 VPWR.n7 VPWR.n6 10.5481
R100 VPWR.n9 VPWR.n8 9.3005
R101 VPWR.n11 VPWR.n3 9.3005
R102 VPWR.n13 VPWR.n12 9.3005
R103 VPWR.n15 VPWR.n14 9.3005
R104 VPWR.n16 VPWR.n0 9.3005
R105 VPWR.n15 VPWR.n2 8.65932
R106 VPWR.n11 VPWR.n10 2.63579
R107 VPWR.n8 VPWR.n7 0.567773
R108 VPWR.n8 VPWR.n3 0.120292
R109 VPWR.n13 VPWR.n3 0.120292
R110 VPWR.n14 VPWR.n13 0.120292
R111 VPWR.n14 VPWR.n0 0.120292
R112 VPWR.n18 VPWR.n0 0.120292
R113 VPWR VPWR.n18 0.0226354
R114 VPB VPB.t4 290.031
R115 VPB.t2 VPB.t3 248.599
R116 VPB.t1 VPB.t2 248.599
R117 VPB.t0 VPB.t1 248.599
R118 VPB.t7 VPB.t0 248.599
R119 VPB.t6 VPB.t7 248.599
R120 VPB.t5 VPB.t6 248.599
R121 VPB.t4 VPB.t5 248.599
R122 VGND.n7 VGND.t0 290.637
R123 VGND.n17 VGND.t5 287.151
R124 VGND.n6 VGND.n5 207.213
R125 VGND.n10 VGND.n4 207.213
R126 VGND.n2 VGND.n1 207.213
R127 VGND.n12 VGND.n11 34.6358
R128 VGND.n16 VGND.n15 34.6358
R129 VGND.n10 VGND.n9 32.0005
R130 VGND.n9 VGND.n6 31.2476
R131 VGND.n12 VGND.n2 25.977
R132 VGND.n5 VGND.t6 24.9236
R133 VGND.n5 VGND.t1 24.9236
R134 VGND.n4 VGND.t7 24.9236
R135 VGND.n4 VGND.t2 24.9236
R136 VGND.n1 VGND.t4 24.9236
R137 VGND.n1 VGND.t3 24.9236
R138 VGND.n17 VGND.n16 13.5534
R139 VGND.n18 VGND.n17 11.1829
R140 VGND.n7 VGND.n6 10.5481
R141 VGND.n9 VGND.n8 9.3005
R142 VGND.n11 VGND.n3 9.3005
R143 VGND.n13 VGND.n12 9.3005
R144 VGND.n15 VGND.n14 9.3005
R145 VGND.n16 VGND.n0 9.3005
R146 VGND.n15 VGND.n2 8.65932
R147 VGND.n11 VGND.n10 2.63579
R148 VGND.n8 VGND.n7 0.567773
R149 VGND.n8 VGND.n3 0.120292
R150 VGND.n13 VGND.n3 0.120292
R151 VGND.n14 VGND.n13 0.120292
R152 VGND.n14 VGND.n0 0.120292
R153 VGND.n18 VGND.n0 0.120292
R154 VGND VGND.n18 0.0226354
R155 VNB VNB.t5 1395.47
R156 VNB.t6 VNB.t0 1196.12
R157 VNB.t1 VNB.t6 1196.12
R158 VNB.t7 VNB.t1 1196.12
R159 VNB.t2 VNB.t7 1196.12
R160 VNB.t4 VNB.t2 1196.12
R161 VNB.t3 VNB.t4 1196.12
R162 VNB.t5 VNB.t3 1196.12
C0 Y VPB 0.034787f
C1 VPWR A 0.127577f
C2 Y VGND 0.574497f
C3 VPB VPWR 0.100209f
C4 VGND VPWR 0.085433f
C5 Y VPWR 0.779949f
C6 VPB A 0.254088f
C7 VGND A 0.116857f
C8 VPB VGND 0.007925f
C9 Y A 0.829319f
C10 VGND VNB 0.51049f
C11 Y VNB 0.126735f
C12 VPWR VNB 0.449913f
C13 A VNB 0.771261f
C14 VPB VNB 0.870552f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 Y.t15 A.t0 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t9 A.t1 Y.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t15 A.t2 Y.t25 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t13 A.t3 VPWR.t8 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t14 A.t4 Y.t18 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t13 A.t5 Y.t17 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t12 A.t6 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t12 A.t7 Y.t16 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t6 A.t8 Y.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t24 A.t9 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR.t15 A.t10 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y.t23 A.t11 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y.t9 A.t12 VPWR.t14 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR.t13 A.t13 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t7 A.t14 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t9 A.t15 Y.t22 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y.t21 A.t16 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND.t7 A.t17 Y.t20 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t6 A.t18 Y.t19 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y.t6 A.t19 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t5 A.t20 Y.t28 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t5 A.t21 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t2 A.t22 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t1 A.t23 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t0 A.t24 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t27 A.t25 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y.t1 A.t26 VPWR.t12 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t26 A.t27 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y.t31 A.t28 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t30 A.t29 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR.t11 A.t30 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y.t29 A.t31 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n2 A.t1 212.081
R1 A.n3 A.t3 212.081
R2 A.n4 A.t8 212.081
R3 A.n5 A.t14 212.081
R4 A.n6 A.t22 212.081
R5 A.n1 A.t21 212.081
R6 A.n10 A.t24 212.081
R7 A.n11 A.t26 212.081
R8 A.n25 A.t30 212.081
R9 A.n24 A.t0 212.081
R10 A.n22 A.t10 212.081
R11 A.n21 A.t12 212.081
R12 A.n12 A.t13 212.081
R13 A.n14 A.t19 212.081
R14 A.n16 A.t23 212.081
R15 A.n15 A.t6 212.081
R16 A.n8 A.n7 196.534
R17 A.n15 A.n13 187.055
R18 A.n9 A.n8 152
R19 A.n27 A.n26 152
R20 A.n23 A.n0 152
R21 A.n20 A.n19 152
R22 A.n18 A.n17 152
R23 A.n2 A.t7 139.78
R24 A.n3 A.t11 139.78
R25 A.n4 A.t5 139.78
R26 A.n5 A.t27 139.78
R27 A.n6 A.t2 139.78
R28 A.n1 A.t31 139.78
R29 A.n10 A.t4 139.78
R30 A.n11 A.t29 139.78
R31 A.n25 A.t20 139.78
R32 A.n24 A.t28 139.78
R33 A.n22 A.t18 139.78
R34 A.n21 A.t25 139.78
R35 A.n12 A.t17 139.78
R36 A.n14 A.t9 139.78
R37 A.n16 A.t15 139.78
R38 A.n15 A.t16 139.78
R39 A.n3 A.n2 61.346
R40 A.n4 A.n3 61.346
R41 A.n5 A.n4 61.346
R42 A.n6 A.n1 61.346
R43 A.n11 A.n10 61.346
R44 A.n25 A.n24 61.346
R45 A.n22 A.n21 61.346
R46 A.n14 A.n12 61.346
R47 A.n16 A.n15 61.346
R48 A.n18 A.n13 46.4005
R49 A.n19 A.n0 45.0672
R50 A.n27 A.n0 44.5338
R51 A A.n18 43.7338
R52 A.n7 A.n5 31.4035
R53 A.n23 A.n22 31.4035
R54 A.n9 A.n1 30.6732
R55 A.n10 A.n9 30.6732
R56 A.n26 A.n11 30.6732
R57 A.n26 A.n25 30.6732
R58 A.n21 A.n20 30.6732
R59 A.n20 A.n12 30.6732
R60 A.n17 A.n14 30.6732
R61 A.n17 A.n16 30.6732
R62 A.n7 A.n6 29.9429
R63 A.n24 A.n23 29.9429
R64 A.n8 A 12.8005
R65 A.n13 A 8.0005
R66 A A.n27 7.46717
R67 A.n19 A 1.06717
R68 VPWR.n14 VPWR.t9 354.187
R69 VPWR.n2 VPWR.n1 320.976
R70 VPWR.n33 VPWR.n4 320.976
R71 VPWR.n6 VPWR.n5 320.976
R72 VPWR.n26 VPWR.n8 320.976
R73 VPWR.n20 VPWR.n19 320.976
R74 VPWR.n17 VPWR.n11 320.976
R75 VPWR.n13 VPWR.n12 320.976
R76 VPWR.n39 VPWR.t7 255.965
R77 VPWR.n21 VPWR.n18 34.6358
R78 VPWR.n25 VPWR.n9 34.6358
R79 VPWR.n28 VPWR.n27 34.6358
R80 VPWR.n32 VPWR.n31 34.6358
R81 VPWR.n38 VPWR.n37 34.6358
R82 VPWR.n16 VPWR.n13 34.2593
R83 VPWR.n34 VPWR.n2 33.5064
R84 VPWR.n34 VPWR.n33 29.7417
R85 VPWR.n17 VPWR.n16 28.9887
R86 VPWR.n1 VPWR.t4 26.5955
R87 VPWR.n1 VPWR.t1 26.5955
R88 VPWR.n4 VPWR.t14 26.5955
R89 VPWR.n4 VPWR.t13 26.5955
R90 VPWR.n5 VPWR.t10 26.5955
R91 VPWR.n5 VPWR.t15 26.5955
R92 VPWR.n8 VPWR.t12 26.5955
R93 VPWR.n8 VPWR.t11 26.5955
R94 VPWR.n19 VPWR.t3 26.5955
R95 VPWR.n19 VPWR.t0 26.5955
R96 VPWR.n11 VPWR.t5 26.5955
R97 VPWR.n11 VPWR.t2 26.5955
R98 VPWR.n12 VPWR.t8 26.5955
R99 VPWR.n12 VPWR.t6 26.5955
R100 VPWR.n31 VPWR.n6 23.7181
R101 VPWR.n21 VPWR.n20 22.9652
R102 VPWR.n39 VPWR.n38 21.0829
R103 VPWR.n27 VPWR.n26 17.6946
R104 VPWR.n26 VPWR.n25 16.9417
R105 VPWR.n20 VPWR.n9 11.6711
R106 VPWR.n28 VPWR.n6 10.9181
R107 VPWR.n16 VPWR.n15 9.3005
R108 VPWR.n18 VPWR.n10 9.3005
R109 VPWR.n22 VPWR.n21 9.3005
R110 VPWR.n23 VPWR.n9 9.3005
R111 VPWR.n25 VPWR.n24 9.3005
R112 VPWR.n27 VPWR.n7 9.3005
R113 VPWR.n29 VPWR.n28 9.3005
R114 VPWR.n31 VPWR.n30 9.3005
R115 VPWR.n32 VPWR.n3 9.3005
R116 VPWR.n35 VPWR.n34 9.3005
R117 VPWR.n37 VPWR.n36 9.3005
R118 VPWR.n38 VPWR.n0 9.3005
R119 VPWR.n40 VPWR.n39 9.3005
R120 VPWR.n14 VPWR.n13 7.57496
R121 VPWR.n18 VPWR.n17 5.64756
R122 VPWR.n33 VPWR.n32 4.89462
R123 VPWR.n37 VPWR.n2 1.12991
R124 VPWR.n15 VPWR.n14 0.534819
R125 VPWR.n15 VPWR.n10 0.120292
R126 VPWR.n22 VPWR.n10 0.120292
R127 VPWR.n23 VPWR.n22 0.120292
R128 VPWR.n24 VPWR.n23 0.120292
R129 VPWR.n24 VPWR.n7 0.120292
R130 VPWR.n29 VPWR.n7 0.120292
R131 VPWR.n30 VPWR.n29 0.120292
R132 VPWR.n30 VPWR.n3 0.120292
R133 VPWR.n35 VPWR.n3 0.120292
R134 VPWR.n36 VPWR.n35 0.120292
R135 VPWR.n36 VPWR.n0 0.120292
R136 VPWR.n40 VPWR.n0 0.120292
R137 VPWR VPWR.n40 0.0226354
R138 Y.n15 Y.n13 243.458
R139 Y.n15 Y.n14 205.059
R140 Y.n17 Y.n16 205.059
R141 Y.n19 Y.n18 205.059
R142 Y.n21 Y.n20 205.059
R143 Y.n23 Y.n22 205.059
R144 Y.n25 Y.n24 205.059
R145 Y.n27 Y.n26 205.059
R146 Y.n2 Y.n0 133.534
R147 Y.n2 Y.n1 99.1759
R148 Y.n4 Y.n3 99.1759
R149 Y.n6 Y.n5 99.1759
R150 Y.n8 Y.n7 99.1759
R151 Y.n10 Y.n9 99.1759
R152 Y.n12 Y.n11 99.1759
R153 Y Y.n29 97.4305
R154 Y.n17 Y.n15 38.4005
R155 Y.n19 Y.n17 38.4005
R156 Y.n21 Y.n19 38.4005
R157 Y.n23 Y.n21 38.4005
R158 Y.n25 Y.n23 38.4005
R159 Y.n27 Y.n25 38.4005
R160 Y.n4 Y.n2 34.3584
R161 Y.n6 Y.n4 34.3584
R162 Y.n8 Y.n6 34.3584
R163 Y.n10 Y.n8 34.3584
R164 Y.n12 Y.n10 34.3584
R165 Y.n28 Y.n12 34.3584
R166 Y.n26 Y.t14 26.5955
R167 Y.n26 Y.t13 26.5955
R168 Y.n13 Y.t3 26.5955
R169 Y.n13 Y.t12 26.5955
R170 Y.n14 Y.t8 26.5955
R171 Y.n14 Y.t6 26.5955
R172 Y.n16 Y.t10 26.5955
R173 Y.n16 Y.t9 26.5955
R174 Y.n18 Y.t0 26.5955
R175 Y.n18 Y.t15 26.5955
R176 Y.n20 Y.t2 26.5955
R177 Y.n20 Y.t1 26.5955
R178 Y.n22 Y.t4 26.5955
R179 Y.n22 Y.t5 26.5955
R180 Y.n24 Y.t11 26.5955
R181 Y.n24 Y.t7 26.5955
R182 Y.n29 Y.t16 24.9236
R183 Y.n29 Y.t23 24.9236
R184 Y.n0 Y.t22 24.9236
R185 Y.n0 Y.t21 24.9236
R186 Y.n1 Y.t20 24.9236
R187 Y.n1 Y.t24 24.9236
R188 Y.n3 Y.t19 24.9236
R189 Y.n3 Y.t27 24.9236
R190 Y.n5 Y.t28 24.9236
R191 Y.n5 Y.t31 24.9236
R192 Y.n7 Y.t18 24.9236
R193 Y.n7 Y.t30 24.9236
R194 Y.n9 Y.t25 24.9236
R195 Y.n9 Y.t29 24.9236
R196 Y.n11 Y.t17 24.9236
R197 Y.n11 Y.t26 24.9236
R198 Y Y.n27 18.4247
R199 Y.n28 Y 11.4429
R200 Y Y.n28 1.74595
R201 VPB.t13 VPB.t14 248.599
R202 VPB.t11 VPB.t13 248.599
R203 VPB.t7 VPB.t11 248.599
R204 VPB.t4 VPB.t7 248.599
R205 VPB.t5 VPB.t4 248.599
R206 VPB.t2 VPB.t5 248.599
R207 VPB.t1 VPB.t2 248.599
R208 VPB.t0 VPB.t1 248.599
R209 VPB.t15 VPB.t0 248.599
R210 VPB.t10 VPB.t15 248.599
R211 VPB.t9 VPB.t10 248.599
R212 VPB.t8 VPB.t9 248.599
R213 VPB.t6 VPB.t8 248.599
R214 VPB.t3 VPB.t6 248.599
R215 VPB.t12 VPB.t3 248.599
R216 VPB VPB.t12 230.841
R217 VGND.n13 VGND.n12 207.213
R218 VGND.n17 VGND.n11 207.213
R219 VGND.n20 VGND.n19 207.213
R220 VGND.n26 VGND.n8 207.213
R221 VGND.n6 VGND.n5 207.213
R222 VGND.n33 VGND.n4 207.213
R223 VGND.n2 VGND.n1 207.213
R224 VGND.n14 VGND.t12 166.852
R225 VGND.n39 VGND.t8 157.567
R226 VGND.n21 VGND.n18 34.6358
R227 VGND.n25 VGND.n9 34.6358
R228 VGND.n28 VGND.n27 34.6358
R229 VGND.n32 VGND.n31 34.6358
R230 VGND.n38 VGND.n37 34.6358
R231 VGND.n16 VGND.n13 34.2593
R232 VGND.n34 VGND.n2 33.5064
R233 VGND.n34 VGND.n33 29.7417
R234 VGND.n17 VGND.n16 28.9887
R235 VGND.n12 VGND.t10 24.9236
R236 VGND.n12 VGND.t13 24.9236
R237 VGND.n11 VGND.t3 24.9236
R238 VGND.n11 VGND.t15 24.9236
R239 VGND.n19 VGND.t0 24.9236
R240 VGND.n19 VGND.t14 24.9236
R241 VGND.n8 VGND.t1 24.9236
R242 VGND.n8 VGND.t5 24.9236
R243 VGND.n5 VGND.t2 24.9236
R244 VGND.n5 VGND.t6 24.9236
R245 VGND.n4 VGND.t4 24.9236
R246 VGND.n4 VGND.t7 24.9236
R247 VGND.n1 VGND.t11 24.9236
R248 VGND.n1 VGND.t9 24.9236
R249 VGND.n31 VGND.n6 23.7181
R250 VGND.n21 VGND.n20 22.9652
R251 VGND.n39 VGND.n38 21.0829
R252 VGND.n27 VGND.n26 17.6946
R253 VGND.n26 VGND.n25 16.9417
R254 VGND.n20 VGND.n9 11.6711
R255 VGND.n28 VGND.n6 10.9181
R256 VGND.n40 VGND.n39 9.3005
R257 VGND.n16 VGND.n15 9.3005
R258 VGND.n18 VGND.n10 9.3005
R259 VGND.n22 VGND.n21 9.3005
R260 VGND.n23 VGND.n9 9.3005
R261 VGND.n25 VGND.n24 9.3005
R262 VGND.n27 VGND.n7 9.3005
R263 VGND.n29 VGND.n28 9.3005
R264 VGND.n31 VGND.n30 9.3005
R265 VGND.n32 VGND.n3 9.3005
R266 VGND.n35 VGND.n34 9.3005
R267 VGND.n37 VGND.n36 9.3005
R268 VGND.n38 VGND.n0 9.3005
R269 VGND.n14 VGND.n13 7.57496
R270 VGND.n18 VGND.n17 5.64756
R271 VGND.n33 VGND.n32 4.89462
R272 VGND.n37 VGND.n2 1.12991
R273 VGND.n15 VGND.n14 0.534819
R274 VGND.n15 VGND.n10 0.120292
R275 VGND.n22 VGND.n10 0.120292
R276 VGND.n23 VGND.n22 0.120292
R277 VGND.n24 VGND.n23 0.120292
R278 VGND.n24 VGND.n7 0.120292
R279 VGND.n29 VGND.n7 0.120292
R280 VGND.n30 VGND.n29 0.120292
R281 VGND.n30 VGND.n3 0.120292
R282 VGND.n35 VGND.n3 0.120292
R283 VGND.n36 VGND.n35 0.120292
R284 VGND.n36 VGND.n0 0.120292
R285 VGND.n40 VGND.n0 0.120292
R286 VGND VGND.n40 0.0226354
R287 VNB.t10 VNB.t12 1196.12
R288 VNB.t13 VNB.t10 1196.12
R289 VNB.t3 VNB.t13 1196.12
R290 VNB.t15 VNB.t3 1196.12
R291 VNB.t0 VNB.t15 1196.12
R292 VNB.t14 VNB.t0 1196.12
R293 VNB.t1 VNB.t14 1196.12
R294 VNB.t5 VNB.t1 1196.12
R295 VNB.t2 VNB.t5 1196.12
R296 VNB.t6 VNB.t2 1196.12
R297 VNB.t4 VNB.t6 1196.12
R298 VNB.t7 VNB.t4 1196.12
R299 VNB.t11 VNB.t7 1196.12
R300 VNB.t9 VNB.t11 1196.12
R301 VNB.t8 VNB.t9 1196.12
R302 VNB VNB.t8 1110.68
C0 VGND VPWR 0.160762f
C1 VGND Y 1.06261f
C2 A VPB 0.525745f
C3 VPWR VPB 0.159316f
C4 Y VPB 0.03049f
C5 VPWR A 0.280261f
C6 Y A 1.4347f
C7 VGND VPB 0.013189f
C8 Y VPWR 1.46621f
C9 VGND A 0.265874f
C10 VGND VNB 0.864536f
C11 Y VNB 0.055057f
C12 VPWR VNB 0.737072f
C13 A VNB 1.54575f
C14 VPB VNB 1.49072f
.ends
