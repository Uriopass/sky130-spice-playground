* NGSPICE file created from sky130_fd_sc_hd__inv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y.t1 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
R0 A.n0 A.t1 230.576
R1 A A.n0 158.667
R2 A.n0 A.t0 158.275
R3 VGND VGND.t0 166.951
R4 Y.n0 Y.t0 235.56
R5 Y Y.t1 152.889
R6 Y Y.n0 2.22659
R7 Y.n0 Y 1.55202
R8 VNB VNB.t0 1612.5
R9 VPWR VPWR.t0 264.904
R10 VPB VPB.t0 350.853
C0 VPWR A 0.037031f
C1 VGND A 0.040045f
C2 A VPB 0.045062f
C3 VGND VPWR 0.033816f
C4 VPWR VPB 0.054478f
C5 Y A 0.047605f
C6 VGND VPB 0.009478f
C7 Y VPWR 0.127579f
C8 VGND Y 0.099841f
C9 Y VPB 0.017744f
C10 VGND VNB 0.251126f
C11 Y VNB 0.096099f
C12 VPWR VNB 0.218922f
C13 A VNB 0.166643f
C14 VPB VNB 0.338976f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t0 A.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n0 A.t3 212.081
R1 A.n1 A.t0 212.081
R2 A A.n1 189.073
R3 A.n0 A.t1 139.78
R4 A.n1 A.t2 139.78
R5 A.n1 A.n0 61.346
R6 VPWR.n0 VPWR.t0 262.851
R7 VPWR.n0 VPWR.t1 259.721
R8 VPWR VPWR.n0 0.491471
R9 Y.n2 Y.n1 208.965
R10 Y Y.n0 96.8352
R11 Y.n1 Y.t0 26.5955
R12 Y.n1 Y.t1 26.5955
R13 Y.n0 Y.t3 24.9236
R14 Y.n0 Y.t2 24.9236
R15 Y.n3 Y 11.2645
R16 Y Y.n3 6.1445
R17 Y.n3 Y 4.65505
R18 Y Y.n2 2.0485
R19 Y.n2 Y 1.55202
R20 VPB.t1 VPB.t0 248.599
R21 VPB VPB.t1 198.287
R22 VGND.n0 VGND.t1 169.418
R23 VGND.n0 VGND.t0 166.787
R24 VGND VGND.n0 0.491471
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 954.045
C0 Y VGND 0.154601f
C1 VPB A 0.074183f
C2 VPB VPWR 0.052063f
C3 A VPWR 0.06305f
C4 VGND VPB 0.006491f
C5 VGND A 0.063754f
C6 VGND VPWR 0.042274f
C7 Y VPB 0.006097f
C8 Y A 0.089386f
C9 Y VPWR 0.209105f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR.t3 A.t0 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t3 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t1 A.t3 Y.t7 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t2 A.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t6 A.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND.t1 A.t6 Y.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t4 A.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n2 A.t1 212.081
R2 A.n7 A.t3 212.081
R3 A.n3 A.t5 212.081
R4 A.n4 A.n3 188.516
R5 A A.n1 154.304
R6 A.n9 A.n8 152
R7 A.n6 A.n5 152
R8 A.n0 A.t6 139.78
R9 A.n2 A.t7 139.78
R10 A.n7 A.t4 139.78
R11 A.n3 A.t2 139.78
R12 A.n1 A.n0 30.6732
R13 A.n2 A.n1 30.6732
R14 A.n8 A.n2 30.6732
R15 A.n8 A.n7 30.6732
R16 A.n7 A.n6 30.6732
R17 A.n6 A.n3 30.6732
R18 A A.n9 19.2005
R19 A.n5 A 17.1525
R20 A A.n4 17.1525
R21 A.n5 A 6.4005
R22 A.n4 A 6.4005
R23 A.n9 A 4.3525
R24 Y.n5 Y.n4 244.069
R25 Y.n2 Y.n0 236.589
R26 Y.n5 Y.n3 204.893
R27 Y.n2 Y.n1 200.321
R28 Y.n3 Y.t1 26.5955
R29 Y.n3 Y.t0 26.5955
R30 Y.n4 Y.t7 26.5955
R31 Y.n4 Y.t6 26.5955
R32 Y.n0 Y.t2 24.9236
R33 Y.n0 Y.t3 24.9236
R34 Y.n1 Y.t5 24.9236
R35 Y.n1 Y.t4 24.9236
R36 Y Y.n5 18.4569
R37 Y.n6 Y 14.008
R38 Y.n6 Y.n2 12.0894
R39 Y Y.n6 2.41559
R40 VPWR.n2 VPWR.t3 884.006
R41 VPWR.n3 VPWR.n1 320.976
R42 VPWR.n5 VPWR.t0 248.843
R43 VPWR.n4 VPWR.n3 34.6358
R44 VPWR.n1 VPWR.t2 26.5955
R45 VPWR.n1 VPWR.t1 26.5955
R46 VPWR.n5 VPWR.n4 22.2123
R47 VPWR.n4 VPWR.n0 9.3005
R48 VPWR.n6 VPWR.n5 9.3005
R49 VPWR.n3 VPWR.n2 7.2029
R50 VPWR.n2 VPWR.n0 0.531054
R51 VPWR.n6 VPWR.n0 0.120292
R52 VPWR VPWR.n6 0.0226354
R53 VPB.t2 VPB.t3 248.599
R54 VPB.t1 VPB.t2 248.599
R55 VPB.t0 VPB.t1 248.599
R56 VPB VPB.t0 221.964
R57 VGND.n2 VGND.t1 292.346
R58 VGND.n5 VGND.t3 286.433
R59 VGND.n3 VGND.n1 207.213
R60 VGND.n4 VGND.n3 34.6358
R61 VGND.n1 VGND.t0 24.9236
R62 VGND.n1 VGND.t2 24.9236
R63 VGND.n5 VGND.n4 22.2123
R64 VGND.n6 VGND.n5 9.3005
R65 VGND.n4 VGND.n0 9.3005
R66 VGND.n3 VGND.n2 7.2029
R67 VGND.n2 VGND.n0 0.531054
R68 VGND.n6 VGND.n0 0.120292
R69 VGND VGND.n6 0.0226354
R70 VNB.t0 VNB.t1 1196.12
R71 VNB.t2 VNB.t0 1196.12
R72 VNB.t3 VNB.t2 1196.12
R73 VNB VNB.t3 1067.96
C0 VPB VPWR 0.065385f
C1 VPWR VGND 0.050092f
C2 A VPB 0.141975f
C3 A VGND 0.081909f
C4 VPB Y 0.015896f
C5 A VPWR 0.098226f
C6 Y VGND 0.262586f
C7 VPWR Y 0.361779f
C8 A Y 0.359887f
C9 VPB VGND 0.006668f
C10 VGND VNB 0.326816f
C11 Y VNB 0.084947f
C12 VPWR VNB 0.296394f
C13 A VNB 0.451855f
C14 VPB VNB 0.516168f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
X0 VPWR.t7 A.t0 Y.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t9 A.t2 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t12 A.t3 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t5 A.t4 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t3 A.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y.t11 A.t6 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR.t3 A.t7 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t10 A.t8 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t7 A.t9 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t1 A.t10 Y.t6 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t3 A.t11 Y.t15 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t2 A.t12 Y.t14 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t1 A.t13 Y.t13 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t5 A.t14 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t0 A.t15 Y.t8 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n1 A.t7 212.081
R1 A.n18 A.t9 212.081
R2 A.n16 A.t10 212.081
R3 A.n2 A.t14 212.081
R4 A.n11 A.t0 212.081
R5 A.n3 A.t1 212.081
R6 A.n6 A.t4 212.081
R7 A.n4 A.t5 212.081
R8 A.n5 A 163.264
R9 A A.n19 152
R10 A.n17 A.n0 152
R11 A.n15 A.n14 152
R12 A.n13 A.n12 152
R13 A.n10 A.n9 152
R14 A.n8 A.n7 152
R15 A.n1 A.t15 139.78
R16 A.n18 A.t3 139.78
R17 A.n16 A.t13 139.78
R18 A.n2 A.t2 139.78
R19 A.n11 A.t12 139.78
R20 A.n3 A.t8 139.78
R21 A.n6 A.t11 139.78
R22 A.n4 A.t6 139.78
R23 A.n19 A.n1 30.6732
R24 A.n19 A.n18 30.6732
R25 A.n18 A.n17 30.6732
R26 A.n17 A.n16 30.6732
R27 A.n16 A.n15 30.6732
R28 A.n15 A.n2 30.6732
R29 A.n12 A.n2 30.6732
R30 A.n12 A.n11 30.6732
R31 A.n11 A.n10 30.6732
R32 A.n10 A.n3 30.6732
R33 A.n7 A.n3 30.6732
R34 A.n7 A.n6 30.6732
R35 A.n6 A.n5 30.6732
R36 A.n5 A.n4 30.6732
R37 A A.n0 21.5045
R38 A.n14 A 19.4565
R39 A A.n13 17.4085
R40 A.n9 A 15.3605
R41 A A.n8 13.3125
R42 A.n8 A 10.2405
R43 A.n9 A 8.1925
R44 A.n13 A 6.1445
R45 A.n14 A 4.0965
R46 A A.n0 2.0485
R47 Y.n1 Y.n0 205.28
R48 Y.n3 Y.n2 205.28
R49 Y.n5 Y.n4 205.28
R50 Y.n7 Y.n6 205.28
R51 Y.n9 Y.n8 99.1759
R52 Y.n11 Y.n10 99.1759
R53 Y.n13 Y.n12 99.1759
R54 Y.n15 Y.n14 99.1759
R55 Y.n3 Y.n1 38.4005
R56 Y.n5 Y.n3 38.4005
R57 Y.n7 Y.n5 38.4005
R58 Y Y.n1 36.4472
R59 Y Y.n7 34.4358
R60 Y.n11 Y.n9 34.3584
R61 Y.n13 Y.n11 34.3584
R62 Y.n15 Y.n13 34.3584
R63 Y Y.n15 27.7875
R64 Y.n0 Y.t4 26.5955
R65 Y.n0 Y.t3 26.5955
R66 Y.n2 Y.t1 26.5955
R67 Y.n2 Y.t0 26.5955
R68 Y.n4 Y.t6 26.5955
R69 Y.n4 Y.t5 26.5955
R70 Y.n6 Y.t2 26.5955
R71 Y.n6 Y.t7 26.5955
R72 Y.n9 Y 25.611
R73 Y.n8 Y.t8 24.9236
R74 Y.n8 Y.t12 24.9236
R75 Y.n10 Y.t13 24.9236
R76 Y.n10 Y.t9 24.9236
R77 Y.n12 Y.t14 24.9236
R78 Y.n12 Y.t10 24.9236
R79 Y.n14 Y.t15 24.9236
R80 Y.n14 Y.t11 24.9236
R81 VPWR.n7 VPWR.t3 345.505
R82 VPWR.n17 VPWR.t4 342.375
R83 VPWR.n2 VPWR.n1 320.976
R84 VPWR.n10 VPWR.n4 320.976
R85 VPWR.n6 VPWR.n5 320.976
R86 VPWR.n12 VPWR.n11 34.6358
R87 VPWR.n16 VPWR.n15 34.6358
R88 VPWR.n10 VPWR.n9 32.0005
R89 VPWR.n9 VPWR.n6 31.2476
R90 VPWR.n1 VPWR.t6 26.5955
R91 VPWR.n1 VPWR.t5 26.5955
R92 VPWR.n4 VPWR.t0 26.5955
R93 VPWR.n4 VPWR.t7 26.5955
R94 VPWR.n5 VPWR.t2 26.5955
R95 VPWR.n5 VPWR.t1 26.5955
R96 VPWR.n12 VPWR.n2 25.977
R97 VPWR.n17 VPWR.n16 13.5534
R98 VPWR.n18 VPWR.n17 11.1829
R99 VPWR.n7 VPWR.n6 10.5481
R100 VPWR.n9 VPWR.n8 9.3005
R101 VPWR.n11 VPWR.n3 9.3005
R102 VPWR.n13 VPWR.n12 9.3005
R103 VPWR.n15 VPWR.n14 9.3005
R104 VPWR.n16 VPWR.n0 9.3005
R105 VPWR.n15 VPWR.n2 8.65932
R106 VPWR.n11 VPWR.n10 2.63579
R107 VPWR.n8 VPWR.n7 0.567773
R108 VPWR.n8 VPWR.n3 0.120292
R109 VPWR.n13 VPWR.n3 0.120292
R110 VPWR.n14 VPWR.n13 0.120292
R111 VPWR.n14 VPWR.n0 0.120292
R112 VPWR.n18 VPWR.n0 0.120292
R113 VPWR VPWR.n18 0.0226354
R114 VPB VPB.t4 290.031
R115 VPB.t2 VPB.t3 248.599
R116 VPB.t1 VPB.t2 248.599
R117 VPB.t0 VPB.t1 248.599
R118 VPB.t7 VPB.t0 248.599
R119 VPB.t6 VPB.t7 248.599
R120 VPB.t5 VPB.t6 248.599
R121 VPB.t4 VPB.t5 248.599
R122 VGND.n7 VGND.t0 290.637
R123 VGND.n17 VGND.t5 287.151
R124 VGND.n6 VGND.n5 207.213
R125 VGND.n10 VGND.n4 207.213
R126 VGND.n2 VGND.n1 207.213
R127 VGND.n12 VGND.n11 34.6358
R128 VGND.n16 VGND.n15 34.6358
R129 VGND.n10 VGND.n9 32.0005
R130 VGND.n9 VGND.n6 31.2476
R131 VGND.n12 VGND.n2 25.977
R132 VGND.n5 VGND.t6 24.9236
R133 VGND.n5 VGND.t1 24.9236
R134 VGND.n4 VGND.t7 24.9236
R135 VGND.n4 VGND.t2 24.9236
R136 VGND.n1 VGND.t4 24.9236
R137 VGND.n1 VGND.t3 24.9236
R138 VGND.n17 VGND.n16 13.5534
R139 VGND.n18 VGND.n17 11.1829
R140 VGND.n7 VGND.n6 10.5481
R141 VGND.n9 VGND.n8 9.3005
R142 VGND.n11 VGND.n3 9.3005
R143 VGND.n13 VGND.n12 9.3005
R144 VGND.n15 VGND.n14 9.3005
R145 VGND.n16 VGND.n0 9.3005
R146 VGND.n15 VGND.n2 8.65932
R147 VGND.n11 VGND.n10 2.63579
R148 VGND.n8 VGND.n7 0.567773
R149 VGND.n8 VGND.n3 0.120292
R150 VGND.n13 VGND.n3 0.120292
R151 VGND.n14 VGND.n13 0.120292
R152 VGND.n14 VGND.n0 0.120292
R153 VGND.n18 VGND.n0 0.120292
R154 VGND VGND.n18 0.0226354
R155 VNB VNB.t5 1395.47
R156 VNB.t6 VNB.t0 1196.12
R157 VNB.t1 VNB.t6 1196.12
R158 VNB.t7 VNB.t1 1196.12
R159 VNB.t2 VNB.t7 1196.12
R160 VNB.t4 VNB.t2 1196.12
R161 VNB.t3 VNB.t4 1196.12
R162 VNB.t5 VNB.t3 1196.12
C0 Y VPB 0.034787f
C1 VPWR A 0.127577f
C2 Y VGND 0.574497f
C3 VPB VPWR 0.100209f
C4 VGND VPWR 0.085433f
C5 Y VPWR 0.779949f
C6 VPB A 0.254088f
C7 VGND A 0.116857f
C8 VPB VGND 0.007925f
C9 Y A 0.829319f
C10 VGND VNB 0.51049f
C11 Y VNB 0.126735f
C12 VPWR VNB 0.449913f
C13 A VNB 0.771261f
C14 VPB VNB 0.870552f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 Y.t15 A.t0 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t9 A.t1 Y.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t15 A.t2 Y.t25 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t13 A.t3 VPWR.t8 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t14 A.t4 Y.t18 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t13 A.t5 Y.t17 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t12 A.t6 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t12 A.t7 Y.t16 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t6 A.t8 Y.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t24 A.t9 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR.t15 A.t10 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y.t23 A.t11 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y.t9 A.t12 VPWR.t14 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR.t13 A.t13 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t7 A.t14 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t9 A.t15 Y.t22 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y.t21 A.t16 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND.t7 A.t17 Y.t20 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t6 A.t18 Y.t19 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y.t6 A.t19 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t5 A.t20 Y.t28 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t5 A.t21 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t2 A.t22 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t1 A.t23 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t0 A.t24 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t27 A.t25 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y.t1 A.t26 VPWR.t12 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t26 A.t27 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y.t31 A.t28 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t30 A.t29 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR.t11 A.t30 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y.t29 A.t31 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n2 A.t1 212.081
R1 A.n3 A.t3 212.081
R2 A.n4 A.t8 212.081
R3 A.n5 A.t14 212.081
R4 A.n6 A.t22 212.081
R5 A.n1 A.t21 212.081
R6 A.n10 A.t24 212.081
R7 A.n11 A.t26 212.081
R8 A.n25 A.t30 212.081
R9 A.n24 A.t0 212.081
R10 A.n22 A.t10 212.081
R11 A.n21 A.t12 212.081
R12 A.n12 A.t13 212.081
R13 A.n14 A.t19 212.081
R14 A.n16 A.t23 212.081
R15 A.n15 A.t6 212.081
R16 A.n8 A.n7 196.534
R17 A.n15 A.n13 187.055
R18 A.n9 A.n8 152
R19 A.n27 A.n26 152
R20 A.n23 A.n0 152
R21 A.n20 A.n19 152
R22 A.n18 A.n17 152
R23 A.n2 A.t7 139.78
R24 A.n3 A.t11 139.78
R25 A.n4 A.t5 139.78
R26 A.n5 A.t27 139.78
R27 A.n6 A.t2 139.78
R28 A.n1 A.t31 139.78
R29 A.n10 A.t4 139.78
R30 A.n11 A.t29 139.78
R31 A.n25 A.t20 139.78
R32 A.n24 A.t28 139.78
R33 A.n22 A.t18 139.78
R34 A.n21 A.t25 139.78
R35 A.n12 A.t17 139.78
R36 A.n14 A.t9 139.78
R37 A.n16 A.t15 139.78
R38 A.n15 A.t16 139.78
R39 A.n3 A.n2 61.346
R40 A.n4 A.n3 61.346
R41 A.n5 A.n4 61.346
R42 A.n6 A.n1 61.346
R43 A.n11 A.n10 61.346
R44 A.n25 A.n24 61.346
R45 A.n22 A.n21 61.346
R46 A.n14 A.n12 61.346
R47 A.n16 A.n15 61.346
R48 A.n18 A.n13 46.4005
R49 A.n19 A.n0 45.0672
R50 A.n27 A.n0 44.5338
R51 A A.n18 43.7338
R52 A.n7 A.n5 31.4035
R53 A.n23 A.n22 31.4035
R54 A.n9 A.n1 30.6732
R55 A.n10 A.n9 30.6732
R56 A.n26 A.n11 30.6732
R57 A.n26 A.n25 30.6732
R58 A.n21 A.n20 30.6732
R59 A.n20 A.n12 30.6732
R60 A.n17 A.n14 30.6732
R61 A.n17 A.n16 30.6732
R62 A.n7 A.n6 29.9429
R63 A.n24 A.n23 29.9429
R64 A.n8 A 12.8005
R65 A.n13 A 8.0005
R66 A A.n27 7.46717
R67 A.n19 A 1.06717
R68 VPWR.n14 VPWR.t9 354.187
R69 VPWR.n2 VPWR.n1 320.976
R70 VPWR.n33 VPWR.n4 320.976
R71 VPWR.n6 VPWR.n5 320.976
R72 VPWR.n26 VPWR.n8 320.976
R73 VPWR.n20 VPWR.n19 320.976
R74 VPWR.n17 VPWR.n11 320.976
R75 VPWR.n13 VPWR.n12 320.976
R76 VPWR.n39 VPWR.t7 255.965
R77 VPWR.n21 VPWR.n18 34.6358
R78 VPWR.n25 VPWR.n9 34.6358
R79 VPWR.n28 VPWR.n27 34.6358
R80 VPWR.n32 VPWR.n31 34.6358
R81 VPWR.n38 VPWR.n37 34.6358
R82 VPWR.n16 VPWR.n13 34.2593
R83 VPWR.n34 VPWR.n2 33.5064
R84 VPWR.n34 VPWR.n33 29.7417
R85 VPWR.n17 VPWR.n16 28.9887
R86 VPWR.n1 VPWR.t4 26.5955
R87 VPWR.n1 VPWR.t1 26.5955
R88 VPWR.n4 VPWR.t14 26.5955
R89 VPWR.n4 VPWR.t13 26.5955
R90 VPWR.n5 VPWR.t10 26.5955
R91 VPWR.n5 VPWR.t15 26.5955
R92 VPWR.n8 VPWR.t12 26.5955
R93 VPWR.n8 VPWR.t11 26.5955
R94 VPWR.n19 VPWR.t3 26.5955
R95 VPWR.n19 VPWR.t0 26.5955
R96 VPWR.n11 VPWR.t5 26.5955
R97 VPWR.n11 VPWR.t2 26.5955
R98 VPWR.n12 VPWR.t8 26.5955
R99 VPWR.n12 VPWR.t6 26.5955
R100 VPWR.n31 VPWR.n6 23.7181
R101 VPWR.n21 VPWR.n20 22.9652
R102 VPWR.n39 VPWR.n38 21.0829
R103 VPWR.n27 VPWR.n26 17.6946
R104 VPWR.n26 VPWR.n25 16.9417
R105 VPWR.n20 VPWR.n9 11.6711
R106 VPWR.n28 VPWR.n6 10.9181
R107 VPWR.n16 VPWR.n15 9.3005
R108 VPWR.n18 VPWR.n10 9.3005
R109 VPWR.n22 VPWR.n21 9.3005
R110 VPWR.n23 VPWR.n9 9.3005
R111 VPWR.n25 VPWR.n24 9.3005
R112 VPWR.n27 VPWR.n7 9.3005
R113 VPWR.n29 VPWR.n28 9.3005
R114 VPWR.n31 VPWR.n30 9.3005
R115 VPWR.n32 VPWR.n3 9.3005
R116 VPWR.n35 VPWR.n34 9.3005
R117 VPWR.n37 VPWR.n36 9.3005
R118 VPWR.n38 VPWR.n0 9.3005
R119 VPWR.n40 VPWR.n39 9.3005
R120 VPWR.n14 VPWR.n13 7.57496
R121 VPWR.n18 VPWR.n17 5.64756
R122 VPWR.n33 VPWR.n32 4.89462
R123 VPWR.n37 VPWR.n2 1.12991
R124 VPWR.n15 VPWR.n14 0.534819
R125 VPWR.n15 VPWR.n10 0.120292
R126 VPWR.n22 VPWR.n10 0.120292
R127 VPWR.n23 VPWR.n22 0.120292
R128 VPWR.n24 VPWR.n23 0.120292
R129 VPWR.n24 VPWR.n7 0.120292
R130 VPWR.n29 VPWR.n7 0.120292
R131 VPWR.n30 VPWR.n29 0.120292
R132 VPWR.n30 VPWR.n3 0.120292
R133 VPWR.n35 VPWR.n3 0.120292
R134 VPWR.n36 VPWR.n35 0.120292
R135 VPWR.n36 VPWR.n0 0.120292
R136 VPWR.n40 VPWR.n0 0.120292
R137 VPWR VPWR.n40 0.0226354
R138 Y.n15 Y.n13 243.458
R139 Y.n15 Y.n14 205.059
R140 Y.n17 Y.n16 205.059
R141 Y.n19 Y.n18 205.059
R142 Y.n21 Y.n20 205.059
R143 Y.n23 Y.n22 205.059
R144 Y.n25 Y.n24 205.059
R145 Y.n27 Y.n26 205.059
R146 Y.n2 Y.n0 133.534
R147 Y.n2 Y.n1 99.1759
R148 Y.n4 Y.n3 99.1759
R149 Y.n6 Y.n5 99.1759
R150 Y.n8 Y.n7 99.1759
R151 Y.n10 Y.n9 99.1759
R152 Y.n12 Y.n11 99.1759
R153 Y Y.n29 97.4305
R154 Y.n17 Y.n15 38.4005
R155 Y.n19 Y.n17 38.4005
R156 Y.n21 Y.n19 38.4005
R157 Y.n23 Y.n21 38.4005
R158 Y.n25 Y.n23 38.4005
R159 Y.n27 Y.n25 38.4005
R160 Y.n4 Y.n2 34.3584
R161 Y.n6 Y.n4 34.3584
R162 Y.n8 Y.n6 34.3584
R163 Y.n10 Y.n8 34.3584
R164 Y.n12 Y.n10 34.3584
R165 Y.n28 Y.n12 34.3584
R166 Y.n26 Y.t14 26.5955
R167 Y.n26 Y.t13 26.5955
R168 Y.n13 Y.t3 26.5955
R169 Y.n13 Y.t12 26.5955
R170 Y.n14 Y.t8 26.5955
R171 Y.n14 Y.t6 26.5955
R172 Y.n16 Y.t10 26.5955
R173 Y.n16 Y.t9 26.5955
R174 Y.n18 Y.t0 26.5955
R175 Y.n18 Y.t15 26.5955
R176 Y.n20 Y.t2 26.5955
R177 Y.n20 Y.t1 26.5955
R178 Y.n22 Y.t4 26.5955
R179 Y.n22 Y.t5 26.5955
R180 Y.n24 Y.t11 26.5955
R181 Y.n24 Y.t7 26.5955
R182 Y.n29 Y.t16 24.9236
R183 Y.n29 Y.t23 24.9236
R184 Y.n0 Y.t22 24.9236
R185 Y.n0 Y.t21 24.9236
R186 Y.n1 Y.t20 24.9236
R187 Y.n1 Y.t24 24.9236
R188 Y.n3 Y.t19 24.9236
R189 Y.n3 Y.t27 24.9236
R190 Y.n5 Y.t28 24.9236
R191 Y.n5 Y.t31 24.9236
R192 Y.n7 Y.t18 24.9236
R193 Y.n7 Y.t30 24.9236
R194 Y.n9 Y.t25 24.9236
R195 Y.n9 Y.t29 24.9236
R196 Y.n11 Y.t17 24.9236
R197 Y.n11 Y.t26 24.9236
R198 Y Y.n27 18.4247
R199 Y.n28 Y 11.4429
R200 Y Y.n28 1.74595
R201 VPB.t13 VPB.t14 248.599
R202 VPB.t11 VPB.t13 248.599
R203 VPB.t7 VPB.t11 248.599
R204 VPB.t4 VPB.t7 248.599
R205 VPB.t5 VPB.t4 248.599
R206 VPB.t2 VPB.t5 248.599
R207 VPB.t1 VPB.t2 248.599
R208 VPB.t0 VPB.t1 248.599
R209 VPB.t15 VPB.t0 248.599
R210 VPB.t10 VPB.t15 248.599
R211 VPB.t9 VPB.t10 248.599
R212 VPB.t8 VPB.t9 248.599
R213 VPB.t6 VPB.t8 248.599
R214 VPB.t3 VPB.t6 248.599
R215 VPB.t12 VPB.t3 248.599
R216 VPB VPB.t12 230.841
R217 VGND.n13 VGND.n12 207.213
R218 VGND.n17 VGND.n11 207.213
R219 VGND.n20 VGND.n19 207.213
R220 VGND.n26 VGND.n8 207.213
R221 VGND.n6 VGND.n5 207.213
R222 VGND.n33 VGND.n4 207.213
R223 VGND.n2 VGND.n1 207.213
R224 VGND.n14 VGND.t12 166.852
R225 VGND.n39 VGND.t8 157.567
R226 VGND.n21 VGND.n18 34.6358
R227 VGND.n25 VGND.n9 34.6358
R228 VGND.n28 VGND.n27 34.6358
R229 VGND.n32 VGND.n31 34.6358
R230 VGND.n38 VGND.n37 34.6358
R231 VGND.n16 VGND.n13 34.2593
R232 VGND.n34 VGND.n2 33.5064
R233 VGND.n34 VGND.n33 29.7417
R234 VGND.n17 VGND.n16 28.9887
R235 VGND.n12 VGND.t10 24.9236
R236 VGND.n12 VGND.t13 24.9236
R237 VGND.n11 VGND.t3 24.9236
R238 VGND.n11 VGND.t15 24.9236
R239 VGND.n19 VGND.t0 24.9236
R240 VGND.n19 VGND.t14 24.9236
R241 VGND.n8 VGND.t1 24.9236
R242 VGND.n8 VGND.t5 24.9236
R243 VGND.n5 VGND.t2 24.9236
R244 VGND.n5 VGND.t6 24.9236
R245 VGND.n4 VGND.t4 24.9236
R246 VGND.n4 VGND.t7 24.9236
R247 VGND.n1 VGND.t11 24.9236
R248 VGND.n1 VGND.t9 24.9236
R249 VGND.n31 VGND.n6 23.7181
R250 VGND.n21 VGND.n20 22.9652
R251 VGND.n39 VGND.n38 21.0829
R252 VGND.n27 VGND.n26 17.6946
R253 VGND.n26 VGND.n25 16.9417
R254 VGND.n20 VGND.n9 11.6711
R255 VGND.n28 VGND.n6 10.9181
R256 VGND.n40 VGND.n39 9.3005
R257 VGND.n16 VGND.n15 9.3005
R258 VGND.n18 VGND.n10 9.3005
R259 VGND.n22 VGND.n21 9.3005
R260 VGND.n23 VGND.n9 9.3005
R261 VGND.n25 VGND.n24 9.3005
R262 VGND.n27 VGND.n7 9.3005
R263 VGND.n29 VGND.n28 9.3005
R264 VGND.n31 VGND.n30 9.3005
R265 VGND.n32 VGND.n3 9.3005
R266 VGND.n35 VGND.n34 9.3005
R267 VGND.n37 VGND.n36 9.3005
R268 VGND.n38 VGND.n0 9.3005
R269 VGND.n14 VGND.n13 7.57496
R270 VGND.n18 VGND.n17 5.64756
R271 VGND.n33 VGND.n32 4.89462
R272 VGND.n37 VGND.n2 1.12991
R273 VGND.n15 VGND.n14 0.534819
R274 VGND.n15 VGND.n10 0.120292
R275 VGND.n22 VGND.n10 0.120292
R276 VGND.n23 VGND.n22 0.120292
R277 VGND.n24 VGND.n23 0.120292
R278 VGND.n24 VGND.n7 0.120292
R279 VGND.n29 VGND.n7 0.120292
R280 VGND.n30 VGND.n29 0.120292
R281 VGND.n30 VGND.n3 0.120292
R282 VGND.n35 VGND.n3 0.120292
R283 VGND.n36 VGND.n35 0.120292
R284 VGND.n36 VGND.n0 0.120292
R285 VGND.n40 VGND.n0 0.120292
R286 VGND VGND.n40 0.0226354
R287 VNB.t10 VNB.t12 1196.12
R288 VNB.t13 VNB.t10 1196.12
R289 VNB.t3 VNB.t13 1196.12
R290 VNB.t15 VNB.t3 1196.12
R291 VNB.t0 VNB.t15 1196.12
R292 VNB.t14 VNB.t0 1196.12
R293 VNB.t1 VNB.t14 1196.12
R294 VNB.t5 VNB.t1 1196.12
R295 VNB.t2 VNB.t5 1196.12
R296 VNB.t6 VNB.t2 1196.12
R297 VNB.t4 VNB.t6 1196.12
R298 VNB.t7 VNB.t4 1196.12
R299 VNB.t11 VNB.t7 1196.12
R300 VNB.t9 VNB.t11 1196.12
R301 VNB.t8 VNB.t9 1196.12
R302 VNB VNB.t8 1110.68
C0 VGND VPWR 0.160762f
C1 VGND Y 1.06261f
C2 A VPB 0.525745f
C3 VPWR VPB 0.159316f
C4 Y VPB 0.03049f
C5 VPWR A 0.280261f
C6 Y A 1.4347f
C7 VGND VPB 0.013189f
C8 Y VPWR 1.46621f
C9 VGND A 0.265874f
C10 VGND VNB 0.864536f
C11 Y VNB 0.055057f
C12 VPWR VNB 0.737072f
C13 A VNB 1.54575f
C14 VPB VNB 1.49072f
.ends


* NGSPICE file created from sky130_fd_sc_hd__or4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4bb_4 VNB VPB VGND VPWR B A X C_N D_N
X0 VPWR.t6 a_315_380.t5 X.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t2 a_315_380.t6 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2 a_315_380.t4 B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t9 C_N.t0 a_27_410.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR.t0 C_N.t1 a_27_410.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR.t2 A.t0 a_583_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t8 a_27_410.t2 a_315_380.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X7 a_583_297.t1 B.t1 a_499_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t3 A.t1 a_315_380.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_397_297.t0 a_205_93.t2 a_315_380.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.257925 ps=2.52 w=1 l=0.15
X10 X.t5 a_315_380.t7 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X.t4 a_315_380.t8 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_499_297.t0 a_27_410.t3 a_397_297.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X13 VPWR.t4 a_315_380.t9 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_205_93.t1 D_N.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X15 a_205_93.t0 D_N.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.11295 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X16 VGND.t5 a_315_380.t10 X.t7 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t4 a_315_380.t11 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_315_380.t1 a_205_93.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X19 X.t0 a_315_380.t12 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 a_315_380.n15 a_315_380.n14 707.908
R1 a_315_380.n4 a_315_380.t9 212.081
R2 a_315_380.n3 a_315_380.t12 212.081
R3 a_315_380.n8 a_315_380.t5 212.081
R4 a_315_380.n10 a_315_380.t6 212.081
R5 a_315_380.n14 a_315_380.n0 197.424
R6 a_315_380.n13 a_315_380.n1 197.424
R7 a_315_380.n6 a_315_380.n5 177.601
R8 a_315_380.n16 a_315_380.n15 162.236
R9 a_315_380.n12 a_315_380.n11 152
R10 a_315_380.n9 a_315_380.n2 152
R11 a_315_380.n7 a_315_380.n6 152
R12 a_315_380.n4 a_315_380.t11 139.78
R13 a_315_380.n3 a_315_380.t8 139.78
R14 a_315_380.n8 a_315_380.t10 139.78
R15 a_315_380.n10 a_315_380.t7 139.78
R16 a_315_380.n13 a_315_380.n12 79.0593
R17 a_315_380.n14 a_315_380.n13 65.5064
R18 a_315_380.n11 a_315_380.n9 49.6611
R19 a_315_380.n8 a_315_380.n7 46.7399
R20 a_315_380.n0 a_315_380.t1 39.6928
R21 a_315_380.n5 a_315_380.n3 35.055
R22 a_315_380.n0 a_315_380.t3 30.462
R23 a_315_380.n5 a_315_380.n4 26.2914
R24 a_315_380.n15 a_315_380.t0 26.2672
R25 a_315_380.n6 a_315_380.n2 25.6005
R26 a_315_380.n12 a_315_380.n2 25.6005
R27 a_315_380.n1 a_315_380.t2 24.9236
R28 a_315_380.n1 a_315_380.t4 24.9236
R29 a_315_380.n7 a_315_380.n3 14.6066
R30 a_315_380.n11 a_315_380.n10 8.76414
R31 a_315_380.n9 a_315_380.n8 2.92171
R32 X.n5 X.n3 252.931
R33 X.n2 X.n0 238.163
R34 X.n5 X.n4 208.507
R35 X.n2 X.n1 98.982
R36 X.n6 X.n5 58.4189
R37 X.n3 X.t3 26.5955
R38 X.n3 X.t2 26.5955
R39 X.n4 X.t1 26.5955
R40 X.n4 X.t0 26.5955
R41 X.n0 X.t7 24.9236
R42 X.n0 X.t5 24.9236
R43 X.n1 X.t6 24.9236
R44 X.n1 X.t4 24.9236
R45 X.n6 X.n2 14.2227
R46 X X.n6 2.78311
R47 VPWR.n19 VPWR.n1 601.679
R48 VPWR.n8 VPWR.t4 351.63
R49 VPWR.n1 VPWR.t1 327.592
R50 VPWR.n11 VPWR.n5 318.293
R51 VPWR.n7 VPWR.n6 318.293
R52 VPWR.n1 VPWR.t0 63.3219
R53 VPWR.n5 VPWR.t5 37.4305
R54 VPWR.n5 VPWR.t2 37.4305
R55 VPWR.n13 VPWR.n12 34.6358
R56 VPWR.n13 VPWR.n2 34.6358
R57 VPWR.n17 VPWR.n2 34.6358
R58 VPWR.n18 VPWR.n17 34.6358
R59 VPWR.n12 VPWR.n11 30.8711
R60 VPWR.n10 VPWR.n7 28.9887
R61 VPWR.n6 VPWR.t3 26.5955
R62 VPWR.n6 VPWR.t6 26.5955
R63 VPWR.n19 VPWR.n18 22.9652
R64 VPWR.n11 VPWR.n10 19.577
R65 VPWR.n10 VPWR.n9 9.3005
R66 VPWR.n11 VPWR.n4 9.3005
R67 VPWR.n12 VPWR.n3 9.3005
R68 VPWR.n14 VPWR.n13 9.3005
R69 VPWR.n15 VPWR.n2 9.3005
R70 VPWR.n17 VPWR.n16 9.3005
R71 VPWR.n18 VPWR.n0 9.3005
R72 VPWR.n20 VPWR.n19 7.12063
R73 VPWR.n8 VPWR.n7 6.48892
R74 VPWR.n9 VPWR.n8 0.663075
R75 VPWR.n20 VPWR.n0 0.148519
R76 VPWR.n9 VPWR.n4 0.120292
R77 VPWR.n4 VPWR.n3 0.120292
R78 VPWR.n14 VPWR.n3 0.120292
R79 VPWR.n15 VPWR.n14 0.120292
R80 VPWR.n16 VPWR.n15 0.120292
R81 VPWR.n16 VPWR.n0 0.120292
R82 VPWR VPWR.n20 0.114842
R83 VPB.t2 VPB.t1 565.265
R84 VPB.t4 VPB.t7 313.707
R85 VPB.t1 VPB.t9 301.87
R86 VPB.t0 VPB.t2 287.072
R87 VPB.t5 VPB.t6 248.599
R88 VPB.t8 VPB.t5 248.599
R89 VPB.t7 VPB.t8 248.599
R90 VPB.t3 VPB.t4 248.599
R91 VPB.t9 VPB.t3 248.599
R92 VPB VPB.t0 192.369
R93 B.n0 B.t1 241.536
R94 B B.n0 183.668
R95 B.n0 B.t0 169.237
R96 VGND.n9 VGND.t4 293.514
R97 VGND.n20 VGND.t0 276.476
R98 VGND.n1 VGND.n0 228.294
R99 VGND.n8 VGND.n7 207.965
R100 VGND.n4 VGND.n3 200.516
R101 VGND.n14 VGND.n13 198.475
R102 VGND.n0 VGND.t9 45.7148
R103 VGND.n13 VGND.t3 43.3851
R104 VGND.n0 VGND.t2 38.5719
R105 VGND.n9 VGND.n8 36.5149
R106 VGND.n12 VGND.n6 34.6358
R107 VGND.n21 VGND.n1 30.8711
R108 VGND.n19 VGND.n4 29.7417
R109 VGND.n15 VGND.n14 27.4829
R110 VGND.n21 VGND.n20 27.4829
R111 VGND.n13 VGND.t7 26.7697
R112 VGND.n7 VGND.t6 24.9236
R113 VGND.n7 VGND.t5 24.9236
R114 VGND.n3 VGND.t1 24.9236
R115 VGND.n3 VGND.t8 24.9236
R116 VGND.n20 VGND.n19 16.9417
R117 VGND.n15 VGND.n4 14.6829
R118 VGND.n14 VGND.n12 13.177
R119 VGND.n23 VGND.n1 11.4238
R120 VGND.n10 VGND.n6 9.3005
R121 VGND.n12 VGND.n11 9.3005
R122 VGND.n14 VGND.n5 9.3005
R123 VGND.n16 VGND.n15 9.3005
R124 VGND.n17 VGND.n4 9.3005
R125 VGND.n19 VGND.n18 9.3005
R126 VGND.n20 VGND.n2 9.3005
R127 VGND.n22 VGND.n21 9.3005
R128 VGND.n8 VGND.n6 3.76521
R129 VGND.n10 VGND.n9 2.15642
R130 VGND.n23 VGND.n22 0.141672
R131 VGND VGND.n23 0.121778
R132 VGND.n11 VGND.n10 0.120292
R133 VGND.n11 VGND.n5 0.120292
R134 VGND.n16 VGND.n5 0.120292
R135 VGND.n17 VGND.n16 0.120292
R136 VGND.n18 VGND.n17 0.120292
R137 VGND.n18 VGND.n2 0.120292
R138 VGND.n22 VGND.n2 0.120292
R139 VNB.t2 VNB.t0 2677.02
R140 VNB.t3 VNB.t7 1509.39
R141 VNB.t0 VNB.t8 1509.39
R142 VNB.t9 VNB.t2 1267.31
R143 VNB.t6 VNB.t4 1196.12
R144 VNB.t5 VNB.t6 1196.12
R145 VNB.t7 VNB.t5 1196.12
R146 VNB.t1 VNB.t3 1196.12
R147 VNB.t8 VNB.t1 1196.12
R148 VNB VNB.t9 1025.24
R149 C_N.n0 C_N.t1 329.902
R150 C_N C_N.n0 153.738
R151 C_N.n0 C_N.t0 132.282
R152 a_27_410.t0 a_27_410.n1 665.061
R153 a_27_410.n1 a_27_410.n0 408.753
R154 a_27_410.n1 a_27_410.t1 312.767
R155 a_27_410.n0 a_27_410.t3 241.536
R156 a_27_410.n0 a_27_410.t2 169.237
R157 A.n0 A.t0 241.536
R158 A A.n0 178.353
R159 A.n0 A.t1 169.237
R160 a_583_297.t0 a_583_297.t1 53.1905
R161 a_499_297.t0 a_499_297.t1 53.1905
R162 a_205_93.n2 a_205_93.n1 636.987
R163 a_205_93.n1 a_205_93.t1 266.481
R164 a_205_93.n0 a_205_93.t2 227.674
R165 a_205_93.n0 a_205_93.t3 155.375
R166 a_205_93.n1 a_205_93.n0 152
R167 a_205_93.n3 a_205_93.n2 59.1005
R168 a_205_93.n2 a_205_93.t0 29.5559
R169 a_397_297.t0 a_397_297.t1 70.9205
R170 D_N D_N.n0 154.429
R171 D_N.n0 D_N.t1 142.994
R172 D_N.n0 D_N.t0 126.927
C0 C_N D_N 0.081313f
C1 VPWR A 0.052577f
C2 VPB B 0.028231f
C3 VPB VGND 0.010456f
C4 X C_N 2.34e-19
C5 D_N B 8.92e-20
C6 D_N VGND 0.018133f
C7 A C_N 5.53e-20
C8 VPWR C_N 0.021171f
C9 X B 0.004605f
C10 X VGND 0.244089f
C11 A B 0.10797f
C12 A VGND 0.018403f
C13 VPWR B 0.082647f
C14 VPB D_N 0.039453f
C15 VPWR VGND 0.110621f
C16 X VPB 0.01233f
C17 C_N B 2.11e-19
C18 C_N VGND 0.031122f
C19 VPB A 0.030992f
C20 VPWR VPB 0.122146f
C21 X D_N 1.03e-19
C22 B VGND 0.017437f
C23 VPWR D_N 0.004101f
C24 VPB C_N 0.093836f
C25 X A 0.015701f
C26 VPWR X 0.357666f
C27 VGND VNB 0.663238f
C28 X VNB 0.058172f
C29 D_N VNB 0.100763f
C30 VPWR VNB 0.542019f
C31 A VNB 0.091075f
C32 B VNB 0.089178f
C33 C_N VNB 0.134167f
C34 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__probe_p_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__probe_p_8 X VPB VNB VGND VPWR A
X0 a_361_47.t10 a_27_47.t6 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_361_47.t9 a_27_47.t7 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_361_47.t8 a_27_47.t8 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t9 a_27_47.t9 a_361_47.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_361_47.t2 a_27_47.t10 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t7 a_27_47.t11 a_361_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t7 a_27_47.t12 a_361_47.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47.t5 A.t1 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_361_47.t0 a_27_47.t13 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47.t1 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_361_47.t6 a_27_47.t14 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t5 a_27_47.t15 a_361_47.t14 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_361_47.t13 a_27_47.t16 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t1 A.t3 a_27_47.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t5 a_27_47.t17 a_361_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t3 a_27_47.t18 a_361_47.t12 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t4 a_27_47.t19 a_361_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t3 a_27_47.t20 a_361_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_361_47.t15 a_27_47.t21 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t1 A.t4 a_27_47.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND.t2 A.t5 a_27_47.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n22 a_27_47.t4 286.348
R1 a_27_47.n24 a_27_47.t3 271.051
R2 a_27_47.n4 a_27_47.t12 221.72
R3 a_27_47.n5 a_27_47.t13 221.72
R4 a_27_47.n3 a_27_47.t15 221.72
R5 a_27_47.n9 a_27_47.t16 221.72
R6 a_27_47.n11 a_27_47.t18 221.72
R7 a_27_47.n1 a_27_47.t21 221.72
R8 a_27_47.n17 a_27_47.t9 221.72
R9 a_27_47.n18 a_27_47.t10 221.72
R10 a_27_47.n25 a_27_47.n24 206.055
R11 a_27_47.n22 a_27_47.n21 198.177
R12 a_27_47.n7 a_27_47.n6 177.601
R13 a_27_47.n20 a_27_47.n19 152
R14 a_27_47.n16 a_27_47.n0 152
R15 a_27_47.n15 a_27_47.n14 152
R16 a_27_47.n13 a_27_47.n12 152
R17 a_27_47.n10 a_27_47.n2 152
R18 a_27_47.n8 a_27_47.n7 152
R19 a_27_47.n4 a_27_47.t11 149.421
R20 a_27_47.n5 a_27_47.t8 149.421
R21 a_27_47.n3 a_27_47.t20 149.421
R22 a_27_47.n9 a_27_47.t7 149.421
R23 a_27_47.n11 a_27_47.t19 149.421
R24 a_27_47.n1 a_27_47.t6 149.421
R25 a_27_47.n17 a_27_47.t17 149.421
R26 a_27_47.n18 a_27_47.t14 149.421
R27 a_27_47.n5 a_27_47.n4 74.9783
R28 a_27_47.n6 a_27_47.n5 66.0523
R29 a_27_47.n16 a_27_47.n15 60.6968
R30 a_27_47.n19 a_27_47.n17 55.3412
R31 a_27_47.n8 a_27_47.n3 51.7709
R32 a_27_47.n12 a_27_47.n1 51.7709
R33 a_27_47.n23 a_27_47.n22 48.9632
R34 a_27_47.n24 a_27_47.n23 38.7339
R35 a_27_47.n10 a_27_47.n9 37.4894
R36 a_27_47.n11 a_27_47.n10 37.4894
R37 a_27_47.t0 a_27_47.n25 26.5955
R38 a_27_47.n25 a_27_47.t5 26.5955
R39 a_27_47.n7 a_27_47.n2 25.6005
R40 a_27_47.n13 a_27_47.n2 25.6005
R41 a_27_47.n14 a_27_47.n13 25.6005
R42 a_27_47.n14 a_27_47.n0 25.6005
R43 a_27_47.n20 a_27_47.n0 25.6005
R44 a_27_47.n21 a_27_47.t2 24.9236
R45 a_27_47.n21 a_27_47.t1 24.9236
R46 a_27_47.n9 a_27_47.n8 23.2079
R47 a_27_47.n12 a_27_47.n11 23.2079
R48 a_27_47.n19 a_27_47.n18 19.6375
R49 a_27_47.n23 a_27_47.n20 18.4476
R50 a_27_47.n6 a_27_47.n3 8.92643
R51 a_27_47.n15 a_27_47.n1 8.92643
R52 a_27_47.n17 a_27_47.n16 5.35606
R53 VGND.n5 VGND.n4 200.516
R54 VGND.n10 VGND.n9 200.516
R55 VGND.n13 VGND.n12 200.516
R56 VGND.n18 VGND.n2 200.516
R57 VGND.n21 VGND.n20 200.516
R58 VGND.n6 VGND.t7 155.156
R59 VGND.n14 VGND.n11 34.6358
R60 VGND.n8 VGND.n5 32.0005
R61 VGND.n18 VGND.n1 28.9887
R62 VGND.n4 VGND.t8 24.9236
R63 VGND.n4 VGND.t3 24.9236
R64 VGND.n9 VGND.t9 24.9236
R65 VGND.n9 VGND.t4 24.9236
R66 VGND.n12 VGND.t10 24.9236
R67 VGND.n12 VGND.t5 24.9236
R68 VGND.n2 VGND.t6 24.9236
R69 VGND.n2 VGND.t1 24.9236
R70 VGND.n20 VGND.t0 24.9236
R71 VGND.n20 VGND.t2 24.9236
R72 VGND.n21 VGND.n19 22.9652
R73 VGND.n19 VGND.n18 15.4358
R74 VGND.n13 VGND.n1 9.41227
R75 VGND.n19 VGND.n0 9.3005
R76 VGND.n18 VGND.n17 9.3005
R77 VGND.n16 VGND.n1 9.3005
R78 VGND.n15 VGND.n14 9.3005
R79 VGND.n11 VGND.n3 9.3005
R80 VGND.n8 VGND.n7 9.3005
R81 VGND.n22 VGND.n21 7.12063
R82 VGND.n10 VGND.n8 6.4005
R83 VGND.n6 VGND.n5 5.79315
R84 VGND.n11 VGND.n10 3.38874
R85 VGND.n7 VGND.n6 0.656787
R86 VGND.n14 VGND.n13 0.376971
R87 VGND.n22 VGND.n0 0.148519
R88 VGND.n7 VGND.n3 0.120292
R89 VGND.n15 VGND.n3 0.120292
R90 VGND.n16 VGND.n15 0.120292
R91 VGND.n17 VGND.n16 0.120292
R92 VGND.n17 VGND.n0 0.120292
R93 VGND VGND.n22 0.11354
R94 a_361_47.n4 a_361_47.n3 374.966
R95 a_361_47.n7 a_361_47.n6 315.985
R96 a_361_47.n5 a_361_47.n1 311.717
R97 a_361_47.n4 a_361_47.n2 311.717
R98 a_361_47.n12 a_361_47.n11 261.425
R99 a_361_47.n9 a_361_47.n8 202.444
R100 a_361_47.n10 a_361_47.n0 198.177
R101 a_361_47.n13 a_361_47.n12 198.177
R102 a_361_47.n5 a_361_47.n4 63.2476
R103 a_361_47.n12 a_361_47.n10 63.2476
R104 a_361_47.n7 a_361_47.n5 50.4476
R105 a_361_47.n10 a_361_47.n9 50.4476
R106 a_361_47.n1 a_361_47.t14 26.5955
R107 a_361_47.n1 a_361_47.t13 26.5955
R108 a_361_47.n2 a_361_47.t12 26.5955
R109 a_361_47.n2 a_361_47.t15 26.5955
R110 a_361_47.n3 a_361_47.t11 26.5955
R111 a_361_47.n3 a_361_47.t2 26.5955
R112 a_361_47.n6 a_361_47.t1 26.5955
R113 a_361_47.n6 a_361_47.t0 26.5955
R114 a_361_47.n8 a_361_47.t7 24.9236
R115 a_361_47.n8 a_361_47.t8 24.9236
R116 a_361_47.n11 a_361_47.t5 24.9236
R117 a_361_47.n11 a_361_47.t6 24.9236
R118 a_361_47.n0 a_361_47.t3 24.9236
R119 a_361_47.n0 a_361_47.t9 24.9236
R120 a_361_47.n13 a_361_47.t4 24.9236
R121 a_361_47.t10 a_361_47.n13 24.9236
R122 a_361_47.n9 a_361_47.n7 22.5887
R123 VNB.t8 VNB.t7 1196.12
R124 VNB.t3 VNB.t8 1196.12
R125 VNB.t9 VNB.t3 1196.12
R126 VNB.t4 VNB.t9 1196.12
R127 VNB.t10 VNB.t4 1196.12
R128 VNB.t5 VNB.t10 1196.12
R129 VNB.t6 VNB.t5 1196.12
R130 VNB.t1 VNB.t6 1196.12
R131 VNB.t0 VNB.t1 1196.12
R132 VNB.t2 VNB.t0 1196.12
R133 VNB VNB.t2 911.327
R134 VPWR.n3 VPWR.n2 320.976
R135 VPWR.n24 VPWR.n1 320.976
R136 VPWR.n17 VPWR.n5 310.502
R137 VPWR.n11 VPWR.n10 310.502
R138 VPWR.n9 VPWR.n8 310.502
R139 VPWR.n7 VPWR.t7 248.906
R140 VPWR.n25 VPWR.n24 43.1829
R141 VPWR.n19 VPWR.n18 34.6358
R142 VPWR.n23 VPWR.n22 34.6358
R143 VPWR.n16 VPWR.n6 34.6358
R144 VPWR.n12 VPWR.n9 32.0005
R145 VPWR.n22 VPWR.n3 27.8593
R146 VPWR.n1 VPWR.t10 26.5955
R147 VPWR.n1 VPWR.t1 26.5955
R148 VPWR.n2 VPWR.t8 26.5955
R149 VPWR.n2 VPWR.t0 26.5955
R150 VPWR.n5 VPWR.t2 26.5955
R151 VPWR.n5 VPWR.t9 26.5955
R152 VPWR.n10 VPWR.t4 26.5955
R153 VPWR.n10 VPWR.t3 26.5955
R154 VPWR.n8 VPWR.t6 26.5955
R155 VPWR.n8 VPWR.t5 26.5955
R156 VPWR.n18 VPWR.n17 9.41227
R157 VPWR.n13 VPWR.n12 9.3005
R158 VPWR.n14 VPWR.n6 9.3005
R159 VPWR.n16 VPWR.n15 9.3005
R160 VPWR.n18 VPWR.n4 9.3005
R161 VPWR.n20 VPWR.n19 9.3005
R162 VPWR.n22 VPWR.n21 9.3005
R163 VPWR.n23 VPWR.n0 9.3005
R164 VPWR.n19 VPWR.n3 6.77697
R165 VPWR.n12 VPWR.n11 6.4005
R166 VPWR.n9 VPWR.n7 5.7932
R167 VPWR.n11 VPWR.n6 3.38874
R168 VPWR.n24 VPWR.n23 0.753441
R169 VPWR.n13 VPWR.n7 0.656729
R170 VPWR.n17 VPWR.n16 0.376971
R171 VPWR.n14 VPWR.n13 0.120292
R172 VPWR.n15 VPWR.n14 0.120292
R173 VPWR.n15 VPWR.n4 0.120292
R174 VPWR.n20 VPWR.n4 0.120292
R175 VPWR.n21 VPWR.n20 0.120292
R176 VPWR.n21 VPWR.n0 0.120292
R177 VPWR.n25 VPWR.n0 0.120292
R178 VPWR VPWR.n25 0.0213333
R179 VPB.t6 VPB.t7 248.599
R180 VPB.t5 VPB.t6 248.599
R181 VPB.t4 VPB.t5 248.599
R182 VPB.t3 VPB.t4 248.599
R183 VPB.t2 VPB.t3 248.599
R184 VPB.t9 VPB.t2 248.599
R185 VPB.t8 VPB.t9 248.599
R186 VPB.t0 VPB.t8 248.599
R187 VPB.t10 VPB.t0 248.599
R188 VPB.t1 VPB.t10 248.599
R189 VPB VPB.t1 189.409
R190 A.n6 A.t4 235.763
R191 A.n1 A.t0 221.72
R192 A.n0 A.t1 221.72
R193 A.n6 A.t5 163.464
R194 A.n3 A.n2 152
R195 A.n5 A.n4 152
R196 A.n7 A.n6 152
R197 A.n1 A.t3 149.421
R198 A.n0 A.t2 149.421
R199 A.n2 A.n1 58.019
R200 A.n5 A.n0 43.7375
R201 A.n4 A.n3 21.7605
R202 A.n7 A 19.5205
R203 A.n6 A.n5 17.8524
R204 A.n2 A.n0 16.9598
R205 A A.n7 9.9205
R206 A.n3 A 5.4405
R207 A.n4 A 2.2405
C0 VPWR X 0.012948f
C1 A X 5.06e-19
C2 VPWR m5_250_389# 9e-20
C3 A VPWR 0.049241f
C4 VPB VGND 0.012473f
C5 A m5_250_389# 8.69e-21
C6 VPB X 6.1e-19
C7 X VGND 6.03e-19
C8 VPWR VPB 0.129645f
C9 VPB m5_250_389# 1.45e-20
C10 A VPB 0.099483f
C11 VPWR VGND 0.093265f
C12 VGND m5_250_389# 1.45e-20
C13 A VGND 0.05431f
C14 X VNB 0.124247f
C15 VGND VNB 0.652926f
C16 VPWR VNB 0.553449f
C17 A VNB 0.321526f
C18 VPB VNB 1.13634f
C19 m5_250_389# VNB 3.44e-19 $ **FLOATING
.ends

* NGSPICE file created from sky130_fd_sc_hd__probec_p_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__probec_p_8 X VPB VNB VGND VPWR A
X0 a_361_47.t7 a_27_47.t6 VGND.t4 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 VPWR m5_872_595# sky130_fd_pr__res_generic_m5 w=0 l=1.2
X1 a_361_47.t6 a_27_47.t7 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_361_47.t5 a_27_47.t8 VGND.t10 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t10 a_27_47.t9 a_361_47.t9 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R1 VGND m5_872_n71# sky130_fd_pr__res_generic_m5 w=0 l=1.2
X4 a_361_47.t8 a_27_47.t10 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t9 a_27_47.t11 a_361_47.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t1 A.t0 a_27_47.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t8 a_27_47.t12 a_361_47.t12 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47.t5 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_361_47.t11 a_27_47.t13 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47.t4 A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_361_47.t3 a_27_47.t14 VGND.t8 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t6 a_27_47.t15 a_361_47.t10 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_361_47.t15 a_27_47.t16 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t0 A.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t7 a_27_47.t17 a_361_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t4 a_27_47.t18 a_361_47.t14 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t6 a_27_47.t19 a_361_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t5 a_27_47.t20 a_361_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_361_47.t13 a_27_47.t21 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t0 A.t4 a_27_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND.t1 A.t5 a_27_47.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R2 a_27_47.n22 a_27_47.t2 286.348
R3 a_27_47.t1 a_27_47.n25 271.051
R4 a_27_47.n4 a_27_47.t12 221.72
R5 a_27_47.n5 a_27_47.t13 221.72
R6 a_27_47.n3 a_27_47.t15 221.72
R7 a_27_47.n9 a_27_47.t16 221.72
R8 a_27_47.n11 a_27_47.t18 221.72
R9 a_27_47.n1 a_27_47.t21 221.72
R10 a_27_47.n17 a_27_47.t9 221.72
R11 a_27_47.n18 a_27_47.t10 221.72
R12 a_27_47.n25 a_27_47.n24 206.056
R13 a_27_47.n22 a_27_47.n21 198.177
R14 a_27_47.n7 a_27_47.n6 177.601
R15 a_27_47.n20 a_27_47.n19 152
R16 a_27_47.n16 a_27_47.n0 152
R17 a_27_47.n15 a_27_47.n14 152
R18 a_27_47.n13 a_27_47.n12 152
R19 a_27_47.n10 a_27_47.n2 152
R20 a_27_47.n8 a_27_47.n7 152
R21 a_27_47.n4 a_27_47.t11 149.421
R22 a_27_47.n5 a_27_47.t8 149.421
R23 a_27_47.n3 a_27_47.t20 149.421
R24 a_27_47.n9 a_27_47.t7 149.421
R25 a_27_47.n11 a_27_47.t19 149.421
R26 a_27_47.n1 a_27_47.t6 149.421
R27 a_27_47.n17 a_27_47.t17 149.421
R28 a_27_47.n18 a_27_47.t14 149.421
R29 a_27_47.n5 a_27_47.n4 74.9783
R30 a_27_47.n6 a_27_47.n5 66.0523
R31 a_27_47.n16 a_27_47.n15 60.6968
R32 a_27_47.n19 a_27_47.n17 55.3412
R33 a_27_47.n8 a_27_47.n3 51.7709
R34 a_27_47.n12 a_27_47.n1 51.7709
R35 a_27_47.n23 a_27_47.n22 48.9632
R36 a_27_47.n25 a_27_47.n23 38.7339
R37 a_27_47.n10 a_27_47.n9 37.4894
R38 a_27_47.n11 a_27_47.n10 37.4894
R39 a_27_47.n24 a_27_47.t3 26.5955
R40 a_27_47.n24 a_27_47.t5 26.5955
R41 a_27_47.n7 a_27_47.n2 25.6005
R42 a_27_47.n13 a_27_47.n2 25.6005
R43 a_27_47.n14 a_27_47.n13 25.6005
R44 a_27_47.n14 a_27_47.n0 25.6005
R45 a_27_47.n20 a_27_47.n0 25.6005
R46 a_27_47.n21 a_27_47.t0 24.9236
R47 a_27_47.n21 a_27_47.t4 24.9236
R48 a_27_47.n9 a_27_47.n8 23.2079
R49 a_27_47.n12 a_27_47.n11 23.2079
R50 a_27_47.n19 a_27_47.n18 19.6375
R51 a_27_47.n23 a_27_47.n20 18.4476
R52 a_27_47.n6 a_27_47.n3 8.92643
R53 a_27_47.n15 a_27_47.n1 8.92643
R54 a_27_47.n17 a_27_47.n16 5.35606
R55 VGND.n5 VGND.n4 200.516
R56 VGND.n10 VGND.n9 200.516
R57 VGND.n13 VGND.n12 200.516
R58 VGND.n18 VGND.n2 200.516
R59 VGND.n21 VGND.n20 200.516
R60 VGND.n6 VGND.t9 155.156
R61 VGND.n14 VGND.n11 34.6358
R62 VGND.n8 VGND.n5 32.0005
R63 VGND.n18 VGND.n1 28.9887
R64 VGND.n4 VGND.t10 24.9236
R65 VGND.n4 VGND.t5 24.9236
R66 VGND.n9 VGND.t3 24.9236
R67 VGND.n9 VGND.t6 24.9236
R68 VGND.n12 VGND.t4 24.9236
R69 VGND.n12 VGND.t7 24.9236
R70 VGND.n2 VGND.t8 24.9236
R71 VGND.n2 VGND.t0 24.9236
R72 VGND.n20 VGND.t2 24.9236
R73 VGND.n20 VGND.t1 24.9236
R74 VGND.n21 VGND.n19 22.9652
R75 VGND.n19 VGND.n18 15.4358
R76 VGND.n13 VGND.n1 9.41227
R77 VGND.n19 VGND.n0 9.3005
R78 VGND.n18 VGND.n17 9.3005
R79 VGND.n16 VGND.n1 9.3005
R80 VGND.n15 VGND.n14 9.3005
R81 VGND.n11 VGND.n3 9.3005
R82 VGND.n8 VGND.n7 9.3005
R83 VGND.n22 VGND.n21 7.12063
R84 VGND.n10 VGND.n8 6.4005
R85 VGND.n6 VGND.n5 5.79315
R86 VGND.n11 VGND.n10 3.38874
R87 VGND.n7 VGND.n6 0.656787
R88 VGND.n14 VGND.n13 0.376971
R89 VGND.n22 VGND.n0 0.148519
R90 VGND.n7 VGND.n3 0.120292
R91 VGND.n15 VGND.n3 0.120292
R92 VGND.n16 VGND.n15 0.120292
R93 VGND.n17 VGND.n16 0.120292
R94 VGND.n17 VGND.n0 0.120292
R95 VGND VGND.n22 0.11354
R96 a_361_47.n4 a_361_47.n3 374.966
R97 a_361_47.n7 a_361_47.n6 315.985
R98 a_361_47.n5 a_361_47.n1 311.717
R99 a_361_47.n4 a_361_47.n2 311.717
R100 a_361_47.n12 a_361_47.n11 261.425
R101 a_361_47.n9 a_361_47.n8 202.444
R102 a_361_47.n10 a_361_47.n0 198.177
R103 a_361_47.n13 a_361_47.n12 198.177
R104 a_361_47.n5 a_361_47.n4 63.2476
R105 a_361_47.n12 a_361_47.n10 63.2476
R106 a_361_47.n7 a_361_47.n5 50.4476
R107 a_361_47.n10 a_361_47.n9 50.4476
R108 a_361_47.n1 a_361_47.t10 26.5955
R109 a_361_47.n1 a_361_47.t15 26.5955
R110 a_361_47.n2 a_361_47.t14 26.5955
R111 a_361_47.n2 a_361_47.t13 26.5955
R112 a_361_47.n3 a_361_47.t9 26.5955
R113 a_361_47.n3 a_361_47.t8 26.5955
R114 a_361_47.n6 a_361_47.t12 26.5955
R115 a_361_47.n6 a_361_47.t11 26.5955
R116 a_361_47.n8 a_361_47.t4 24.9236
R117 a_361_47.n8 a_361_47.t5 24.9236
R118 a_361_47.n11 a_361_47.t2 24.9236
R119 a_361_47.n11 a_361_47.t3 24.9236
R120 a_361_47.n0 a_361_47.t0 24.9236
R121 a_361_47.n0 a_361_47.t6 24.9236
R122 a_361_47.n13 a_361_47.t1 24.9236
R123 a_361_47.t7 a_361_47.n13 24.9236
R124 a_361_47.n9 a_361_47.n7 22.5887
R125 VNB VNB.t7 48835.8
R126 VNB.t7 VNB.t8 746.668
R127 VNB.t8 VNB.t3 746.668
R128 VNB.t3 VNB.t9 746.668
R129 VNB.t9 VNB.t4 746.668
R130 VNB.t4 VNB.t10 746.668
R131 VNB.t10 VNB.t5 746.668
R132 VNB.t5 VNB.t6 746.668
R133 VNB.t6 VNB.t0 746.668
R134 VNB.t0 VNB.t2 746.668
R135 VNB.t2 VNB.t1 746.668
R136 VNB VNB.t1 568.889
R137 VPWR.n3 VPWR.n2 320.976
R138 VPWR.n24 VPWR.n1 320.976
R139 VPWR.n17 VPWR.n5 310.502
R140 VPWR.n11 VPWR.n10 310.502
R141 VPWR.n9 VPWR.n8 310.502
R142 VPWR.n7 VPWR.t8 248.906
R143 VPWR.n25 VPWR.n24 43.1829
R144 VPWR.n19 VPWR.n18 34.6358
R145 VPWR.n23 VPWR.n22 34.6358
R146 VPWR.n16 VPWR.n6 34.6358
R147 VPWR.n12 VPWR.n9 32.0005
R148 VPWR.n22 VPWR.n3 27.8593
R149 VPWR.n1 VPWR.t2 26.5955
R150 VPWR.n1 VPWR.t0 26.5955
R151 VPWR.n2 VPWR.t9 26.5955
R152 VPWR.n2 VPWR.t1 26.5955
R153 VPWR.n5 VPWR.t3 26.5955
R154 VPWR.n5 VPWR.t10 26.5955
R155 VPWR.n10 VPWR.t5 26.5955
R156 VPWR.n10 VPWR.t4 26.5955
R157 VPWR.n8 VPWR.t7 26.5955
R158 VPWR.n8 VPWR.t6 26.5955
R159 VPWR.n18 VPWR.n17 9.41227
R160 VPWR.n13 VPWR.n12 9.3005
R161 VPWR.n14 VPWR.n6 9.3005
R162 VPWR.n16 VPWR.n15 9.3005
R163 VPWR.n18 VPWR.n4 9.3005
R164 VPWR.n20 VPWR.n19 9.3005
R165 VPWR.n22 VPWR.n21 9.3005
R166 VPWR.n23 VPWR.n0 9.3005
R167 VPWR.n19 VPWR.n3 6.77697
R168 VPWR.n12 VPWR.n11 6.4005
R169 VPWR.n9 VPWR.n7 5.7932
R170 VPWR.n11 VPWR.n6 3.38874
R171 VPWR.n24 VPWR.n23 0.753441
R172 VPWR.n13 VPWR.n7 0.656729
R173 VPWR.n17 VPWR.n16 0.376971
R174 VPWR.n14 VPWR.n13 0.120292
R175 VPWR.n15 VPWR.n14 0.120292
R176 VPWR.n15 VPWR.n4 0.120292
R177 VPWR.n20 VPWR.n4 0.120292
R178 VPWR.n21 VPWR.n20 0.120292
R179 VPWR.n21 VPWR.n0 0.120292
R180 VPWR.n25 VPWR.n0 0.120292
R181 VPWR VPWR.n25 0.0213333
R182 VPB.t7 VPB.t8 248.599
R183 VPB.t6 VPB.t7 248.599
R184 VPB.t5 VPB.t6 248.599
R185 VPB.t4 VPB.t5 248.599
R186 VPB.t3 VPB.t4 248.599
R187 VPB.t10 VPB.t3 248.599
R188 VPB.t9 VPB.t10 248.599
R189 VPB.t1 VPB.t9 248.599
R190 VPB.t2 VPB.t1 248.599
R191 VPB.t0 VPB.t2 248.599
R192 VPB VPB.t0 189.409
R193 A.n6 A.t4 235.763
R194 A.n1 A.t0 221.72
R195 A.n0 A.t1 221.72
R196 A.n6 A.t5 163.464
R197 A.n3 A.n2 152
R198 A.n5 A.n4 152
R199 A.n7 A.n6 152
R200 A.n1 A.t3 149.421
R201 A.n0 A.t2 149.421
R202 A.n2 A.n1 58.019
R203 A.n5 A.n0 43.7375
R204 A.n4 A.n3 21.7605
R205 A.n7 A 19.5205
R206 A.n6 A.n5 17.8524
R207 A.n2 A.n0 16.9598
R208 A A.n7 9.9205
R209 A.n3 A 5.4405
R210 A.n4 A 2.2405
C0 VPWR m5_872_575# 9.28e-19
C1 A m5_212_112# 2.85e-19
C2 VGND m5_212_112# 4.68e-19
C3 VPWR A 0.049241f
C4 VGND VPWR 0.321008f
C5 m5_872_595# VPWR 1.49e-20
C6 VGND m5_872_n71# 1.49e-20
C7 VPB X 0.003532f
C8 VGND A 0.05431f
C9 VPB m5_212_112# 8.85e-20
C10 VPWR VPB 0.140712f
C11 X m5_212_112# 1.91e-19
C12 VPWR X 0.007108f
C13 VPWR m5_212_112# 4.68e-19
C14 VPB A 0.099483f
C15 VGND m5_872_n91# 9.28e-19
C16 VGND VPB 0.018545f
C17 A X 0.010266f
C18 VGND X 0.006466f
C19 X VNB 0.462652f
C20 VGND VNB 1.09844f
C21 VPWR VNB 0.994271f
C22 A VNB 0.321526f
C23 VPB VNB 1.13634f
C24 m5_872_n71# VNB 5.57e-19
C25 m5_872_n91# VNB 7.76e-19 $ **FLOATING
C26 m5_872_595# VNB 5.57e-19
C27 m5_872_575# VNB 7.76e-19 $ **FLOATING
C28 m5_212_112# VNB 0.007354f $ **FLOATING
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbn_1 VGND VPWR VPB VNB CLK_N SCD SCE D SET_B RESET_B
+ Q_N Q
X0 a_381_363.t0 SCD.t0 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_1102_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2 VPWR.t10 a_1396_21.t2 a_2122_329.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X3 Q.t1 a_2596_47.t2 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X4 a_917_47.t3 a_27_47.t2 a_453_47.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07035 ps=0.755 w=0.42 l=0.15
X5 VPWR.t12 SCE.t0 a_423_315.t1 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND.t1 SCE.t1 a_423_315.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_1614_47.t1 a_1102_21# VGND.t9 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.098 pd=0.99 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_1030_47.t0 a_27_47.t3 a_917_47.t2 VNB.t15 sky130_fd_pr__special_nfet_01v8 ad=0.07335 pd=0.78 as=0.0747 ps=0.775 w=0.36 l=0.15
X9 VPWR.t2 RESET_B.t0 a_1396_21.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1539 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 VPWR.t11 CLK_N.t0 a_27_47.t0 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_1572_329.t1 a_1102_21# VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1743 pd=1.41 as=0.2247 ps=1.375 w=0.84 l=0.15
X12 a_2122_329.t1 a_1714_47.t4 a_1887_21.t2 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.12285 ps=1.17 w=0.84 l=0.15
X13 VGND.t3 a_1887_21.t4 a_1822_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.066 ps=0.745 w=0.42 l=0.15
X14 VPWR.t7 a_1102_21# a_1017_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X15 VPWR.t0 a_1887_21.t5 a_1800_413.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X16 a_1887_21.t1 a_1714_47.t5 a_2004_47.t1 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.11885 ps=1.075 w=0.64 l=0.15
X17 a_1887_21.t3 SET_B.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X18 a_1800_413.t0 a_27_47.t4 a_1714_47.t2 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1102_21# a_917_47.t4 a_1241_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.10205 ps=0.995 w=0.64 l=0.15
X20 a_193_47.t0 a_27_47.t5 VGND.t6 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 a_453_47.t1 D.t0 a_735_47.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.05985 ps=0.705 w=0.42 l=0.15
X22 a_1714_47.t3 a_193_47.t2 a_1572_329.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1743 ps=1.41 w=0.42 l=0.15
X23 a_2004_47.t0 a_1396_21.t3 a_1887_21.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 Q.t0 a_2596_47.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X25 VGND.t4 a_1887_21.t6 a_2596_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 a_193_47.t1 a_27_47.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_1241_47.t2 SET_B.t1 VGND.t13 VNB.t23 sky130_fd_pr__nfet_01v8 ad=0.10205 pd=0.995 as=0.08295 ps=0.815 w=0.42 l=0.15
X28 a_1241_47.t1 a_1396_21.t4 a_1102_21# VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X29 a_1017_413.t0 a_193_47.t3 a_917_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X30 VGND.t10 a_1102_21# a_1030_47.t1 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08295 pd=0.815 as=0.07335 ps=0.78 w=0.42 l=0.15
X31 a_735_47.t0 a_423_315.t2 VGND.t8 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.05985 ps=0.705 w=0.42 l=0.15
X32 VPWR.t3 a_1887_21.t7 a_2596_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X33 a_453_47.t5 a_423_315.t3 a_381_363.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X34 a_381_47.t1 SCD.t1 VGND.t7 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_1822_47.t0 a_193_47.t4 a_1714_47.t0 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0702 ps=0.75 w=0.36 l=0.15
X36 Q_N.t0 a_1887_21.t8 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X37 Q_N.t1 a_1887_21.t9 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1539 ps=1.335 w=1 l=0.15
X38 a_1714_47.t1 a_27_47.t7 a_1614_47.t0 VNB.t13 sky130_fd_pr__special_nfet_01v8 ad=0.0702 pd=0.75 as=0.098 ps=0.99 w=0.36 l=0.15
X39 a_453_47.t2 D.t1 a_752_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X40 a_917_47.t1 a_193_47.t5 a_453_47.t0 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.0747 pd=0.775 as=0.066 ps=0.745 w=0.36 l=0.15
X41 a_2004_47.t2 SET_B.t2 VGND.t12 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.11885 pd=1.075 as=0.05985 ps=0.705 w=0.42 l=0.15
X42 a_752_413.t0 SCE.t2 VPWR.t13 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 VGND.t11 CLK_N.t1 a_27_47.t1 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X44 a_453_47.t4 SCE.t3 a_381_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1239 pd=1.43 as=0.0441 ps=0.63 w=0.42 l=0.15
X45 VGND.t0 RESET_B.t1 a_1396_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 SCD.n0 SCD.t1 301.533
R1 SCD.n0 SCD.t0 197.62
R2 SCD SCD.n0 154.058
R3 VPWR.n22 VPWR.t10 793.365
R4 VPWR.n16 VPWR.n15 732.75
R5 VPWR.n43 VPWR.t7 686.259
R6 VPWR.n58 VPWR.n1 604.394
R7 VPWR.n50 VPWR.n5 601.292
R8 VPWR.n29 VPWR.n28 585
R9 VPWR.n37 VPWR.t8 397.274
R10 VPWR.n56 VPWR.t6 374.75
R11 VPWR.n18 VPWR.n17 321.776
R12 VPWR.n28 VPWR.t4 91.4648
R13 VPWR.n28 VPWR.t0 91.4648
R14 VPWR.n5 VPWR.t13 63.3219
R15 VPWR.n5 VPWR.t12 63.3219
R16 VPWR.n15 VPWR.t2 63.1021
R17 VPWR.n17 VPWR.t3 57.7247
R18 VPWR.n1 VPWR.t1 41.5552
R19 VPWR.n1 VPWR.t11 41.5552
R20 VPWR.n51 VPWR.n3 34.6358
R21 VPWR.n55 VPWR.n3 34.6358
R22 VPWR.n45 VPWR.n44 34.6358
R23 VPWR.n45 VPWR.n6 34.6358
R24 VPWR.n49 VPWR.n6 34.6358
R25 VPWR.n38 VPWR.n9 34.6358
R26 VPWR.n42 VPWR.n9 34.6358
R27 VPWR.n31 VPWR.n30 34.6358
R28 VPWR.n31 VPWR.n11 34.6358
R29 VPWR.n35 VPWR.n11 34.6358
R30 VPWR.n36 VPWR.n35 34.6358
R31 VPWR.n23 VPWR.n13 34.6358
R32 VPWR.n17 VPWR.t9 32.5902
R33 VPWR.n44 VPWR.n43 31.2476
R34 VPWR.n27 VPWR.n13 28.9134
R35 VPWR.n15 VPWR.t5 28.0332
R36 VPWR.n51 VPWR.n50 24.0946
R37 VPWR.n58 VPWR.n57 22.9652
R38 VPWR.n56 VPWR.n55 21.4593
R39 VPWR.n57 VPWR.n56 21.0829
R40 VPWR.n50 VPWR.n49 20.3299
R41 VPWR.n30 VPWR.n29 18.1464
R42 VPWR.n23 VPWR.n22 13.6287
R43 VPWR.n21 VPWR.n20 10.706
R44 VPWR.n20 VPWR.n16 10.1241
R45 VPWR.n43 VPWR.n42 9.41227
R46 VPWR.n20 VPWR.n19 9.3005
R47 VPWR.n21 VPWR.n14 9.3005
R48 VPWR.n24 VPWR.n23 9.3005
R49 VPWR.n25 VPWR.n13 9.3005
R50 VPWR.n27 VPWR.n26 9.3005
R51 VPWR.n30 VPWR.n12 9.3005
R52 VPWR.n32 VPWR.n31 9.3005
R53 VPWR.n33 VPWR.n11 9.3005
R54 VPWR.n35 VPWR.n34 9.3005
R55 VPWR.n36 VPWR.n10 9.3005
R56 VPWR.n39 VPWR.n38 9.3005
R57 VPWR.n40 VPWR.n9 9.3005
R58 VPWR.n42 VPWR.n41 9.3005
R59 VPWR.n43 VPWR.n8 9.3005
R60 VPWR.n44 VPWR.n7 9.3005
R61 VPWR.n46 VPWR.n45 9.3005
R62 VPWR.n47 VPWR.n6 9.3005
R63 VPWR.n49 VPWR.n48 9.3005
R64 VPWR.n50 VPWR.n4 9.3005
R65 VPWR.n52 VPWR.n51 9.3005
R66 VPWR.n53 VPWR.n3 9.3005
R67 VPWR.n55 VPWR.n54 9.3005
R68 VPWR.n56 VPWR.n2 9.3005
R69 VPWR.n57 VPWR.n0 9.3005
R70 VPWR.n18 VPWR.n16 7.8441
R71 VPWR.n59 VPWR.n58 7.12063
R72 VPWR.n37 VPWR.n36 6.4005
R73 VPWR.n22 VPWR.n21 3.8405
R74 VPWR.n38 VPWR.n37 3.38874
R75 VPWR.n29 VPWR.n27 2.44414
R76 VPWR.n19 VPWR.n18 0.21101
R77 VPWR.n59 VPWR.n0 0.148519
R78 VPWR.n19 VPWR.n14 0.120292
R79 VPWR.n24 VPWR.n14 0.120292
R80 VPWR.n25 VPWR.n24 0.120292
R81 VPWR.n26 VPWR.n25 0.120292
R82 VPWR.n26 VPWR.n12 0.120292
R83 VPWR.n32 VPWR.n12 0.120292
R84 VPWR.n33 VPWR.n32 0.120292
R85 VPWR.n34 VPWR.n33 0.120292
R86 VPWR.n34 VPWR.n10 0.120292
R87 VPWR.n39 VPWR.n10 0.120292
R88 VPWR.n40 VPWR.n39 0.120292
R89 VPWR.n41 VPWR.n40 0.120292
R90 VPWR.n41 VPWR.n8 0.120292
R91 VPWR.n8 VPWR.n7 0.120292
R92 VPWR.n46 VPWR.n7 0.120292
R93 VPWR.n47 VPWR.n46 0.120292
R94 VPWR.n48 VPWR.n47 0.120292
R95 VPWR.n48 VPWR.n4 0.120292
R96 VPWR.n52 VPWR.n4 0.120292
R97 VPWR.n53 VPWR.n52 0.120292
R98 VPWR.n54 VPWR.n53 0.120292
R99 VPWR.n54 VPWR.n2 0.120292
R100 VPWR.n2 VPWR.n0 0.120292
R101 VPWR VPWR.n59 0.114842
R102 a_381_363.t0 a_381_363.t1 64.6411
R103 VPB.t11 VPB.t12 1287.38
R104 VPB.t13 VPB.t19 636.293
R105 VPB.t15 VPB.t2 588.942
R106 VPB.t8 VPB.t4 556.386
R107 VPB.t1 VPB.t10 556.386
R108 VPB.t12 VPB.t9 426.168
R109 VPB.t3 VPB.t11 355.14
R110 VPB.t17 VPB.t0 349.221
R111 VPB.t0 VPB.t6 319.627
R112 VPB.t2 VPB.t8 287.072
R113 VPB.t7 VPB.t5 287.072
R114 VPB.t6 VPB.t16 284.113
R115 VPB.t4 VPB.t14 281.154
R116 VPB.t9 VPB.t17 248.599
R117 VPB.t5 VPB.t3 248.599
R118 VPB.t20 VPB.t7 248.599
R119 VPB.t19 VPB.t20 248.599
R120 VPB.t18 VPB.t1 248.599
R121 VPB.t16 VPB.t15 213.084
R122 VPB.t10 VPB.t13 213.084
R123 VPB VPB.t18 142.056
R124 SET_B.n1 SET_B.n0 438.599
R125 SET_B.n2 SET_B.t0 386.848
R126 SET_B.n3 SET_B.n2 178.222
R127 SET_B.n3 SET_B.n1 156.823
R128 SET_B.n1 SET_B.t1 142.635
R129 SET_B.n2 SET_B.t2 142.635
R130 SET_B SET_B.n3 5.0092
R131 SET_B.n3 SET_B 3.15412
R132 a_1396_21.t1 a_1396_21.n4 740.542
R133 a_1396_21.n1 a_1396_21.t0 286.716
R134 a_1396_21.n3 a_1396_21.t4 212.989
R135 a_1396_21.n4 a_1396_21.n3 211.846
R136 a_1396_21.n0 a_1396_21.t3 211.513
R137 a_1396_21.n0 a_1396_21.t2 206.935
R138 a_1396_21.n3 a_1396_21.n2 204.869
R139 a_1396_21.n1 a_1396_21.n0 152
R140 a_1396_21.n4 a_1396_21.n1 9.77505
R141 a_2122_329.t0 a_2122_329.t1 49.2505
R142 a_2596_47.t1 a_2596_47.n1 384.125
R143 a_2596_47.n1 a_2596_47.t0 243.28
R144 a_2596_47.n0 a_2596_47.t2 239.505
R145 a_2596_47.n1 a_2596_47.n0 175.079
R146 a_2596_47.n0 a_2596_47.t3 167.204
R147 Q.n1 Q.t1 353.606
R148 Q.n0 Q.t0 209.923
R149 Q Q.n0 68.3375
R150 Q.n1 Q 9.10538
R151 Q Q.n1 7.47898
R152 Q.n0 Q 6.64665
R153 a_27_47.n1 a_27_47.t2 493.933
R154 a_27_47.t0 a_27_47.n5 420.808
R155 a_27_47.n0 a_27_47.t4 343.399
R156 a_27_47.n0 a_27_47.t7 283.659
R157 a_27_47.n4 a_27_47.t6 262.945
R158 a_27_47.n3 a_27_47.t1 261.135
R159 a_27_47.n4 a_27_47.t5 227.597
R160 a_27_47.n2 a_27_47.n1 164.404
R161 a_27_47.n5 a_27_47.n4 152
R162 a_27_47.n1 a_27_47.t3 138.977
R163 a_27_47.n5 a_27_47.n3 21.4266
R164 a_27_47.n3 a_27_47.n2 13.2617
R165 a_27_47.n2 a_27_47.n0 12.1899
R166 a_453_47.n2 a_453_47.n0 663.077
R167 a_453_47.t5 a_453_47.n3 424.159
R168 a_453_47.n3 a_453_47.t4 291.046
R169 a_453_47.n2 a_453_47.n1 256.082
R170 a_453_47.n0 a_453_47.t3 93.81
R171 a_453_47.n1 a_453_47.t0 63.3338
R172 a_453_47.n0 a_453_47.t2 63.3219
R173 a_453_47.n3 a_453_47.n2 34.6156
R174 a_453_47.n1 a_453_47.t1 29.7268
R175 a_917_47.n4 a_917_47.n3 704.789
R176 a_917_47.n3 a_917_47.n0 293.938
R177 a_917_47.n2 a_917_47.t4 220.706
R178 a_917_47.n3 a_917_47.n2 220.218
R179 a_917_47.n2 a_917_47.n1 214.135
R180 a_917_47.n0 a_917_47.t2 93.3338
R181 a_917_47.t0 a_917_47.n4 63.3219
R182 a_917_47.n4 a_917_47.t3 63.3219
R183 a_917_47.n0 a_917_47.t1 45.0005
R184 SCE.n2 SCE.n1 285.988
R185 SCE.n3 SCE.n2 266.591
R186 SCE.n1 SCE.t2 228.148
R187 SCE.n4 SCE.n3 152
R188 SCE.n3 SCE.t3 97.8329
R189 SCE.n2 SCE.t1 93.1872
R190 SCE.n1 SCE.t0 93.1872
R191 SCE SCE.n4 28.4177
R192 SCE.n0 SCE 17.1641
R193 SCE.n4 SCE 4.04261
R194 SCE.n0 SCE 2.61868
R195 SCE SCE.n0 1.51629
R196 a_423_315.n0 a_423_315.t1 678.063
R197 a_423_315.n0 a_423_315.t3 478.704
R198 a_423_315.n1 a_423_315.t2 284.283
R199 a_423_315.t0 a_423_315.n1 284.104
R200 a_423_315.n1 a_423_315.n0 76.2817
R201 VGND.n31 VGND.t9 279.471
R202 VGND.n56 VGND.t7 245.448
R203 VGND.n14 VGND.n13 207.882
R204 VGND.n39 VGND.n38 205.707
R205 VGND.n24 VGND.n23 202.724
R206 VGND.n59 VGND.n58 199.739
R207 VGND.n50 VGND.n4 198.964
R208 VGND.n16 VGND.n15 110.672
R209 VGND.n38 VGND.t10 74.2862
R210 VGND.n15 VGND.t0 57.8264
R211 VGND.n13 VGND.t4 54.2862
R212 VGND.n23 VGND.t3 42.8576
R213 VGND.n4 VGND.t1 42.8576
R214 VGND.n23 VGND.t12 38.5719
R215 VGND.n38 VGND.t13 38.5719
R216 VGND.n4 VGND.t8 38.5719
R217 VGND.n58 VGND.t6 38.5719
R218 VGND.n58 VGND.t11 38.5719
R219 VGND.n17 VGND.n12 34.6358
R220 VGND.n21 VGND.n12 34.6358
R221 VGND.n22 VGND.n21 34.6358
R222 VGND.n25 VGND.n22 34.6358
R223 VGND.n29 VGND.n10 34.6358
R224 VGND.n30 VGND.n29 34.6358
R225 VGND.n32 VGND.n30 34.6358
R226 VGND.n36 VGND.n8 34.6358
R227 VGND.n37 VGND.n36 34.6358
R228 VGND.n40 VGND.n37 34.6358
R229 VGND.n44 VGND.n6 34.6358
R230 VGND.n45 VGND.n44 34.6358
R231 VGND.n46 VGND.n45 34.6358
R232 VGND.n46 VGND.n3 34.6358
R233 VGND.n52 VGND.n51 34.6358
R234 VGND.n52 VGND.n1 34.6358
R235 VGND.n56 VGND.n1 27.4829
R236 VGND.n50 VGND.n3 26.7299
R237 VGND.n13 VGND.t2 25.9346
R238 VGND.n15 VGND.t5 24.7418
R239 VGND.n59 VGND.n57 22.9652
R240 VGND.n40 VGND.n39 21.8358
R241 VGND.n57 VGND.n56 21.0829
R242 VGND.n17 VGND.n16 20.3299
R243 VGND.n51 VGND.n50 17.6946
R244 VGND.n39 VGND.n6 12.8005
R245 VGND.n24 VGND.n10 9.78874
R246 VGND.n57 VGND.n0 9.3005
R247 VGND.n56 VGND.n55 9.3005
R248 VGND.n54 VGND.n1 9.3005
R249 VGND.n53 VGND.n52 9.3005
R250 VGND.n51 VGND.n2 9.3005
R251 VGND.n50 VGND.n49 9.3005
R252 VGND.n48 VGND.n3 9.3005
R253 VGND.n47 VGND.n46 9.3005
R254 VGND.n45 VGND.n5 9.3005
R255 VGND.n44 VGND.n43 9.3005
R256 VGND.n42 VGND.n6 9.3005
R257 VGND.n41 VGND.n40 9.3005
R258 VGND.n37 VGND.n7 9.3005
R259 VGND.n36 VGND.n35 9.3005
R260 VGND.n34 VGND.n8 9.3005
R261 VGND.n33 VGND.n32 9.3005
R262 VGND.n30 VGND.n9 9.3005
R263 VGND.n29 VGND.n28 9.3005
R264 VGND.n27 VGND.n10 9.3005
R265 VGND.n26 VGND.n25 9.3005
R266 VGND.n22 VGND.n11 9.3005
R267 VGND.n21 VGND.n20 9.3005
R268 VGND.n19 VGND.n12 9.3005
R269 VGND.n18 VGND.n17 9.3005
R270 VGND.n60 VGND.n59 7.12063
R271 VGND.n16 VGND.n14 7.10092
R272 VGND.n32 VGND.n31 5.64756
R273 VGND.n25 VGND.n24 5.27109
R274 VGND.n31 VGND.n8 2.25932
R275 VGND.n18 VGND.n14 0.218009
R276 VGND.n60 VGND.n0 0.148519
R277 VGND.n19 VGND.n18 0.120292
R278 VGND.n20 VGND.n19 0.120292
R279 VGND.n20 VGND.n11 0.120292
R280 VGND.n26 VGND.n11 0.120292
R281 VGND.n27 VGND.n26 0.120292
R282 VGND.n28 VGND.n27 0.120292
R283 VGND.n28 VGND.n9 0.120292
R284 VGND.n33 VGND.n9 0.120292
R285 VGND.n34 VGND.n33 0.120292
R286 VGND.n35 VGND.n34 0.120292
R287 VGND.n35 VGND.n7 0.120292
R288 VGND.n41 VGND.n7 0.120292
R289 VGND.n42 VGND.n41 0.120292
R290 VGND.n43 VGND.n42 0.120292
R291 VGND.n43 VGND.n5 0.120292
R292 VGND.n47 VGND.n5 0.120292
R293 VGND.n48 VGND.n47 0.120292
R294 VGND.n49 VGND.n48 0.120292
R295 VGND.n49 VGND.n2 0.120292
R296 VGND.n53 VGND.n2 0.120292
R297 VGND.n54 VGND.n53 0.120292
R298 VGND.n55 VGND.n54 0.120292
R299 VGND.n55 VGND.n0 0.120292
R300 VGND VGND.n60 0.114842
R301 VNB.t2 VNB.t3 2776.7
R302 VNB.t11 VNB.t10 2677.02
R303 VNB.t7 VNB.t1 2677.02
R304 VNB.t6 VNB.t19 2677.02
R305 VNB.t14 VNB.t16 2677.02
R306 VNB.t22 VNB.t20 1666.02
R307 VNB.t9 VNB.t15 1609.06
R308 VNB.t18 VNB.t23 1552.1
R309 VNB.t13 VNB.t8 1537.86
R310 VNB.t15 VNB.t18 1452.43
R311 VNB.t23 VNB.t0 1438.19
R312 VNB.t19 VNB.t13 1423.95
R313 VNB.t1 VNB.t11 1381.23
R314 VNB.t10 VNB.t4 1352.75
R315 VNB.t8 VNB.t5 1352.75
R316 VNB.t12 VNB.t9 1352.75
R317 VNB.t5 VNB.t22 1238.83
R318 VNB.t17 VNB.t12 1238.83
R319 VNB.t3 VNB.t17 1238.83
R320 VNB.t20 VNB.t7 1196.12
R321 VNB.t0 VNB.t6 1196.12
R322 VNB.t21 VNB.t14 1196.12
R323 VNB.t16 VNB.t2 1025.24
R324 VNB VNB.t21 683.495
R325 a_1614_47.n0 a_1614_47.t0 75.0005
R326 a_1614_47.n1 a_1614_47.n0 67.2005
R327 a_1614_47.n0 a_1614_47.t1 13.144
R328 a_1030_47.t1 a_1030_47.t0 99.0472
R329 RESET_B.n0 RESET_B.t1 203.042
R330 RESET_B.n0 RESET_B.t0 174.123
R331 RESET_B RESET_B.n0 154.111
R332 CLK_N.n0 CLK_N.t0 272.062
R333 CLK_N.n0 CLK_N.t1 236.716
R334 CLK_N.n1 CLK_N.n0 152
R335 CLK_N CLK_N.n1 7.6805
R336 CLK_N.n1 CLK_N 4.75479
R337 a_1572_329.t1 a_1572_329.t0 236.869
R338 a_1714_47.n3 a_1714_47.n2 692.294
R339 a_1714_47.n2 a_1714_47.n0 275.937
R340 a_1714_47.n1 a_1714_47.t4 241.536
R341 a_1714_47.n2 a_1714_47.n1 235.919
R342 a_1714_47.n1 a_1714_47.t5 196.549
R343 a_1714_47.n0 a_1714_47.t1 70.0005
R344 a_1714_47.t2 a_1714_47.n3 63.3219
R345 a_1714_47.n3 a_1714_47.t3 63.3219
R346 a_1714_47.n0 a_1714_47.t0 60.0005
R347 a_1887_21.n7 a_1887_21.n6 594.413
R348 a_1887_21.n5 a_1887_21.t4 386.848
R349 a_1887_21.n4 a_1887_21.n2 305.288
R350 a_1887_21.n1 a_1887_21.t9 292.413
R351 a_1887_21.n4 a_1887_21.n3 278.113
R352 a_1887_21.n0 a_1887_21.t7 231.945
R353 a_1887_21.n1 a_1887_21.t8 220.113
R354 a_1887_21.n6 a_1887_21.n5 204.841
R355 a_1887_21.n0 a_1887_21.t6 164.464
R356 a_1887_21.n2 a_1887_21.n0 151.742
R357 a_1887_21.n5 a_1887_21.t5 142.635
R358 a_1887_21.n7 a_1887_21.t3 91.4648
R359 a_1887_21.t2 a_1887_21.n7 32.8338
R360 a_1887_21.n6 a_1887_21.n4 30.4946
R361 a_1887_21.n3 a_1887_21.t0 25.313
R362 a_1887_21.n3 a_1887_21.t1 25.313
R363 a_1887_21.n2 a_1887_21.n1 2.67828
R364 a_1822_47.t1 a_1822_47.t0 93.0601
R365 a_1017_413.t0 a_1017_413.t1 211.071
R366 a_1800_413.t0 a_1800_413.t1 206.381
R367 a_2004_47.t0 a_2004_47.n0 455.964
R368 a_2004_47.n0 a_2004_47.t2 64.2862
R369 a_2004_47.n0 a_2004_47.t1 47.7237
R370 a_1241_47.n0 a_1241_47.t1 465.606
R371 a_1241_47.n0 a_1241_47.t2 62.8576
R372 a_1241_47.t0 a_1241_47.n0 26.2951
R373 a_193_47.n0 a_193_47.t4 524.309
R374 a_193_47.t1 a_193_47.n3 367.062
R375 a_193_47.n1 a_193_47.t5 321.067
R376 a_193_47.n1 a_193_47.t3 307.325
R377 a_193_47.n3 a_193_47.t0 302.7
R378 a_193_47.n2 a_193_47.n0 171.565
R379 a_193_47.n0 a_193_47.t2 148.35
R380 a_193_47.n3 a_193_47.n2 12.4849
R381 a_193_47.n2 a_193_47.n1 9.3005
R382 D.n0 D.t0 308.481
R383 D.n0 D.t1 224.934
R384 D.n1 D.n0 152
R385 D D.n1 24.5111
R386 D.n1 D 5.45235
R387 a_735_47.t0 a_735_47.t1 81.4291
R388 a_381_47.t0 a_381_47.t1 60.0005
R389 Q_N.n1 Q_N.t1 353.795
R390 Q_N.n0 Q_N.t0 209.923
R391 Q_N Q_N.n0 79.4391
R392 Q_N.n1 Q_N 8.2361
R393 Q_N Q_N.n1 6.90173
R394 Q_N.n0 Q_N 5.61454
R395 a_752_413.t0 a_752_413.t1 126.644
C0 VGND Q 0.064261f
C1 Q RESET_B 6.25e-20
C2 Q_N RESET_B 0.001681f
C3 Q_N VGND 0.086192f
C4 VPWR Q 0.098264f
C5 Q_N VPWR 0.061416f
C6 VGND RESET_B 0.028485f
C7 VPWR RESET_B 0.009854f
C8 VGND VPWR 0.081614f
C9 SET_B Q 1.23e-19
C10 Q_N SET_B 3.62e-19
C11 SET_B RESET_B 0.002263f
C12 VGND SET_B 0.294482f
C13 D RESET_B 4.17e-21
C14 VGND D 0.010765f
C15 VPWR SET_B 0.025481f
C16 VGND SCE 0.073258f
C17 VGND SCD 0.033229f
C18 VPWR D 0.049441f
C19 VPWR SCE 0.038617f
C20 VPWR SCD 0.042428f
C21 CLK_N VGND 0.01748f
C22 VPB Q 0.012264f
C23 CLK_N VPWR 0.017689f
C24 Q_N VPB 0.010238f
C25 D SCE 0.05245f
C26 VPB RESET_B 0.047075f
C27 VGND VPB 0.015537f
C28 SCD SCE 0.10264f
C29 VPWR VPB 0.307265f
C30 VPB SET_B 0.145752f
C31 VPB D 0.086957f
C32 VPB SCE 0.138182f
C33 SCD VPB 0.077422f
C34 CLK_N VPB 0.069967f
C35 VPWR a_1351_329# 0.009837f
C36 a_1102_21# RESET_B 6.51e-21
C37 VGND a_1102_21# 0.054252f
C38 VPWR a_1102_21# 0.160129f
C39 SET_B a_1102_21# 0.1761f
C40 VPB a_1102_21# 0.142801f
C41 a_1351_329# a_1102_21# 0.010395f
C42 Q VNB 0.094533f
C43 Q_N VNB 0.013509f
C44 RESET_B VNB 0.132569f
C45 VGND VNB 1.54739f
C46 VPWR VNB 1.24599f
C47 SET_B VNB 0.265114f
C48 D VNB 0.115683f
C49 SCE VNB 0.301733f
C50 SCD VNB 0.139433f
C51 CLK_N VNB 0.196032f
C52 VPB VNB 2.81966f
C53 a_1102_21# VNB 0.241075f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfsbp_2 SCD CLK Q_N D SET_B SCE Q VPWR VGND VPB VNB
X0 a_1006_47.t1 a_818_47.t2 a_181_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_1781_295.t1 a_1597_329.t4 VPWR.t13 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND.t0 a_328_21.t2 a_265_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 Q_N.t1 a_1597_329.t5 VGND.t14 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_818_47.t0 a_652_47.t2 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VPWR.t3 a_2501_47.t2 Q.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 a_1090_47.t0 a_818_47.t3 a_1006_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR.t0 SCD.t0 a_27_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 Q.t2 a_2501_47.t3 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X9 VPWR.t9 SET_B.t0 a_1132_21.t1 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.27 as=0.0714 ps=0.76 w=0.42 l=0.15
X10 a_1517_47.t1 a_1006_47.t4 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.2336 pd=1.37 as=0.09575 ps=0.965 w=0.64 l=0.15
X11 VGND.t10 a_1132_21.t2 a_1090_47.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 VGND.t11 a_1597_329.t6 a_2501_47.t0 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_181_47.t3 SCE.t0 a_109_47.t0 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 VGND.t9 SCE.t1 a_328_21.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1006_47.t3 a_652_47.t3 a_181_47.t2 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 VGND.t6 a_2501_47.t4 Q.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_818_47.t1 a_652_47.t4 VPWR.t8 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X18 VGND.t8 SET_B.t1 a_1885_47.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0735 ps=0.77 w=0.42 l=0.15
X19 VPWR.t1 SCE.t2 a_328_21.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.162825 ps=1.8 w=0.64 l=0.15
X20 a_1597_329.t0 a_818_47.t4 a_1517_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.09 as=0.2336 ps=1.37 w=0.64 l=0.15
X21 a_181_47.t4 D.t0 a_193_369.t1 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.1056 pd=0.97 as=0.0672 ps=0.85 w=0.64 l=0.15
X22 a_27_369.t0 a_328_21.t3 a_181_47.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.162825 pd=1.8 as=0.1056 ps=0.97 w=0.64 l=0.15
X23 a_1597_329.t3 a_652_47.t5 a_1525_329.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.32 as=0.0882 ps=1.05 w=0.84 l=0.15
X24 a_265_47.t1 D.t1 a_181_47.t5 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X25 a_1781_295.t0 a_1597_329.t7 VGND.t12 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 a_1813_47.t0 a_652_47.t6 a_1597_329.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.09 w=0.42 l=0.15
X27 a_1350_47.t0 a_1006_47.t5 a_1132_21.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 Q.t0 a_2501_47.t5 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X29 a_193_369.t0 SCE.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 a_1525_329.t0 a_1006_47.t6 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.1428 ps=1.27 w=0.84 l=0.15
X31 a_1885_47.t1 a_1781_295.t2 a_1813_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X32 VPWR.t12 a_1597_329.t8 Q_N.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.325 pd=2.65 as=0.135 ps=1.27 w=1 l=0.15
X33 VGND.t5 CLK.t0 a_652_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X34 VPWR.t7 CLK.t1 a_652_47.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X35 VPWR.t10 a_1132_21.t3 a_1102_413.t0 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.09345 pd=0.865 as=0.063 ps=0.72 w=0.42 l=0.15
X36 VGND.t2 SET_B.t2 a_1350_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.09575 pd=0.965 as=0.0441 ps=0.63 w=0.42 l=0.15
X37 VGND.t13 a_1597_329.t9 Q_N.t0 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.21125 pd=1.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 a_1102_413.t1 a_652_47.t7 a_1006_47.t2 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.06825 ps=0.745 w=0.42 l=0.15
X39 Q_N.t2 a_1597_329.t10 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR.t14 a_1597_329.t11 a_2501_47.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X41 a_1597_329.t1 SET_B.t3 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08505 ps=0.825 w=0.42 l=0.15
X42 a_109_47.t1 SCD.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_818_47.t1 a_818_47.n4 673.492
R1 a_818_47.n1 a_818_47.t4 385.065
R2 a_818_47.n3 a_818_47.t3 383.315
R3 a_818_47.n3 a_818_47.t2 319.728
R4 a_818_47.n2 a_818_47.t0 274.921
R5 a_818_47.n2 a_818_47.n1 204.853
R6 a_818_47.n4 a_818_47.n3 190.707
R7 a_818_47.n1 a_818_47.n0 148.35
R8 a_818_47.n4 a_818_47.n2 2.5605
R9 a_181_47.n1 a_181_47.t0 691.576
R10 a_181_47.n3 a_181_47.n2 610.928
R11 a_181_47.n1 a_181_47.t2 285.824
R12 a_181_47.n2 a_181_47.n0 268.38
R13 a_181_47.n3 a_181_47.t4 60.0239
R14 a_181_47.t1 a_181_47.n3 41.5552
R15 a_181_47.n0 a_181_47.t5 38.5719
R16 a_181_47.n0 a_181_47.t3 38.5719
R17 a_181_47.n2 a_181_47.n1 21.7005
R18 a_1006_47.n5 a_1006_47.n0 659.918
R19 a_1006_47.n3 a_1006_47.n2 312.132
R20 a_1006_47.n1 a_1006_47.t6 263.863
R21 a_1006_47.n3 a_1006_47.t5 243.046
R22 a_1006_47.n6 a_1006_47.n5 242.078
R23 a_1006_47.n4 a_1006_47.n1 201.111
R24 a_1006_47.n1 a_1006_47.t4 167.463
R25 a_1006_47.n4 a_1006_47.n3 152
R26 a_1006_47.n0 a_1006_47.t1 89.1195
R27 a_1006_47.n0 a_1006_47.t2 63.3219
R28 a_1006_47.n5 a_1006_47.n4 50.0711
R29 a_1006_47.t0 a_1006_47.n6 38.5719
R30 a_1006_47.n6 a_1006_47.t3 38.5719
R31 VPB.t16 VPB.t8 961.838
R32 VPB.t18 VPB.t17 642.212
R33 VPB.t13 VPB.t12 594.861
R34 VPB.t0 VPB.t11 556.386
R35 VPB.t8 VPB.t0 556.386
R36 VPB.t15 VPB.t6 556.386
R37 VPB.t2 VPB.t10 556.386
R38 VPB.t7 VPB.t2 550.467
R39 VPB.t17 VPB.t9 343.303
R40 VPB.t19 VPB.t7 284.113
R41 VPB.t12 VPB.t5 281.154
R42 VPB.t6 VPB.t14 281.154
R43 VPB.t14 VPB.t18 266.356
R44 VPB.t5 VPB.t4 248.599
R45 VPB.t11 VPB.t13 248.599
R46 VPB.t10 VPB.t15 248.599
R47 VPB.t1 VPB.t3 248.599
R48 VPB.t9 VPB.t16 213.084
R49 VPB.t3 VPB.t19 213.084
R50 VPB VPB.t1 192.369
R51 a_1597_329.t3 a_1597_329.n7 774.99
R52 a_1597_329.n7 a_1597_329.t1 662.782
R53 a_1597_329.n4 a_1597_329.n3 469.707
R54 a_1597_329.n0 a_1597_329.t11 249.034
R55 a_1597_329.n1 a_1597_329.t8 212.081
R56 a_1597_329.n2 a_1597_329.t10 212.081
R57 a_1597_329.n0 a_1597_329.t6 176.733
R58 a_1597_329.n7 a_1597_329.n6 176.599
R59 a_1597_329.n6 a_1597_329.t4 167.038
R60 a_1597_329.n5 a_1597_329.n2 147.522
R61 a_1597_329.n1 a_1597_329.n0 146.792
R62 a_1597_329.n1 a_1597_329.t9 139.78
R63 a_1597_329.n2 a_1597_329.t5 139.78
R64 a_1597_329.n4 a_1597_329.t7 132.282
R65 a_1597_329.n3 a_1597_329.t2 81.4291
R66 a_1597_329.n2 a_1597_329.n1 61.346
R67 a_1597_329.n6 a_1597_329.n5 60.666
R68 a_1597_329.n3 a_1597_329.t0 34.8666
R69 a_1597_329.n5 a_1597_329.n4 13.0648
R70 VPWR.n53 VPWR.t1 717.596
R71 VPWR.n41 VPWR.t10 695.119
R72 VPWR.n28 VPWR.t13 663.062
R73 VPWR.n30 VPWR.t5 662.285
R74 VPWR.n60 VPWR.n1 598.965
R75 VPWR.n5 VPWR.n4 598.965
R76 VPWR.n10 VPWR.n9 585
R77 VPWR.n18 VPWR.n17 311.579
R78 VPWR.n19 VPWR.t3 265.658
R79 VPWR.n22 VPWR.t12 259.317
R80 VPWR.n15 VPWR.t11 255.905
R81 VPWR.n9 VPWR.t6 87.9469
R82 VPWR.n9 VPWR.t9 84.4291
R83 VPWR.n17 VPWR.t14 56.9458
R84 VPWR.n1 VPWR.t2 41.5552
R85 VPWR.n1 VPWR.t0 41.5552
R86 VPWR.n4 VPWR.t8 41.5552
R87 VPWR.n4 VPWR.t7 41.5552
R88 VPWR.n54 VPWR.n2 34.6358
R89 VPWR.n58 VPWR.n2 34.6358
R90 VPWR.n59 VPWR.n58 34.6358
R91 VPWR.n45 VPWR.n7 34.6358
R92 VPWR.n46 VPWR.n45 34.6358
R93 VPWR.n47 VPWR.n46 34.6358
R94 VPWR.n34 VPWR.n12 34.6358
R95 VPWR.n35 VPWR.n34 34.6358
R96 VPWR.n23 VPWR.n15 33.1299
R97 VPWR.n17 VPWR.t4 33.1097
R98 VPWR.n40 VPWR.n39 30.6829
R99 VPWR.n30 VPWR.n29 30.1181
R100 VPWR.n47 VPWR.n5 29.7417
R101 VPWR.n28 VPWR.n27 28.6123
R102 VPWR.n52 VPWR.n51 28.4707
R103 VPWR.n41 VPWR.n40 25.6005
R104 VPWR.n22 VPWR.n21 25.224
R105 VPWR.n60 VPWR.n59 22.9652
R106 VPWR.n23 VPWR.n22 22.2123
R107 VPWR.n27 VPWR.n15 20.3299
R108 VPWR.n41 VPWR.n7 18.824
R109 VPWR.n21 VPWR.n18 17.6946
R110 VPWR.n54 VPWR.n53 16.3529
R111 VPWR.n29 VPWR.n28 15.8123
R112 VPWR.n51 VPWR.n5 14.6829
R113 VPWR.n30 VPWR.n12 14.3064
R114 VPWR.n36 VPWR.n35 10.6358
R115 VPWR.n21 VPWR.n20 9.3005
R116 VPWR.n22 VPWR.n16 9.3005
R117 VPWR.n24 VPWR.n23 9.3005
R118 VPWR.n25 VPWR.n15 9.3005
R119 VPWR.n27 VPWR.n26 9.3005
R120 VPWR.n28 VPWR.n14 9.3005
R121 VPWR.n29 VPWR.n13 9.3005
R122 VPWR.n31 VPWR.n30 9.3005
R123 VPWR.n32 VPWR.n12 9.3005
R124 VPWR.n34 VPWR.n33 9.3005
R125 VPWR.n35 VPWR.n11 9.3005
R126 VPWR.n37 VPWR.n36 9.3005
R127 VPWR.n39 VPWR.n38 9.3005
R128 VPWR.n40 VPWR.n8 9.3005
R129 VPWR.n42 VPWR.n41 9.3005
R130 VPWR.n43 VPWR.n7 9.3005
R131 VPWR.n45 VPWR.n44 9.3005
R132 VPWR.n46 VPWR.n6 9.3005
R133 VPWR.n48 VPWR.n47 9.3005
R134 VPWR.n49 VPWR.n5 9.3005
R135 VPWR.n51 VPWR.n50 9.3005
R136 VPWR.n52 VPWR.n3 9.3005
R137 VPWR.n55 VPWR.n54 9.3005
R138 VPWR.n56 VPWR.n2 9.3005
R139 VPWR.n58 VPWR.n57 9.3005
R140 VPWR.n59 VPWR.n0 9.3005
R141 VPWR.n61 VPWR.n60 7.12063
R142 VPWR.n36 VPWR.n10 6.87109
R143 VPWR.n19 VPWR.n18 6.75413
R144 VPWR.n53 VPWR.n52 2.31027
R145 VPWR.n39 VPWR.n10 1.78874
R146 VPWR.n20 VPWR.n19 0.589392
R147 VPWR.n61 VPWR.n0 0.148519
R148 VPWR.n20 VPWR.n16 0.120292
R149 VPWR.n24 VPWR.n16 0.120292
R150 VPWR.n25 VPWR.n24 0.120292
R151 VPWR.n26 VPWR.n25 0.120292
R152 VPWR.n26 VPWR.n14 0.120292
R153 VPWR.n14 VPWR.n13 0.120292
R154 VPWR.n31 VPWR.n13 0.120292
R155 VPWR.n32 VPWR.n31 0.120292
R156 VPWR.n33 VPWR.n32 0.120292
R157 VPWR.n33 VPWR.n11 0.120292
R158 VPWR.n37 VPWR.n11 0.120292
R159 VPWR.n38 VPWR.n37 0.120292
R160 VPWR.n38 VPWR.n8 0.120292
R161 VPWR.n42 VPWR.n8 0.120292
R162 VPWR.n43 VPWR.n42 0.120292
R163 VPWR.n44 VPWR.n43 0.120292
R164 VPWR.n44 VPWR.n6 0.120292
R165 VPWR.n48 VPWR.n6 0.120292
R166 VPWR.n49 VPWR.n48 0.120292
R167 VPWR.n50 VPWR.n49 0.120292
R168 VPWR.n50 VPWR.n3 0.120292
R169 VPWR.n55 VPWR.n3 0.120292
R170 VPWR.n56 VPWR.n55 0.120292
R171 VPWR.n57 VPWR.n56 0.120292
R172 VPWR.n57 VPWR.n0 0.120292
R173 VPWR VPWR.n61 0.114842
R174 a_1781_295.n2 a_1781_295.t1 696.909
R175 a_1781_295.n1 a_1781_295.n0 448.372
R176 a_1781_295.t0 a_1781_295.n2 285.67
R177 a_1781_295.n2 a_1781_295.n1 256.642
R178 a_1781_295.n1 a_1781_295.t2 159.172
R179 a_328_21.n2 a_328_21.n1 628.706
R180 a_328_21.n0 a_328_21.t3 269.921
R181 a_328_21.n1 a_328_21.t1 260.365
R182 a_328_21.n1 a_328_21.n0 200.93
R183 a_328_21.n0 a_328_21.t2 178.924
R184 a_328_21.n2 a_328_21.t0 129.492
R185 a_328_21.n3 a_328_21.n2 3.78896
R186 a_265_47.t0 a_265_47.t1 90.0005
R187 VGND.n59 VGND.t0 243.028
R188 VGND.n65 VGND.t1 223.571
R189 VGND.n57 VGND.t9 223.571
R190 VGND.n44 VGND.t10 223.571
R191 VGND.n28 VGND.n27 203.433
R192 VGND.n52 VGND.n51 200.361
R193 VGND.n15 VGND.n14 197.981
R194 VGND.n37 VGND.n36 185
R195 VGND.n21 VGND.t14 160.222
R196 VGND.n16 VGND.t6 155.905
R197 VGND.n19 VGND.t13 149.802
R198 VGND.n27 VGND.t8 55.7148
R199 VGND.n14 VGND.t11 45.7148
R200 VGND.n36 VGND.t3 42.0094
R201 VGND.n27 VGND.t12 40.0005
R202 VGND.n36 VGND.t2 38.5719
R203 VGND.n51 VGND.t4 38.5719
R204 VGND.n51 VGND.t5 38.5719
R205 VGND.n22 VGND.n20 34.6358
R206 VGND.n26 VGND.n11 34.6358
R207 VGND.n30 VGND.n29 34.6358
R208 VGND.n30 VGND.n9 34.6358
R209 VGND.n34 VGND.n9 34.6358
R210 VGND.n35 VGND.n34 34.6358
R211 VGND.n43 VGND.n42 34.6358
R212 VGND.n49 VGND.n5 34.6358
R213 VGND.n50 VGND.n49 34.6358
R214 VGND.n63 VGND.n1 34.6358
R215 VGND.n14 VGND.t7 34.506
R216 VGND.n64 VGND.n63 34.0711
R217 VGND.n59 VGND.n58 33.1299
R218 VGND.n52 VGND.n50 32.377
R219 VGND.n45 VGND.n5 30.214
R220 VGND.n21 VGND.n11 29.7417
R221 VGND.n56 VGND.n3 28.5534
R222 VGND.n38 VGND.n35 27.6309
R223 VGND.n19 VGND.n13 25.224
R224 VGND.n20 VGND.n19 22.2123
R225 VGND.n15 VGND.n13 17.6946
R226 VGND.n59 VGND.n1 17.3181
R227 VGND.n58 VGND.n57 16.1005
R228 VGND.n52 VGND.n3 14.3064
R229 VGND.n29 VGND.n28 10.9181
R230 VGND.n66 VGND.n65 9.86521
R231 VGND.n42 VGND.n7 9.66183
R232 VGND.n64 VGND.n0 9.3005
R233 VGND.n63 VGND.n62 9.3005
R234 VGND.n61 VGND.n1 9.3005
R235 VGND.n60 VGND.n59 9.3005
R236 VGND.n58 VGND.n2 9.3005
R237 VGND.n56 VGND.n55 9.3005
R238 VGND.n54 VGND.n3 9.3005
R239 VGND.n53 VGND.n52 9.3005
R240 VGND.n50 VGND.n4 9.3005
R241 VGND.n49 VGND.n48 9.3005
R242 VGND.n47 VGND.n5 9.3005
R243 VGND.n46 VGND.n45 9.3005
R244 VGND.n43 VGND.n6 9.3005
R245 VGND.n42 VGND.n41 9.3005
R246 VGND.n40 VGND.n7 9.3005
R247 VGND.n39 VGND.n38 9.3005
R248 VGND.n35 VGND.n8 9.3005
R249 VGND.n34 VGND.n33 9.3005
R250 VGND.n32 VGND.n9 9.3005
R251 VGND.n31 VGND.n30 9.3005
R252 VGND.n29 VGND.n10 9.3005
R253 VGND.n26 VGND.n25 9.3005
R254 VGND.n24 VGND.n11 9.3005
R255 VGND.n23 VGND.n22 9.3005
R256 VGND.n20 VGND.n12 9.3005
R257 VGND.n19 VGND.n18 9.3005
R258 VGND.n17 VGND.n13 9.3005
R259 VGND.n44 VGND.n43 8.50873
R260 VGND.n65 VGND.n64 8.09462
R261 VGND.n16 VGND.n15 6.75413
R262 VGND.n38 VGND.n37 4.9623
R263 VGND.n22 VGND.n21 4.89462
R264 VGND.n28 VGND.n26 4.89462
R265 VGND.n45 VGND.n44 4.53868
R266 VGND.n57 VGND.n56 2.5005
R267 VGND.n37 VGND.n7 1.65443
R268 VGND.n17 VGND.n16 0.589392
R269 VGND.n18 VGND.n17 0.120292
R270 VGND.n18 VGND.n12 0.120292
R271 VGND.n23 VGND.n12 0.120292
R272 VGND.n24 VGND.n23 0.120292
R273 VGND.n25 VGND.n24 0.120292
R274 VGND.n25 VGND.n10 0.120292
R275 VGND.n31 VGND.n10 0.120292
R276 VGND.n32 VGND.n31 0.120292
R277 VGND.n33 VGND.n32 0.120292
R278 VGND.n33 VGND.n8 0.120292
R279 VGND.n39 VGND.n8 0.120292
R280 VGND.n40 VGND.n39 0.120292
R281 VGND.n41 VGND.n40 0.120292
R282 VGND.n41 VGND.n6 0.120292
R283 VGND.n46 VGND.n6 0.120292
R284 VGND.n47 VGND.n46 0.120292
R285 VGND.n48 VGND.n47 0.120292
R286 VGND.n48 VGND.n4 0.120292
R287 VGND.n53 VGND.n4 0.120292
R288 VGND.n54 VGND.n53 0.120292
R289 VGND.n55 VGND.n54 0.120292
R290 VGND.n55 VGND.n2 0.120292
R291 VGND.n60 VGND.n2 0.120292
R292 VGND.n61 VGND.n60 0.120292
R293 VGND.n62 VGND.n61 0.120292
R294 VGND.n62 VGND.n0 0.120292
R295 VGND.n66 VGND.n0 0.120292
R296 VGND VGND.n66 0.0226354
R297 VNB.t19 VNB.t21 3075.73
R298 VNB.t18 VNB.t20 2862.14
R299 VNB.t17 VNB.t5 2677.02
R300 VNB.t7 VNB.t13 2677.02
R301 VNB.t16 VNB.t8 2677.02
R302 VNB.t0 VNB.t16 2677.02
R303 VNB.t6 VNB.t1 2506.15
R304 VNB.t1 VNB.t10 1708.74
R305 VNB.t9 VNB.t14 1423.95
R306 VNB.t14 VNB.t19 1381.23
R307 VNB.t20 VNB.t12 1352.75
R308 VNB.t4 VNB.t6 1352.75
R309 VNB.t22 VNB.t0 1324.27
R310 VNB.t12 VNB.t11 1196.12
R311 VNB.t21 VNB.t18 1196.12
R312 VNB.t13 VNB.t2 1196.12
R313 VNB.t8 VNB.t7 1196.12
R314 VNB.t15 VNB.t22 1196.12
R315 VNB.t10 VNB.t9 1025.24
R316 VNB.t5 VNB.t4 1025.24
R317 VNB.t2 VNB.t17 1025.24
R318 VNB.t3 VNB.t15 1025.24
R319 VNB VNB.t3 925.567
R320 Q_N.n1 Q_N 591.806
R321 Q_N.n1 Q_N.n0 585
R322 Q_N.n2 Q_N.n1 585
R323 Q_N Q_N.n4 186.458
R324 Q_N.n4 Q_N.n3 185
R325 Q_N.n1 Q_N.t3 26.5955
R326 Q_N.n1 Q_N.t2 26.5955
R327 Q_N.n4 Q_N.t0 24.9236
R328 Q_N.n4 Q_N.t1 24.9236
R329 Q_N Q_N.n3 9.55999
R330 Q_N.n0 Q_N 6.80556
R331 Q_N Q_N.n2 6.80556
R332 Q_N.n0 Q_N 4.21316
R333 Q_N.n2 Q_N 4.21316
R334 Q_N.n3 Q_N 1.45873
R335 a_652_47.t0 a_652_47.n5 663.644
R336 a_652_47.n3 a_652_47.t6 429.212
R337 a_652_47.n3 a_652_47.t5 419.243
R338 a_652_47.n0 a_652_47.t3 393.634
R339 a_652_47.n4 a_652_47.t7 316.05
R340 a_652_47.n2 a_652_47.t1 288.964
R341 a_652_47.n1 a_652_47.t4 249.397
R342 a_652_47.n2 a_652_47.n1 152
R343 a_652_47.n1 a_652_47.n0 105.025
R344 a_652_47.n0 a_652_47.t2 91.5805
R345 a_652_47.n4 a_652_47.n3 68.928
R346 a_652_47.n5 a_652_47.n2 30.2774
R347 a_652_47.n5 a_652_47.n4 10.4804
R348 a_2501_47.t1 a_2501_47.n2 404.825
R349 a_2501_47.n2 a_2501_47.t0 261.971
R350 a_2501_47.n0 a_2501_47.t2 212.081
R351 a_2501_47.n1 a_2501_47.t3 212.081
R352 a_2501_47.n2 a_2501_47.n1 184.858
R353 a_2501_47.n0 a_2501_47.t4 139.78
R354 a_2501_47.n1 a_2501_47.t5 139.78
R355 a_2501_47.n1 a_2501_47.n0 61.346
R356 Q.n0 Q 591.207
R357 Q.n1 Q.n0 585
R358 Q.n5 Q.n4 185
R359 Q.n0 Q.t3 26.5955
R360 Q.n0 Q.t2 26.5955
R361 Q.n4 Q.t1 24.9236
R362 Q.n4 Q.t0 24.9236
R363 Q.n3 Q 15.9294
R364 Q Q.n5 12.6066
R365 Q.n2 Q 11.249
R366 Q.n1 Q 6.98232
R367 Q Q.n1 6.20656
R368 Q.n3 Q 3.41383
R369 Q Q.n2 2.84494
R370 Q Q.n3 2.32777
R371 Q.n2 Q 1.93989
R372 Q.n5 Q 0.582318
R373 a_1090_47.t0 a_1090_47.t1 60.0005
R374 SCD.n0 SCD.t0 299.433
R375 SCD.n0 SCD.t1 206.245
R376 SCD.n1 SCD.n0 152
R377 SCD.n1 SCD 19.828
R378 SCD SCD.n1 14.3064
R379 a_27_369.n0 a_27_369.t1 1323.74
R380 a_27_369.n0 a_27_369.t0 123.291
R381 a_27_369.n1 a_27_369.n0 3.78896
R382 SET_B.n1 SET_B.t1 358.397
R383 SET_B.n0 SET_B.t2 357.659
R384 SET_B.n2 SET_B.n1 219.648
R385 SET_B.n1 SET_B.t3 170.196
R386 SET_B.n0 SET_B.t0 166.577
R387 SET_B.n2 SET_B.n0 159
R388 SET_B SET_B.n2 3.4005
R389 a_1132_21.n0 a_1132_21.t1 892.923
R390 a_1132_21.t0 a_1132_21.n1 419.579
R391 a_1132_21.n1 a_1132_21.n0 201.407
R392 a_1132_21.n0 a_1132_21.t3 139.55
R393 a_1132_21.n1 a_1132_21.t2 129.338
R394 a_1517_47.t0 a_1517_47.t1 136.875
R395 SCE.n1 SCE.t2 296.43
R396 SCE.n0 SCE.t3 263.18
R397 SCE.n0 SCE.t0 231.73
R398 SCE.n1 SCE.t1 203.244
R399 SCE.n2 SCE.n1 173.137
R400 SCE.n2 SCE.n0 154.744
R401 SCE SCE.n2 3.88621
R402 a_109_47.t0 a_109_47.t1 60.0005
R403 a_1885_47.t0 a_1885_47.t1 100.001
R404 D.n0 D.t0 373.283
R405 D.n1 D.n0 152
R406 D.n0 D.t1 132.282
R407 D.n1 D 23.1303
R408 D D.n1 7.41103
R409 a_193_369.t0 a_193_369.t1 64.6411
R410 a_1525_329.t0 a_1525_329.t1 49.2505
R411 a_1813_47.t0 a_1813_47.t1 60.0005
R412 a_1350_47.t0 a_1350_47.t1 60.0005
R413 CLK.n0 CLK.t1 248.458
R414 CLK.n0 CLK.t0 216.869
R415 CLK.n1 CLK.n0 152
R416 CLK.n1 CLK 18.1413
R417 CLK CLK.n1 2.90959
R418 a_1102_413.t0 a_1102_413.t1 140.714
C0 Q VGND 0.142748f
C1 Q VPWR 0.196711f
C2 Q_N VGND 0.162855f
C3 Q SET_B 6.54e-20
C4 VGND VPWR 0.159441f
C5 Q_N VPWR 0.222201f
C6 SET_B VGND 0.043001f
C7 SET_B Q_N 2.38e-19
C8 D VGND 0.00863f
C9 SET_B VPWR 0.101852f
C10 D VPWR 0.008091f
C11 CLK VGND 0.040824f
C12 CLK VPWR 0.038784f
C13 VGND SCE 0.1436f
C14 VPWR SCE 0.065329f
C15 VPB Q 0.005913f
C16 D SCE 0.202134f
C17 SCD VGND 0.045183f
C18 VPB Q_N 0.00554f
C19 SCD VPWR 0.016342f
C20 CLK SCE 0.095776f
C21 VPB VGND 0.024942f
C22 VPB VPWR 0.329773f
C23 VPB SET_B 0.203809f
C24 VPB D 0.045769f
C25 VPB CLK 0.082276f
C26 SCD SCE 0.170177f
C27 VPB SCE 0.129094f
C28 VPB SCD 0.070898f
C29 a_1723_413# VPWR 8.96e-19
C30 SET_B a_1723_413# 2.84e-19
C31 Q VNB 0.024421f
C32 Q_N VNB 0.003971f
C33 VGND VNB 1.59881f
C34 VPWR VNB 1.27614f
C35 SET_B VNB 0.221463f
C36 CLK VNB 0.139079f
C37 D VNB 0.106116f
C38 SCE VNB 0.252516f
C39 SCD VNB 0.205442f
C40 VPB VNB 2.81966f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfsbp_1 SCD CLK Q_N D SET_B SCE Q VPWR VGND VPB VNB
X0 Q.t1 a_2412_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 a_1129_21.t1 a_997_413.t4 VPWR.t11 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.0924 ps=0.86 w=0.42 l=0.15
X2 VPWR.t10 SCD.t0 a_27_369.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_1081_413# a_643_369.t2 a_997_413.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1587_329# SET_B.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.10395 ps=0.915 w=0.42 l=0.15
X5 a_809_369.t1 a_643_369.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_997_413.t2 a_809_369.t2 a_181_47.t3 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_1770_295.t0 a_1587_329# VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 Q_N.t0 a_1587_329# VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 VPWR.t8 SET_B.t1 a_1129_21.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.27 as=0.07035 ps=0.755 w=0.42 l=0.15
X10 Q_N.t1 a_1587_329# VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_181_47.t4 SCE.t0 a_109_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 a_1514_47# a_997_413.t5 VGND.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.2224 pd=1.335 as=0.09575 ps=0.965 w=0.64 l=0.15
X13 VPWR.t1 a_1770_295.t2 a_1712_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.10395 pd=0.915 as=0.0609 ps=0.71 w=0.42 l=0.15
X14 VGND SET_B a_1347_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09575 pd=0.965 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 Q.t0 a_2412_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X16 a_27_369.t0 a_319_21.t2 a_181_47.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X17 VGND.t0 SCE.t1 a_319_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_181_47.t1 D.t0 a_193_369.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X19 a_265_47.t1 D.t1 a_181_47.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_997_413.t0 a_643_369.t4 a_181_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VGND.t5 a_1587_329# a_2412_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X22 a_1087_47# a_809_369.t3 a_997_413.t3 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_369.t0 SCE.t2 VPWR.t13 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_809_369.t0 a_643_369.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 VPWR.t2 SCE.t3 a_319_21.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 VGND SET_B a_1879_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08505 pd=0.825 as=0.1029 ps=0.91 w=0.42 l=0.15
X27 VPWR.t5 a_1587_329# a_2412_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 VPWR.t9 CLK.t0 a_643_369.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 a_1514_329# a_997_413.t6 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0903 pd=1.055 as=0.1428 ps=1.27 w=0.84 l=0.15
X30 a_1712_413.t1 a_809_369.t4 a_1587_329# VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.15225 ps=1.315 w=0.42 l=0.15
X31 VGND.t1 a_319_21.t3 a_265_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 VGND.t9 CLK.t1 a_643_369.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 a_1770_295.t1 a_1587_329# VGND.t7 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08505 ps=0.825 w=0.42 l=0.15
X34 a_109_47.t1 SCD.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_2412_47.t0 a_2412_47.n1 398.825
R1 a_2412_47.n1 a_2412_47.t1 257.401
R2 a_2412_47.n0 a_2412_47.t3 241.536
R3 a_2412_47.n1 a_2412_47.n0 177.213
R4 a_2412_47.n0 a_2412_47.t2 169.237
R5 VGND.n46 VGND.t1 259.166
R6 VGND.n18 VGND.t7 244.278
R7 VGND.n44 VGND.t0 237.877
R8 VGND.n53 VGND.t4 237.506
R9 VGND.n26 VGND.t8 227.01
R10 VGND.n14 VGND.n12 218.172
R11 VGND.n40 VGND.n39 199.865
R12 VGND.n13 VGND.t6 160.014
R13 VGND.n12 VGND.t5 54.2862
R14 VGND.n39 VGND.t3 38.5719
R15 VGND.n39 VGND.t9 38.5719
R16 VGND.n17 VGND.n11 34.6358
R17 VGND.n20 VGND.n19 34.6358
R18 VGND.n20 VGND.n9 34.6358
R19 VGND.n24 VGND.n9 34.6358
R20 VGND.n25 VGND.n24 34.6358
R21 VGND.n32 VGND.n31 34.6358
R22 VGND.n37 VGND.n5 34.6358
R23 VGND.n38 VGND.n37 34.6358
R24 VGND.n47 VGND.n45 34.6358
R25 VGND.n51 VGND.n1 34.6358
R26 VGND.n52 VGND.n51 34.6358
R27 VGND.n40 VGND.n38 32.377
R28 VGND.n27 VGND.n25 32.1993
R29 VGND.n44 VGND.n3 31.624
R30 VGND.n19 VGND.n18 31.2476
R31 VGND.n33 VGND.n5 27.3528
R32 VGND.n12 VGND.t2 25.9346
R33 VGND.n13 VGND.n11 23.3417
R34 VGND.n33 VGND.n32 16.6884
R35 VGND.n46 VGND.n1 16.1887
R36 VGND.n53 VGND.n52 15.8123
R37 VGND.n40 VGND.n3 13.5534
R38 VGND.n45 VGND.n44 12.0476
R39 VGND.n31 VGND.n7 10.5755
R40 VGND.n54 VGND.n53 9.3005
R41 VGND.n52 VGND.n0 9.3005
R42 VGND.n51 VGND.n50 9.3005
R43 VGND.n49 VGND.n1 9.3005
R44 VGND.n48 VGND.n47 9.3005
R45 VGND.n45 VGND.n2 9.3005
R46 VGND.n44 VGND.n43 9.3005
R47 VGND.n42 VGND.n3 9.3005
R48 VGND.n41 VGND.n40 9.3005
R49 VGND.n38 VGND.n4 9.3005
R50 VGND.n37 VGND.n36 9.3005
R51 VGND.n35 VGND.n5 9.3005
R52 VGND.n34 VGND.n33 9.3005
R53 VGND.n32 VGND.n6 9.3005
R54 VGND.n31 VGND.n30 9.3005
R55 VGND.n29 VGND.n7 9.3005
R56 VGND.n28 VGND.n27 9.3005
R57 VGND.n25 VGND.n8 9.3005
R58 VGND.n24 VGND.n23 9.3005
R59 VGND.n22 VGND.n9 9.3005
R60 VGND.n21 VGND.n20 9.3005
R61 VGND.n19 VGND.n10 9.3005
R62 VGND.n17 VGND.n16 9.3005
R63 VGND.n15 VGND.n11 9.3005
R64 VGND.n14 VGND.n13 7.38075
R65 VGND.n27 VGND.n26 5.17803
R66 VGND.n47 VGND.n46 4.89462
R67 VGND.n18 VGND.n17 3.38874
R68 VGND.n26 VGND.n7 1.4387
R69 VGND.n15 VGND.n14 0.206847
R70 VGND.n16 VGND.n15 0.120292
R71 VGND.n16 VGND.n10 0.120292
R72 VGND.n21 VGND.n10 0.120292
R73 VGND.n22 VGND.n21 0.120292
R74 VGND.n23 VGND.n22 0.120292
R75 VGND.n23 VGND.n8 0.120292
R76 VGND.n28 VGND.n8 0.120292
R77 VGND.n29 VGND.n28 0.120292
R78 VGND.n30 VGND.n29 0.120292
R79 VGND.n30 VGND.n6 0.120292
R80 VGND.n34 VGND.n6 0.120292
R81 VGND.n35 VGND.n34 0.120292
R82 VGND.n36 VGND.n35 0.120292
R83 VGND.n36 VGND.n4 0.120292
R84 VGND.n41 VGND.n4 0.120292
R85 VGND.n42 VGND.n41 0.120292
R86 VGND.n43 VGND.n42 0.120292
R87 VGND.n43 VGND.n2 0.120292
R88 VGND.n48 VGND.n2 0.120292
R89 VGND.n49 VGND.n48 0.120292
R90 VGND.n50 VGND.n49 0.120292
R91 VGND.n50 VGND.n0 0.120292
R92 VGND.n54 VGND.n0 0.120292
R93 VGND VGND.n54 0.0213333
R94 Q.n1 Q 593.095
R95 Q.n1 Q.n0 585
R96 Q.n2 Q.n1 585
R97 Q.n5 Q.t1 129.036
R98 Q.n1 Q.t0 26.5955
R99 Q.n4 Q 19.3735
R100 Q.n0 Q 8.09462
R101 Q Q.n5 6.83238
R102 Q.n3 Q.n2 6.21226
R103 Q.n5 Q 5.70906
R104 Q.n0 Q 4.70638
R105 Q.n2 Q 4.70638
R106 Q.n4 Q 4.15185
R107 Q Q.n3 3.45996
R108 Q Q.n4 2.25932
R109 Q.n3 Q 1.88285
R110 VNB.t9 VNB.t6 8600.65
R111 VNB.t13 VNB.t9 6080.26
R112 VNB.t2 VNB.t1 2762.46
R113 VNB.t8 VNB.t7 2677.02
R114 VNB.t6 VNB.t8 2677.02
R115 VNB.t4 VNB.t0 2677.02
R116 VNB.t1 VNB.t10 2677.02
R117 VNB.t7 VNB.t3 1352.75
R118 VNB.t0 VNB.t13 1196.12
R119 VNB.t10 VNB.t4 1196.12
R120 VNB.t12 VNB.t2 1196.12
R121 VNB.t11 VNB.t12 1196.12
R122 VNB.t5 VNB.t11 1025.24
R123 VNB VNB.t5 911.327
R124 a_997_413.n5 a_997_413.n0 662.052
R125 a_997_413.n3 a_997_413.t4 583.074
R126 a_997_413.n1 a_997_413.t6 267.243
R127 a_997_413.n3 a_997_413.n2 251.078
R128 a_997_413.n6 a_997_413.n5 234.409
R129 a_997_413.n4 a_997_413.n1 196.618
R130 a_997_413.n1 a_997_413.t5 170.843
R131 a_997_413.n4 a_997_413.n3 152
R132 a_997_413.n0 a_997_413.t1 63.3219
R133 a_997_413.n0 a_997_413.t2 63.3219
R134 a_997_413.n5 a_997_413.n4 46.7187
R135 a_997_413.n6 a_997_413.t3 38.5719
R136 a_997_413.t0 a_997_413.n6 38.5719
R137 VPWR.n45 VPWR.t2 731.903
R138 VPWR.n34 VPWR.t11 713.88
R139 VPWR.n21 VPWR.t6 663.062
R140 VPWR.n52 VPWR.n1 603.433
R141 VPWR.n5 VPWR.n4 598.965
R142 VPWR.n23 VPWR.n14 598.965
R143 VPWR.n10 VPWR.n9 585
R144 VPWR.n18 VPWR.n17 335.767
R145 VPWR.n16 VPWR.t7 255.905
R146 VPWR.n14 VPWR.t1 168.857
R147 VPWR.n9 VPWR.t12 87.9469
R148 VPWR.n9 VPWR.t8 84.4291
R149 VPWR.n14 VPWR.t4 63.3219
R150 VPWR.n17 VPWR.t5 58.4849
R151 VPWR.n1 VPWR.t13 41.5552
R152 VPWR.n1 VPWR.t10 41.5552
R153 VPWR.n4 VPWR.t0 41.5552
R154 VPWR.n4 VPWR.t9 41.5552
R155 VPWR.n46 VPWR.n2 34.6358
R156 VPWR.n50 VPWR.n2 34.6358
R157 VPWR.n51 VPWR.n50 34.6358
R158 VPWR.n38 VPWR.n7 34.6358
R159 VPWR.n39 VPWR.n38 34.6358
R160 VPWR.n40 VPWR.n39 34.6358
R161 VPWR.n27 VPWR.n12 34.6358
R162 VPWR.n28 VPWR.n27 34.6358
R163 VPWR.n40 VPWR.n5 33.5064
R164 VPWR.n17 VPWR.t3 31.663
R165 VPWR.n45 VPWR.n44 31.624
R166 VPWR.n34 VPWR.n33 29.7417
R167 VPWR.n52 VPWR.n51 28.9887
R168 VPWR.n33 VPWR.n32 27.577
R169 VPWR.n23 VPWR.n22 27.4829
R170 VPWR.n21 VPWR.n20 25.977
R171 VPWR.n20 VPWR.n16 23.3417
R172 VPWR.n22 VPWR.n21 18.4476
R173 VPWR.n23 VPWR.n12 16.9417
R174 VPWR.n34 VPWR.n7 14.6829
R175 VPWR.n29 VPWR.n28 13.7417
R176 VPWR.n46 VPWR.n45 12.0476
R177 VPWR.n44 VPWR.n5 10.9181
R178 VPWR.n20 VPWR.n19 9.3005
R179 VPWR.n21 VPWR.n15 9.3005
R180 VPWR.n22 VPWR.n13 9.3005
R181 VPWR.n24 VPWR.n23 9.3005
R182 VPWR.n25 VPWR.n12 9.3005
R183 VPWR.n27 VPWR.n26 9.3005
R184 VPWR.n28 VPWR.n11 9.3005
R185 VPWR.n30 VPWR.n29 9.3005
R186 VPWR.n32 VPWR.n31 9.3005
R187 VPWR.n33 VPWR.n8 9.3005
R188 VPWR.n35 VPWR.n34 9.3005
R189 VPWR.n36 VPWR.n7 9.3005
R190 VPWR.n38 VPWR.n37 9.3005
R191 VPWR.n39 VPWR.n6 9.3005
R192 VPWR.n41 VPWR.n40 9.3005
R193 VPWR.n42 VPWR.n5 9.3005
R194 VPWR.n44 VPWR.n43 9.3005
R195 VPWR.n45 VPWR.n3 9.3005
R196 VPWR.n47 VPWR.n46 9.3005
R197 VPWR.n48 VPWR.n2 9.3005
R198 VPWR.n50 VPWR.n49 9.3005
R199 VPWR.n51 VPWR.n0 9.3005
R200 VPWR.n29 VPWR.n10 7.90638
R201 VPWR.n18 VPWR.n16 7.39033
R202 VPWR.n53 VPWR.n52 7.12063
R203 VPWR.n32 VPWR.n10 0.753441
R204 VPWR.n19 VPWR.n18 0.197686
R205 VPWR.n53 VPWR.n0 0.148519
R206 VPWR.n19 VPWR.n15 0.120292
R207 VPWR.n15 VPWR.n13 0.120292
R208 VPWR.n24 VPWR.n13 0.120292
R209 VPWR.n25 VPWR.n24 0.120292
R210 VPWR.n26 VPWR.n25 0.120292
R211 VPWR.n26 VPWR.n11 0.120292
R212 VPWR.n30 VPWR.n11 0.120292
R213 VPWR.n31 VPWR.n30 0.120292
R214 VPWR.n31 VPWR.n8 0.120292
R215 VPWR.n35 VPWR.n8 0.120292
R216 VPWR.n36 VPWR.n35 0.120292
R217 VPWR.n37 VPWR.n36 0.120292
R218 VPWR.n37 VPWR.n6 0.120292
R219 VPWR.n41 VPWR.n6 0.120292
R220 VPWR.n42 VPWR.n41 0.120292
R221 VPWR.n43 VPWR.n42 0.120292
R222 VPWR.n43 VPWR.n3 0.120292
R223 VPWR.n47 VPWR.n3 0.120292
R224 VPWR.n48 VPWR.n47 0.120292
R225 VPWR.n49 VPWR.n48 0.120292
R226 VPWR.n49 VPWR.n0 0.120292
R227 VPWR VPWR.n53 0.11354
R228 a_1129_21.n3 a_1129_21.n2 808.119
R229 a_1129_21.n2 a_1129_21.n1 336.712
R230 a_1129_21.n2 a_1129_21.n0 139.822
R231 a_1129_21.t0 a_1129_21.n3 84.4291
R232 a_1129_21.n3 a_1129_21.t1 72.7029
R233 VPB.t4 VPB.t17 651.091
R234 VPB.t16 VPB.t13 585.981
R235 VPB.t10 VPB.t9 559.346
R236 VPB.t9 VPB.t8 556.386
R237 VPB.t5 VPB.t10 556.386
R238 VPB.t0 VPB.t15 556.386
R239 VPB.t2 VPB.t12 556.386
R240 VPB.t7 VPB.t2 556.386
R241 VPB.t1 VPB.t5 381.776
R242 VPB.t11 VPB.t16 343.303
R243 VPB.t17 VPB.t11 287.072
R244 VPB.t8 VPB.t3 281.154
R245 VPB.t13 VPB.t1 260.437
R246 VPB.t15 VPB.t4 248.599
R247 VPB.t12 VPB.t0 248.599
R248 VPB.t6 VPB.t7 248.599
R249 VPB.t14 VPB.t18 248.599
R250 VPB.t18 VPB.t6 213.084
R251 VPB VPB.t14 189.409
R252 SCD.n0 SCD.t0 297.825
R253 SCD.n0 SCD.t1 204.639
R254 SCD.n1 SCD.n0 152
R255 SCD.n1 SCD 19.4467
R256 SCD SCD.n1 14.0313
R257 a_27_369.t0 a_27_369.t1 1468.53
R258 a_643_369.t0 a_643_369.n7 670.08
R259 a_643_369.n2 a_643_369.n0 424.721
R260 a_643_369.n2 a_643_369.n1 419.243
R261 a_643_369.n4 a_643_369.t4 393.634
R262 a_643_369.n3 a_643_369.t2 317.574
R263 a_643_369.n6 a_643_369.t1 291.962
R264 a_643_369.n5 a_643_369.t5 267.3
R265 a_643_369.n6 a_643_369.n5 152
R266 a_643_369.n5 a_643_369.n4 100.206
R267 a_643_369.n4 a_643_369.t3 91.5805
R268 a_643_369.n3 a_643_369.n2 42.3659
R269 a_643_369.n7 a_643_369.n6 30.0313
R270 a_643_369.n7 a_643_369.n3 10.6775
R271 SET_B.n1 SET_B.n0 352.901
R272 SET_B.n3 SET_B.n2 350.789
R273 SET_B.n4 SET_B.n3 228.845
R274 SET_B.n3 SET_B.t0 209.403
R275 SET_B.n1 SET_B.t1 167.094
R276 SET_B.n4 SET_B.n1 157.12
R277 SET_B SET_B.n4 2.90183
R278 a_809_369.t0 a_809_369.n4 672.456
R279 a_809_369.n3 a_809_369.t3 433.509
R280 a_809_369.n1 a_809_369.n0 383.459
R281 a_809_369.n3 a_809_369.t2 321.334
R282 a_809_369.n2 a_809_369.t1 274.921
R283 a_809_369.n2 a_809_369.n1 204.804
R284 a_809_369.n4 a_809_369.n3 182.673
R285 a_809_369.n1 a_809_369.t4 148.35
R286 a_809_369.n4 a_809_369.n2 2.5605
R287 a_181_47.n1 a_181_47.t3 692.5
R288 a_181_47.n3 a_181_47.n2 616.648
R289 a_181_47.n2 a_181_47.n0 415.272
R290 a_181_47.n1 a_181_47.t0 288.805
R291 a_181_47.n3 a_181_47.t2 41.5552
R292 a_181_47.t1 a_181_47.n3 41.5552
R293 a_181_47.n0 a_181_47.t5 38.5719
R294 a_181_47.n0 a_181_47.t4 38.5719
R295 a_181_47.n2 a_181_47.n1 22.626
R296 a_1770_295.t0 a_1770_295.n2 698.292
R297 a_1770_295.n1 a_1770_295.t2 458.437
R298 a_1770_295.n2 a_1770_295.t1 278.209
R299 a_1770_295.n2 a_1770_295.n1 258.38
R300 a_1770_295.n1 a_1770_295.n0 161.202
R301 Q_N.n1 Q_N 593.145
R302 Q_N.n1 Q_N.n0 585
R303 Q_N.n2 Q_N.n1 585
R304 Q_N.n3 Q_N.t1 129.312
R305 Q_N.n1 Q_N.t0 26.5955
R306 Q_N.n0 Q_N 8.14595
R307 Q_N Q_N.n2 8.14595
R308 Q_N.n3 Q_N 7.23019
R309 Q_N Q_N.n3 5.71727
R310 Q_N.n0 Q_N 5.04292
R311 Q_N.n2 Q_N 5.04292
R312 SCE.n1 SCE.t3 295.168
R313 SCE.n0 SCE.t2 263.493
R314 SCE.n0 SCE.t0 232.163
R315 SCE.n1 SCE.t1 201.982
R316 SCE.n2 SCE.n1 173.302
R317 SCE.n2 SCE.n0 154.744
R318 SCE SCE.n2 3.88621
R319 a_109_47.t0 a_109_47.t1 60.0005
R320 a_1712_413.t0 a_1712_413.t1 136.024
R321 a_319_21.t0 a_319_21.n1 754.953
R322 a_319_21.n0 a_319_21.t2 284.38
R323 a_319_21.n1 a_319_21.t1 259.56
R324 a_319_21.n0 a_319_21.t3 191.194
R325 a_319_21.n1 a_319_21.n0 152
R326 D.n0 D.t0 373.283
R327 D.n1 D.n0 152
R328 D.n0 D.t1 132.282
R329 D.n1 D 23.5434
R330 D D.n1 7.54336
R331 a_193_369.t0 a_193_369.t1 64.6411
R332 a_265_47.t0 a_265_47.t1 77.1434
R333 CLK.n0 CLK.t0 255.077
R334 CLK.n0 CLK.t1 218.642
R335 CLK.n1 CLK.n0 152
R336 CLK.n1 CLK 20.3641
R337 CLK CLK.n1 2.90959
C0 D SCE 0.201502f
C1 a_1587_329# Q_N 0.060734f
C2 a_1587_329# a_1514_47# 0.003753f
C3 a_1347_47# VGND 0.004877f
C4 VPB VPWR 0.299408f
C5 a_1807_47# VPWR 2.14e-19
C6 SCE VPWR 0.06207f
C7 CLK VPWR 0.03214f
C8 a_1587_329# a_1514_329# 4.67e-19
C9 SCE VPB 0.130323f
C10 VGND Q_N 0.099586f
C11 VGND a_1514_47# 0.022344f
C12 CLK VPB 0.079477f
C13 VGND SCD 0.046163f
C14 CLK SCE 0.090278f
C15 SET_B Q_N 1.89e-19
C16 a_1587_329# Q 0.004035f
C17 VGND a_1587_329# 0.276178f
C18 SET_B a_1587_329# 0.28381f
C19 Q_N VPWR 0.128905f
C20 SCD VPWR 0.017446f
C21 a_1587_329# VPWR 0.379027f
C22 a_1587_329# a_1879_47# 0.011245f
C23 a_1081_413# VPWR 9.08e-19
C24 SET_B a_1514_329# 1.44e-19
C25 VGND Q 0.090879f
C26 Q_N VPB 0.010465f
C27 VGND a_1087_47# 0.005178f
C28 SCD VPB 0.070598f
C29 SCD SCE 0.170067f
C30 a_1514_329# VPWR 0.005944f
C31 SET_B Q 7.09e-20
C32 VGND SET_B 0.046474f
C33 a_1587_329# VPB 0.288699f
C34 VGND D 0.008969f
C35 a_1587_329# a_1807_47# 0.004624f
C36 Q VPWR 0.119664f
C37 VGND VPWR 0.11403f
C38 VGND a_1879_47# 0.003135f
C39 SET_B VPWR 0.102581f
C40 D VPWR 0.007833f
C41 Q VPB 0.012103f
C42 VGND VPB 0.022743f
C43 VGND SCE 0.130889f
C44 VGND a_1807_47# 0.001719f
C45 a_1879_47# VPWR 6.22e-19
C46 VGND CLK 0.037001f
C47 SET_B VPB 0.210906f
C48 SET_B a_1807_47# 9.13e-19
C49 D VPB 0.043598f
C50 Q VNB 0.091437f
C51 Q_N VNB 0.007215f
C52 VGND VNB 1.47853f
C53 VPWR VNB 1.17013f
C54 SET_B VNB 0.233014f
C55 CLK VNB 0.137461f
C56 D VNB 0.104074f
C57 SCE VNB 0.254717f
C58 SCD VNB 0.204781f
C59 VPB VNB 2.64247f
C60 a_1587_329# VNB 0.478914f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtp_4 VPB VNB VPWR VGND SCE SCD D RESET_B CLK Q
X0 a_193_47.t0 a_27_47.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_780_389.t1 a_299_66.t2 a_620_389.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.82 as=0.1755 ps=1.19 w=0.54 l=0.15
X2 a_1245_303.t2 a_1079_413# VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.2184 ps=2.2 w=0.84 l=0.15
X3 VPWR.t11 a_1592_47.t4 a_1767_21.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VGND.t3 a_1767_21.t3 a_1701_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06705 ps=0.75 w=0.42 l=0.15
X5 a_1758_413.t1 a_193_47.t2 a_1592_47.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0546 pd=0.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1767_21.t2 a_1592_47.t5 a_1946_47.t1 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.05145 ps=0.665 w=0.42 l=0.15
X7 VGND.t0 SCD.t0 a_817_66.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.18
X8 a_538_389.t0 SCE.t0 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0702 pd=0.8 as=0.0729 ps=0.81 w=0.54 l=0.15
X9 VPWR.t1 SCD.t1 a_780_389.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.64 as=0.0756 ps=0.82 w=0.54 l=0.15
X10 VPWR.t5 SCE.t1 a_299_66.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.189 ps=1.78 w=0.54 l=0.15
X11 a_1767_21.t0 RESET_B.t0 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X12 a_193_47.t1 a_27_47.t3 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_620_389.t3 D.t0 a_569_119.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.110275 pd=1.065 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 VGND.t4 a_1767_21.t4 Q.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_1293_47.t1 a_1245_303.t4 a_1187_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0759 ps=0.8 w=0.42 l=0.15
X16 VPWR.t8 a_1767_21.t5 Q.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X17 a_620_389.t4 D.t1 a_538_389.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1755 pd=1.19 as=0.0702 ps=0.8 w=0.54 l=0.15
X18 Q.t4 a_1767_21.t6 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X19 a_569_119.t0 a_299_66.t3 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 VPWR.t4 a_1767_21.t7 a_1758_413.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0546 ps=0.68 w=0.42 l=0.15
X21 VGND.t8 RESET_B.t1 a_1293_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 Q.t1 a_1767_21.t8 VPWR.t12 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 Q.t3 a_1767_21.t9 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_1191_413.t0 RESET_B.t2 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1007 ps=0.94 w=0.42 l=0.15
X25 a_1079_413# a_27_47.t4 a_620_389.t0 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.063 pd=0.71 as=0.0936 ps=1.24 w=0.36 l=0.15
X26 a_1946_47.t0 RESET_B.t3 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.05145 pd=0.665 as=0.12495 ps=1.015 w=0.42 l=0.15
X27 a_1701_47.t1 a_27_47.t5 a_1592_47.t0 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X28 Q.t0 a_1767_21.t10 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X29 a_1592_47.t3 a_193_47.t3 a_1245_303.t1 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X30 VGND.t7 SCE.t2 a_299_66.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_1592_47.t1 a_27_47.t6 a_1245_303.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12075 ps=1.165 w=0.42 l=0.15
X32 a_1245_303.t3 a_1079_413# VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1346 ps=1.15 w=0.64 l=0.15
X33 a_1079_413# a_193_47.t4 a_620_389.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0861 pd=0.83 as=0.1533 ps=1.57 w=0.42 l=0.15
X34 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X35 a_817_66.t0 SCE.t3 a_620_389.t5 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.110275 ps=1.065 w=0.42 l=0.5
X36 VGND.t11 CLK.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n4 a_27_47.n3 532.726
R1 a_27_47.n2 a_27_47.t6 496.003
R2 a_27_47.t0 a_27_47.n0 391.175
R3 a_27_47.n4 a_27_47.t4 279.101
R4 a_27_47.n0 a_27_47.t1 271.212
R5 a_27_47.n1 a_27_47.t2 241.536
R6 a_27_47.n2 a_27_47.t5 199.762
R7 a_27_47.n5 a_27_47.n2 170.347
R8 a_27_47.n1 a_27_47.t3 169.237
R9 a_27_47.n5 a_27_47.n4 164.312
R10 a_27_47.n0 a_27_47.n1 152
R11 a_27_47.n0 a_27_47.n5 14.0789
R12 VPWR.n8 VPWR.t7 806.511
R13 VPWR.n36 VPWR.t1 700.982
R14 VPWR.n29 VPWR.t3 688.191
R15 VPWR.n16 VPWR.t11 663.062
R16 VPWR.n43 VPWR.n42 615.871
R17 VPWR.n50 VPWR.n1 604.394
R18 VPWR.n11 VPWR.n10 603.433
R19 VPWR.n15 VPWR.t12 250.464
R20 VPWR.n14 VPWR.n13 229.496
R21 VPWR.n10 VPWR.t4 114.918
R22 VPWR.n10 VPWR.t6 63.3219
R23 VPWR.n42 VPWR.t9 49.2505
R24 VPWR.n42 VPWR.t5 49.2505
R25 VPWR.n40 VPWR.n4 34.6358
R26 VPWR.n41 VPWR.n40 34.6358
R27 VPWR.n44 VPWR.n41 34.6358
R28 VPWR.n48 VPWR.n2 34.6358
R29 VPWR.n49 VPWR.n48 34.6358
R30 VPWR.n30 VPWR.n6 34.6358
R31 VPWR.n34 VPWR.n6 34.6358
R32 VPWR.n35 VPWR.n34 34.6358
R33 VPWR.n22 VPWR.n21 34.6358
R34 VPWR.n23 VPWR.n22 34.6358
R35 VPWR.n28 VPWR.n27 31.3563
R36 VPWR.n1 VPWR.t0 29.5505
R37 VPWR.n36 VPWR.n4 29.3652
R38 VPWR.n21 VPWR.n11 29.3652
R39 VPWR.n13 VPWR.t8 28.5655
R40 VPWR.n1 VPWR.t2 26.5955
R41 VPWR.n13 VPWR.t10 26.5955
R42 VPWR.n43 VPWR.n2 25.224
R43 VPWR.n23 VPWR.n8 22.9652
R44 VPWR.n50 VPWR.n49 21.8358
R45 VPWR.n17 VPWR.n11 21.0829
R46 VPWR.n16 VPWR.n15 20.3299
R47 VPWR.n30 VPWR.n29 19.7527
R48 VPWR.n27 VPWR.n8 18.4476
R49 VPWR.n17 VPWR.n16 17.3181
R50 VPWR.n36 VPWR.n35 15.0593
R51 VPWR.n44 VPWR.n43 9.41227
R52 VPWR.n16 VPWR.n12 9.3005
R53 VPWR.n18 VPWR.n17 9.3005
R54 VPWR.n19 VPWR.n11 9.3005
R55 VPWR.n21 VPWR.n20 9.3005
R56 VPWR.n22 VPWR.n9 9.3005
R57 VPWR.n24 VPWR.n23 9.3005
R58 VPWR.n25 VPWR.n8 9.3005
R59 VPWR.n27 VPWR.n26 9.3005
R60 VPWR.n28 VPWR.n7 9.3005
R61 VPWR.n31 VPWR.n30 9.3005
R62 VPWR.n32 VPWR.n6 9.3005
R63 VPWR.n34 VPWR.n33 9.3005
R64 VPWR.n35 VPWR.n5 9.3005
R65 VPWR.n37 VPWR.n36 9.3005
R66 VPWR.n38 VPWR.n4 9.3005
R67 VPWR.n40 VPWR.n39 9.3005
R68 VPWR.n41 VPWR.n3 9.3005
R69 VPWR.n45 VPWR.n44 9.3005
R70 VPWR.n46 VPWR.n2 9.3005
R71 VPWR.n48 VPWR.n47 9.3005
R72 VPWR.n49 VPWR.n0 9.3005
R73 VPWR.n51 VPWR.n50 7.18025
R74 VPWR.n15 VPWR.n14 6.64175
R75 VPWR.n29 VPWR.n28 2.70272
R76 VPWR.n14 VPWR.n12 0.568643
R77 VPWR.n51 VPWR.n0 0.147761
R78 VPWR.n18 VPWR.n12 0.120292
R79 VPWR.n19 VPWR.n18 0.120292
R80 VPWR.n20 VPWR.n19 0.120292
R81 VPWR.n20 VPWR.n9 0.120292
R82 VPWR.n24 VPWR.n9 0.120292
R83 VPWR.n25 VPWR.n24 0.120292
R84 VPWR.n26 VPWR.n25 0.120292
R85 VPWR.n26 VPWR.n7 0.120292
R86 VPWR.n31 VPWR.n7 0.120292
R87 VPWR.n32 VPWR.n31 0.120292
R88 VPWR.n33 VPWR.n32 0.120292
R89 VPWR.n33 VPWR.n5 0.120292
R90 VPWR.n37 VPWR.n5 0.120292
R91 VPWR.n38 VPWR.n37 0.120292
R92 VPWR.n39 VPWR.n38 0.120292
R93 VPWR.n39 VPWR.n3 0.120292
R94 VPWR.n45 VPWR.n3 0.120292
R95 VPWR.n46 VPWR.n45 0.120292
R96 VPWR.n47 VPWR.n46 0.120292
R97 VPWR.n47 VPWR.n0 0.120292
R98 VPWR VPWR.n51 0.113006
R99 a_193_47.n0 a_193_47.t3 342.533
R100 a_193_47.n2 a_193_47.n1 338.877
R101 a_193_47.t0 a_193_47.n4 332.233
R102 a_193_47.n0 a_193_47.t2 307.817
R103 a_193_47.n4 a_193_47.t1 302.798
R104 a_193_47.n2 a_193_47.t4 300.252
R105 a_193_47.n3 a_193_47.n2 15.9565
R106 a_193_47.n4 a_193_47.n3 13.0278
R107 a_193_47.n3 a_193_47.n0 11.9849
R108 VPB.t8 VPB.t5 917.446
R109 VPB.t3 VPB.t7 774.313
R110 VPB.t1 VPB.t8 637.548
R111 VPB.t16 VPB.t17 556.386
R112 VPB.t5 VPB.t11 556.386
R113 VPB.t15 VPB.t4 511.784
R114 VPB.t6 VPB.t10 313.707
R115 VPB.t11 VPB.t2 281.154
R116 VPB.t4 VPB.t1 275.084
R117 VPB.t7 VPB.t13 268.688
R118 VPB.t13 VPB.t15 262.291
R119 VPB.t0 VPB.t3 257.478
R120 VPB.t12 VPB.t14 254.518
R121 VPB.t2 VPB.t9 254.518
R122 VPB.t17 VPB.t12 248.599
R123 VPB.t10 VPB.t16 248.599
R124 VPB.t9 VPB.t6 242.679
R125 VPB VPB.t0 177.571
R126 a_299_66.n0 a_299_66.t2 1108.99
R127 a_299_66.t1 a_299_66.n0 700.674
R128 a_299_66.n0 a_299_66.t3 346.219
R129 a_299_66.n0 a_299_66.t0 288.474
R130 a_620_389.n0 a_620_389.t2 686.09
R131 a_620_389.n3 a_620_389.n2 599.683
R132 a_620_389.n0 a_620_389.t0 360.05
R133 a_620_389.n2 a_620_389.n1 276.555
R134 a_620_389.n3 a_620_389.t4 162.344
R135 a_620_389.n1 a_620_389.t5 106.636
R136 a_620_389.n2 a_620_389.n0 83.2005
R137 a_620_389.t1 a_620_389.n3 74.7875
R138 a_620_389.n1 a_620_389.t3 38.5724
R139 a_780_389.t0 a_780_389.t1 102.148
R140 a_1245_303.n4 a_1245_303.n3 644.628
R141 a_1245_303.n1 a_1245_303.t4 365.918
R142 a_1245_303.n3 a_1245_303.n2 269.793
R143 a_1245_303.n3 a_1245_303.n1 227.672
R144 a_1245_303.n1 a_1245_303.n0 158.392
R145 a_1245_303.n4 a_1245_303.t0 72.7029
R146 a_1245_303.n2 a_1245_303.t1 63.3338
R147 a_1245_303.t2 a_1245_303.n4 50.4231
R148 a_1245_303.n2 a_1245_303.t3 26.7713
R149 a_1592_47.n1 a_1592_47.t5 1025.84
R150 a_1592_47.n3 a_1592_47.n2 635.218
R151 a_1592_47.n1 a_1592_47.t4 412.283
R152 a_1592_47.n2 a_1592_47.n0 302.889
R153 a_1592_47.n2 a_1592_47.n1 220.894
R154 a_1592_47.n0 a_1592_47.t3 70.0005
R155 a_1592_47.t1 a_1592_47.n3 68.0124
R156 a_1592_47.n3 a_1592_47.t2 63.3219
R157 a_1592_47.n0 a_1592_47.t0 61.6672
R158 a_1767_21.n6 a_1767_21.t7 1015.03
R159 a_1767_21.n9 a_1767_21.n8 783.903
R160 a_1767_21.n7 a_1767_21.n6 257.036
R161 a_1767_21.n7 a_1767_21.t2 223.571
R162 a_1767_21.n2 a_1767_21.n0 212.081
R163 a_1767_21.n3 a_1767_21.t10 212.081
R164 a_1767_21.n4 a_1767_21.t5 212.081
R165 a_1767_21.n5 a_1767_21.t8 212.081
R166 a_1767_21.n6 a_1767_21.t3 178.585
R167 a_1767_21.n8 a_1767_21.n5 173.925
R168 a_1767_21.n2 a_1767_21.n1 139.78
R169 a_1767_21.n3 a_1767_21.t6 139.78
R170 a_1767_21.n4 a_1767_21.t4 139.78
R171 a_1767_21.n5 a_1767_21.t9 139.78
R172 a_1767_21.n8 a_1767_21.n7 64.0131
R173 a_1767_21.n9 a_1767_21.t1 63.3219
R174 a_1767_21.t0 a_1767_21.n9 63.3219
R175 a_1767_21.n4 a_1767_21.n3 62.8066
R176 a_1767_21.n3 a_1767_21.n2 61.346
R177 a_1767_21.n5 a_1767_21.n4 61.346
R178 a_1701_47.t0 a_1701_47.t1 93.5174
R179 VGND.n13 VGND.t2 290.289
R180 VGND.n43 VGND.t6 252.274
R181 VGND.n1 VGND.t7 241.996
R182 VGND.n36 VGND.t0 241.22
R183 VGND.n15 VGND.n14 216.678
R184 VGND.n11 VGND.n10 205.707
R185 VGND.n28 VGND.n8 199.739
R186 VGND.n50 VGND.n49 199.739
R187 VGND.n10 VGND.t9 117.144
R188 VGND.n8 VGND.t8 72.8576
R189 VGND.n8 VGND.t10 60.5809
R190 VGND.n10 VGND.t3 52.8576
R191 VGND.n18 VGND.n17 34.6358
R192 VGND.n19 VGND.n18 34.6358
R193 VGND.n23 VGND.n22 34.6358
R194 VGND.n24 VGND.n23 34.6358
R195 VGND.n24 VGND.n7 34.6358
R196 VGND.n30 VGND.n29 34.6358
R197 VGND.n30 VGND.n5 34.6358
R198 VGND.n34 VGND.n5 34.6358
R199 VGND.n35 VGND.n34 34.6358
R200 VGND.n37 VGND.n3 34.6358
R201 VGND.n41 VGND.n3 34.6358
R202 VGND.n42 VGND.n41 34.6358
R203 VGND.n48 VGND.n47 34.6358
R204 VGND.n17 VGND.n13 34.2593
R205 VGND.n14 VGND.t4 26.7697
R206 VGND.n28 VGND.n7 25.977
R207 VGND.n14 VGND.t1 24.9236
R208 VGND.n49 VGND.t5 24.9236
R209 VGND.n49 VGND.t11 24.9236
R210 VGND.n50 VGND.n48 22.9652
R211 VGND.n43 VGND.n42 19.9534
R212 VGND.n47 VGND.n1 19.9534
R213 VGND.n19 VGND.n11 19.577
R214 VGND.n29 VGND.n28 18.4476
R215 VGND.n22 VGND.n11 15.0593
R216 VGND.n43 VGND.n1 14.3064
R217 VGND.n48 VGND.n0 9.3005
R218 VGND.n47 VGND.n46 9.3005
R219 VGND.n45 VGND.n1 9.3005
R220 VGND.n44 VGND.n43 9.3005
R221 VGND.n17 VGND.n16 9.3005
R222 VGND.n18 VGND.n12 9.3005
R223 VGND.n20 VGND.n19 9.3005
R224 VGND.n22 VGND.n21 9.3005
R225 VGND.n23 VGND.n9 9.3005
R226 VGND.n25 VGND.n24 9.3005
R227 VGND.n26 VGND.n7 9.3005
R228 VGND.n28 VGND.n27 9.3005
R229 VGND.n29 VGND.n6 9.3005
R230 VGND.n31 VGND.n30 9.3005
R231 VGND.n32 VGND.n5 9.3005
R232 VGND.n34 VGND.n33 9.3005
R233 VGND.n35 VGND.n4 9.3005
R234 VGND.n38 VGND.n37 9.3005
R235 VGND.n39 VGND.n3 9.3005
R236 VGND.n41 VGND.n40 9.3005
R237 VGND.n42 VGND.n2 9.3005
R238 VGND.n15 VGND.n13 7.54862
R239 VGND.n51 VGND.n50 7.12063
R240 VGND.n37 VGND.n36 5.64756
R241 VGND.n36 VGND.n35 4.14168
R242 VGND.n16 VGND.n15 0.576163
R243 VGND.n51 VGND.n0 0.148519
R244 VGND.n16 VGND.n12 0.120292
R245 VGND.n20 VGND.n12 0.120292
R246 VGND.n21 VGND.n20 0.120292
R247 VGND.n21 VGND.n9 0.120292
R248 VGND.n25 VGND.n9 0.120292
R249 VGND.n26 VGND.n25 0.120292
R250 VGND.n27 VGND.n26 0.120292
R251 VGND.n27 VGND.n6 0.120292
R252 VGND.n31 VGND.n6 0.120292
R253 VGND.n32 VGND.n31 0.120292
R254 VGND.n33 VGND.n32 0.120292
R255 VGND.n33 VGND.n4 0.120292
R256 VGND.n38 VGND.n4 0.120292
R257 VGND.n39 VGND.n38 0.120292
R258 VGND.n40 VGND.n39 0.120292
R259 VGND.n40 VGND.n2 0.120292
R260 VGND.n44 VGND.n2 0.120292
R261 VGND.n45 VGND.n44 0.120292
R262 VGND.n46 VGND.n45 0.120292
R263 VGND.n46 VGND.n0 0.120292
R264 VGND VGND.n51 0.101821
R265 VNB.t6 VNB.t11 2933.33
R266 VNB.t18 VNB.t1 2748.22
R267 VNB.t0 VNB.t6 2747.16
R268 VNB.t7 VNB.t9 2677.02
R269 VNB.t9 VNB.t8 2512.82
R270 VNB.t4 VNB.t13 2121.68
R271 VNB.t10 VNB.t14 1879.61
R272 VNB.t16 VNB.t17 1863.06
R273 VNB.t12 VNB.t5 1552.1
R274 VNB.t17 VNB.t0 1453.45
R275 VNB.t5 VNB.t4 1366.99
R276 VNB.t14 VNB.t12 1352.75
R277 VNB.t3 VNB.t2 1224.6
R278 VNB.t1 VNB.t3 1196.12
R279 VNB.t15 VNB.t7 1196.12
R280 VNB.t13 VNB.t18 1124.92
R281 VNB.t11 VNB.t10 1025.24
R282 VNB.t8 VNB.t16 951.351
R283 VNB VNB.t15 726.215
R284 a_1758_413.t0 a_1758_413.t1 121.953
R285 a_1946_47.t0 a_1946_47.t1 70.0005
R286 SCD.n0 SCD.t0 248.767
R287 SCD.n0 SCD.t1 191.998
R288 SCD SCD.n0 155.072
R289 a_817_66.t1 a_817_66.t0 60.0005
R290 SCE.t2 SCE.t3 729.321
R291 SCE.n0 SCE.t0 273.134
R292 SCE.n1 SCE.t2 215.901
R293 SCE SCE.n1 159.054
R294 SCE.n1 SCE.n0 145.296
R295 SCE.n0 SCE.t1 138.173
R296 a_538_389.t0 a_538_389.t1 94.8524
R297 Q Q.n0 586.723
R298 Q.n6 Q.n0 585
R299 Q.n3 Q.t0 384.11
R300 Q.n3 Q.t4 228.612
R301 Q.n2 Q.n1 185
R302 Q.n5 Q 89.6005
R303 Q.n4 Q.n3 31.8066
R304 Q.n0 Q.t2 26.5955
R305 Q.n0 Q.t1 26.5955
R306 Q.n1 Q.t5 24.9236
R307 Q.n1 Q.t3 24.9236
R308 Q.n5 Q.n4 24.3815
R309 Q.n4 Q.n2 20.3141
R310 Q Q.n5 16.0005
R311 Q Q.n6 15.0159
R312 Q.n2 Q 10.0928
R313 Q.n6 Q 1.72358
R314 Q.n5 Q 0.738962
R315 RESET_B.n1 RESET_B.t0 2026.37
R316 RESET_B.n0 RESET_B.t2 398.99
R317 RESET_B.n1 RESET_B.t3 204.458
R318 RESET_B.n3 RESET_B.n0 163.06
R319 RESET_B.n2 RESET_B.n1 157.826
R320 RESET_B.n0 RESET_B.t1 136.21
R321 RESET_B.n4 RESET_B 11.2557
R322 RESET_B.n3 RESET_B.n2 9.43939
R323 RESET_B.n4 RESET_B.n3 9.30982
R324 RESET_B.n2 RESET_B 5.91708
R325 RESET_B RESET_B.n4 3.75222
R326 D.n0 D.t0 234.942
R327 D.n0 D.t1 164.25
R328 D D.n0 157.819
R329 a_569_119.t0 a_569_119.t1 60.0005
R330 a_1187_47.n0 a_1187_47.t0 9.47418
R331 a_1293_47.t0 a_1293_47.t1 60.0005
R332 CLK.n0 CLK.t0 428.579
R333 CLK.n0 CLK.t1 426.168
R334 CLK.n1 CLK.n0 152
R335 CLK.n1 CLK 10.4234
R336 CLK CLK.n1 2.01193
C0 VPWR VGND 0.086439f
C1 D VGND 0.001786f
C2 CLK VGND 0.017295f
C3 VPWR D 0.062452f
C4 CLK VPWR 0.01885f
C5 RESET_B Q 0.002838f
C6 SCD Q 5.45e-21
C7 VPB Q 0.010601f
C8 RESET_B SCD 4.26e-19
C9 RESET_B VPB 0.152772f
C10 SCE SCD 0.033759f
C11 SCE RESET_B 1.82e-19
C12 SCD VPB 0.06936f
C13 SCE VPB 0.182158f
C14 RESET_B a_1079_413# 0.146062f
C15 SCD a_1079_413# 2.16e-19
C16 VPB a_1079_413# 0.09595f
C17 VGND Q 0.192016f
C18 VPWR Q 0.370166f
C19 RESET_B VGND 0.27163f
C20 SCD VGND 0.069739f
C21 D Q 1.13e-21
C22 VPB VGND 0.012251f
C23 SCE VGND 0.086893f
C24 VPWR RESET_B 0.07406f
C25 VPWR SCD 0.01224f
C26 RESET_B D 8.56e-20
C27 D SCD 0.005659f
C28 VPWR VPB 0.285878f
C29 CLK RESET_B 2.16e-20
C30 D VPB 0.068911f
C31 SCE VPWR 0.066374f
C32 a_1079_413# VGND 0.126685f
C33 SCE D 0.051599f
C34 CLK VPB 0.040886f
C35 CLK SCE 2.38e-19
C36 VPWR a_1079_413# 0.068775f
C37 D a_1079_413# 2.79e-20
C38 Q VNB 0.045447f
C39 VGND VNB 1.42023f
C40 RESET_B VNB 0.269536f
C41 VPWR VNB 1.16632f
C42 SCD VNB 0.13368f
C43 D VNB 0.093585f
C44 SCE VNB 0.51427f
C45 CLK VNB 0.15698f
C46 VPB VNB 2.51881f
C47 a_1079_413# VNB 0.150381f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtp_2 VPB VNB VPWR VGND SCE SCD D RESET_B CLK Q
X0 a_193_47.t0 a_27_47.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_780_389.t1 a_299_66.t2 a_620_389.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.82 as=0.1755 ps=1.19 w=0.54 l=0.15
X2 a_1245_303.t1 a_1079_413# VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.2184 ps=2.2 w=0.84 l=0.15
X3 VPWR.t10 a_1592_47.t4 a_1767_21.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VGND.t10 a_1767_21.t3 a_1701_47.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06705 ps=0.75 w=0.42 l=0.15
X5 a_1758_413.t0 a_193_47.t2 a_1592_47.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0546 pd=0.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1767_21.t2 a_1592_47.t5 a_1946_47.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.05145 ps=0.665 w=0.42 l=0.15
X7 VGND.t1 SCD.t0 a_817_66.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.18
X8 a_538_389.t0 SCE.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0702 pd=0.8 as=0.0729 ps=0.81 w=0.54 l=0.15
X9 VPWR.t1 SCD.t1 a_780_389.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.64 as=0.0756 ps=0.82 w=0.54 l=0.15
X10 VPWR.t6 SCE.t1 a_299_66.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.189 ps=1.78 w=0.54 l=0.15
X11 a_1767_21.t0 RESET_B.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X12 a_193_47.t1 a_27_47.t3 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_620_389.t0 D.t0 a_569_119.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.110275 pd=1.065 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 VGND.t9 a_1767_21.t4 Q.t3 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_1293_47.t0 a_1245_303.t4 a_1187_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0759 ps=0.8 w=0.42 l=0.15
X16 VPWR.t8 a_1767_21.t5 Q.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X17 a_620_389.t5 D.t1 a_538_389.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1755 pd=1.19 as=0.0702 ps=0.8 w=0.54 l=0.15
X18 a_569_119.t0 a_299_66.t3 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 VPWR.t9 a_1767_21.t6 a_1758_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0546 ps=0.68 w=0.42 l=0.15
X20 VGND.t7 RESET_B.t1 a_1293_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 Q.t0 a_1767_21.t7 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 Q.t2 a_1767_21.t8 VGND.t8 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_1191_413# RESET_B.t2 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1007 ps=0.94 w=0.42 l=0.15
X24 a_1079_413# a_27_47.t4 a_620_389.t3 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.063 pd=0.71 as=0.0936 ps=1.24 w=0.36 l=0.15
X25 a_1946_47.t0 RESET_B.t3 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.05145 pd=0.665 as=0.12495 ps=1.015 w=0.42 l=0.15
X26 a_1701_47.t0 a_27_47.t5 a_1592_47.t1 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X27 a_1592_47.t2 a_193_47.t3 a_1245_303.t3 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X28 VGND.t2 SCE.t2 a_299_66.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_1592_47.t0 a_27_47.t6 a_1245_303.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12075 ps=1.165 w=0.42 l=0.15
X30 a_1245_303.t0 a_1079_413# VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1346 ps=1.15 w=0.64 l=0.15
X31 a_1079_413# a_193_47.t4 a_620_389.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0861 pd=0.83 as=0.1533 ps=1.57 w=0.42 l=0.15
X32 VPWR.t5 CLK.t0 a_27_47.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X33 a_817_66.t1 SCE.t3 a_620_389.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.110275 ps=1.065 w=0.42 l=0.5
X34 VGND.t5 CLK.t1 a_27_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n4 a_27_47.n3 532.726
R1 a_27_47.n2 a_27_47.t6 496.003
R2 a_27_47.t0 a_27_47.n0 391.175
R3 a_27_47.n4 a_27_47.t4 279.101
R4 a_27_47.n0 a_27_47.t1 271.212
R5 a_27_47.n1 a_27_47.t2 241.536
R6 a_27_47.n2 a_27_47.t5 199.762
R7 a_27_47.n5 a_27_47.n2 170.347
R8 a_27_47.n1 a_27_47.t3 169.237
R9 a_27_47.n5 a_27_47.n4 164.312
R10 a_27_47.n0 a_27_47.n1 152
R11 a_27_47.n0 a_27_47.n5 14.0789
R12 VPWR.n8 VPWR.t0 806.511
R13 VPWR.n35 VPWR.t1 700.982
R14 VPWR.n28 VPWR.t11 688.191
R15 VPWR.n15 VPWR.t10 663.062
R16 VPWR.n42 VPWR.n41 615.871
R17 VPWR.n49 VPWR.n1 604.394
R18 VPWR.n11 VPWR.n10 603.433
R19 VPWR.n13 VPWR.t8 259.166
R20 VPWR.n14 VPWR.t7 250.464
R21 VPWR.n10 VPWR.t9 114.918
R22 VPWR.n10 VPWR.t3 63.3219
R23 VPWR.n41 VPWR.t2 49.2505
R24 VPWR.n41 VPWR.t6 49.2505
R25 VPWR.n39 VPWR.n4 34.6358
R26 VPWR.n40 VPWR.n39 34.6358
R27 VPWR.n43 VPWR.n40 34.6358
R28 VPWR.n47 VPWR.n2 34.6358
R29 VPWR.n48 VPWR.n47 34.6358
R30 VPWR.n29 VPWR.n6 34.6358
R31 VPWR.n33 VPWR.n6 34.6358
R32 VPWR.n34 VPWR.n33 34.6358
R33 VPWR.n21 VPWR.n20 34.6358
R34 VPWR.n22 VPWR.n21 34.6358
R35 VPWR.n27 VPWR.n26 31.3563
R36 VPWR.n1 VPWR.t5 29.5505
R37 VPWR.n35 VPWR.n4 29.3652
R38 VPWR.n20 VPWR.n11 29.3652
R39 VPWR.n1 VPWR.t4 26.5955
R40 VPWR.n42 VPWR.n2 25.224
R41 VPWR.n22 VPWR.n8 22.9652
R42 VPWR.n49 VPWR.n48 21.8358
R43 VPWR.n16 VPWR.n11 21.0829
R44 VPWR.n15 VPWR.n14 20.3299
R45 VPWR.n29 VPWR.n28 19.7527
R46 VPWR.n26 VPWR.n8 18.4476
R47 VPWR.n16 VPWR.n15 17.3181
R48 VPWR.n35 VPWR.n34 15.0593
R49 VPWR.n43 VPWR.n42 9.41227
R50 VPWR.n15 VPWR.n12 9.3005
R51 VPWR.n17 VPWR.n16 9.3005
R52 VPWR.n18 VPWR.n11 9.3005
R53 VPWR.n20 VPWR.n19 9.3005
R54 VPWR.n21 VPWR.n9 9.3005
R55 VPWR.n23 VPWR.n22 9.3005
R56 VPWR.n24 VPWR.n8 9.3005
R57 VPWR.n26 VPWR.n25 9.3005
R58 VPWR.n27 VPWR.n7 9.3005
R59 VPWR.n30 VPWR.n29 9.3005
R60 VPWR.n31 VPWR.n6 9.3005
R61 VPWR.n33 VPWR.n32 9.3005
R62 VPWR.n34 VPWR.n5 9.3005
R63 VPWR.n36 VPWR.n35 9.3005
R64 VPWR.n37 VPWR.n4 9.3005
R65 VPWR.n39 VPWR.n38 9.3005
R66 VPWR.n40 VPWR.n3 9.3005
R67 VPWR.n44 VPWR.n43 9.3005
R68 VPWR.n45 VPWR.n2 9.3005
R69 VPWR.n47 VPWR.n46 9.3005
R70 VPWR.n48 VPWR.n0 9.3005
R71 VPWR.n50 VPWR.n49 7.18025
R72 VPWR.n14 VPWR.n13 6.56401
R73 VPWR.n28 VPWR.n27 2.70272
R74 VPWR.n13 VPWR.n12 0.652261
R75 VPWR.n50 VPWR.n0 0.147761
R76 VPWR.n17 VPWR.n12 0.120292
R77 VPWR.n18 VPWR.n17 0.120292
R78 VPWR.n19 VPWR.n18 0.120292
R79 VPWR.n19 VPWR.n9 0.120292
R80 VPWR.n23 VPWR.n9 0.120292
R81 VPWR.n24 VPWR.n23 0.120292
R82 VPWR.n25 VPWR.n24 0.120292
R83 VPWR.n25 VPWR.n7 0.120292
R84 VPWR.n30 VPWR.n7 0.120292
R85 VPWR.n31 VPWR.n30 0.120292
R86 VPWR.n32 VPWR.n31 0.120292
R87 VPWR.n32 VPWR.n5 0.120292
R88 VPWR.n36 VPWR.n5 0.120292
R89 VPWR.n37 VPWR.n36 0.120292
R90 VPWR.n38 VPWR.n37 0.120292
R91 VPWR.n38 VPWR.n3 0.120292
R92 VPWR.n44 VPWR.n3 0.120292
R93 VPWR.n45 VPWR.n44 0.120292
R94 VPWR.n46 VPWR.n45 0.120292
R95 VPWR.n46 VPWR.n0 0.120292
R96 VPWR VPWR.n50 0.113006
R97 a_193_47.n0 a_193_47.t3 342.533
R98 a_193_47.n2 a_193_47.n1 338.877
R99 a_193_47.t0 a_193_47.n4 332.233
R100 a_193_47.n0 a_193_47.t2 307.817
R101 a_193_47.n4 a_193_47.t1 302.798
R102 a_193_47.n2 a_193_47.t4 300.252
R103 a_193_47.n3 a_193_47.n2 15.9565
R104 a_193_47.n4 a_193_47.n3 13.0278
R105 a_193_47.n3 a_193_47.n0 11.9849
R106 VPB.t9 VPB.t16 917.446
R107 VPB.t6 VPB.t8 774.313
R108 VPB.t1 VPB.t9 637.548
R109 VPB.t14 VPB.t11 556.386
R110 VPB.t16 VPB.t0 556.386
R111 VPB.t15 VPB.t4 511.784
R112 VPB.t13 VPB.t3 313.707
R113 VPB.t0 VPB.t5 281.154
R114 VPB.t4 VPB.t1 275.084
R115 VPB.t8 VPB.t2 268.688
R116 VPB.t2 VPB.t15 262.291
R117 VPB.t7 VPB.t6 257.478
R118 VPB.t5 VPB.t10 254.518
R119 VPB.t11 VPB.t12 248.599
R120 VPB.t3 VPB.t14 248.599
R121 VPB.t10 VPB.t13 242.679
R122 VPB VPB.t7 177.571
R123 a_299_66.n0 a_299_66.t2 1108.99
R124 a_299_66.t1 a_299_66.n0 700.674
R125 a_299_66.n0 a_299_66.t3 346.219
R126 a_299_66.n0 a_299_66.t0 288.474
R127 a_620_389.n0 a_620_389.t4 686.09
R128 a_620_389.n3 a_620_389.n2 599.683
R129 a_620_389.n0 a_620_389.t3 360.05
R130 a_620_389.n2 a_620_389.n1 276.555
R131 a_620_389.n3 a_620_389.t5 162.344
R132 a_620_389.n1 a_620_389.t1 106.636
R133 a_620_389.n2 a_620_389.n0 83.2005
R134 a_620_389.t2 a_620_389.n3 74.7875
R135 a_620_389.n1 a_620_389.t0 38.5724
R136 a_780_389.t0 a_780_389.t1 102.148
R137 a_1245_303.n4 a_1245_303.n3 644.628
R138 a_1245_303.n1 a_1245_303.t4 365.918
R139 a_1245_303.n3 a_1245_303.n2 269.793
R140 a_1245_303.n3 a_1245_303.n1 227.672
R141 a_1245_303.n1 a_1245_303.n0 158.392
R142 a_1245_303.n4 a_1245_303.t2 72.7029
R143 a_1245_303.n2 a_1245_303.t3 63.3338
R144 a_1245_303.t1 a_1245_303.n4 50.4231
R145 a_1245_303.n2 a_1245_303.t0 26.7713
R146 a_1592_47.n1 a_1592_47.t5 1025.84
R147 a_1592_47.n3 a_1592_47.n2 635.218
R148 a_1592_47.n1 a_1592_47.t4 412.283
R149 a_1592_47.n2 a_1592_47.n0 302.889
R150 a_1592_47.n2 a_1592_47.n1 220.894
R151 a_1592_47.n0 a_1592_47.t2 70.0005
R152 a_1592_47.t0 a_1592_47.n3 68.0124
R153 a_1592_47.n3 a_1592_47.t3 63.3219
R154 a_1592_47.n0 a_1592_47.t1 61.6672
R155 a_1767_21.n2 a_1767_21.t6 1015.03
R156 a_1767_21.n5 a_1767_21.n4 783.903
R157 a_1767_21.n3 a_1767_21.n2 257.036
R158 a_1767_21.n3 a_1767_21.t2 223.571
R159 a_1767_21.n0 a_1767_21.t5 212.081
R160 a_1767_21.n1 a_1767_21.t7 212.081
R161 a_1767_21.n2 a_1767_21.t3 178.585
R162 a_1767_21.n4 a_1767_21.n1 173.925
R163 a_1767_21.n0 a_1767_21.t4 139.78
R164 a_1767_21.n1 a_1767_21.t8 139.78
R165 a_1767_21.n4 a_1767_21.n3 64.0131
R166 a_1767_21.n5 a_1767_21.t1 63.3219
R167 a_1767_21.t0 a_1767_21.n5 63.3219
R168 a_1767_21.n1 a_1767_21.n0 61.346
R169 a_1701_47.t1 a_1701_47.t0 93.5174
R170 VGND.n14 VGND.t9 297.507
R171 VGND.n13 VGND.t8 290.289
R172 VGND.n42 VGND.t3 252.274
R173 VGND.n1 VGND.t2 241.996
R174 VGND.n35 VGND.t1 241.22
R175 VGND.n11 VGND.n10 205.707
R176 VGND.n27 VGND.n8 199.739
R177 VGND.n49 VGND.n48 199.739
R178 VGND.n10 VGND.t6 117.144
R179 VGND.n8 VGND.t7 72.8576
R180 VGND.n8 VGND.t0 60.5809
R181 VGND.n10 VGND.t10 52.8576
R182 VGND.n17 VGND.n16 34.6358
R183 VGND.n18 VGND.n17 34.6358
R184 VGND.n22 VGND.n21 34.6358
R185 VGND.n23 VGND.n22 34.6358
R186 VGND.n23 VGND.n7 34.6358
R187 VGND.n29 VGND.n28 34.6358
R188 VGND.n29 VGND.n5 34.6358
R189 VGND.n33 VGND.n5 34.6358
R190 VGND.n34 VGND.n33 34.6358
R191 VGND.n36 VGND.n3 34.6358
R192 VGND.n40 VGND.n3 34.6358
R193 VGND.n41 VGND.n40 34.6358
R194 VGND.n47 VGND.n46 34.6358
R195 VGND.n16 VGND.n13 34.2593
R196 VGND.n27 VGND.n7 25.977
R197 VGND.n48 VGND.t4 24.9236
R198 VGND.n48 VGND.t5 24.9236
R199 VGND.n49 VGND.n47 22.9652
R200 VGND.n42 VGND.n41 19.9534
R201 VGND.n46 VGND.n1 19.9534
R202 VGND.n18 VGND.n11 19.577
R203 VGND.n28 VGND.n27 18.4476
R204 VGND.n21 VGND.n11 15.0593
R205 VGND.n42 VGND.n1 14.3064
R206 VGND.n47 VGND.n0 9.3005
R207 VGND.n46 VGND.n45 9.3005
R208 VGND.n44 VGND.n1 9.3005
R209 VGND.n43 VGND.n42 9.3005
R210 VGND.n16 VGND.n15 9.3005
R211 VGND.n17 VGND.n12 9.3005
R212 VGND.n19 VGND.n18 9.3005
R213 VGND.n21 VGND.n20 9.3005
R214 VGND.n22 VGND.n9 9.3005
R215 VGND.n24 VGND.n23 9.3005
R216 VGND.n25 VGND.n7 9.3005
R217 VGND.n27 VGND.n26 9.3005
R218 VGND.n28 VGND.n6 9.3005
R219 VGND.n30 VGND.n29 9.3005
R220 VGND.n31 VGND.n5 9.3005
R221 VGND.n33 VGND.n32 9.3005
R222 VGND.n34 VGND.n4 9.3005
R223 VGND.n37 VGND.n36 9.3005
R224 VGND.n38 VGND.n3 9.3005
R225 VGND.n40 VGND.n39 9.3005
R226 VGND.n41 VGND.n2 9.3005
R227 VGND.n14 VGND.n13 7.51197
R228 VGND.n50 VGND.n49 7.12063
R229 VGND.n36 VGND.n35 5.64756
R230 VGND.n35 VGND.n34 4.14168
R231 VGND.n15 VGND.n14 0.614509
R232 VGND.n50 VGND.n0 0.148519
R233 VGND.n15 VGND.n12 0.120292
R234 VGND.n19 VGND.n12 0.120292
R235 VGND.n20 VGND.n19 0.120292
R236 VGND.n20 VGND.n9 0.120292
R237 VGND.n24 VGND.n9 0.120292
R238 VGND.n25 VGND.n24 0.120292
R239 VGND.n26 VGND.n25 0.120292
R240 VGND.n26 VGND.n6 0.120292
R241 VGND.n30 VGND.n6 0.120292
R242 VGND.n31 VGND.n30 0.120292
R243 VGND.n32 VGND.n31 0.120292
R244 VGND.n32 VGND.n4 0.120292
R245 VGND.n37 VGND.n4 0.120292
R246 VGND.n38 VGND.n37 0.120292
R247 VGND.n39 VGND.n38 0.120292
R248 VGND.n39 VGND.n2 0.120292
R249 VGND.n43 VGND.n2 0.120292
R250 VGND.n44 VGND.n43 0.120292
R251 VGND.n45 VGND.n44 0.120292
R252 VGND.n45 VGND.n0 0.120292
R253 VGND VGND.n50 0.101821
R254 VNB.t8 VNB.t3 2933.33
R255 VNB.t17 VNB.t14 2748.22
R256 VNB.t4 VNB.t8 2747.16
R257 VNB.t9 VNB.t5 2677.02
R258 VNB.t5 VNB.t6 2512.82
R259 VNB.t16 VNB.t11 2121.68
R260 VNB.t13 VNB.t1 1879.61
R261 VNB.t0 VNB.t2 1863.06
R262 VNB.t12 VNB.t7 1552.1
R263 VNB.t2 VNB.t4 1453.45
R264 VNB.t7 VNB.t16 1366.99
R265 VNB.t1 VNB.t12 1352.75
R266 VNB.t14 VNB.t15 1196.12
R267 VNB.t10 VNB.t9 1196.12
R268 VNB.t11 VNB.t17 1124.92
R269 VNB.t3 VNB.t13 1025.24
R270 VNB.t6 VNB.t0 951.351
R271 VNB VNB.t10 726.215
R272 a_1758_413.t0 a_1758_413.t1 121.953
R273 a_1946_47.t0 a_1946_47.t1 70.0005
R274 SCD.n0 SCD.t0 248.767
R275 SCD.n0 SCD.t1 191.998
R276 SCD SCD.n0 155.072
R277 a_817_66.t0 a_817_66.t1 60.0005
R278 SCE.t2 SCE.t3 729.321
R279 SCE.n0 SCE.t0 273.134
R280 SCE.n1 SCE.t2 215.901
R281 SCE SCE.n1 159.054
R282 SCE.n1 SCE.n0 145.296
R283 SCE.n0 SCE.t1 138.173
R284 a_538_389.t0 a_538_389.t1 94.8524
R285 RESET_B.n1 RESET_B.t0 2026.37
R286 RESET_B.n0 RESET_B.t2 398.99
R287 RESET_B.n1 RESET_B.t3 204.458
R288 RESET_B.n3 RESET_B.n0 163.06
R289 RESET_B.n2 RESET_B.n1 157.826
R290 RESET_B.n0 RESET_B.t1 136.21
R291 RESET_B.n4 RESET_B 11.2557
R292 RESET_B.n3 RESET_B.n2 9.43939
R293 RESET_B.n4 RESET_B.n3 9.30982
R294 RESET_B.n2 RESET_B 5.91708
R295 RESET_B RESET_B.n4 3.75222
R296 D.n0 D.t0 234.942
R297 D.n0 D.t1 164.25
R298 D D.n0 157.819
R299 a_569_119.t0 a_569_119.t1 60.0005
R300 Q Q.n0 586.723
R301 Q.n4 Q.n0 585
R302 Q.n2 Q.n1 185
R303 Q.n3 Q 89.6005
R304 Q.n3 Q.n2 64.8093
R305 Q.n0 Q.t1 26.5955
R306 Q.n0 Q.t0 26.5955
R307 Q.n1 Q.t3 24.9236
R308 Q.n1 Q.t2 24.9236
R309 Q Q.n3 16.0005
R310 Q Q.n4 15.0159
R311 Q.n2 Q 10.0928
R312 Q.n4 Q 1.72358
R313 Q.n3 Q 0.738962
R314 a_1187_47.n0 a_1187_47.t0 9.47418
R315 a_1293_47.t0 a_1293_47.t1 60.0005
R316 CLK.n0 CLK.t0 428.579
R317 CLK.n0 CLK.t1 426.168
R318 CLK.n1 CLK.n0 152
R319 CLK.n1 CLK 10.4234
R320 CLK CLK.n1 2.01193
C0 RESET_B a_1079_413# 0.146062f
C1 a_1079_413# SCD 2.16e-19
C2 Q VGND 0.08411f
C3 Q VPWR 0.170606f
C4 RESET_B VGND 0.271407f
C5 RESET_B VPWR 0.07406f
C6 VGND SCD 0.069738f
C7 Q D 1.13e-21
C8 SCD VPWR 0.01224f
C9 RESET_B D 8.56e-20
C10 VGND SCE 0.086893f
C11 SCE VPWR 0.066374f
C12 D SCD 0.005659f
C13 SCE D 0.051599f
C14 VPB CLK 0.040886f
C15 VPB a_1191_413# 0.011156f
C16 Q RESET_B 0.001328f
C17 Q SCD 3.09e-21
C18 RESET_B SCD 4.26e-19
C19 RESET_B SCE 1.82e-19
C20 SCE SCD 0.033759f
C21 CLK VGND 0.017295f
C22 CLK VPWR 0.01885f
C23 a_1079_413# a_1191_413# 0.04854f
C24 VPB a_1079_413# 0.09595f
C25 a_1191_413# VPWR 0.110782f
C26 CLK RESET_B 2.16e-20
C27 VPB VGND 0.011009f
C28 VPB VPWR 0.266658f
C29 CLK SCE 2.38e-19
C30 VPB D 0.068911f
C31 RESET_B a_1191_413# 0.011249f
C32 VGND a_1079_413# 0.126685f
C33 a_1079_413# VPWR 0.068775f
C34 a_1079_413# D 2.79e-20
C35 Q VPB 0.005349f
C36 VPB RESET_B 0.152772f
C37 VGND VPWR 0.066677f
C38 VPB SCD 0.06936f
C39 VPB SCE 0.182158f
C40 VGND D 0.001786f
C41 D VPWR 0.062452f
C42 Q VNB 0.03888f
C43 VGND VNB 1.32382f
C44 RESET_B VNB 0.272421f
C45 VPWR VNB 1.08933f
C46 SCD VNB 0.13368f
C47 D VNB 0.093585f
C48 SCE VNB 0.51427f
C49 CLK VNB 0.15698f
C50 VPB VNB 2.34162f
C51 a_1191_413# VNB 0.00653f
C52 a_1079_413# VNB 0.150381f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtp_1 VPB VNB VPWR VGND SCE SCD D RESET_B CLK Q
X0 a_193_47.t1 a_27_47.t2 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_780_389.t1 a_299_66.t2 a_620_389.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.82 as=0.1755 ps=1.19 w=0.54 l=0.15
X2 a_1245_303.t2 a_1079_413# VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.2184 ps=2.2 w=0.84 l=0.15
X3 VPWR.t4 a_1592_47.t4 a_1767_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VGND.t4 a_1767_21.t3 a_1701_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06705 ps=0.75 w=0.42 l=0.15
X5 a_1758_413.t1 a_193_47.t2 a_1592_47.t3 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0546 pd=0.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1767_21.t0 a_1592_47.t5 a_1946_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.05145 ps=0.665 w=0.42 l=0.15
X7 VGND.t1 SCD.t0 a_817_66.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.18
X8 a_538_389.t0 SCE.t0 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0702 pd=0.8 as=0.0729 ps=0.81 w=0.54 l=0.15
X9 VPWR.t6 SCD.t1 a_780_389.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.64 as=0.0756 ps=0.82 w=0.54 l=0.15
X10 VPWR.t8 SCE.t1 a_299_66.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.189 ps=1.78 w=0.54 l=0.15
X11 a_1767_21.t2 RESET_B.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X12 a_193_47.t0 a_27_47.t3 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_620_389.t1 D.t0 a_569_119.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.110275 pd=1.065 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 a_1293_47.t0 a_1245_303.t4 a_1187_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0759 ps=0.8 w=0.42 l=0.15
X15 a_620_389.t4 D.t1 a_538_389.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1755 pd=1.19 as=0.0702 ps=0.8 w=0.54 l=0.15
X16 a_569_119.t1 a_299_66.t3 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VPWR.t1 a_1767_21.t4 a_1758_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0546 ps=0.68 w=0.42 l=0.15
X18 VGND.t2 RESET_B.t1 a_1293_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 Q.t1 a_1767_21.t5 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X20 Q.t0 a_1767_21.t6 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_1191_413# RESET_B.t2 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1007 ps=0.94 w=0.42 l=0.15
X22 a_1079_413# a_27_47.t4 a_620_389.t2 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.063 pd=0.71 as=0.0936 ps=1.24 w=0.36 l=0.15
X23 a_1946_47.t1 RESET_B.t3 VGND.t9 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.05145 pd=0.665 as=0.12495 ps=1.015 w=0.42 l=0.15
X24 a_1701_47.t1 a_27_47.t5 a_1592_47.t1 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X25 a_1592_47.t2 a_193_47.t3 a_1245_303.t3 VNB.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X26 VGND.t0 SCE.t2 a_299_66.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_1592_47.t0 a_27_47.t6 a_1245_303.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12075 ps=1.165 w=0.42 l=0.15
X28 a_1245_303.t1 a_1079_413# VGND.t6 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1346 ps=1.15 w=0.64 l=0.15
X29 a_1079_413# a_193_47.t4 a_620_389.t5 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0861 pd=0.83 as=0.1533 ps=1.57 w=0.42 l=0.15
X30 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X31 a_817_66.t1 SCE.t3 a_620_389.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.110275 ps=1.065 w=0.42 l=0.5
X32 VGND.t8 CLK.t1 a_27_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n4 a_27_47.n3 532.726
R1 a_27_47.n2 a_27_47.t6 496.003
R2 a_27_47.t0 a_27_47.n0 391.175
R3 a_27_47.n4 a_27_47.t4 279.101
R4 a_27_47.n0 a_27_47.t1 271.212
R5 a_27_47.n1 a_27_47.t2 241.536
R6 a_27_47.n2 a_27_47.t5 199.762
R7 a_27_47.n5 a_27_47.n2 170.347
R8 a_27_47.n1 a_27_47.t3 169.237
R9 a_27_47.n5 a_27_47.n4 164.312
R10 a_27_47.n0 a_27_47.n1 152
R11 a_27_47.n0 a_27_47.n5 14.0789
R12 VPWR.n8 VPWR.t10 806.511
R13 VPWR.n33 VPWR.t6 700.982
R14 VPWR.n26 VPWR.t3 688.191
R15 VPWR.n13 VPWR.t4 663.062
R16 VPWR.n40 VPWR.n39 615.871
R17 VPWR.n47 VPWR.n1 604.394
R18 VPWR.n11 VPWR.n10 603.433
R19 VPWR.n12 VPWR.t2 254.494
R20 VPWR.n10 VPWR.t1 114.918
R21 VPWR.n10 VPWR.t5 63.3219
R22 VPWR.n39 VPWR.t9 49.2505
R23 VPWR.n39 VPWR.t8 49.2505
R24 VPWR.n37 VPWR.n4 34.6358
R25 VPWR.n38 VPWR.n37 34.6358
R26 VPWR.n41 VPWR.n38 34.6358
R27 VPWR.n45 VPWR.n2 34.6358
R28 VPWR.n46 VPWR.n45 34.6358
R29 VPWR.n27 VPWR.n6 34.6358
R30 VPWR.n31 VPWR.n6 34.6358
R31 VPWR.n32 VPWR.n31 34.6358
R32 VPWR.n19 VPWR.n18 34.6358
R33 VPWR.n20 VPWR.n19 34.6358
R34 VPWR.n25 VPWR.n24 31.3563
R35 VPWR.n1 VPWR.t0 29.5505
R36 VPWR.n33 VPWR.n4 29.3652
R37 VPWR.n18 VPWR.n11 29.3652
R38 VPWR.n1 VPWR.t7 26.5955
R39 VPWR.n40 VPWR.n2 25.224
R40 VPWR.n20 VPWR.n8 22.9652
R41 VPWR.n47 VPWR.n46 21.8358
R42 VPWR.n14 VPWR.n11 21.0829
R43 VPWR.n27 VPWR.n26 19.7527
R44 VPWR.n24 VPWR.n8 18.4476
R45 VPWR.n14 VPWR.n13 17.3181
R46 VPWR.n33 VPWR.n32 15.0593
R47 VPWR.n41 VPWR.n40 9.41227
R48 VPWR.n15 VPWR.n14 9.3005
R49 VPWR.n16 VPWR.n11 9.3005
R50 VPWR.n18 VPWR.n17 9.3005
R51 VPWR.n19 VPWR.n9 9.3005
R52 VPWR.n21 VPWR.n20 9.3005
R53 VPWR.n22 VPWR.n8 9.3005
R54 VPWR.n24 VPWR.n23 9.3005
R55 VPWR.n25 VPWR.n7 9.3005
R56 VPWR.n28 VPWR.n27 9.3005
R57 VPWR.n29 VPWR.n6 9.3005
R58 VPWR.n31 VPWR.n30 9.3005
R59 VPWR.n32 VPWR.n5 9.3005
R60 VPWR.n34 VPWR.n33 9.3005
R61 VPWR.n35 VPWR.n4 9.3005
R62 VPWR.n37 VPWR.n36 9.3005
R63 VPWR.n38 VPWR.n3 9.3005
R64 VPWR.n42 VPWR.n41 9.3005
R65 VPWR.n43 VPWR.n2 9.3005
R66 VPWR.n45 VPWR.n44 9.3005
R67 VPWR.n46 VPWR.n0 9.3005
R68 VPWR.n48 VPWR.n47 7.18025
R69 VPWR.n13 VPWR.n12 5.11699
R70 VPWR.n26 VPWR.n25 2.70272
R71 VPWR.n15 VPWR.n12 1.96442
R72 VPWR.n48 VPWR.n0 0.147761
R73 VPWR.n16 VPWR.n15 0.120292
R74 VPWR.n17 VPWR.n16 0.120292
R75 VPWR.n17 VPWR.n9 0.120292
R76 VPWR.n21 VPWR.n9 0.120292
R77 VPWR.n22 VPWR.n21 0.120292
R78 VPWR.n23 VPWR.n22 0.120292
R79 VPWR.n23 VPWR.n7 0.120292
R80 VPWR.n28 VPWR.n7 0.120292
R81 VPWR.n29 VPWR.n28 0.120292
R82 VPWR.n30 VPWR.n29 0.120292
R83 VPWR.n30 VPWR.n5 0.120292
R84 VPWR.n34 VPWR.n5 0.120292
R85 VPWR.n35 VPWR.n34 0.120292
R86 VPWR.n36 VPWR.n35 0.120292
R87 VPWR.n36 VPWR.n3 0.120292
R88 VPWR.n42 VPWR.n3 0.120292
R89 VPWR.n43 VPWR.n42 0.120292
R90 VPWR.n44 VPWR.n43 0.120292
R91 VPWR.n44 VPWR.n0 0.120292
R92 VPWR VPWR.n48 0.113006
R93 a_193_47.n0 a_193_47.t3 342.533
R94 a_193_47.n2 a_193_47.n1 338.877
R95 a_193_47.t1 a_193_47.n4 332.233
R96 a_193_47.n0 a_193_47.t2 307.817
R97 a_193_47.n4 a_193_47.t0 302.798
R98 a_193_47.n2 a_193_47.t4 300.252
R99 a_193_47.n3 a_193_47.n2 15.9565
R100 a_193_47.n4 a_193_47.n3 13.0278
R101 a_193_47.n3 a_193_47.n0 11.9849
R102 VPB.t14 VPB.t4 917.446
R103 VPB.t9 VPB.t10 774.313
R104 VPB.t7 VPB.t14 637.548
R105 VPB.t5 VPB.t3 556.386
R106 VPB.t4 VPB.t12 556.386
R107 VPB.t13 VPB.t0 511.784
R108 VPB.t2 VPB.t6 313.707
R109 VPB.t12 VPB.t8 281.154
R110 VPB.t0 VPB.t7 275.084
R111 VPB.t10 VPB.t11 268.688
R112 VPB.t11 VPB.t13 262.291
R113 VPB.t1 VPB.t9 257.478
R114 VPB.t8 VPB.t15 254.518
R115 VPB.t6 VPB.t5 248.599
R116 VPB.t15 VPB.t2 242.679
R117 VPB VPB.t1 177.571
R118 a_299_66.n0 a_299_66.t2 1108.99
R119 a_299_66.t1 a_299_66.n0 700.674
R120 a_299_66.n0 a_299_66.t3 346.219
R121 a_299_66.n0 a_299_66.t0 288.474
R122 a_620_389.n0 a_620_389.t5 686.09
R123 a_620_389.n3 a_620_389.n2 599.683
R124 a_620_389.n0 a_620_389.t2 360.05
R125 a_620_389.n2 a_620_389.n1 276.555
R126 a_620_389.n3 a_620_389.t4 162.344
R127 a_620_389.n1 a_620_389.t0 106.636
R128 a_620_389.n2 a_620_389.n0 83.2005
R129 a_620_389.t3 a_620_389.n3 74.7875
R130 a_620_389.n1 a_620_389.t1 38.5724
R131 a_780_389.t0 a_780_389.t1 102.148
R132 a_1245_303.n4 a_1245_303.n3 644.628
R133 a_1245_303.n1 a_1245_303.t4 365.918
R134 a_1245_303.n3 a_1245_303.n2 269.793
R135 a_1245_303.n3 a_1245_303.n1 227.672
R136 a_1245_303.n1 a_1245_303.n0 158.392
R137 a_1245_303.n4 a_1245_303.t0 72.7029
R138 a_1245_303.n2 a_1245_303.t3 63.3338
R139 a_1245_303.t2 a_1245_303.n4 50.4231
R140 a_1245_303.n2 a_1245_303.t1 26.7713
R141 a_1592_47.n1 a_1592_47.t5 1025.84
R142 a_1592_47.n3 a_1592_47.n2 635.218
R143 a_1592_47.n1 a_1592_47.t4 412.283
R144 a_1592_47.n2 a_1592_47.n0 302.889
R145 a_1592_47.n2 a_1592_47.n1 220.894
R146 a_1592_47.n0 a_1592_47.t2 70.0005
R147 a_1592_47.t0 a_1592_47.n3 68.0124
R148 a_1592_47.n3 a_1592_47.t3 63.3219
R149 a_1592_47.n0 a_1592_47.t1 61.6672
R150 a_1767_21.n3 a_1767_21.t4 1015.03
R151 a_1767_21.n2 a_1767_21.n0 783.903
R152 a_1767_21.n4 a_1767_21.n3 257.036
R153 a_1767_21.n1 a_1767_21.t5 239.505
R154 a_1767_21.t0 a_1767_21.n4 223.571
R155 a_1767_21.n3 a_1767_21.t3 178.585
R156 a_1767_21.n1 a_1767_21.t6 167.204
R157 a_1767_21.n2 a_1767_21.n1 162.24
R158 a_1767_21.n4 a_1767_21.n2 64.0131
R159 a_1767_21.n0 a_1767_21.t1 63.3219
R160 a_1767_21.n0 a_1767_21.t2 63.3219
R161 a_1701_47.t0 a_1701_47.t1 93.5174
R162 VGND.n12 VGND.t3 297.289
R163 VGND.n35 VGND.t7 252.274
R164 VGND.n1 VGND.t0 241.996
R165 VGND.n28 VGND.t1 241.22
R166 VGND.n11 VGND.n10 205.707
R167 VGND.n20 VGND.n8 199.739
R168 VGND.n42 VGND.n41 199.739
R169 VGND.n10 VGND.t9 117.144
R170 VGND.n8 VGND.t2 72.8576
R171 VGND.n8 VGND.t6 60.5809
R172 VGND.n10 VGND.t4 52.8576
R173 VGND.n15 VGND.n14 34.6358
R174 VGND.n16 VGND.n15 34.6358
R175 VGND.n16 VGND.n7 34.6358
R176 VGND.n22 VGND.n21 34.6358
R177 VGND.n22 VGND.n5 34.6358
R178 VGND.n26 VGND.n5 34.6358
R179 VGND.n27 VGND.n26 34.6358
R180 VGND.n29 VGND.n3 34.6358
R181 VGND.n33 VGND.n3 34.6358
R182 VGND.n34 VGND.n33 34.6358
R183 VGND.n40 VGND.n39 34.6358
R184 VGND.n12 VGND.n11 27.1309
R185 VGND.n20 VGND.n7 25.977
R186 VGND.n41 VGND.t5 24.9236
R187 VGND.n41 VGND.t8 24.9236
R188 VGND.n42 VGND.n40 22.9652
R189 VGND.n35 VGND.n34 19.9534
R190 VGND.n39 VGND.n1 19.9534
R191 VGND.n21 VGND.n20 18.4476
R192 VGND.n14 VGND.n11 15.0593
R193 VGND.n35 VGND.n1 14.3064
R194 VGND.n40 VGND.n0 9.3005
R195 VGND.n39 VGND.n38 9.3005
R196 VGND.n37 VGND.n1 9.3005
R197 VGND.n36 VGND.n35 9.3005
R198 VGND.n14 VGND.n13 9.3005
R199 VGND.n15 VGND.n9 9.3005
R200 VGND.n17 VGND.n16 9.3005
R201 VGND.n18 VGND.n7 9.3005
R202 VGND.n20 VGND.n19 9.3005
R203 VGND.n21 VGND.n6 9.3005
R204 VGND.n23 VGND.n22 9.3005
R205 VGND.n24 VGND.n5 9.3005
R206 VGND.n26 VGND.n25 9.3005
R207 VGND.n27 VGND.n4 9.3005
R208 VGND.n30 VGND.n29 9.3005
R209 VGND.n31 VGND.n3 9.3005
R210 VGND.n33 VGND.n32 9.3005
R211 VGND.n34 VGND.n2 9.3005
R212 VGND.n43 VGND.n42 7.12063
R213 VGND.n29 VGND.n28 5.64756
R214 VGND.n28 VGND.n27 4.14168
R215 VGND.n13 VGND.n12 0.193917
R216 VGND.n43 VGND.n0 0.148519
R217 VGND.n13 VGND.n9 0.120292
R218 VGND.n17 VGND.n9 0.120292
R219 VGND.n18 VGND.n17 0.120292
R220 VGND.n19 VGND.n18 0.120292
R221 VGND.n19 VGND.n6 0.120292
R222 VGND.n23 VGND.n6 0.120292
R223 VGND.n24 VGND.n23 0.120292
R224 VGND.n25 VGND.n24 0.120292
R225 VGND.n25 VGND.n4 0.120292
R226 VGND.n30 VGND.n4 0.120292
R227 VGND.n31 VGND.n30 0.120292
R228 VGND.n32 VGND.n31 0.120292
R229 VGND.n32 VGND.n2 0.120292
R230 VGND.n36 VGND.n2 0.120292
R231 VGND.n37 VGND.n36 0.120292
R232 VGND.n38 VGND.n37 0.120292
R233 VGND.n38 VGND.n0 0.120292
R234 VGND VGND.n43 0.101821
R235 VNB.t10 VNB.t2 2933.33
R236 VNB.t1 VNB.t5 2748.22
R237 VNB.t3 VNB.t10 2747.16
R238 VNB.t11 VNB.t0 2677.02
R239 VNB.t0 VNB.t13 2512.82
R240 VNB.t6 VNB.t16 2121.68
R241 VNB.t4 VNB.t12 1879.61
R242 VNB.t8 VNB.t7 1863.06
R243 VNB.t15 VNB.t9 1552.1
R244 VNB.t7 VNB.t3 1453.45
R245 VNB.t9 VNB.t6 1366.99
R246 VNB.t12 VNB.t15 1352.75
R247 VNB.t14 VNB.t11 1196.12
R248 VNB.t16 VNB.t1 1124.92
R249 VNB.t2 VNB.t4 1025.24
R250 VNB.t13 VNB.t8 951.351
R251 VNB VNB.t14 726.215
R252 a_1758_413.t0 a_1758_413.t1 121.953
R253 a_1946_47.t0 a_1946_47.t1 70.0005
R254 SCD.n0 SCD.t0 248.767
R255 SCD.n0 SCD.t1 191.998
R256 SCD SCD.n0 155.072
R257 a_817_66.t0 a_817_66.t1 60.0005
R258 SCE.t2 SCE.t3 729.321
R259 SCE.n0 SCE.t0 273.134
R260 SCE.n1 SCE.t2 215.901
R261 SCE SCE.n1 159.054
R262 SCE.n1 SCE.n0 145.296
R263 SCE.n0 SCE.t1 138.173
R264 a_538_389.t0 a_538_389.t1 94.8524
R265 RESET_B.n1 RESET_B.t0 2026.37
R266 RESET_B.n0 RESET_B.t2 398.99
R267 RESET_B.n1 RESET_B.t3 204.458
R268 RESET_B.n3 RESET_B.n0 163.06
R269 RESET_B.n2 RESET_B.n1 157.826
R270 RESET_B.n0 RESET_B.t1 136.21
R271 RESET_B.n4 RESET_B 11.2557
R272 RESET_B.n3 RESET_B.n2 9.43939
R273 RESET_B.n4 RESET_B.n3 9.30982
R274 RESET_B.n2 RESET_B 5.91708
R275 RESET_B RESET_B.n4 3.75222
R276 D.n0 D.t0 234.942
R277 D.n0 D.t1 164.25
R278 D D.n0 157.819
R279 a_569_119.t0 a_569_119.t1 60.0005
R280 a_1187_47.n0 a_1187_47.t0 9.47418
R281 a_1293_47.t0 a_1293_47.t1 60.0005
R282 Q.n2 Q.t1 353.606
R283 Q.n0 Q.t0 209.923
R284 Q.n1 Q 89.6005
R285 Q.n1 Q.n0 64.8093
R286 Q Q.n1 16.0005
R287 Q.n0 Q 10.0928
R288 Q.n2 Q 9.10538
R289 Q Q.n2 7.47898
R290 Q.n1 Q 0.738962
R291 CLK.n0 CLK.t0 428.579
R292 CLK.n0 CLK.t1 426.168
R293 CLK.n1 CLK.n0 152
R294 CLK.n1 CLK 10.4234
R295 CLK CLK.n1 2.01193
C0 Q RESET_B 0.001328f
C1 SCD Q 3.09e-21
C2 Q VPB 0.011159f
C3 RESET_B SCE 1.82e-19
C4 SCD RESET_B 4.26e-19
C5 SCD SCE 0.033759f
C6 RESET_B VPB 0.152772f
C7 SCE VPB 0.182158f
C8 SCD VPB 0.06936f
C9 RESET_B a_1079_413# 0.146062f
C10 SCD a_1079_413# 2.16e-19
C11 VPB a_1079_413# 0.09595f
C12 VGND D 0.001786f
C13 VPWR VGND 0.046151f
C14 VGND CLK 0.017295f
C15 VPWR D 0.062452f
C16 VPWR CLK 0.01885f
C17 VPWR a_1191_413# 0.110782f
C18 Q VGND 0.057668f
C19 Q D 1.13e-21
C20 VPWR Q 0.100202f
C21 RESET_B VGND 0.271028f
C22 RESET_B D 8.56e-20
C23 VGND SCE 0.086893f
C24 SCD VGND 0.069735f
C25 VPWR RESET_B 0.07406f
C26 SCE D 0.051599f
C27 VGND VPB 0.00922f
C28 RESET_B CLK 2.16e-20
C29 SCD VPWR 0.01224f
C30 SCD D 0.005659f
C31 VPWR SCE 0.066374f
C32 SCE CLK 2.38e-19
C33 VPWR VPB 0.249451f
C34 D VPB 0.068911f
C35 VPB CLK 0.040886f
C36 RESET_B a_1191_413# 0.011249f
C37 VGND a_1079_413# 0.126685f
C38 D a_1079_413# 2.79e-20
C39 VPWR a_1079_413# 0.068775f
C40 VPB a_1191_413# 0.011156f
C41 a_1079_413# a_1191_413# 0.04854f
C42 Q VNB 0.089262f
C43 VGND VNB 1.2607f
C44 RESET_B VNB 0.273601f
C45 VPWR VNB 1.01734f
C46 SCD VNB 0.13368f
C47 D VNB 0.093585f
C48 SCE VNB 0.51427f
C49 CLK VNB 0.15698f
C50 VPB VNB 2.25302f
C51 a_1191_413# VNB 0.00653f
C52 a_1079_413# VNB 0.150381f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtn_1 VPB VNB VPWR VGND SCE SCD D RESET_B CLK_N Q
X0 a_193_47.t1 a_27_47.t2 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_780_389.t0 a_299_66.t2 a_620_389.t2 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.82 as=0.1755 ps=1.19 w=0.54 l=0.15
X2 a_1245_303.t1 a_1079_413# VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.2184 ps=2.2 w=0.84 l=0.15
X3 VPWR.t3 a_1592_47.t4 a_1767_21.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VGND.t8 a_1767_21.t3 a_1701_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06705 ps=0.75 w=0.42 l=0.15
X5 a_1758_413.t0 a_27_47.t3 a_1592_47.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0546 pd=0.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1767_21.t1 a_1592_47.t5 a_1946_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.05145 ps=0.665 w=0.42 l=0.15
X7 VGND.t9 SCD.t0 a_817_66.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.18
X8 a_538_389.t1 SCE.t0 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0702 pd=0.8 as=0.0729 ps=0.81 w=0.54 l=0.15
X9 VPWR.t9 SCD.t1 a_780_389.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.64 as=0.0756 ps=0.82 w=0.54 l=0.15
X10 VPWR.t0 SCE.t1 a_299_66.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.189 ps=1.78 w=0.54 l=0.15
X11 a_1767_21.t2 RESET_B.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X12 a_193_47.t0 a_27_47.t4 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_620_389.t1 D.t0 a_569_119.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.110275 pd=1.065 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 a_1293_47.t1 a_1245_303.t4 a_1187_47.t0 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0759 ps=0.8 w=0.42 l=0.15
X15 a_620_389.t0 D.t1 a_538_389.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1755 pd=1.19 as=0.0702 ps=0.8 w=0.54 l=0.15
X16 a_569_119.t1 a_299_66.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VPWR.t5 a_1767_21.t4 a_1758_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0546 ps=0.68 w=0.42 l=0.15
X18 VGND.t4 RESET_B.t1 a_1293_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 Q.t0 a_1767_21.t5 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X20 Q.t1 a_1767_21.t6 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_1191_413.t0 RESET_B.t2 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1007 ps=0.94 w=0.42 l=0.15
X22 a_1079_413# a_193_47.t2 a_620_389.t4 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.063 pd=0.71 as=0.0936 ps=1.24 w=0.36 l=0.15
X23 a_1946_47.t1 RESET_B.t3 VGND.t6 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.05145 pd=0.665 as=0.12495 ps=1.015 w=0.42 l=0.15
X24 a_1701_47.t0 a_193_47.t3 a_1592_47.t0 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X25 a_1592_47.t3 a_27_47.t5 a_1245_303.t3 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X26 VGND.t2 SCE.t2 a_299_66.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_1592_47.t1 a_193_47.t4 a_1245_303.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12075 ps=1.165 w=0.42 l=0.15
X28 a_1245_303.t0 a_1079_413# VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1346 ps=1.15 w=0.64 l=0.15
X29 a_1079_413# a_27_47.t6 a_620_389.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0861 pd=0.83 as=0.1533 ps=1.57 w=0.42 l=0.15
X30 VPWR.t2 CLK_N.t0 a_27_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X31 a_817_66.t0 SCE.t3 a_620_389.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.110275 ps=1.065 w=0.42 l=0.5
X32 VGND.t0 CLK_N.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t1 a_27_47.n6 351.659
R1 a_27_47.n2 a_27_47.t5 342.533
R2 a_27_47.n4 a_27_47.n3 338.877
R3 a_27_47.n2 a_27_47.t3 307.817
R4 a_27_47.n4 a_27_47.t6 300.252
R5 a_27_47.n1 a_27_47.t0 271.212
R6 a_27_47.n0 a_27_47.t2 241.536
R7 a_27_47.n0 a_27_47.t4 169.237
R8 a_27_47.n1 a_27_47.n0 152
R9 a_27_47.n6 a_27_47.n1 40.7345
R10 a_27_47.n5 a_27_47.n4 15.9565
R11 a_27_47.n6 a_27_47.n5 13.3475
R12 a_27_47.n5 a_27_47.n2 11.9849
R13 VPWR.n8 VPWR.t1 806.511
R14 VPWR.n33 VPWR.t9 700.982
R15 VPWR.n26 VPWR.t8 688.191
R16 VPWR.n13 VPWR.t3 663.062
R17 VPWR.n40 VPWR.n39 615.871
R18 VPWR.n47 VPWR.n1 604.394
R19 VPWR.n11 VPWR.n10 603.433
R20 VPWR.n12 VPWR.t6 254.494
R21 VPWR.n10 VPWR.t5 114.918
R22 VPWR.n10 VPWR.t4 63.3219
R23 VPWR.n39 VPWR.t10 49.2505
R24 VPWR.n39 VPWR.t0 49.2505
R25 VPWR.n37 VPWR.n4 34.6358
R26 VPWR.n38 VPWR.n37 34.6358
R27 VPWR.n41 VPWR.n38 34.6358
R28 VPWR.n45 VPWR.n2 34.6358
R29 VPWR.n46 VPWR.n45 34.6358
R30 VPWR.n27 VPWR.n6 34.6358
R31 VPWR.n31 VPWR.n6 34.6358
R32 VPWR.n32 VPWR.n31 34.6358
R33 VPWR.n19 VPWR.n18 34.6358
R34 VPWR.n20 VPWR.n19 34.6358
R35 VPWR.n25 VPWR.n24 31.3563
R36 VPWR.n1 VPWR.t2 29.5505
R37 VPWR.n33 VPWR.n4 29.3652
R38 VPWR.n18 VPWR.n11 29.3652
R39 VPWR.n1 VPWR.t7 26.5955
R40 VPWR.n40 VPWR.n2 25.224
R41 VPWR.n20 VPWR.n8 22.9652
R42 VPWR.n47 VPWR.n46 21.8358
R43 VPWR.n14 VPWR.n11 21.0829
R44 VPWR.n27 VPWR.n26 19.7527
R45 VPWR.n24 VPWR.n8 18.4476
R46 VPWR.n14 VPWR.n13 17.3181
R47 VPWR.n33 VPWR.n32 15.0593
R48 VPWR.n41 VPWR.n40 9.41227
R49 VPWR.n15 VPWR.n14 9.3005
R50 VPWR.n16 VPWR.n11 9.3005
R51 VPWR.n18 VPWR.n17 9.3005
R52 VPWR.n19 VPWR.n9 9.3005
R53 VPWR.n21 VPWR.n20 9.3005
R54 VPWR.n22 VPWR.n8 9.3005
R55 VPWR.n24 VPWR.n23 9.3005
R56 VPWR.n25 VPWR.n7 9.3005
R57 VPWR.n28 VPWR.n27 9.3005
R58 VPWR.n29 VPWR.n6 9.3005
R59 VPWR.n31 VPWR.n30 9.3005
R60 VPWR.n32 VPWR.n5 9.3005
R61 VPWR.n34 VPWR.n33 9.3005
R62 VPWR.n35 VPWR.n4 9.3005
R63 VPWR.n37 VPWR.n36 9.3005
R64 VPWR.n38 VPWR.n3 9.3005
R65 VPWR.n42 VPWR.n41 9.3005
R66 VPWR.n43 VPWR.n2 9.3005
R67 VPWR.n45 VPWR.n44 9.3005
R68 VPWR.n46 VPWR.n0 9.3005
R69 VPWR.n48 VPWR.n47 7.18025
R70 VPWR.n13 VPWR.n12 5.11699
R71 VPWR.n26 VPWR.n25 2.70272
R72 VPWR.n15 VPWR.n12 1.96442
R73 VPWR.n48 VPWR.n0 0.147761
R74 VPWR.n16 VPWR.n15 0.120292
R75 VPWR.n17 VPWR.n16 0.120292
R76 VPWR.n17 VPWR.n9 0.120292
R77 VPWR.n21 VPWR.n9 0.120292
R78 VPWR.n22 VPWR.n21 0.120292
R79 VPWR.n23 VPWR.n22 0.120292
R80 VPWR.n23 VPWR.n7 0.120292
R81 VPWR.n28 VPWR.n7 0.120292
R82 VPWR.n29 VPWR.n28 0.120292
R83 VPWR.n30 VPWR.n29 0.120292
R84 VPWR.n30 VPWR.n5 0.120292
R85 VPWR.n34 VPWR.n5 0.120292
R86 VPWR.n35 VPWR.n34 0.120292
R87 VPWR.n36 VPWR.n35 0.120292
R88 VPWR.n36 VPWR.n3 0.120292
R89 VPWR.n42 VPWR.n3 0.120292
R90 VPWR.n43 VPWR.n42 0.120292
R91 VPWR.n44 VPWR.n43 0.120292
R92 VPWR.n44 VPWR.n0 0.120292
R93 VPWR VPWR.n48 0.113006
R94 a_193_47.n2 a_193_47.n1 532.726
R95 a_193_47.n0 a_193_47.t4 496.003
R96 a_193_47.t1 a_193_47.n4 379.293
R97 a_193_47.n2 a_193_47.t2 279.101
R98 a_193_47.n4 a_193_47.t0 255.74
R99 a_193_47.n0 a_193_47.t3 199.762
R100 a_193_47.n3 a_193_47.n0 170.347
R101 a_193_47.n3 a_193_47.n2 164.312
R102 a_193_47.n4 a_193_47.n3 12.5563
R103 VPB.t9 VPB.t12 917.446
R104 VPB.t11 VPB.t0 774.313
R105 VPB.t14 VPB.t9 637.548
R106 VPB.t4 VPB.t8 556.386
R107 VPB.t12 VPB.t2 556.386
R108 VPB.t1 VPB.t13 511.784
R109 VPB.t7 VPB.t6 313.707
R110 VPB.t2 VPB.t5 281.154
R111 VPB.t13 VPB.t14 275.084
R112 VPB.t0 VPB.t15 268.688
R113 VPB.t15 VPB.t1 262.291
R114 VPB.t3 VPB.t11 257.478
R115 VPB.t5 VPB.t10 254.518
R116 VPB.t6 VPB.t4 248.599
R117 VPB.t10 VPB.t7 242.679
R118 VPB VPB.t3 177.571
R119 a_299_66.n0 a_299_66.t2 1108.99
R120 a_299_66.t0 a_299_66.n0 700.674
R121 a_299_66.n0 a_299_66.t3 346.219
R122 a_299_66.n0 a_299_66.t1 288.474
R123 a_620_389.n0 a_620_389.t5 686.09
R124 a_620_389.n3 a_620_389.n2 599.683
R125 a_620_389.n0 a_620_389.t4 360.05
R126 a_620_389.n2 a_620_389.n1 276.555
R127 a_620_389.t0 a_620_389.n3 162.344
R128 a_620_389.n1 a_620_389.t3 106.636
R129 a_620_389.n2 a_620_389.n0 83.2005
R130 a_620_389.n3 a_620_389.t2 74.7875
R131 a_620_389.n1 a_620_389.t1 38.5724
R132 a_780_389.t0 a_780_389.t1 102.148
R133 a_1245_303.n4 a_1245_303.n3 644.628
R134 a_1245_303.n1 a_1245_303.t4 365.918
R135 a_1245_303.n3 a_1245_303.n2 269.793
R136 a_1245_303.n3 a_1245_303.n1 227.672
R137 a_1245_303.n1 a_1245_303.n0 158.392
R138 a_1245_303.n4 a_1245_303.t2 72.7029
R139 a_1245_303.n2 a_1245_303.t3 63.3338
R140 a_1245_303.t1 a_1245_303.n4 50.4231
R141 a_1245_303.n2 a_1245_303.t0 26.7713
R142 a_1592_47.n1 a_1592_47.t5 1025.84
R143 a_1592_47.n3 a_1592_47.n2 635.218
R144 a_1592_47.n1 a_1592_47.t4 412.283
R145 a_1592_47.n2 a_1592_47.n0 302.889
R146 a_1592_47.n2 a_1592_47.n1 220.894
R147 a_1592_47.n0 a_1592_47.t3 70.0005
R148 a_1592_47.t1 a_1592_47.n3 68.0124
R149 a_1592_47.n3 a_1592_47.t2 63.3219
R150 a_1592_47.n0 a_1592_47.t0 61.6672
R151 a_1767_21.n1 a_1767_21.t4 1015.03
R152 a_1767_21.n4 a_1767_21.n3 783.903
R153 a_1767_21.n2 a_1767_21.n1 257.036
R154 a_1767_21.n0 a_1767_21.t5 239.505
R155 a_1767_21.n2 a_1767_21.t1 223.571
R156 a_1767_21.n1 a_1767_21.t3 178.585
R157 a_1767_21.n0 a_1767_21.t6 167.204
R158 a_1767_21.n3 a_1767_21.n0 162.24
R159 a_1767_21.n3 a_1767_21.n2 64.0131
R160 a_1767_21.t0 a_1767_21.n4 63.3219
R161 a_1767_21.n4 a_1767_21.t2 63.3219
R162 a_1701_47.t1 a_1701_47.t0 93.5174
R163 VGND.n12 VGND.t7 297.289
R164 VGND.n35 VGND.t3 252.274
R165 VGND.n1 VGND.t2 241.996
R166 VGND.n28 VGND.t9 241.22
R167 VGND.n11 VGND.n10 205.707
R168 VGND.n20 VGND.n8 199.739
R169 VGND.n42 VGND.n41 199.739
R170 VGND.n10 VGND.t6 117.144
R171 VGND.n8 VGND.t4 72.8576
R172 VGND.n8 VGND.t1 60.5809
R173 VGND.n10 VGND.t8 52.8576
R174 VGND.n15 VGND.n14 34.6358
R175 VGND.n16 VGND.n15 34.6358
R176 VGND.n16 VGND.n7 34.6358
R177 VGND.n22 VGND.n21 34.6358
R178 VGND.n22 VGND.n5 34.6358
R179 VGND.n26 VGND.n5 34.6358
R180 VGND.n27 VGND.n26 34.6358
R181 VGND.n29 VGND.n3 34.6358
R182 VGND.n33 VGND.n3 34.6358
R183 VGND.n34 VGND.n33 34.6358
R184 VGND.n40 VGND.n39 34.6358
R185 VGND.n12 VGND.n11 27.1309
R186 VGND.n20 VGND.n7 25.977
R187 VGND.n41 VGND.t5 24.9236
R188 VGND.n41 VGND.t0 24.9236
R189 VGND.n42 VGND.n40 22.9652
R190 VGND.n35 VGND.n34 19.9534
R191 VGND.n39 VGND.n1 19.9534
R192 VGND.n21 VGND.n20 18.4476
R193 VGND.n14 VGND.n11 15.0593
R194 VGND.n35 VGND.n1 14.3064
R195 VGND.n40 VGND.n0 9.3005
R196 VGND.n39 VGND.n38 9.3005
R197 VGND.n37 VGND.n1 9.3005
R198 VGND.n36 VGND.n35 9.3005
R199 VGND.n14 VGND.n13 9.3005
R200 VGND.n15 VGND.n9 9.3005
R201 VGND.n17 VGND.n16 9.3005
R202 VGND.n18 VGND.n7 9.3005
R203 VGND.n20 VGND.n19 9.3005
R204 VGND.n21 VGND.n6 9.3005
R205 VGND.n23 VGND.n22 9.3005
R206 VGND.n24 VGND.n5 9.3005
R207 VGND.n26 VGND.n25 9.3005
R208 VGND.n27 VGND.n4 9.3005
R209 VGND.n30 VGND.n29 9.3005
R210 VGND.n31 VGND.n3 9.3005
R211 VGND.n33 VGND.n32 9.3005
R212 VGND.n34 VGND.n2 9.3005
R213 VGND.n43 VGND.n42 7.12063
R214 VGND.n29 VGND.n28 5.64756
R215 VGND.n28 VGND.n27 4.14168
R216 VGND.n13 VGND.n12 0.193917
R217 VGND.n43 VGND.n0 0.148519
R218 VGND.n13 VGND.n9 0.120292
R219 VGND.n17 VGND.n9 0.120292
R220 VGND.n18 VGND.n17 0.120292
R221 VGND.n19 VGND.n18 0.120292
R222 VGND.n19 VGND.n6 0.120292
R223 VGND.n23 VGND.n6 0.120292
R224 VGND.n24 VGND.n23 0.120292
R225 VGND.n25 VGND.n24 0.120292
R226 VGND.n25 VGND.n4 0.120292
R227 VGND.n30 VGND.n4 0.120292
R228 VGND.n31 VGND.n30 0.120292
R229 VGND.n32 VGND.n31 0.120292
R230 VGND.n32 VGND.n2 0.120292
R231 VGND.n36 VGND.n2 0.120292
R232 VGND.n37 VGND.n36 0.120292
R233 VGND.n38 VGND.n37 0.120292
R234 VGND.n38 VGND.n0 0.120292
R235 VGND VGND.n43 0.101821
R236 VNB.t9 VNB.t16 2933.33
R237 VNB.t7 VNB.t13 2748.22
R238 VNB.t15 VNB.t9 2747.16
R239 VNB.t11 VNB.t3 2677.02
R240 VNB.t3 VNB.t4 2512.82
R241 VNB.t14 VNB.t12 2121.68
R242 VNB.t6 VNB.t1 1879.61
R243 VNB.t2 VNB.t5 1863.06
R244 VNB.t10 VNB.t8 1552.1
R245 VNB.t5 VNB.t15 1453.45
R246 VNB.t8 VNB.t14 1366.99
R247 VNB.t1 VNB.t10 1352.75
R248 VNB.t0 VNB.t11 1196.12
R249 VNB.t12 VNB.t7 1124.92
R250 VNB.t16 VNB.t6 1025.24
R251 VNB.t4 VNB.t2 951.351
R252 VNB VNB.t0 726.215
R253 a_1758_413.t0 a_1758_413.t1 121.953
R254 a_1946_47.t0 a_1946_47.t1 70.0005
R255 SCD.n0 SCD.t0 248.767
R256 SCD.n0 SCD.t1 191.998
R257 SCD SCD.n0 155.072
R258 a_817_66.t1 a_817_66.t0 60.0005
R259 SCE.t2 SCE.t3 729.321
R260 SCE.n0 SCE.t0 273.134
R261 SCE.n1 SCE.t2 215.901
R262 SCE SCE.n1 159.054
R263 SCE.n1 SCE.n0 145.296
R264 SCE.n0 SCE.t1 138.173
R265 a_538_389.t0 a_538_389.t1 94.8524
R266 RESET_B.n1 RESET_B.t0 2026.37
R267 RESET_B.n0 RESET_B.t2 398.99
R268 RESET_B.n1 RESET_B.t3 204.458
R269 RESET_B.n3 RESET_B.n0 163.06
R270 RESET_B.n2 RESET_B.n1 157.826
R271 RESET_B.n0 RESET_B.t1 136.21
R272 RESET_B.n4 RESET_B 11.2557
R273 RESET_B.n3 RESET_B.n2 9.43939
R274 RESET_B.n4 RESET_B.n3 9.30982
R275 RESET_B.n2 RESET_B 5.91708
R276 RESET_B RESET_B.n4 3.75222
R277 D.n0 D.t0 234.942
R278 D.n0 D.t1 164.25
R279 D D.n0 157.819
R280 a_569_119.t0 a_569_119.t1 60.0005
R281 a_1187_47.n0 a_1187_47.t0 9.47418
R282 a_1293_47.t0 a_1293_47.t1 60.0005
R283 Q.n2 Q.t0 353.606
R284 Q.n0 Q.t1 209.923
R285 Q.n1 Q 89.6005
R286 Q.n1 Q.n0 64.8093
R287 Q Q.n1 16.0005
R288 Q.n0 Q 10.0928
R289 Q.n2 Q 9.10538
R290 Q Q.n2 7.47898
R291 Q.n1 Q 0.738962
R292 CLK_N.n0 CLK_N.t0 428.579
R293 CLK_N.n0 CLK_N.t1 426.168
R294 CLK_N.n1 CLK_N.n0 152
R295 CLK_N.n1 CLK_N 10.4234
R296 CLK_N CLK_N.n1 2.01193
C0 SCD Q 3.09e-21
C1 RESET_B Q 0.001328f
C2 D Q 1.13e-21
C3 Q VPB 0.011159f
C4 SCD SCE 0.033759f
C5 SCE RESET_B 1.82e-19
C6 SCE D 0.051599f
C7 SCE VPB 0.182158f
C8 VPWR VGND 0.043221f
C9 VPWR CLK_N 0.01885f
C10 VGND CLK_N 0.017295f
C11 SCD VPWR 0.01224f
C12 VPWR RESET_B 0.07406f
C13 VPWR D 0.062452f
C14 SCD VGND 0.069735f
C15 RESET_B VGND 0.271028f
C16 D VGND 0.001786f
C17 VPWR VPB 0.249383f
C18 RESET_B CLK_N 2.16e-20
C19 VGND VPB 0.009396f
C20 VPB CLK_N 0.040886f
C21 VPWR a_1079_413# 0.068775f
C22 VGND a_1079_413# 0.126685f
C23 VPWR Q 0.100202f
C24 VGND Q 0.057668f
C25 SCD RESET_B 4.26e-19
C26 VPWR SCE 0.066374f
C27 SCD D 0.005659f
C28 D RESET_B 8.56e-20
C29 SCD VPB 0.06936f
C30 SCE VGND 0.086893f
C31 RESET_B VPB 0.152772f
C32 SCE CLK_N 2.38e-19
C33 D VPB 0.068911f
C34 SCD a_1079_413# 2.16e-19
C35 RESET_B a_1079_413# 0.146062f
C36 D a_1079_413# 2.79e-20
C37 a_1079_413# VPB 0.09595f
C38 Q VNB 0.089262f
C39 VGND VNB 1.26076f
C40 RESET_B VNB 0.273601f
C41 VPWR VNB 1.01821f
C42 SCD VNB 0.13368f
C43 D VNB 0.093585f
C44 SCE VNB 0.51427f
C45 CLK_N VNB 0.15698f
C46 VPB VNB 2.25302f
C47 a_1079_413# VNB 0.150381f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrbp_2 VPB VNB VPWR VGND Q_N Q SCE SCD D RESET_B CLK
X0 a_193_47.t0 a_27_47.t2 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_780_389.t1 a_299_66.t2 a_620_389.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.82 as=0.1755 ps=1.19 w=0.54 l=0.15
X2 a_1245_303.t2 a_1079_413# VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.2184 ps=2.2 w=0.84 l=0.15
X3 VPWR.t10 a_1592_47.t4 a_1767_21.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VGND.t4 a_1767_21.t3 Q.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.10075 ps=0.96 w=0.65 l=0.15
X5 VGND.t1 a_1767_21.t4 a_1701_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06705 ps=0.75 w=0.42 l=0.15
X6 a_1758_413.t1 a_193_47.t2 a_1592_47.t2 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0546 pd=0.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 a_1767_21.t1 a_1592_47.t5 a_1946_47.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.05145 ps=0.665 w=0.42 l=0.15
X8 VPWR.t12 a_1767_21.t5 a_2135_47.t0 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 VGND.t8 SCD.t0 a_817_66.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.18
X10 a_538_389.t1 SCE.t0 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0702 pd=0.8 as=0.0729 ps=0.81 w=0.54 l=0.15
X11 VPWR.t2 SCD.t1 a_780_389.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.64 as=0.0756 ps=0.82 w=0.54 l=0.15
X12 VPWR.t1 SCE.t1 a_299_66.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.189 ps=1.78 w=0.54 l=0.15
X13 a_1767_21.t2 RESET_B.t0 VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X14 a_193_47.t1 a_27_47.t3 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_620_389.t5 D.t0 a_569_119.t0 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.110275 pd=1.065 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 Q.t1 a_1767_21.t6 VPWR.t13 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.149 ps=1.325 w=1 l=0.15
X17 a_1293_47.t1 a_1245_303.t4 a_1187_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0759 ps=0.8 w=0.42 l=0.15
X18 Q.t3 a_1767_21.t7 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.098625 ps=0.98 w=0.65 l=0.15
X19 a_620_389.t1 D.t1 a_538_389.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1755 pd=1.19 as=0.0702 ps=0.8 w=0.54 l=0.15
X20 Q_N.t3 a_2135_47.t2 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X21 a_569_119.t1 a_299_66.t3 VGND.t10 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X22 VPWR.t0 a_1767_21.t8 a_1758_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0546 ps=0.68 w=0.42 l=0.15
X23 VGND.t9 RESET_B.t1 a_1293_47.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 VPWR.t3 a_2135_47.t3 Q_N.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND.t2 a_1767_21.t9 a_2135_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 a_1191_413.t0 RESET_B.t2 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1007 ps=0.94 w=0.42 l=0.15
X27 a_1079_413# a_27_47.t4 a_620_389.t2 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.063 pd=0.71 as=0.0936 ps=1.24 w=0.36 l=0.15
X28 Q_N.t0 a_2135_47.t4 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X29 a_1946_47.t1 RESET_B.t3 VGND.t13 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.05145 pd=0.665 as=0.12495 ps=1.015 w=0.42 l=0.15
X30 a_1701_47.t1 a_27_47.t5 a_1592_47.t1 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X31 VPWR.t14 a_1767_21.t10 Q.t0 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.155 ps=1.31 w=1 l=0.15
X32 a_1592_47.t3 a_193_47.t3 a_1245_303.t1 VNB.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X33 VGND.t12 SCE.t2 a_299_66.t1 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X34 a_1592_47.t0 a_27_47.t6 a_1245_303.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12075 ps=1.165 w=0.42 l=0.15
X35 a_1245_303.t3 a_1079_413# VGND.t11 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1346 ps=1.15 w=0.64 l=0.15
X36 a_1079_413# a_193_47.t4 a_620_389.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0861 pd=0.83 as=0.1533 ps=1.57 w=0.42 l=0.15
X37 VGND.t6 a_2135_47.t5 Q_N.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 VPWR.t8 CLK.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X39 a_817_66.t1 SCE.t3 a_620_389.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.110275 ps=1.065 w=0.42 l=0.5
X40 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n4 a_27_47.n3 532.726
R1 a_27_47.n2 a_27_47.t6 496.003
R2 a_27_47.t1 a_27_47.n0 391.175
R3 a_27_47.n4 a_27_47.t4 279.101
R4 a_27_47.n0 a_27_47.t0 271.212
R5 a_27_47.n1 a_27_47.t2 241.536
R6 a_27_47.n2 a_27_47.t5 199.762
R7 a_27_47.n5 a_27_47.n2 170.347
R8 a_27_47.n1 a_27_47.t3 169.237
R9 a_27_47.n5 a_27_47.n4 164.312
R10 a_27_47.n0 a_27_47.n1 152
R11 a_27_47.n0 a_27_47.n5 14.0789
R12 VPWR.n8 VPWR.t9 806.511
R13 VPWR.n43 VPWR.t2 700.982
R14 VPWR.n36 VPWR.t6 688.191
R15 VPWR.n23 VPWR.t10 663.062
R16 VPWR.n50 VPWR.n49 615.871
R17 VPWR.n57 VPWR.n1 604.394
R18 VPWR.n11 VPWR.n10 603.433
R19 VPWR.n14 VPWR.n13 601.679
R20 VPWR.n17 VPWR.n16 599.74
R21 VPWR.n15 VPWR.t3 267.262
R22 VPWR.n10 VPWR.t0 114.918
R23 VPWR.n10 VPWR.t11 63.3219
R24 VPWR.n13 VPWR.t12 50.7896
R25 VPWR.n49 VPWR.t7 49.2505
R26 VPWR.n49 VPWR.t1 49.2505
R27 VPWR.n13 VPWR.t13 38.7078
R28 VPWR.n47 VPWR.n4 34.6358
R29 VPWR.n48 VPWR.n47 34.6358
R30 VPWR.n51 VPWR.n48 34.6358
R31 VPWR.n55 VPWR.n2 34.6358
R32 VPWR.n56 VPWR.n55 34.6358
R33 VPWR.n37 VPWR.n6 34.6358
R34 VPWR.n41 VPWR.n6 34.6358
R35 VPWR.n42 VPWR.n41 34.6358
R36 VPWR.n29 VPWR.n28 34.6358
R37 VPWR.n30 VPWR.n29 34.6358
R38 VPWR.n16 VPWR.t14 32.5055
R39 VPWR.n35 VPWR.n34 31.3563
R40 VPWR.n1 VPWR.t8 29.5505
R41 VPWR.n43 VPWR.n4 29.3652
R42 VPWR.n28 VPWR.n11 29.3652
R43 VPWR.n23 VPWR.n22 27.1064
R44 VPWR.n1 VPWR.t5 26.5955
R45 VPWR.n16 VPWR.t4 26.5955
R46 VPWR.n50 VPWR.n2 25.224
R47 VPWR.n18 VPWR.n14 23.3417
R48 VPWR.n30 VPWR.n8 22.9652
R49 VPWR.n18 VPWR.n17 22.2123
R50 VPWR.n57 VPWR.n56 21.8358
R51 VPWR.n24 VPWR.n11 21.0829
R52 VPWR.n22 VPWR.n14 21.0829
R53 VPWR.n37 VPWR.n36 19.7527
R54 VPWR.n34 VPWR.n8 18.4476
R55 VPWR.n24 VPWR.n23 17.3181
R56 VPWR.n43 VPWR.n42 15.0593
R57 VPWR.n51 VPWR.n50 9.41227
R58 VPWR.n19 VPWR.n18 9.3005
R59 VPWR.n20 VPWR.n14 9.3005
R60 VPWR.n22 VPWR.n21 9.3005
R61 VPWR.n23 VPWR.n12 9.3005
R62 VPWR.n25 VPWR.n24 9.3005
R63 VPWR.n26 VPWR.n11 9.3005
R64 VPWR.n28 VPWR.n27 9.3005
R65 VPWR.n29 VPWR.n9 9.3005
R66 VPWR.n31 VPWR.n30 9.3005
R67 VPWR.n32 VPWR.n8 9.3005
R68 VPWR.n34 VPWR.n33 9.3005
R69 VPWR.n35 VPWR.n7 9.3005
R70 VPWR.n38 VPWR.n37 9.3005
R71 VPWR.n39 VPWR.n6 9.3005
R72 VPWR.n41 VPWR.n40 9.3005
R73 VPWR.n42 VPWR.n5 9.3005
R74 VPWR.n44 VPWR.n43 9.3005
R75 VPWR.n45 VPWR.n4 9.3005
R76 VPWR.n47 VPWR.n46 9.3005
R77 VPWR.n48 VPWR.n3 9.3005
R78 VPWR.n52 VPWR.n51 9.3005
R79 VPWR.n53 VPWR.n2 9.3005
R80 VPWR.n55 VPWR.n54 9.3005
R81 VPWR.n56 VPWR.n0 9.3005
R82 VPWR.n58 VPWR.n57 7.18025
R83 VPWR.n17 VPWR.n15 6.58707
R84 VPWR.n36 VPWR.n35 2.70272
R85 VPWR.n19 VPWR.n15 0.61689
R86 VPWR.n58 VPWR.n0 0.147761
R87 VPWR.n20 VPWR.n19 0.120292
R88 VPWR.n21 VPWR.n20 0.120292
R89 VPWR.n21 VPWR.n12 0.120292
R90 VPWR.n25 VPWR.n12 0.120292
R91 VPWR.n26 VPWR.n25 0.120292
R92 VPWR.n27 VPWR.n26 0.120292
R93 VPWR.n27 VPWR.n9 0.120292
R94 VPWR.n31 VPWR.n9 0.120292
R95 VPWR.n32 VPWR.n31 0.120292
R96 VPWR.n33 VPWR.n32 0.120292
R97 VPWR.n33 VPWR.n7 0.120292
R98 VPWR.n38 VPWR.n7 0.120292
R99 VPWR.n39 VPWR.n38 0.120292
R100 VPWR.n40 VPWR.n39 0.120292
R101 VPWR.n40 VPWR.n5 0.120292
R102 VPWR.n44 VPWR.n5 0.120292
R103 VPWR.n45 VPWR.n44 0.120292
R104 VPWR.n46 VPWR.n45 0.120292
R105 VPWR.n46 VPWR.n3 0.120292
R106 VPWR.n52 VPWR.n3 0.120292
R107 VPWR.n53 VPWR.n52 0.120292
R108 VPWR.n54 VPWR.n53 0.120292
R109 VPWR.n54 VPWR.n0 0.120292
R110 VPWR VPWR.n58 0.113006
R111 a_193_47.n0 a_193_47.t3 342.533
R112 a_193_47.n2 a_193_47.n1 338.877
R113 a_193_47.t0 a_193_47.n4 332.233
R114 a_193_47.n0 a_193_47.t2 307.817
R115 a_193_47.n4 a_193_47.t1 302.798
R116 a_193_47.n2 a_193_47.t4 300.252
R117 a_193_47.n3 a_193_47.n2 15.9565
R118 a_193_47.n4 a_193_47.n3 13.0278
R119 a_193_47.n3 a_193_47.n0 11.9849
R120 VPB.t12 VPB.t9 917.446
R121 VPB.t8 VPB.t2 774.313
R122 VPB.t4 VPB.t12 637.548
R123 VPB.t15 VPB.t17 556.386
R124 VPB.t9 VPB.t14 556.386
R125 VPB.t3 VPB.t0 511.784
R126 VPB.t1 VPB.t16 313.707
R127 VPB.t17 VPB.t18 281.154
R128 VPB.t14 VPB.t7 281.154
R129 VPB.t0 VPB.t4 275.084
R130 VPB.t18 VPB.t19 272.274
R131 VPB.t2 VPB.t10 268.688
R132 VPB.t19 VPB.t6 266.356
R133 VPB.t10 VPB.t3 262.291
R134 VPB.t11 VPB.t8 257.478
R135 VPB.t7 VPB.t13 254.518
R136 VPB.t6 VPB.t5 248.599
R137 VPB.t16 VPB.t15 248.599
R138 VPB.t13 VPB.t1 242.679
R139 VPB VPB.t11 177.571
R140 a_299_66.n0 a_299_66.t2 1108.99
R141 a_299_66.t0 a_299_66.n0 700.674
R142 a_299_66.n0 a_299_66.t3 346.219
R143 a_299_66.n0 a_299_66.t1 288.474
R144 a_620_389.n0 a_620_389.t3 686.09
R145 a_620_389.n3 a_620_389.n2 599.683
R146 a_620_389.n0 a_620_389.t2 360.05
R147 a_620_389.n2 a_620_389.n1 276.555
R148 a_620_389.t1 a_620_389.n3 162.344
R149 a_620_389.n1 a_620_389.t0 106.636
R150 a_620_389.n2 a_620_389.n0 83.2005
R151 a_620_389.n3 a_620_389.t4 74.7875
R152 a_620_389.n1 a_620_389.t5 38.5724
R153 a_780_389.t0 a_780_389.t1 102.148
R154 a_1245_303.n4 a_1245_303.n3 644.628
R155 a_1245_303.n1 a_1245_303.t4 365.918
R156 a_1245_303.n3 a_1245_303.n2 269.793
R157 a_1245_303.n3 a_1245_303.n1 227.672
R158 a_1245_303.n1 a_1245_303.n0 158.392
R159 a_1245_303.n4 a_1245_303.t0 72.7029
R160 a_1245_303.n2 a_1245_303.t1 63.3338
R161 a_1245_303.t2 a_1245_303.n4 50.4231
R162 a_1245_303.n2 a_1245_303.t3 26.7713
R163 a_1592_47.n1 a_1592_47.t5 1025.84
R164 a_1592_47.n3 a_1592_47.n2 635.218
R165 a_1592_47.n1 a_1592_47.t4 412.283
R166 a_1592_47.n2 a_1592_47.n0 302.889
R167 a_1592_47.n2 a_1592_47.n1 220.894
R168 a_1592_47.n0 a_1592_47.t3 70.0005
R169 a_1592_47.t0 a_1592_47.n3 68.0124
R170 a_1592_47.n3 a_1592_47.t2 63.3219
R171 a_1592_47.n0 a_1592_47.t1 61.6672
R172 a_1767_21.n3 a_1767_21.t8 1015.03
R173 a_1767_21.n6 a_1767_21.n5 792.436
R174 a_1767_21.n0 a_1767_21.t5 257.067
R175 a_1767_21.n4 a_1767_21.n3 257.036
R176 a_1767_21.n4 a_1767_21.t1 223.571
R177 a_1767_21.n1 a_1767_21.t10 212.081
R178 a_1767_21.n2 a_1767_21.t6 212.081
R179 a_1767_21.n3 a_1767_21.t4 178.585
R180 a_1767_21.n5 a_1767_21.n0 178.398
R181 a_1767_21.n0 a_1767_21.t9 176.733
R182 a_1767_21.n1 a_1767_21.t3 139.78
R183 a_1767_21.n2 a_1767_21.t7 139.78
R184 a_1767_21.n5 a_1767_21.n4 72.424
R185 a_1767_21.n0 a_1767_21.n2 70.1096
R186 a_1767_21.n2 a_1767_21.n1 67.1884
R187 a_1767_21.t0 a_1767_21.n6 63.3219
R188 a_1767_21.n6 a_1767_21.t2 63.3219
R189 Q Q.n0 603.287
R190 Q Q.n1 202.554
R191 Q.n0 Q.t1 34.4755
R192 Q.n1 Q.t3 32.3082
R193 Q.n0 Q.t0 26.5955
R194 Q.n1 Q.t2 24.9236
R195 VGND.n50 VGND.t10 252.274
R196 VGND.n1 VGND.t12 241.996
R197 VGND.n43 VGND.t8 241.22
R198 VGND.n17 VGND.n15 221.142
R199 VGND.n11 VGND.n10 205.707
R200 VGND.n20 VGND.n19 202.688
R201 VGND.n35 VGND.n8 199.739
R202 VGND.n57 VGND.n56 199.739
R203 VGND.n16 VGND.t6 165.125
R204 VGND.n10 VGND.t13 117.144
R205 VGND.n8 VGND.t9 72.8576
R206 VGND.n8 VGND.t11 60.5809
R207 VGND.n10 VGND.t1 52.8576
R208 VGND.n19 VGND.t2 48.5719
R209 VGND.n18 VGND.n17 34.6358
R210 VGND.n24 VGND.n13 34.6358
R211 VGND.n25 VGND.n24 34.6358
R212 VGND.n26 VGND.n25 34.6358
R213 VGND.n30 VGND.n29 34.6358
R214 VGND.n31 VGND.n30 34.6358
R215 VGND.n31 VGND.n7 34.6358
R216 VGND.n37 VGND.n36 34.6358
R217 VGND.n37 VGND.n5 34.6358
R218 VGND.n41 VGND.n5 34.6358
R219 VGND.n42 VGND.n41 34.6358
R220 VGND.n44 VGND.n3 34.6358
R221 VGND.n48 VGND.n3 34.6358
R222 VGND.n49 VGND.n48 34.6358
R223 VGND.n55 VGND.n54 34.6358
R224 VGND.n19 VGND.t3 32.5719
R225 VGND.n15 VGND.t4 30.462
R226 VGND.n20 VGND.n18 27.4829
R227 VGND.n35 VGND.n7 25.977
R228 VGND.n15 VGND.t5 24.9236
R229 VGND.n56 VGND.t7 24.9236
R230 VGND.n56 VGND.t0 24.9236
R231 VGND.n57 VGND.n55 22.9652
R232 VGND.n20 VGND.n13 21.0829
R233 VGND.n50 VGND.n49 19.9534
R234 VGND.n54 VGND.n1 19.9534
R235 VGND.n26 VGND.n11 19.577
R236 VGND.n36 VGND.n35 18.4476
R237 VGND.n29 VGND.n11 15.0593
R238 VGND.n50 VGND.n1 14.3064
R239 VGND.n55 VGND.n0 9.3005
R240 VGND.n54 VGND.n53 9.3005
R241 VGND.n52 VGND.n1 9.3005
R242 VGND.n51 VGND.n50 9.3005
R243 VGND.n18 VGND.n14 9.3005
R244 VGND.n21 VGND.n20 9.3005
R245 VGND.n22 VGND.n13 9.3005
R246 VGND.n24 VGND.n23 9.3005
R247 VGND.n25 VGND.n12 9.3005
R248 VGND.n27 VGND.n26 9.3005
R249 VGND.n29 VGND.n28 9.3005
R250 VGND.n30 VGND.n9 9.3005
R251 VGND.n32 VGND.n31 9.3005
R252 VGND.n33 VGND.n7 9.3005
R253 VGND.n35 VGND.n34 9.3005
R254 VGND.n36 VGND.n6 9.3005
R255 VGND.n38 VGND.n37 9.3005
R256 VGND.n39 VGND.n5 9.3005
R257 VGND.n41 VGND.n40 9.3005
R258 VGND.n42 VGND.n4 9.3005
R259 VGND.n45 VGND.n44 9.3005
R260 VGND.n46 VGND.n3 9.3005
R261 VGND.n48 VGND.n47 9.3005
R262 VGND.n49 VGND.n2 9.3005
R263 VGND.n17 VGND.n16 7.24166
R264 VGND.n58 VGND.n57 7.12063
R265 VGND.n44 VGND.n43 5.64756
R266 VGND.n43 VGND.n42 4.14168
R267 VGND.n16 VGND.n14 0.508344
R268 VGND.n58 VGND.n0 0.148519
R269 VGND.n21 VGND.n14 0.120292
R270 VGND.n22 VGND.n21 0.120292
R271 VGND.n23 VGND.n22 0.120292
R272 VGND.n23 VGND.n12 0.120292
R273 VGND.n27 VGND.n12 0.120292
R274 VGND.n28 VGND.n27 0.120292
R275 VGND.n28 VGND.n9 0.120292
R276 VGND.n32 VGND.n9 0.120292
R277 VGND.n33 VGND.n32 0.120292
R278 VGND.n34 VGND.n33 0.120292
R279 VGND.n34 VGND.n6 0.120292
R280 VGND.n38 VGND.n6 0.120292
R281 VGND.n39 VGND.n38 0.120292
R282 VGND.n40 VGND.n39 0.120292
R283 VGND.n40 VGND.n4 0.120292
R284 VGND.n45 VGND.n4 0.120292
R285 VGND.n46 VGND.n45 0.120292
R286 VGND.n47 VGND.n46 0.120292
R287 VGND.n47 VGND.n2 0.120292
R288 VGND.n51 VGND.n2 0.120292
R289 VGND.n52 VGND.n51 0.120292
R290 VGND.n53 VGND.n52 0.120292
R291 VGND.n53 VGND.n0 0.120292
R292 VGND VGND.n58 0.101821
R293 VNB.t10 VNB.t6 2933.33
R294 VNB.t13 VNB.t10 2747.16
R295 VNB.t12 VNB.t1 2733.98
R296 VNB.t11 VNB.t19 2677.02
R297 VNB.t19 VNB.t16 2512.82
R298 VNB.t3 VNB.t20 2121.68
R299 VNB.t14 VNB.t17 1879.61
R300 VNB.t18 VNB.t5 1863.06
R301 VNB.t15 VNB.t9 1552.1
R302 VNB.t5 VNB.t13 1453.45
R303 VNB.t1 VNB.t2 1366.99
R304 VNB.t9 VNB.t3 1366.99
R305 VNB.t17 VNB.t15 1352.75
R306 VNB.t2 VNB.t4 1310.03
R307 VNB.t4 VNB.t7 1281.55
R308 VNB.t7 VNB.t8 1196.12
R309 VNB.t0 VNB.t11 1196.12
R310 VNB.t20 VNB.t12 1124.92
R311 VNB.t6 VNB.t14 1025.24
R312 VNB.t16 VNB.t18 951.351
R313 VNB VNB.t0 726.215
R314 a_1701_47.t0 a_1701_47.t1 93.5174
R315 a_1758_413.t0 a_1758_413.t1 121.953
R316 a_1946_47.t0 a_1946_47.t1 70.0005
R317 a_2135_47.t0 a_2135_47.n2 388.889
R318 a_2135_47.n2 a_2135_47.t1 344.161
R319 a_2135_47.n2 a_2135_47.n1 253.565
R320 a_2135_47.n1 a_2135_47.t4 212.081
R321 a_2135_47.n0 a_2135_47.t3 212.081
R322 a_2135_47.n1 a_2135_47.t2 139.78
R323 a_2135_47.n0 a_2135_47.t5 139.78
R324 a_2135_47.n1 a_2135_47.n0 61.346
R325 SCD.n0 SCD.t0 248.767
R326 SCD.n0 SCD.t1 191.998
R327 SCD SCD.n0 155.072
R328 a_817_66.t0 a_817_66.t1 60.0005
R329 SCE.t2 SCE.t3 729.321
R330 SCE.n0 SCE.t0 273.134
R331 SCE.n1 SCE.t2 215.901
R332 SCE SCE.n1 159.054
R333 SCE.n1 SCE.n0 145.296
R334 SCE.n0 SCE.t1 138.173
R335 a_538_389.t0 a_538_389.t1 94.8524
R336 RESET_B.n1 RESET_B.t0 2026.37
R337 RESET_B.n0 RESET_B.t2 398.99
R338 RESET_B.n1 RESET_B.t3 204.458
R339 RESET_B.n3 RESET_B.n0 163.06
R340 RESET_B.n2 RESET_B.n1 157.826
R341 RESET_B.n0 RESET_B.t1 136.21
R342 RESET_B.n4 RESET_B 11.2557
R343 RESET_B.n3 RESET_B.n2 9.43939
R344 RESET_B.n4 RESET_B.n3 9.30982
R345 RESET_B.n2 RESET_B 5.91708
R346 RESET_B RESET_B.n4 3.75222
R347 D.n0 D.t0 234.942
R348 D.n0 D.t1 164.25
R349 D D.n0 157.819
R350 a_569_119.t0 a_569_119.t1 60.0005
R351 a_1187_47.n0 a_1187_47.t0 9.47418
R352 a_1293_47.t0 a_1293_47.t1 60.0005
R353 Q_N Q_N.n0 239.123
R354 Q_N Q_N.n1 116.588
R355 Q_N.n0 Q_N.t1 26.5955
R356 Q_N.n0 Q_N.t0 26.5955
R357 Q_N.n1 Q_N.t2 24.9236
R358 Q_N.n1 Q_N.t3 24.9236
R359 CLK.n0 CLK.t0 428.579
R360 CLK.n0 CLK.t1 426.168
R361 CLK.n1 CLK.n0 152
R362 CLK.n1 CLK 10.4234
R363 CLK CLK.n1 2.01193
C0 a_1079_413# RESET_B 0.146062f
C1 SCD a_1079_413# 2.16e-19
C2 VGND Q 0.117924f
C3 VGND RESET_B 0.270701f
C4 Q VPWR 0.013756f
C5 VGND SCE 0.086893f
C6 VPWR RESET_B 0.07406f
C7 SCE VPWR 0.066374f
C8 CLK RESET_B 2.16e-20
C9 CLK SCE 2.38e-19
C10 VGND SCD 0.069739f
C11 SCD VPWR 0.01224f
C12 D RESET_B 8.56e-20
C13 D SCE 0.051599f
C14 D SCD 0.005659f
C15 VGND a_1079_413# 0.126685f
C16 a_1079_413# VPWR 0.068775f
C17 D a_1079_413# 2.79e-20
C18 VGND VPWR 0.092871f
C19 VGND CLK 0.017295f
C20 CLK VPWR 0.01885f
C21 VGND D 0.001786f
C22 D VPWR 0.062452f
C23 Q_N VPB 0.004363f
C24 Q VPB 0.002075f
C25 VPB RESET_B 0.152772f
C26 VPB SCE 0.182158f
C27 SCD VPB 0.06936f
C28 Q Q_N 0.005911f
C29 Q_N RESET_B 3.23e-19
C30 Q_N SCD 7.96e-23
C31 VPB a_1079_413# 0.09595f
C32 VGND VPB 0.012136f
C33 VPB VPWR 0.287728f
C34 VPB CLK 0.040886f
C35 D VPB 0.068911f
C36 Q RESET_B 0.001081f
C37 SCE RESET_B 1.82e-19
C38 Q SCD 3.64e-21
C39 SCD RESET_B 4.26e-19
C40 SCD SCE 0.033759f
C41 VGND Q_N 0.14259f
C42 Q_N VPWR 0.152099f
C43 Q_N VNB 0.026888f
C44 Q VNB 0.004144f
C45 VGND VNB 1.47394f
C46 RESET_B VNB 0.268513f
C47 VPWR VNB 1.20019f
C48 SCD VNB 0.13368f
C49 D VNB 0.093585f
C50 SCE VNB 0.51427f
C51 CLK VNB 0.15698f
C52 VPB VNB 2.60741f
C53 a_1079_413# VNB 0.150381f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrbp_1 VPB VNB VPWR VGND Q_N SCE SCD D RESET_B CLK Q
X0 a_193_47.t1 a_27_47.t2 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_780_389.t0 a_299_66.t2 a_620_389.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.82 as=0.1755 ps=1.19 w=0.54 l=0.15
X2 VGND.t10 a_1767_21.t3 a_2324_47.t0 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3 a_1245_303.t3 a_1079_413# VPWR.t11 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.2184 ps=2.2 w=0.84 l=0.15
X4 VPWR.t2 a_1592_47.t4 a_1767_21.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND.t9 a_1767_21.t4 a_1701_47.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06705 ps=0.75 w=0.42 l=0.15
X6 a_1758_413.t0 a_193_47.t2 a_1592_47.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0546 pd=0.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR.t4 a_1767_21.t5 a_2324_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8 a_1767_21.t1 a_1592_47.t5 a_1946_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.05145 ps=0.665 w=0.42 l=0.15
X9 VGND.t3 SCD.t0 a_817_66.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.18
X10 a_538_389.t0 SCE.t0 VPWR.t12 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0702 pd=0.8 as=0.0729 ps=0.81 w=0.54 l=0.15
X11 VPWR.t7 SCD.t1 a_780_389.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.64 as=0.0756 ps=0.82 w=0.54 l=0.15
X12 VPWR.t1 SCE.t1 a_299_66.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.189 ps=1.78 w=0.54 l=0.15
X13 a_1767_21.t2 RESET_B.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X14 a_193_47.t0 a_27_47.t3 VGND.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_620_389.t1 D.t0 a_569_119.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.110275 pd=1.065 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_1293_47.t1 a_1245_303.t4 a_1187_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0759 ps=0.8 w=0.42 l=0.15
X17 a_620_389.t5 D.t1 a_538_389.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1755 pd=1.19 as=0.0702 ps=0.8 w=0.54 l=0.15
X18 a_569_119.t0 a_299_66.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 VPWR.t9 a_1767_21.t6 a_1758_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0546 ps=0.68 w=0.42 l=0.15
X20 VGND.t1 RESET_B.t1 a_1293_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 Q.t1 a_1767_21.t7 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 Q.t0 a_1767_21.t8 VGND.t11 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X23 Q_N.t0 a_2324_47.t2 VGND.t8 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X24 a_1191_413.t0 RESET_B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1007 ps=0.94 w=0.42 l=0.15
X25 a_1079_413# a_27_47.t4 a_620_389.t3 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.063 pd=0.71 as=0.0936 ps=1.24 w=0.36 l=0.15
X26 a_1946_47.t0 RESET_B.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.05145 pd=0.665 as=0.12495 ps=1.015 w=0.42 l=0.15
X27 Q_N.t1 a_2324_47.t3 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X28 a_1701_47.t0 a_27_47.t5 a_1592_47.t0 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X29 a_1592_47.t2 a_193_47.t3 a_1245_303.t1 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X30 VGND.t0 SCE.t2 a_299_66.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_1592_47.t1 a_27_47.t6 a_1245_303.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12075 ps=1.165 w=0.42 l=0.15
X32 a_1245_303.t2 a_1079_413# VGND.t7 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1346 ps=1.15 w=0.64 l=0.15
X33 a_1079_413# a_193_47.t4 a_620_389.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0861 pd=0.83 as=0.1533 ps=1.57 w=0.42 l=0.15
X34 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X35 a_817_66.t1 SCE.t3 a_620_389.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.110275 ps=1.065 w=0.42 l=0.5
X36 VGND.t6 CLK.t1 a_27_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n4 a_27_47.n3 532.726
R1 a_27_47.n2 a_27_47.t6 496.003
R2 a_27_47.t0 a_27_47.n0 391.175
R3 a_27_47.n4 a_27_47.t4 279.101
R4 a_27_47.n0 a_27_47.t1 271.212
R5 a_27_47.n1 a_27_47.t2 241.536
R6 a_27_47.n2 a_27_47.t5 199.762
R7 a_27_47.n5 a_27_47.n2 170.347
R8 a_27_47.n1 a_27_47.t3 169.237
R9 a_27_47.n5 a_27_47.n4 164.312
R10 a_27_47.n0 a_27_47.n1 152
R11 a_27_47.n0 a_27_47.n5 14.0789
R12 VPWR.n8 VPWR.t11 806.511
R13 VPWR.n36 VPWR.t7 700.982
R14 VPWR.n29 VPWR.t0 688.191
R15 VPWR.n16 VPWR.t2 663.062
R16 VPWR.n43 VPWR.n42 615.871
R17 VPWR.n50 VPWR.n1 604.394
R18 VPWR.n11 VPWR.n10 603.433
R19 VPWR.n14 VPWR.n13 318.031
R20 VPWR.n15 VPWR.t10 250.464
R21 VPWR.n10 VPWR.t9 114.918
R22 VPWR.n10 VPWR.t5 63.3219
R23 VPWR.n42 VPWR.t12 49.2505
R24 VPWR.n42 VPWR.t1 49.2505
R25 VPWR.n13 VPWR.t6 36.1587
R26 VPWR.n13 VPWR.t4 36.1587
R27 VPWR.n40 VPWR.n4 34.6358
R28 VPWR.n41 VPWR.n40 34.6358
R29 VPWR.n44 VPWR.n41 34.6358
R30 VPWR.n48 VPWR.n2 34.6358
R31 VPWR.n49 VPWR.n48 34.6358
R32 VPWR.n30 VPWR.n6 34.6358
R33 VPWR.n34 VPWR.n6 34.6358
R34 VPWR.n35 VPWR.n34 34.6358
R35 VPWR.n22 VPWR.n21 34.6358
R36 VPWR.n23 VPWR.n22 34.6358
R37 VPWR.n28 VPWR.n27 31.3563
R38 VPWR.n1 VPWR.t3 29.5505
R39 VPWR.n36 VPWR.n4 29.3652
R40 VPWR.n21 VPWR.n11 29.3652
R41 VPWR.n1 VPWR.t8 26.5955
R42 VPWR.n43 VPWR.n2 25.224
R43 VPWR.n23 VPWR.n8 22.9652
R44 VPWR.n50 VPWR.n49 21.8358
R45 VPWR.n17 VPWR.n11 21.0829
R46 VPWR.n16 VPWR.n15 20.3299
R47 VPWR.n30 VPWR.n29 19.7527
R48 VPWR.n27 VPWR.n8 18.4476
R49 VPWR.n17 VPWR.n16 17.3181
R50 VPWR.n36 VPWR.n35 15.0593
R51 VPWR.n44 VPWR.n43 9.41227
R52 VPWR.n16 VPWR.n12 9.3005
R53 VPWR.n18 VPWR.n17 9.3005
R54 VPWR.n19 VPWR.n11 9.3005
R55 VPWR.n21 VPWR.n20 9.3005
R56 VPWR.n22 VPWR.n9 9.3005
R57 VPWR.n24 VPWR.n23 9.3005
R58 VPWR.n25 VPWR.n8 9.3005
R59 VPWR.n27 VPWR.n26 9.3005
R60 VPWR.n28 VPWR.n7 9.3005
R61 VPWR.n31 VPWR.n30 9.3005
R62 VPWR.n32 VPWR.n6 9.3005
R63 VPWR.n34 VPWR.n33 9.3005
R64 VPWR.n35 VPWR.n5 9.3005
R65 VPWR.n37 VPWR.n36 9.3005
R66 VPWR.n38 VPWR.n4 9.3005
R67 VPWR.n40 VPWR.n39 9.3005
R68 VPWR.n41 VPWR.n3 9.3005
R69 VPWR.n45 VPWR.n44 9.3005
R70 VPWR.n46 VPWR.n2 9.3005
R71 VPWR.n48 VPWR.n47 9.3005
R72 VPWR.n49 VPWR.n0 9.3005
R73 VPWR.n51 VPWR.n50 7.18025
R74 VPWR.n15 VPWR.n14 7.0068
R75 VPWR.n29 VPWR.n28 2.70272
R76 VPWR.n14 VPWR.n12 0.231742
R77 VPWR.n51 VPWR.n0 0.147761
R78 VPWR.n18 VPWR.n12 0.120292
R79 VPWR.n19 VPWR.n18 0.120292
R80 VPWR.n20 VPWR.n19 0.120292
R81 VPWR.n20 VPWR.n9 0.120292
R82 VPWR.n24 VPWR.n9 0.120292
R83 VPWR.n25 VPWR.n24 0.120292
R84 VPWR.n26 VPWR.n25 0.120292
R85 VPWR.n26 VPWR.n7 0.120292
R86 VPWR.n31 VPWR.n7 0.120292
R87 VPWR.n32 VPWR.n31 0.120292
R88 VPWR.n33 VPWR.n32 0.120292
R89 VPWR.n33 VPWR.n5 0.120292
R90 VPWR.n37 VPWR.n5 0.120292
R91 VPWR.n38 VPWR.n37 0.120292
R92 VPWR.n39 VPWR.n38 0.120292
R93 VPWR.n39 VPWR.n3 0.120292
R94 VPWR.n45 VPWR.n3 0.120292
R95 VPWR.n46 VPWR.n45 0.120292
R96 VPWR.n47 VPWR.n46 0.120292
R97 VPWR.n47 VPWR.n0 0.120292
R98 VPWR VPWR.n51 0.113006
R99 a_193_47.n0 a_193_47.t3 342.533
R100 a_193_47.n2 a_193_47.n1 338.877
R101 a_193_47.t1 a_193_47.n4 332.233
R102 a_193_47.n0 a_193_47.t2 307.817
R103 a_193_47.n4 a_193_47.t0 302.798
R104 a_193_47.n2 a_193_47.t4 300.252
R105 a_193_47.n3 a_193_47.n2 15.9565
R106 a_193_47.n4 a_193_47.n3 13.0278
R107 a_193_47.n3 a_193_47.n0 11.9849
R108 VPB.t11 VPB.t0 917.446
R109 VPB.t10 VPB.t1 774.313
R110 VPB.t8 VPB.t11 637.548
R111 VPB.t2 VPB.t14 556.386
R112 VPB.t0 VPB.t16 556.386
R113 VPB.t15 VPB.t7 511.784
R114 VPB.t14 VPB 414.33
R115 VPB.t13 VPB.t5 313.707
R116 VPB.t16 VPB.t9 281.154
R117 VPB.t7 VPB.t8 275.084
R118 VPB.t1 VPB.t17 268.688
R119 VPB.t17 VPB.t15 262.291
R120 VPB.t4 VPB.t6 260.437
R121 VPB.t3 VPB.t10 257.478
R122 VPB.t9 VPB.t12 254.518
R123 VPB.t5 VPB.t2 248.599
R124 VPB.t12 VPB.t13 242.679
R125 VPB VPB.t3 177.571
R126 VPB VPB.t4 142.056
R127 a_299_66.n0 a_299_66.t2 1108.99
R128 a_299_66.t0 a_299_66.n0 700.674
R129 a_299_66.n0 a_299_66.t3 346.219
R130 a_299_66.n0 a_299_66.t1 288.474
R131 a_620_389.n0 a_620_389.t4 686.09
R132 a_620_389.n3 a_620_389.n2 599.683
R133 a_620_389.n0 a_620_389.t3 360.05
R134 a_620_389.n2 a_620_389.n1 276.555
R135 a_620_389.n3 a_620_389.t5 162.344
R136 a_620_389.n1 a_620_389.t2 106.636
R137 a_620_389.n2 a_620_389.n0 83.2005
R138 a_620_389.t0 a_620_389.n3 74.7875
R139 a_620_389.n1 a_620_389.t1 38.5724
R140 a_780_389.t0 a_780_389.t1 102.148
R141 a_1767_21.n2 a_1767_21.t6 1015.03
R142 a_1767_21.n5 a_1767_21.n4 783.903
R143 a_1767_21.n3 a_1767_21.n2 257.036
R144 a_1767_21.n0 a_1767_21.t5 239.393
R145 a_1767_21.n3 a_1767_21.t1 223.571
R146 a_1767_21.n1 a_1767_21.t7 212.081
R147 a_1767_21.n2 a_1767_21.t4 178.585
R148 a_1767_21.n4 a_1767_21.n1 173.925
R149 a_1767_21.n0 a_1767_21.t3 154.24
R150 a_1767_21.n1 a_1767_21.t8 139.78
R151 a_1767_21.n1 a_1767_21.n0 132.916
R152 a_1767_21.n4 a_1767_21.n3 64.0131
R153 a_1767_21.t0 a_1767_21.n5 63.3219
R154 a_1767_21.n5 a_1767_21.t2 63.3219
R155 a_2324_47.t1 a_2324_47.n1 405.735
R156 a_2324_47.n1 a_2324_47.t0 294.611
R157 a_2324_47.n0 a_2324_47.t3 254.389
R158 a_2324_47.n0 a_2324_47.t2 211.01
R159 a_2324_47.n1 a_2324_47.n0 152
R160 VGND.n13 VGND.t11 290.289
R161 VGND.n43 VGND.t2 252.274
R162 VGND.n1 VGND.t0 241.996
R163 VGND.n36 VGND.t3 241.22
R164 VGND.n15 VGND.n14 205.746
R165 VGND.n11 VGND.n10 205.707
R166 VGND.n28 VGND.n8 199.739
R167 VGND.n50 VGND.n49 199.739
R168 VGND.n10 VGND.t4 117.144
R169 VGND.n8 VGND.t1 72.8576
R170 VGND.n8 VGND.t7 60.5809
R171 VGND.n10 VGND.t9 52.8576
R172 VGND.n18 VGND.n17 34.6358
R173 VGND.n19 VGND.n18 34.6358
R174 VGND.n23 VGND.n22 34.6358
R175 VGND.n24 VGND.n23 34.6358
R176 VGND.n24 VGND.n7 34.6358
R177 VGND.n30 VGND.n29 34.6358
R178 VGND.n30 VGND.n5 34.6358
R179 VGND.n34 VGND.n5 34.6358
R180 VGND.n35 VGND.n34 34.6358
R181 VGND.n37 VGND.n3 34.6358
R182 VGND.n41 VGND.n3 34.6358
R183 VGND.n42 VGND.n41 34.6358
R184 VGND.n48 VGND.n47 34.6358
R185 VGND.n17 VGND.n13 34.2593
R186 VGND.n14 VGND.t8 33.462
R187 VGND.n14 VGND.t10 33.462
R188 VGND.n28 VGND.n7 25.977
R189 VGND.n49 VGND.t5 24.9236
R190 VGND.n49 VGND.t6 24.9236
R191 VGND.n50 VGND.n48 22.9652
R192 VGND.n43 VGND.n42 19.9534
R193 VGND.n47 VGND.n1 19.9534
R194 VGND.n19 VGND.n11 19.577
R195 VGND.n29 VGND.n28 18.4476
R196 VGND.n22 VGND.n11 15.0593
R197 VGND.n43 VGND.n1 14.3064
R198 VGND.n48 VGND.n0 9.3005
R199 VGND.n47 VGND.n46 9.3005
R200 VGND.n45 VGND.n1 9.3005
R201 VGND.n44 VGND.n43 9.3005
R202 VGND.n17 VGND.n16 9.3005
R203 VGND.n18 VGND.n12 9.3005
R204 VGND.n20 VGND.n19 9.3005
R205 VGND.n22 VGND.n21 9.3005
R206 VGND.n23 VGND.n9 9.3005
R207 VGND.n25 VGND.n24 9.3005
R208 VGND.n26 VGND.n7 9.3005
R209 VGND.n28 VGND.n27 9.3005
R210 VGND.n29 VGND.n6 9.3005
R211 VGND.n31 VGND.n30 9.3005
R212 VGND.n32 VGND.n5 9.3005
R213 VGND.n34 VGND.n33 9.3005
R214 VGND.n35 VGND.n4 9.3005
R215 VGND.n38 VGND.n37 9.3005
R216 VGND.n39 VGND.n3 9.3005
R217 VGND.n41 VGND.n40 9.3005
R218 VGND.n42 VGND.n2 9.3005
R219 VGND.n15 VGND.n13 7.91825
R220 VGND.n51 VGND.n50 7.12063
R221 VGND.n37 VGND.n36 5.64756
R222 VGND.n36 VGND.n35 4.14168
R223 VGND.n16 VGND.n15 0.205869
R224 VGND.n51 VGND.n0 0.148519
R225 VGND.n16 VGND.n12 0.120292
R226 VGND.n20 VGND.n12 0.120292
R227 VGND.n21 VGND.n20 0.120292
R228 VGND.n21 VGND.n9 0.120292
R229 VGND.n25 VGND.n9 0.120292
R230 VGND.n26 VGND.n25 0.120292
R231 VGND.n27 VGND.n26 0.120292
R232 VGND.n27 VGND.n6 0.120292
R233 VGND.n31 VGND.n6 0.120292
R234 VGND.n32 VGND.n31 0.120292
R235 VGND.n33 VGND.n32 0.120292
R236 VGND.n33 VGND.n4 0.120292
R237 VGND.n38 VGND.n4 0.120292
R238 VGND.n39 VGND.n38 0.120292
R239 VGND.n40 VGND.n39 0.120292
R240 VGND.n40 VGND.n2 0.120292
R241 VGND.n44 VGND.n2 0.120292
R242 VGND.n45 VGND.n44 0.120292
R243 VGND.n46 VGND.n45 0.120292
R244 VGND.n46 VGND.n0 0.120292
R245 VGND VGND.n51 0.101821
R246 VNB.t10 VNB.t0 2933.33
R247 VNB.t1 VNB.t16 2748.22
R248 VNB.t5 VNB.t10 2747.16
R249 VNB.t11 VNB.t2 2677.02
R250 VNB.t2 VNB.t4 2512.82
R251 VNB.t17 VNB.t6 2121.68
R252 VNB.t16 VNB 1993.53
R253 VNB.t3 VNB.t14 1879.61
R254 VNB.t7 VNB.t8 1863.06
R255 VNB.t12 VNB.t9 1552.1
R256 VNB.t8 VNB.t5 1453.45
R257 VNB.t9 VNB.t17 1366.99
R258 VNB.t14 VNB.t12 1352.75
R259 VNB.t18 VNB.t15 1253.07
R260 VNB.t13 VNB.t11 1196.12
R261 VNB.t6 VNB.t1 1124.92
R262 VNB.t0 VNB.t3 1025.24
R263 VNB.t4 VNB.t7 951.351
R264 VNB VNB.t13 726.215
R265 VNB VNB.t18 683.495
R266 a_1245_303.n4 a_1245_303.n3 644.628
R267 a_1245_303.n1 a_1245_303.t4 365.918
R268 a_1245_303.n3 a_1245_303.n2 269.793
R269 a_1245_303.n3 a_1245_303.n1 227.672
R270 a_1245_303.n1 a_1245_303.n0 158.392
R271 a_1245_303.n4 a_1245_303.t0 72.7029
R272 a_1245_303.n2 a_1245_303.t1 63.3338
R273 a_1245_303.t3 a_1245_303.n4 50.4231
R274 a_1245_303.n2 a_1245_303.t2 26.7713
R275 a_1592_47.n1 a_1592_47.t5 1025.84
R276 a_1592_47.n3 a_1592_47.n2 635.218
R277 a_1592_47.n1 a_1592_47.t4 412.283
R278 a_1592_47.n2 a_1592_47.n0 302.889
R279 a_1592_47.n2 a_1592_47.n1 220.894
R280 a_1592_47.n0 a_1592_47.t2 70.0005
R281 a_1592_47.t1 a_1592_47.n3 68.0124
R282 a_1592_47.n3 a_1592_47.t3 63.3219
R283 a_1592_47.n0 a_1592_47.t0 61.6672
R284 a_1701_47.t1 a_1701_47.t0 93.5174
R285 a_1758_413.t0 a_1758_413.t1 121.953
R286 a_1946_47.t0 a_1946_47.t1 70.0005
R287 SCD.n0 SCD.t0 248.767
R288 SCD.n0 SCD.t1 191.998
R289 SCD SCD.n0 155.072
R290 a_817_66.t0 a_817_66.t1 60.0005
R291 SCE.t2 SCE.t3 729.321
R292 SCE.n0 SCE.t0 273.134
R293 SCE.n1 SCE.t2 215.901
R294 SCE SCE.n1 159.054
R295 SCE.n1 SCE.n0 145.296
R296 SCE.n0 SCE.t1 138.173
R297 a_538_389.t0 a_538_389.t1 94.8524
R298 RESET_B.n1 RESET_B.t0 2026.37
R299 RESET_B.n0 RESET_B.t2 398.99
R300 RESET_B.n1 RESET_B.t3 204.458
R301 RESET_B.n3 RESET_B.n0 163.06
R302 RESET_B.n2 RESET_B.n1 157.826
R303 RESET_B.n0 RESET_B.t1 136.21
R304 RESET_B.n4 RESET_B 11.2557
R305 RESET_B.n3 RESET_B.n2 9.43939
R306 RESET_B.n4 RESET_B.n3 9.30982
R307 RESET_B.n2 RESET_B 5.91708
R308 RESET_B RESET_B.n4 3.75222
R309 D.n0 D.t0 234.942
R310 D.n0 D.t1 164.25
R311 D D.n0 157.819
R312 a_569_119.t0 a_569_119.t1 60.0005
R313 a_1187_47.n0 a_1187_47.t0 9.47418
R314 a_1293_47.t0 a_1293_47.t1 60.0005
R315 Q.n2 Q.t1 353.606
R316 Q.n0 Q.t0 209.923
R317 Q.n1 Q 89.6005
R318 Q.n1 Q.n0 64.8093
R319 Q Q.n1 16.0005
R320 Q.n0 Q 10.0928
R321 Q.n2 Q 9.10538
R322 Q Q.n2 7.47898
R323 Q.n1 Q 0.738962
R324 Q_N Q_N.t1 382.396
R325 Q_N Q_N.t0 291.714
R326 CLK.n0 CLK.t0 428.579
R327 CLK.n0 CLK.t1 426.168
R328 CLK.n1 CLK.n0 152
R329 CLK.n1 CLK 10.4234
R330 CLK CLK.n1 2.01193
C0 Q_N VPWR 0.089681f
C1 VPWR D 0.062452f
C2 VPWR CLK 0.01885f
C3 SCD VPWR 0.01224f
C4 VPWR VGND 0.075715f
C5 Q VPWR 0.100294f
C6 Q_N VGND 0.054631f
C7 VPWR SCE 0.066374f
C8 VGND D 0.001786f
C9 Q D 1.13e-21
C10 SCD D 0.005659f
C11 VPWR VPB 0.282335f
C12 CLK VGND 0.017295f
C13 Q_N VPB 0.013082f
C14 SCE D 0.051599f
C15 VPB D 0.068911f
C16 CLK SCE 2.38e-19
C17 VPB CLK 0.040886f
C18 VPWR a_1079_413# 0.068775f
C19 a_1079_413# D 2.79e-20
C20 SCD VGND 0.06974f
C21 VPWR RESET_B 0.07406f
C22 Q SCD 3.09e-21
C23 Q VGND 0.05776f
C24 Q_N RESET_B 2.46e-19
C25 VGND SCE 0.086893f
C26 RESET_B D 8.56e-20
C27 SCD SCE 0.033759f
C28 VPB VGND 0.014605f
C29 CLK RESET_B 2.16e-20
C30 SCD VPB 0.06936f
C31 Q VPB 0.011015f
C32 VPB SCE 0.182158f
C33 SCD a_1079_413# 2.16e-19
C34 VGND a_1079_413# 0.126685f
C35 VPB a_1079_413# 0.09595f
C36 SCD RESET_B 4.26e-19
C37 RESET_B VGND 0.271028f
C38 Q RESET_B 0.001328f
C39 RESET_B SCE 1.82e-19
C40 VPB RESET_B 0.152772f
C41 RESET_B a_1079_413# 0.146062f
C42 Q_N VNB 0.093794f
C43 Q VNB 0.012452f
C44 VGND VNB 1.40475f
C45 RESET_B VNB 0.269957f
C46 VPWR VNB 1.12848f
C47 SCD VNB 0.13368f
C48 D VNB 0.093585f
C49 SCE VNB 0.51427f
C50 CLK VNB 0.15698f
C51 VPB VNB 2.51881f
C52 a_1079_413# VNB 0.150381f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfbbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbp_1 VGND VPWR VPB VNB CLK SCD SCE D SET_B RESET_B Q_N
+ Q
X0 a_381_363.t1 SCD.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_1107_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2 VPWR.t9 a_1400_21.t2 a_2122_329.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X3 Q.t0 a_2596_47.t2 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X4 a_931_47.t2 a_193_47.t2 a_453_363.t5 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07035 ps=0.755 w=0.42 l=0.15
X5 a_1251_47.t0 a_1400_21.t3 a_1107_21# VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 VPWR.t11 SCE.t0 a_423_315.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1407 ps=1.51 w=0.42 l=0.15
X7 VPWR.t7 RESET_B.t0 a_1400_21.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1539 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 VPWR.t12 CLK.t0 a_27_47.t0 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_1572_329.t1 a_1107_21# VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1743 pd=1.41 as=0.2247 ps=1.375 w=0.84 l=0.15
X10 a_2122_329.t1 a_1714_47.t4 a_1887_21.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.12285 ps=1.17 w=0.84 l=0.15
X11 a_2026_47.t2 SET_B.t0 VGND.t12 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.09575 pd=0.965 as=0.08295 ps=0.815 w=0.42 l=0.15
X12 VGND.t10 a_1887_21.t4 a_1822_47.t1 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08295 pd=0.815 as=0.066 ps=0.745 w=0.42 l=0.15
X13 a_1041_47.t1 a_193_47.t3 a_931_47.t3 VNB.t21 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X14 VPWR.t4 a_1107_21# a_1017_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X15 a_1107_21# a_931_47.t4 a_1251_47.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.09575 ps=0.965 w=0.64 l=0.15
X16 VPWR.t13 a_1887_21.t5 a_1800_413.t0 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X17 a_764_47.t1 a_423_315.t2 VGND.t8 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.07245 ps=0.765 w=0.42 l=0.15
X18 a_1887_21.t1 a_1714_47.t5 a_2026_47.t0 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.09575 ps=0.965 w=0.64 l=0.15
X19 a_1887_21.t3 SET_B.t1 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X20 a_1800_413.t1 a_193_47.t4 a_1714_47.t2 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 a_931_47.t1 a_27_47.t2 a_453_363.t2 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X22 a_193_47.t1 a_27_47.t3 VGND.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_453_363.t3 D.t0 a_764_47.t0 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 VGND.t7 SCE.t1 a_423_315.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.07245 pd=0.765 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_1714_47.t0 a_27_47.t4 a_1572_329.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1743 ps=1.41 w=0.42 l=0.15
X26 VGND.t5 a_1107_21# a_1041_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X27 a_2026_47.t1 a_1400_21.t4 a_1887_21.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 Q.t1 a_2596_47.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X29 VGND.t9 a_1887_21.t6 a_2596_47.t1 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 a_193_47.t0 a_27_47.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X31 a_1017_413.t0 a_27_47.t6 a_931_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 a_453_363.t1 SCE.t2 a_381_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0504 ps=0.66 w=0.42 l=0.15
X33 VPWR.t1 a_1887_21.t7 a_2596_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X34 a_453_363.t0 a_423_315.t3 a_381_363.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X35 a_381_47.t0 SCD.t1 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X36 a_1822_47.t0 a_27_47.t7 a_1714_47.t1 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0702 ps=0.75 w=0.36 l=0.15
X37 Q_N.t0 a_1887_21.t8 VGND.t11 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X38 Q_N.t1 a_1887_21.t9 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1539 ps=1.335 w=1 l=0.15
X39 a_1714_47.t3 a_193_47.t5 a_1618_47.t1 VNB.t20 sky130_fd_pr__special_nfet_01v8 ad=0.0702 pd=0.75 as=0.0944 ps=0.97 w=0.36 l=0.15
X40 a_453_363.t4 D.t1 a_752_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X41 a_1618_47.t0 a_1107_21# VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0944 pd=0.97 as=0.1664 ps=1.8 w=0.64 l=0.15
X42 a_752_413.t0 SCE.t3 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 VGND.t2 CLK.t1 a_27_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X44 VGND.t3 RESET_B.t1 a_1400_21.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 SCD.n0 SCD.t1 302.411
R1 SCD.n0 SCD.t0 173.877
R2 SCD SCD.n0 154.058
R3 VPWR.n22 VPWR.t9 793.365
R4 VPWR.n16 VPWR.n15 732.75
R5 VPWR.n43 VPWR.t4 686.259
R6 VPWR.n58 VPWR.n1 604.394
R7 VPWR.n50 VPWR.n5 601.292
R8 VPWR.n29 VPWR.n28 585
R9 VPWR.n37 VPWR.t5 397.274
R10 VPWR.n56 VPWR.t3 376.099
R11 VPWR.n18 VPWR.n17 321.339
R12 VPWR.n28 VPWR.t10 91.4648
R13 VPWR.n28 VPWR.t13 91.4648
R14 VPWR.n5 VPWR.t2 63.3219
R15 VPWR.n5 VPWR.t11 63.3219
R16 VPWR.n15 VPWR.t7 63.1021
R17 VPWR.n17 VPWR.t1 58.4849
R18 VPWR.n1 VPWR.t0 41.5552
R19 VPWR.n1 VPWR.t12 41.5552
R20 VPWR.n51 VPWR.n3 34.6358
R21 VPWR.n55 VPWR.n3 34.6358
R22 VPWR.n45 VPWR.n44 34.6358
R23 VPWR.n45 VPWR.n6 34.6358
R24 VPWR.n49 VPWR.n6 34.6358
R25 VPWR.n38 VPWR.n9 34.6358
R26 VPWR.n42 VPWR.n9 34.6358
R27 VPWR.n31 VPWR.n30 34.6358
R28 VPWR.n31 VPWR.n11 34.6358
R29 VPWR.n35 VPWR.n11 34.6358
R30 VPWR.n36 VPWR.n35 34.6358
R31 VPWR.n23 VPWR.n13 34.6358
R32 VPWR.n17 VPWR.t6 31.831
R33 VPWR.n44 VPWR.n43 31.2476
R34 VPWR.n27 VPWR.n13 28.9134
R35 VPWR.n15 VPWR.t8 28.0332
R36 VPWR.n51 VPWR.n50 24.0946
R37 VPWR.n57 VPWR.n56 22.9652
R38 VPWR.n58 VPWR.n57 22.9652
R39 VPWR.n56 VPWR.n55 21.4593
R40 VPWR.n50 VPWR.n49 20.3299
R41 VPWR.n30 VPWR.n29 18.1464
R42 VPWR.n23 VPWR.n22 13.6287
R43 VPWR.n21 VPWR.n20 10.706
R44 VPWR.n20 VPWR.n16 10.1241
R45 VPWR.n43 VPWR.n42 9.41227
R46 VPWR.n20 VPWR.n19 9.3005
R47 VPWR.n21 VPWR.n14 9.3005
R48 VPWR.n24 VPWR.n23 9.3005
R49 VPWR.n25 VPWR.n13 9.3005
R50 VPWR.n27 VPWR.n26 9.3005
R51 VPWR.n30 VPWR.n12 9.3005
R52 VPWR.n32 VPWR.n31 9.3005
R53 VPWR.n33 VPWR.n11 9.3005
R54 VPWR.n35 VPWR.n34 9.3005
R55 VPWR.n36 VPWR.n10 9.3005
R56 VPWR.n39 VPWR.n38 9.3005
R57 VPWR.n40 VPWR.n9 9.3005
R58 VPWR.n42 VPWR.n41 9.3005
R59 VPWR.n43 VPWR.n8 9.3005
R60 VPWR.n44 VPWR.n7 9.3005
R61 VPWR.n46 VPWR.n45 9.3005
R62 VPWR.n47 VPWR.n6 9.3005
R63 VPWR.n49 VPWR.n48 9.3005
R64 VPWR.n50 VPWR.n4 9.3005
R65 VPWR.n52 VPWR.n51 9.3005
R66 VPWR.n53 VPWR.n3 9.3005
R67 VPWR.n55 VPWR.n54 9.3005
R68 VPWR.n56 VPWR.n2 9.3005
R69 VPWR.n57 VPWR.n0 9.3005
R70 VPWR.n18 VPWR.n16 7.84364
R71 VPWR.n59 VPWR.n58 7.12063
R72 VPWR.n37 VPWR.n36 6.4005
R73 VPWR.n22 VPWR.n21 3.8405
R74 VPWR.n38 VPWR.n37 3.38874
R75 VPWR.n29 VPWR.n27 2.44414
R76 VPWR.n19 VPWR.n18 0.211436
R77 VPWR.n59 VPWR.n0 0.148519
R78 VPWR.n19 VPWR.n14 0.120292
R79 VPWR.n24 VPWR.n14 0.120292
R80 VPWR.n25 VPWR.n24 0.120292
R81 VPWR.n26 VPWR.n25 0.120292
R82 VPWR.n26 VPWR.n12 0.120292
R83 VPWR.n32 VPWR.n12 0.120292
R84 VPWR.n33 VPWR.n32 0.120292
R85 VPWR.n34 VPWR.n33 0.120292
R86 VPWR.n34 VPWR.n10 0.120292
R87 VPWR.n39 VPWR.n10 0.120292
R88 VPWR.n40 VPWR.n39 0.120292
R89 VPWR.n41 VPWR.n40 0.120292
R90 VPWR.n41 VPWR.n8 0.120292
R91 VPWR.n8 VPWR.n7 0.120292
R92 VPWR.n46 VPWR.n7 0.120292
R93 VPWR.n47 VPWR.n46 0.120292
R94 VPWR.n48 VPWR.n47 0.120292
R95 VPWR.n48 VPWR.n4 0.120292
R96 VPWR.n52 VPWR.n4 0.120292
R97 VPWR.n53 VPWR.n52 0.120292
R98 VPWR.n54 VPWR.n53 0.120292
R99 VPWR.n54 VPWR.n2 0.120292
R100 VPWR.n2 VPWR.n0 0.120292
R101 VPWR VPWR.n59 0.114842
R102 a_381_363.t0 a_381_363.t1 64.6411
R103 VPB.t7 VPB.t8 1287.38
R104 VPB.t3 VPB.t16 636.293
R105 VPB.t12 VPB.t10 588.942
R106 VPB.t11 VPB.t4 556.386
R107 VPB.t1 VPB.t6 556.386
R108 VPB.t8 VPB.t0 426.168
R109 VPB.t2 VPB.t7 355.14
R110 VPB.t20 VPB.t18 349.221
R111 VPB.t18 VPB.t15 319.627
R112 VPB.t10 VPB.t11 287.072
R113 VPB.t13 VPB.t19 287.072
R114 VPB.t15 VPB.t14 284.113
R115 VPB.t4 VPB.t9 281.154
R116 VPB.t0 VPB.t20 248.599
R117 VPB.t19 VPB.t2 248.599
R118 VPB.t5 VPB.t13 248.599
R119 VPB.t16 VPB.t5 248.599
R120 VPB.t17 VPB.t1 248.599
R121 VPB.t14 VPB.t12 213.084
R122 VPB.t6 VPB.t3 213.084
R123 VPB VPB.t17 142.056
R124 SET_B.n2 SET_B.n0 389.618
R125 SET_B.n3 SET_B.t1 386.848
R126 SET_B.n4 SET_B.n3 178.222
R127 SET_B.n4 SET_B.n2 157.042
R128 SET_B.n3 SET_B.t0 142.635
R129 SET_B.n2 SET_B.n1 142.569
R130 SET_B SET_B.n4 5.0092
R131 SET_B.n4 SET_B 3.29747
R132 a_1400_21.t1 a_1400_21.n4 740.542
R133 a_1400_21.n1 a_1400_21.t0 287.966
R134 a_1400_21.n4 a_1400_21.n3 211.846
R135 a_1400_21.n0 a_1400_21.t4 211.513
R136 a_1400_21.n0 a_1400_21.t2 206.935
R137 a_1400_21.n3 a_1400_21.n2 204.869
R138 a_1400_21.n3 a_1400_21.t3 204.411
R139 a_1400_21.n1 a_1400_21.n0 152
R140 a_1400_21.n4 a_1400_21.n1 9.77505
R141 a_2122_329.t0 a_2122_329.t1 49.2505
R142 a_2596_47.t0 a_2596_47.n1 384.125
R143 a_2596_47.n1 a_2596_47.t1 243.28
R144 a_2596_47.n0 a_2596_47.t2 238.59
R145 a_2596_47.n1 a_2596_47.n0 175.079
R146 a_2596_47.n0 a_2596_47.t3 166.291
R147 Q.n1 Q.t0 353.606
R148 Q.n0 Q.t1 209.923
R149 Q Q.n0 69.451
R150 Q.n1 Q 9.10538
R151 Q Q.n1 7.47898
R152 Q.n0 Q 6.64665
R153 a_193_47.n1 a_193_47.t2 533.949
R154 a_193_47.t0 a_193_47.n3 424.863
R155 a_193_47.n0 a_193_47.t4 343.399
R156 a_193_47.n0 a_193_47.t5 283.659
R157 a_193_47.n3 a_193_47.t1 242.915
R158 a_193_47.n2 a_193_47.n1 164.76
R159 a_193_47.n1 a_193_47.t3 141.923
R160 a_193_47.n3 a_193_47.n2 12.8956
R161 a_193_47.n2 a_193_47.n0 12.1452
R162 a_453_363.n2 a_453_363.n0 648.148
R163 a_453_363.t0 a_453_363.n3 404.389
R164 a_453_363.n3 a_453_363.t1 270.257
R165 a_453_363.n2 a_453_363.n1 225.96
R166 a_453_363.n0 a_453_363.t5 93.81
R167 a_453_363.n1 a_453_363.t2 63.3338
R168 a_453_363.n0 a_453_363.t4 63.3219
R169 a_453_363.n3 a_453_363.n2 33.8555
R170 a_453_363.n1 a_453_363.t3 29.7268
R171 a_931_47.n4 a_931_47.n3 707.533
R172 a_931_47.n3 a_931_47.n0 288.925
R173 a_931_47.n2 a_931_47.t4 216.9
R174 a_931_47.n3 a_931_47.n2 216.829
R175 a_931_47.n2 a_931_47.n1 210.474
R176 a_931_47.n0 a_931_47.t1 70.0005
R177 a_931_47.n0 a_931_47.t3 63.3338
R178 a_931_47.t0 a_931_47.n4 63.3219
R179 a_931_47.n4 a_931_47.t2 63.3219
R180 a_1251_47.t0 a_1251_47.t1 509.728
R181 VNB.t10 VNB.t17 2976.05
R182 VNB.t6 VNB.t4 2933.33
R183 VNB.t14 VNB.t18 2677.02
R184 VNB.t2 VNB.t8 2677.02
R185 VNB.t3 VNB.t9 2677.02
R186 VNB.t12 VNB.t7 2677.02
R187 VNB.t11 VNB.t21 1566.34
R188 VNB.t19 VNB.t22 1552.1
R189 VNB.t20 VNB.t0 1537.86
R190 VNB.t4 VNB.t5 1409.71
R191 VNB.t8 VNB.t14 1381.23
R192 VNB.t9 VNB.t20 1366.99
R193 VNB.t21 VNB.t10 1366.99
R194 VNB.t18 VNB.t1 1352.75
R195 VNB.t22 VNB.t16 1352.75
R196 VNB.t0 VNB.t19 1352.75
R197 VNB.t15 VNB.t11 1352.75
R198 VNB.t16 VNB.t2 1196.12
R199 VNB.t17 VNB.t3 1196.12
R200 VNB.t13 VNB.t12 1196.12
R201 VNB.t7 VNB.t6 1110.68
R202 VNB.t5 VNB.t15 1025.24
R203 VNB VNB.t13 683.495
R204 SCE.n1 SCE.n0 310.087
R205 SCE.n2 SCE.n1 296.029
R206 SCE.n0 SCE.t3 228.148
R207 SCE.n3 SCE.n2 157.272
R208 SCE.n2 SCE.t2 97.2038
R209 SCE.n0 SCE.t0 93.1872
R210 SCE.n1 SCE.t1 93.1872
R211 SCE SCE.n3 29.3823
R212 SCE.n3 SCE 10.1823
R213 a_423_315.t0 a_423_315.n1 719.841
R214 a_423_315.n1 a_423_315.t3 467.93
R215 a_423_315.n0 a_423_315.t2 285.834
R216 a_423_315.n0 a_423_315.t1 281.849
R217 a_423_315.n1 a_423_315.n0 89.0358
R218 RESET_B.n0 RESET_B.t1 203.042
R219 RESET_B.n0 RESET_B.t0 174.123
R220 RESET_B RESET_B.n0 154.111
R221 CLK.n0 CLK.t0 272.062
R222 CLK.n0 CLK.t1 236.716
R223 CLK.n1 CLK.n0 152
R224 CLK CLK.n1 7.6805
R225 CLK.n1 CLK 4.75479
R226 a_27_47.n2 a_27_47.t7 524.309
R227 a_27_47.t0 a_27_47.n5 389.055
R228 a_27_47.n3 a_27_47.t2 312.796
R229 a_27_47.n3 a_27_47.t6 307.325
R230 a_27_47.n1 a_27_47.t1 287.17
R231 a_27_47.n0 a_27_47.t5 262.945
R232 a_27_47.n0 a_27_47.t3 227.597
R233 a_27_47.n4 a_27_47.n2 171.565
R234 a_27_47.n1 a_27_47.n0 152
R235 a_27_47.n2 a_27_47.t4 148.35
R236 a_27_47.n5 a_27_47.n1 35.3396
R237 a_27_47.n5 a_27_47.n4 12.8956
R238 a_27_47.n4 a_27_47.n3 9.3005
R239 a_1572_329.t1 a_1572_329.t0 236.869
R240 a_1714_47.n3 a_1714_47.n2 692.294
R241 a_1714_47.n2 a_1714_47.n0 275.937
R242 a_1714_47.n1 a_1714_47.t4 241.536
R243 a_1714_47.n2 a_1714_47.n1 235.919
R244 a_1714_47.n1 a_1714_47.t5 196.549
R245 a_1714_47.n0 a_1714_47.t3 70.0005
R246 a_1714_47.n3 a_1714_47.t2 63.3219
R247 a_1714_47.t0 a_1714_47.n3 63.3219
R248 a_1714_47.n0 a_1714_47.t1 60.0005
R249 a_1887_21.n6 a_1887_21.n5 594.413
R250 a_1887_21.n4 a_1887_21.t4 386.848
R251 a_1887_21.n3 a_1887_21.n1 305.288
R252 a_1887_21.n3 a_1887_21.n2 277.892
R253 a_1887_21.n1 a_1887_21.t9 268.313
R254 a_1887_21.n0 a_1887_21.t7 231.945
R255 a_1887_21.n5 a_1887_21.n4 204.841
R256 a_1887_21.n1 a_1887_21.t8 196.013
R257 a_1887_21.n0 a_1887_21.t6 164.464
R258 a_1887_21.n1 a_1887_21.n0 151.742
R259 a_1887_21.n4 a_1887_21.t5 142.635
R260 a_1887_21.n6 a_1887_21.t3 91.4648
R261 a_1887_21.t0 a_1887_21.n6 32.8338
R262 a_1887_21.n5 a_1887_21.n3 30.4946
R263 a_1887_21.n2 a_1887_21.t2 25.313
R264 a_1887_21.n2 a_1887_21.t1 25.313
R265 VGND.n38 VGND.t5 287.135
R266 VGND.n31 VGND.t6 280.289
R267 VGND.n55 VGND.t4 247.636
R268 VGND.n14 VGND.n13 207.882
R269 VGND.n24 VGND.n23 202.724
R270 VGND.n58 VGND.n57 199.739
R271 VGND.n49 VGND.n4 198.964
R272 VGND.n16 VGND.n15 110.672
R273 VGND.n23 VGND.t12 70.0005
R274 VGND.n4 VGND.t7 60.0005
R275 VGND.n15 VGND.t3 57.8264
R276 VGND.n13 VGND.t9 54.2862
R277 VGND.n23 VGND.t10 42.8576
R278 VGND.n4 VGND.t8 38.5719
R279 VGND.n57 VGND.t1 38.5719
R280 VGND.n57 VGND.t2 38.5719
R281 VGND.n17 VGND.n12 34.6358
R282 VGND.n21 VGND.n12 34.6358
R283 VGND.n22 VGND.n21 34.6358
R284 VGND.n25 VGND.n22 34.6358
R285 VGND.n29 VGND.n10 34.6358
R286 VGND.n30 VGND.n29 34.6358
R287 VGND.n32 VGND.n30 34.6358
R288 VGND.n36 VGND.n8 34.6358
R289 VGND.n37 VGND.n36 34.6358
R290 VGND.n39 VGND.n37 34.6358
R291 VGND.n43 VGND.n6 34.6358
R292 VGND.n44 VGND.n43 34.6358
R293 VGND.n45 VGND.n44 34.6358
R294 VGND.n45 VGND.n3 34.6358
R295 VGND.n51 VGND.n50 34.6358
R296 VGND.n51 VGND.n1 34.6358
R297 VGND.n50 VGND.n49 28.6123
R298 VGND.n55 VGND.n1 27.4829
R299 VGND.n13 VGND.t0 25.9346
R300 VGND.n15 VGND.t11 24.7418
R301 VGND.n56 VGND.n55 22.9652
R302 VGND.n58 VGND.n56 22.9652
R303 VGND.n17 VGND.n16 20.3299
R304 VGND.n39 VGND.n38 18.0711
R305 VGND.n38 VGND.n6 16.5652
R306 VGND.n49 VGND.n3 15.8123
R307 VGND.n24 VGND.n10 9.78874
R308 VGND.n56 VGND.n0 9.3005
R309 VGND.n55 VGND.n54 9.3005
R310 VGND.n53 VGND.n1 9.3005
R311 VGND.n52 VGND.n51 9.3005
R312 VGND.n50 VGND.n2 9.3005
R313 VGND.n49 VGND.n48 9.3005
R314 VGND.n47 VGND.n3 9.3005
R315 VGND.n46 VGND.n45 9.3005
R316 VGND.n44 VGND.n5 9.3005
R317 VGND.n43 VGND.n42 9.3005
R318 VGND.n41 VGND.n6 9.3005
R319 VGND.n40 VGND.n39 9.3005
R320 VGND.n37 VGND.n7 9.3005
R321 VGND.n36 VGND.n35 9.3005
R322 VGND.n34 VGND.n8 9.3005
R323 VGND.n33 VGND.n32 9.3005
R324 VGND.n30 VGND.n9 9.3005
R325 VGND.n29 VGND.n28 9.3005
R326 VGND.n27 VGND.n10 9.3005
R327 VGND.n26 VGND.n25 9.3005
R328 VGND.n22 VGND.n11 9.3005
R329 VGND.n21 VGND.n20 9.3005
R330 VGND.n19 VGND.n12 9.3005
R331 VGND.n18 VGND.n17 9.3005
R332 VGND.n59 VGND.n58 7.12063
R333 VGND.n16 VGND.n14 7.10092
R334 VGND.n32 VGND.n31 5.64756
R335 VGND.n25 VGND.n24 5.27109
R336 VGND.n31 VGND.n8 3.76521
R337 VGND.n18 VGND.n14 0.218009
R338 VGND.n59 VGND.n0 0.148519
R339 VGND.n19 VGND.n18 0.120292
R340 VGND.n20 VGND.n19 0.120292
R341 VGND.n20 VGND.n11 0.120292
R342 VGND.n26 VGND.n11 0.120292
R343 VGND.n27 VGND.n26 0.120292
R344 VGND.n28 VGND.n27 0.120292
R345 VGND.n28 VGND.n9 0.120292
R346 VGND.n33 VGND.n9 0.120292
R347 VGND.n34 VGND.n33 0.120292
R348 VGND.n35 VGND.n34 0.120292
R349 VGND.n35 VGND.n7 0.120292
R350 VGND.n40 VGND.n7 0.120292
R351 VGND.n41 VGND.n40 0.120292
R352 VGND.n42 VGND.n41 0.120292
R353 VGND.n42 VGND.n5 0.120292
R354 VGND.n46 VGND.n5 0.120292
R355 VGND.n47 VGND.n46 0.120292
R356 VGND.n48 VGND.n47 0.120292
R357 VGND.n48 VGND.n2 0.120292
R358 VGND.n52 VGND.n2 0.120292
R359 VGND.n53 VGND.n52 0.120292
R360 VGND.n54 VGND.n53 0.120292
R361 VGND.n54 VGND.n0 0.120292
R362 VGND VGND.n59 0.114842
R363 a_2026_47.n0 a_2026_47.t1 457.231
R364 a_2026_47.t0 a_2026_47.n0 42.0094
R365 a_2026_47.n0 a_2026_47.t2 38.5719
R366 a_1822_47.t1 a_1822_47.t0 93.0601
R367 a_1041_47.t0 a_1041_47.t1 93.5174
R368 a_1017_413.t0 a_1017_413.t1 211.071
R369 a_1800_413.t0 a_1800_413.t1 206.381
R370 a_764_47.t0 a_764_47.t1 60.0005
R371 D.n0 D.t0 308.481
R372 D.n0 D.t1 224.934
R373 D.n1 D.n0 152
R374 D.n1 D 40.6405
R375 D D.n1 2.8805
R376 a_381_47.t0 a_381_47.t1 68.5719
R377 Q_N.n1 Q_N.t1 353.795
R378 Q_N.n0 Q_N.t0 209.923
R379 Q_N Q_N.n0 79.4391
R380 Q_N.n1 Q_N 8.2361
R381 Q_N Q_N.n1 6.90173
R382 Q_N.n0 Q_N 5.61454
R383 a_1618_47.n0 a_1618_47.t1 68.3338
R384 a_1618_47.n1 a_1618_47.n0 67.2005
R385 a_1618_47.n0 a_1618_47.t0 13.144
R386 a_752_413.t0 a_752_413.t1 126.644
C0 RESET_B Q 6.25e-20
C1 VPWR Q 0.099121f
C2 VPWR RESET_B 0.009858f
C3 VPB Q 0.012264f
C4 VPB RESET_B 0.047075f
C5 VPB VPWR 0.306924f
C6 RESET_B D 3.53e-21
C7 VPWR SCD 0.042724f
C8 VPWR D 0.04608f
C9 VPB SCD 0.07562f
C10 VPB D 0.086201f
C11 VGND a_1107_21# 0.052207f
C12 SET_B a_1107_21# 0.174486f
C13 VPWR a_1351_329# 0.009837f
C14 RESET_B a_1107_21# 6.51e-21
C15 VPWR a_1107_21# 0.15986f
C16 VPB a_1107_21# 0.14068f
C17 a_1351_329# a_1107_21# 0.010422f
C18 VGND Q_N 0.086192f
C19 CLK VGND 0.01947f
C20 Q_N SET_B 3.62e-19
C21 VGND SCE 0.072336f
C22 VGND SET_B 0.295728f
C23 RESET_B Q_N 0.001681f
C24 VGND Q 0.064306f
C25 VGND RESET_B 0.028707f
C26 VPWR Q_N 0.061427f
C27 VPWR VGND 0.084754f
C28 VPB Q_N 0.010224f
C29 CLK VPWR 0.019459f
C30 VPB VGND 0.016647f
C31 Q SET_B 1.21e-19
C32 RESET_B SET_B 0.002334f
C33 VGND SCD 0.029712f
C34 VPWR SCE 0.038333f
C35 VPWR SET_B 0.025404f
C36 VGND D 0.01764f
C37 VPB CLK 0.070599f
C38 VPB SCE 0.131544f
C39 SCD SCE 0.10925f
C40 VPB SET_B 0.144895f
C41 SCE D 0.052343f
C42 Q VNB 0.09443f
C43 Q_N VNB 0.013507f
C44 RESET_B VNB 0.132613f
C45 VGND VNB 1.54697f
C46 VPWR VNB 1.24623f
C47 SET_B VNB 0.265223f
C48 D VNB 0.112806f
C49 SCE VNB 0.304916f
C50 SCD VNB 0.129448f
C51 CLK VNB 0.196677f
C52 VPB VNB 2.81966f
C53 a_1107_21# VNB 0.239078f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbn_2 VGND VPWR VPB VNB CLK_N SCD SCE D SET_B RESET_B
+ Q_N Q
X0 a_381_363.t0 SCD.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_1107_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X2 VPWR.t11 a_1401_21.t2 a_2122_329.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X3 a_931_47.t1 a_27_47.t2 a_453_47.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07035 ps=0.755 w=0.42 l=0.15
X4 VPWR.t12 SCE.t0 a_423_315.t1 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1407 ps=1.51 w=0.42 l=0.15
X5 VPWR.t0 CLK_N.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_1572_329.t0 a_1107_21# VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1743 pd=1.41 as=0.2247 ps=1.375 w=0.84 l=0.15
X7 a_2122_329.t1 a_1714_47.t3 a_1888_21.t1 VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.12285 ps=1.17 w=0.84 l=0.15
X8 VGND.t10 a_1888_21.t4 a_1823_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X9 a_1041_47.t1 a_27_47.t3 a_931_47.t2 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X10 VPWR.t9 a_1107_21# a_1017_413.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X11 VPWR.t7 a_1888_21.t5 a_1800_413.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 a_1888_21.t0 a_1714_47.t4 a_2004_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.1199 ps=1.08 w=0.64 l=0.15
X13 a_764_47.t0 a_423_315.t2 VGND.t2 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.07245 ps=0.765 w=0.42 l=0.15
X14 Q.t1 a_2696_47.t2 VGND.t4 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X15 a_1888_21.t3 SET_B.t0 VPWR.t14 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X16 a_1800_413.t1 a_27_47.t4 a_1714_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_931_47.t3 a_193_47.t2 a_453_47.t5 VNB.t20 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X18 VGND.t9 a_1888_21.t6 a_2696_47.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 a_193_47.t0 a_27_47.t5 VGND.t12 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR.t13 a_1888_21.t7 a_2696_47.t1 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X21 a_453_47.t4 D.t0 a_764_47.t1 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 VGND.t11 SCE.t1 a_423_315.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.07245 pd=0.765 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 a_1714_47.t2 a_193_47.t3 a_1572_329.t1 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1743 ps=1.41 w=0.42 l=0.15
X24 VPWR.t6 a_1888_21.t8 Q_N.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 a_2004_47.t1 a_1401_21.t3 a_1888_21.t2 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.83 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 VGND.t6 a_1107_21# a_1041_47.t0 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X27 VGND.t7 a_1888_21.t9 Q_N.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VGND.t0 a_2696_47.t3 Q.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VPWR.t8 a_2696_47.t4 Q.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 Q_N.t2 a_1888_21.t10 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X31 a_193_47.t1 a_27_47.t6 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 Q.t2 a_2696_47.t5 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X33 a_1017_413.t1 a_193_47.t4 a_931_47.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X34 Q_N.t0 a_1888_21.t11 VGND.t8 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X35 a_453_47.t1 a_423_315.t3 a_381_363.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X36 a_381_47.t0 SCD.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 a_1714_47.t0 a_27_47.t7 a_1619_47# VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X38 a_453_47.t0 D.t1 a_752_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 a_1251_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0968 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X40 a_1619_47# a_1107_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X41 a_2004_47.t2 SET_B.t1 VGND.t13 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.1199 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X42 VPWR.t15 RESET_B.t0 a_1401_21.t1 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X43 VGND.t3 RESET_B.t1 a_1401_21.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X44 a_752_413.t0 SCE.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 VGND.t5 CLK_N.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X46 a_453_47.t2 SCE.t3 a_381_47.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
R0 SCD.n0 SCD.t1 301.269
R1 SCD.n0 SCD.t0 172.736
R2 SCD SCD.n0 154.058
R3 VPWR.n31 VPWR.t11 793.365
R4 VPWR.n24 VPWR.n23 732.75
R5 VPWR.n52 VPWR.t9 686.259
R6 VPWR.n67 VPWR.n1 604.394
R7 VPWR.n59 VPWR.n5 600.583
R8 VPWR.n38 VPWR.n37 585
R9 VPWR.n46 VPWR.t10 397.274
R10 VPWR.n65 VPWR.t1 374.75
R11 VPWR.n18 VPWR.n17 315.236
R12 VPWR.n19 VPWR.t8 258.538
R13 VPWR.n22 VPWR.t6 252.288
R14 VPWR.n37 VPWR.t14 91.4648
R15 VPWR.n37 VPWR.t7 91.4648
R16 VPWR.n5 VPWR.t2 63.3219
R17 VPWR.n5 VPWR.t12 63.3219
R18 VPWR.n23 VPWR.t15 63.1021
R19 VPWR.n17 VPWR.t13 58.4849
R20 VPWR.n1 VPWR.t4 41.5552
R21 VPWR.n1 VPWR.t0 41.5552
R22 VPWR.n60 VPWR.n3 34.6358
R23 VPWR.n64 VPWR.n3 34.6358
R24 VPWR.n54 VPWR.n53 34.6358
R25 VPWR.n54 VPWR.n6 34.6358
R26 VPWR.n58 VPWR.n6 34.6358
R27 VPWR.n47 VPWR.n9 34.6358
R28 VPWR.n51 VPWR.n9 34.6358
R29 VPWR.n40 VPWR.n39 34.6358
R30 VPWR.n40 VPWR.n11 34.6358
R31 VPWR.n44 VPWR.n11 34.6358
R32 VPWR.n45 VPWR.n44 34.6358
R33 VPWR.n32 VPWR.n13 34.6358
R34 VPWR.n17 VPWR.t5 31.831
R35 VPWR.n53 VPWR.n52 31.2476
R36 VPWR.n36 VPWR.n13 28.9134
R37 VPWR.n21 VPWR.n18 28.6123
R38 VPWR.n23 VPWR.t3 27.7871
R39 VPWR.n25 VPWR.n22 26.3534
R40 VPWR.n22 VPWR.n21 25.224
R41 VPWR.n67 VPWR.n66 22.9652
R42 VPWR.n60 VPWR.n59 22.9652
R43 VPWR.n25 VPWR.n24 21.9111
R44 VPWR.n65 VPWR.n64 21.4593
R45 VPWR.n66 VPWR.n65 21.0829
R46 VPWR.n59 VPWR.n58 20.3299
R47 VPWR.n39 VPWR.n38 18.1464
R48 VPWR.n32 VPWR.n31 13.6287
R49 VPWR.n29 VPWR.n15 10.706
R50 VPWR.n30 VPWR.n29 10.706
R51 VPWR.n52 VPWR.n51 9.41227
R52 VPWR.n21 VPWR.n20 9.3005
R53 VPWR.n22 VPWR.n16 9.3005
R54 VPWR.n26 VPWR.n25 9.3005
R55 VPWR.n27 VPWR.n15 9.3005
R56 VPWR.n29 VPWR.n28 9.3005
R57 VPWR.n30 VPWR.n14 9.3005
R58 VPWR.n33 VPWR.n32 9.3005
R59 VPWR.n34 VPWR.n13 9.3005
R60 VPWR.n36 VPWR.n35 9.3005
R61 VPWR.n39 VPWR.n12 9.3005
R62 VPWR.n41 VPWR.n40 9.3005
R63 VPWR.n42 VPWR.n11 9.3005
R64 VPWR.n44 VPWR.n43 9.3005
R65 VPWR.n45 VPWR.n10 9.3005
R66 VPWR.n48 VPWR.n47 9.3005
R67 VPWR.n49 VPWR.n9 9.3005
R68 VPWR.n51 VPWR.n50 9.3005
R69 VPWR.n52 VPWR.n8 9.3005
R70 VPWR.n53 VPWR.n7 9.3005
R71 VPWR.n55 VPWR.n54 9.3005
R72 VPWR.n56 VPWR.n6 9.3005
R73 VPWR.n58 VPWR.n57 9.3005
R74 VPWR.n59 VPWR.n4 9.3005
R75 VPWR.n61 VPWR.n60 9.3005
R76 VPWR.n62 VPWR.n3 9.3005
R77 VPWR.n64 VPWR.n63 9.3005
R78 VPWR.n65 VPWR.n2 9.3005
R79 VPWR.n66 VPWR.n0 9.3005
R80 VPWR.n68 VPWR.n67 7.12063
R81 VPWR.n46 VPWR.n45 6.4005
R82 VPWR.n19 VPWR.n18 6.29708
R83 VPWR.n31 VPWR.n30 3.8405
R84 VPWR.n47 VPWR.n46 3.38874
R85 VPWR.n38 VPWR.n36 2.44414
R86 VPWR.n24 VPWR.n15 1.2805
R87 VPWR.n20 VPWR.n19 0.669899
R88 VPWR.n68 VPWR.n0 0.148519
R89 VPWR.n20 VPWR.n16 0.120292
R90 VPWR.n26 VPWR.n16 0.120292
R91 VPWR.n27 VPWR.n26 0.120292
R92 VPWR.n28 VPWR.n27 0.120292
R93 VPWR.n28 VPWR.n14 0.120292
R94 VPWR.n33 VPWR.n14 0.120292
R95 VPWR.n34 VPWR.n33 0.120292
R96 VPWR.n35 VPWR.n34 0.120292
R97 VPWR.n35 VPWR.n12 0.120292
R98 VPWR.n41 VPWR.n12 0.120292
R99 VPWR.n42 VPWR.n41 0.120292
R100 VPWR.n43 VPWR.n42 0.120292
R101 VPWR.n43 VPWR.n10 0.120292
R102 VPWR.n48 VPWR.n10 0.120292
R103 VPWR.n49 VPWR.n48 0.120292
R104 VPWR.n50 VPWR.n49 0.120292
R105 VPWR.n50 VPWR.n8 0.120292
R106 VPWR.n8 VPWR.n7 0.120292
R107 VPWR.n55 VPWR.n7 0.120292
R108 VPWR.n56 VPWR.n55 0.120292
R109 VPWR.n57 VPWR.n56 0.120292
R110 VPWR.n57 VPWR.n4 0.120292
R111 VPWR.n61 VPWR.n4 0.120292
R112 VPWR.n62 VPWR.n61 0.120292
R113 VPWR.n63 VPWR.n62 0.120292
R114 VPWR.n63 VPWR.n2 0.120292
R115 VPWR.n2 VPWR.n0 0.120292
R116 VPWR VPWR.n68 0.114842
R117 a_381_363.t0 a_381_363.t1 64.6411
R118 VPB.t13 VPB.t14 1287.38
R119 VPB.t16 VPB.t21 636.293
R120 VPB.t12 VPB.t17 636.293
R121 VPB.t8 VPB.t18 556.386
R122 VPB.t6 VPB.t1 556.386
R123 VPB.t14 VPB.t19 426.168
R124 VPB.t15 VPB.t13 355.14
R125 VPB.t5 VPB.t9 349.221
R126 VPB.t9 VPB.t20 319.627
R127 VPB.t21 VPB.t3 287.072
R128 VPB.t11 VPB.t4 287.072
R129 VPB.t20 VPB.t22 284.113
R130 VPB.t18 VPB.t7 281.154
R131 VPB.t7 VPB.t10 248.599
R132 VPB.t3 VPB.t8 248.599
R133 VPB.t19 VPB.t5 248.599
R134 VPB.t4 VPB.t15 248.599
R135 VPB.t2 VPB.t11 248.599
R136 VPB.t17 VPB.t2 248.599
R137 VPB.t0 VPB.t6 248.599
R138 VPB.t22 VPB.t16 213.084
R139 VPB.t1 VPB.t12 213.084
R140 VPB VPB.t0 142.056
R141 SET_B.n2 SET_B.n0 389.618
R142 SET_B.n3 SET_B.t0 387.207
R143 SET_B.n4 SET_B.n3 178.222
R144 SET_B.n4 SET_B.n2 157.042
R145 SET_B.n3 SET_B.t1 142.994
R146 SET_B.n2 SET_B.n1 142.569
R147 SET_B SET_B.n4 5.0092
R148 SET_B.n4 SET_B 3.29747
R149 a_1401_21.t1 a_1401_21.n5 746.564
R150 a_1401_21.n1 a_1401_21.t0 289.192
R151 a_1401_21.n5 a_1401_21.n4 211.846
R152 a_1401_21.n0 a_1401_21.t3 211.737
R153 a_1401_21.n0 a_1401_21.t2 207.404
R154 a_1401_21.n4 a_1401_21.n3 205.625
R155 a_1401_21.n4 a_1401_21.n2 204.869
R156 a_1401_21.n1 a_1401_21.n0 152
R157 a_1401_21.n5 a_1401_21.n1 9.77505
R158 a_2122_329.t0 a_2122_329.t1 49.2505
R159 VNB.t15 VNB.t10 8216.18
R160 VNB.t17 VNB.t12 3018.77
R161 VNB.t10 VNB.t5 2904.85
R162 VNB.t16 VNB.t6 2890.61
R163 VNB.t4 VNB.t14 2677.02
R164 VNB.t9 VNB.t1 2677.02
R165 VNB.t19 VNB.t7 1680.26
R166 VNB.t20 VNB.t8 1566.34
R167 VNB.t12 VNB.t13 1409.71
R168 VNB.t6 VNB.t3 1381.23
R169 VNB.t8 VNB.t15 1366.99
R170 VNB.t14 VNB.t11 1352.75
R171 VNB.t18 VNB.t20 1352.75
R172 VNB.t5 VNB.t19 1224.6
R173 VNB.t11 VNB.t0 1196.12
R174 VNB.t3 VNB.t4 1196.12
R175 VNB.t7 VNB.t16 1196.12
R176 VNB.t2 VNB.t9 1196.12
R177 VNB.t13 VNB.t18 1025.24
R178 VNB.t1 VNB.t17 1025.24
R179 VNB VNB.t2 683.495
R180 a_27_47.n1 a_27_47.t2 533.949
R181 a_27_47.t0 a_27_47.n5 424.394
R182 a_27_47.n0 a_27_47.t4 343.399
R183 a_27_47.n0 a_27_47.t7 283.3
R184 a_27_47.n3 a_27_47.t1 265.743
R185 a_27_47.n4 a_27_47.t6 262.945
R186 a_27_47.n4 a_27_47.t5 227.597
R187 a_27_47.n2 a_27_47.n1 164.76
R188 a_27_47.n5 a_27_47.n4 152
R189 a_27_47.n1 a_27_47.t3 141.923
R190 a_27_47.n5 a_27_47.n3 21.4266
R191 a_27_47.n3 a_27_47.n2 13.3063
R192 a_27_47.n2 a_27_47.n0 12.1452
R193 a_453_47.n2 a_453_47.n0 648.148
R194 a_453_47.t1 a_453_47.n3 471.418
R195 a_453_47.n3 a_453_47.t2 282.817
R196 a_453_47.n2 a_453_47.n1 225.96
R197 a_453_47.n0 a_453_47.t3 93.81
R198 a_453_47.n1 a_453_47.t5 63.3338
R199 a_453_47.n0 a_453_47.t0 63.3219
R200 a_453_47.n3 a_453_47.n2 33.7313
R201 a_453_47.n1 a_453_47.t4 29.7268
R202 a_931_47.n5 a_931_47.n4 707.533
R203 a_931_47.n4 a_931_47.n0 288.925
R204 a_931_47.n3 a_931_47.n2 216.9
R205 a_931_47.n4 a_931_47.n3 216.829
R206 a_931_47.n3 a_931_47.n1 210.474
R207 a_931_47.n0 a_931_47.t3 70.0005
R208 a_931_47.n0 a_931_47.t2 63.3338
R209 a_931_47.t0 a_931_47.n5 63.3219
R210 a_931_47.n5 a_931_47.t1 63.3219
R211 SCE.n1 SCE.n0 310.087
R212 SCE.n2 SCE.n1 290.406
R213 SCE.n0 SCE.t2 228.148
R214 SCE.n3 SCE.n2 152
R215 SCE.n2 SCE.t3 101.221
R216 SCE.n0 SCE.t0 93.1872
R217 SCE.n1 SCE.t1 93.1872
R218 SCE.n3 SCE 26.0043
R219 SCE SCE.n3 5.86232
R220 a_423_315.n0 a_423_315.t1 719.841
R221 a_423_315.n0 a_423_315.t3 467.93
R222 a_423_315.n1 a_423_315.t2 285.834
R223 a_423_315.t0 a_423_315.n1 284.56
R224 a_423_315.n1 a_423_315.n0 89.0358
R225 CLK_N.n0 CLK_N.t0 272.062
R226 CLK_N.n0 CLK_N.t1 236.716
R227 CLK_N.n1 CLK_N.n0 152
R228 CLK_N CLK_N.n1 7.6805
R229 CLK_N.n1 CLK_N 4.75479
R230 a_1572_329.t0 a_1572_329.t1 236.869
R231 a_1714_47.n2 a_1714_47.n1 692.294
R232 a_1714_47.n1 a_1714_47.t0 345.937
R233 a_1714_47.n0 a_1714_47.t3 241.536
R234 a_1714_47.n1 a_1714_47.n0 235.919
R235 a_1714_47.n0 a_1714_47.t4 196.549
R236 a_1714_47.t1 a_1714_47.n2 63.3219
R237 a_1714_47.n2 a_1714_47.t2 63.3219
R238 a_1888_21.n7 a_1888_21.n6 594.413
R239 a_1888_21.n5 a_1888_21.t4 387.207
R240 a_1888_21.n4 a_1888_21.n2 311.765
R241 a_1888_21.n2 a_1888_21.t10 308.481
R242 a_1888_21.n4 a_1888_21.n3 275.635
R243 a_1888_21.n2 a_1888_21.t11 236.18
R244 a_1888_21.n0 a_1888_21.t7 231.476
R245 a_1888_21.n1 a_1888_21.t8 221.72
R246 a_1888_21.n6 a_1888_21.n5 204.841
R247 a_1888_21.n0 a_1888_21.t6 163.995
R248 a_1888_21.n1 a_1888_21.t9 149.421
R249 a_1888_21.n1 a_1888_21.n0 144.601
R250 a_1888_21.n5 a_1888_21.t5 142.994
R251 a_1888_21.n7 a_1888_21.t3 91.4648
R252 a_1888_21.n2 a_1888_21.n1 85.6894
R253 a_1888_21.t1 a_1888_21.n7 32.8338
R254 a_1888_21.n6 a_1888_21.n4 30.4946
R255 a_1888_21.n3 a_1888_21.t2 25.313
R256 a_1888_21.n3 a_1888_21.t0 25.313
R257 a_1823_47.n0 a_1823_47.t0 11.0774
R258 VGND.n45 VGND.t6 287.135
R259 VGND.n62 VGND.t1 245.448
R260 VGND.n32 VGND.n31 202.724
R261 VGND.n17 VGND.n16 201.488
R262 VGND.n65 VGND.n64 199.739
R263 VGND.n56 VGND.n4 198.964
R264 VGND.n15 VGND.t0 163.38
R265 VGND.n14 VGND.t7 157.02
R266 VGND.n24 VGND.n23 110.672
R267 VGND.n4 VGND.t11 60.0005
R268 VGND.n23 VGND.t3 57.8264
R269 VGND.n16 VGND.t9 54.2862
R270 VGND.n31 VGND.t10 41.4291
R271 VGND.n31 VGND.t13 38.5719
R272 VGND.n4 VGND.t2 38.5719
R273 VGND.n64 VGND.t12 38.5719
R274 VGND.n64 VGND.t5 38.5719
R275 VGND.n25 VGND.n12 34.6358
R276 VGND.n29 VGND.n12 34.6358
R277 VGND.n30 VGND.n29 34.6358
R278 VGND.n33 VGND.n30 34.6358
R279 VGND.n37 VGND.n10 34.6358
R280 VGND.n38 VGND.n37 34.6358
R281 VGND.n39 VGND.n38 34.6358
R282 VGND.n43 VGND.n8 34.6358
R283 VGND.n44 VGND.n43 34.6358
R284 VGND.n46 VGND.n44 34.6358
R285 VGND.n50 VGND.n6 34.6358
R286 VGND.n51 VGND.n50 34.6358
R287 VGND.n52 VGND.n51 34.6358
R288 VGND.n52 VGND.n3 34.6358
R289 VGND.n58 VGND.n57 34.6358
R290 VGND.n58 VGND.n1 34.6358
R291 VGND.n18 VGND.n17 28.6123
R292 VGND.n57 VGND.n56 28.6123
R293 VGND.n62 VGND.n1 27.4829
R294 VGND.n22 VGND.n14 26.3534
R295 VGND.n25 VGND.n24 26.3534
R296 VGND.n16 VGND.t4 25.9346
R297 VGND.n18 VGND.n14 25.224
R298 VGND.n23 VGND.t8 24.7418
R299 VGND.n65 VGND.n63 22.9652
R300 VGND.n63 VGND.n62 21.0829
R301 VGND.n24 VGND.n22 18.0711
R302 VGND.n46 VGND.n45 18.0711
R303 VGND.n45 VGND.n6 16.5652
R304 VGND.n56 VGND.n3 15.8123
R305 VGND.n32 VGND.n10 9.78874
R306 VGND.n39 VGND.n8 9.78873
R307 VGND.n63 VGND.n0 9.3005
R308 VGND.n62 VGND.n61 9.3005
R309 VGND.n60 VGND.n1 9.3005
R310 VGND.n59 VGND.n58 9.3005
R311 VGND.n57 VGND.n2 9.3005
R312 VGND.n56 VGND.n55 9.3005
R313 VGND.n54 VGND.n3 9.3005
R314 VGND.n53 VGND.n52 9.3005
R315 VGND.n51 VGND.n5 9.3005
R316 VGND.n50 VGND.n49 9.3005
R317 VGND.n48 VGND.n6 9.3005
R318 VGND.n47 VGND.n46 9.3005
R319 VGND.n44 VGND.n7 9.3005
R320 VGND.n43 VGND.n42 9.3005
R321 VGND.n41 VGND.n8 9.3005
R322 VGND.n40 VGND.n39 9.3005
R323 VGND.n38 VGND.n9 9.3005
R324 VGND.n37 VGND.n36 9.3005
R325 VGND.n35 VGND.n10 9.3005
R326 VGND.n34 VGND.n33 9.3005
R327 VGND.n30 VGND.n11 9.3005
R328 VGND.n29 VGND.n28 9.3005
R329 VGND.n27 VGND.n12 9.3005
R330 VGND.n26 VGND.n25 9.3005
R331 VGND.n24 VGND.n13 9.3005
R332 VGND.n22 VGND.n21 9.3005
R333 VGND.n20 VGND.n14 9.3005
R334 VGND.n19 VGND.n18 9.3005
R335 VGND.n66 VGND.n65 7.12063
R336 VGND.n17 VGND.n15 6.29708
R337 VGND.n33 VGND.n32 5.27109
R338 VGND.n19 VGND.n15 0.669899
R339 VGND.n66 VGND.n0 0.148519
R340 VGND.n20 VGND.n19 0.120292
R341 VGND.n21 VGND.n20 0.120292
R342 VGND.n21 VGND.n13 0.120292
R343 VGND.n26 VGND.n13 0.120292
R344 VGND.n27 VGND.n26 0.120292
R345 VGND.n28 VGND.n27 0.120292
R346 VGND.n28 VGND.n11 0.120292
R347 VGND.n34 VGND.n11 0.120292
R348 VGND.n35 VGND.n34 0.120292
R349 VGND.n36 VGND.n35 0.120292
R350 VGND.n36 VGND.n9 0.120292
R351 VGND.n40 VGND.n9 0.120292
R352 VGND.n41 VGND.n40 0.120292
R353 VGND.n42 VGND.n41 0.120292
R354 VGND.n42 VGND.n7 0.120292
R355 VGND.n47 VGND.n7 0.120292
R356 VGND.n48 VGND.n47 0.120292
R357 VGND.n49 VGND.n48 0.120292
R358 VGND.n49 VGND.n5 0.120292
R359 VGND.n53 VGND.n5 0.120292
R360 VGND.n54 VGND.n53 0.120292
R361 VGND.n55 VGND.n54 0.120292
R362 VGND.n55 VGND.n2 0.120292
R363 VGND.n59 VGND.n2 0.120292
R364 VGND.n60 VGND.n59 0.120292
R365 VGND.n61 VGND.n60 0.120292
R366 VGND.n61 VGND.n0 0.120292
R367 VGND VGND.n66 0.114842
R368 a_1041_47.t0 a_1041_47.t1 93.5174
R369 a_1017_413.t0 a_1017_413.t1 211.071
R370 a_1800_413.t0 a_1800_413.t1 206.381
R371 a_2004_47.n0 a_2004_47.t1 459.442
R372 a_2004_47.n0 a_2004_47.t2 64.2862
R373 a_2004_47.t0 a_2004_47.n0 49.1523
R374 a_764_47.t0 a_764_47.t1 60.0005
R375 a_2696_47.t1 a_2696_47.n2 384.125
R376 a_2696_47.n2 a_2696_47.t0 243.28
R377 a_2696_47.n0 a_2696_47.t4 212.081
R378 a_2696_47.n1 a_2696_47.t5 212.081
R379 a_2696_47.n2 a_2696_47.n1 187.494
R380 a_2696_47.n0 a_2696_47.t3 139.78
R381 a_2696_47.n1 a_2696_47.t2 139.78
R382 a_2696_47.n1 a_2696_47.n0 61.346
R383 Q Q.n0 586.793
R384 Q.n3 Q.n0 585
R385 Q.n2 Q.n1 185
R386 Q Q.n2 69.6887
R387 Q.n0 Q.t3 26.5955
R388 Q.n0 Q.t2 26.5955
R389 Q.n1 Q.t0 24.9236
R390 Q.n1 Q.t1 24.9236
R391 Q Q.n3 15.6165
R392 Q.n2 Q 6.9125
R393 Q.n3 Q 1.7925
R394 a_193_47.n1 a_193_47.n0 525.917
R395 a_193_47.t1 a_193_47.n4 367.062
R396 a_193_47.n2 a_193_47.t2 312.796
R397 a_193_47.n2 a_193_47.t4 307.325
R398 a_193_47.n4 a_193_47.t0 302.7
R399 a_193_47.n3 a_193_47.n1 171.565
R400 a_193_47.n1 a_193_47.t3 148.35
R401 a_193_47.n4 a_193_47.n3 12.4849
R402 a_193_47.n3 a_193_47.n2 9.3005
R403 D.n0 D.t0 308.481
R404 D.n0 D.t1 224.934
R405 D.n1 D.n0 152
R406 D.n1 D 40.6405
R407 D D.n1 2.8805
R408 Q_N Q_N.n0 586.537
R409 Q_N.n3 Q_N.n0 585
R410 Q_N.n2 Q_N.n1 185
R411 Q_N Q_N.n2 85.2786
R412 Q_N.n0 Q_N.t3 26.5955
R413 Q_N.n0 Q_N.t2 26.5955
R414 Q_N.n1 Q_N.t1 24.9236
R415 Q_N.n1 Q_N.t0 24.9236
R416 Q_N Q_N.n3 15.8725
R417 Q_N.n2 Q_N 6.4005
R418 Q_N.n3 Q_N 1.5365
R419 a_381_47.t0 a_381_47.t1 60.0005
R420 a_752_413.t0 a_752_413.t1 126.644
R421 RESET_B.n0 RESET_B.t1 201.874
R422 RESET_B.n0 RESET_B.t0 172.953
R423 RESET_B RESET_B.n0 154
C0 VGND Q_N 0.134412f
C1 SET_B Q_N 3.06e-19
C2 SET_B VGND 0.292237f
C3 VGND SCD 0.030148f
C4 VPWR CLK_N 0.019459f
C5 CLK_N VPB 0.070599f
C6 VGND a_1251_47# 0.162848f
C7 VPWR a_1351_329# 0.009837f
C8 SET_B a_1251_47# 0.029124f
C9 VGND CLK_N 0.01947f
C10 RESET_B a_1107_21# 6.32e-21
C11 VPWR a_1107_21# 0.15986f
C12 D RESET_B 2.27e-21
C13 a_1107_21# VPB 0.140705f
C14 D VPWR 0.04608f
C15 D VPB 0.086201f
C16 a_1619_47# a_1107_21# 9.75e-19
C17 RESET_B Q 4.25e-20
C18 VPWR Q 0.179079f
C19 Q VPB 0.005707f
C20 VPWR RESET_B 0.01025f
C21 RESET_B VPB 0.049182f
C22 VPWR VPB 0.340272f
C23 a_1619_47# VPWR 6.2e-19
C24 SCE D 0.052343f
C25 VGND a_1107_21# 0.052419f
C26 D VGND 0.01764f
C27 SET_B a_1107_21# 0.174513f
C28 SCE VPWR 0.038339f
C29 SCE VPB 0.133044f
C30 a_1251_47# a_1107_21# 0.069647f
C31 VGND Q 0.115695f
C32 RESET_B Q_N 0.001648f
C33 VPWR Q_N 0.136109f
C34 SET_B Q 9.31e-20
C35 Q_N VPB 0.004297f
C36 VGND RESET_B 0.029382f
C37 VPWR VGND 0.127775f
C38 SET_B RESET_B 0.00216f
C39 VGND VPB 0.020125f
C40 SET_B VPWR 0.025494f
C41 VPWR SCD 0.043231f
C42 SET_B VPB 0.144946f
C43 SCD VPB 0.077138f
C44 a_1619_47# VGND 0.009148f
C45 a_1619_47# SET_B 0.00383f
C46 a_1619_47# a_1251_47# 3.34e-19
C47 SCE VGND 0.073066f
C48 SCE SCD 0.112623f
C49 a_1107_21# a_1351_329# 0.010433f
C50 Q VNB 0.027092f
C51 Q_N VNB 0.010034f
C52 RESET_B VNB 0.136415f
C53 VGND VNB 1.67416f
C54 VPWR VNB 1.35967f
C55 SET_B VNB 0.263389f
C56 D VNB 0.112806f
C57 SCE VNB 0.3013f
C58 SCD VNB 0.130547f
C59 CLK_N VNB 0.196677f
C60 VPB VNB 2.99686f
C61 a_1251_47# VNB 0.013628f
C62 a_1107_21# VNB 0.239034f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfstp_1 SCD CLK D SET_B SCE Q VPWR VGND VPB VNB
X0 VPWR.t6 a_1597_329.t3 a_2227_47.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1506 pd=1.33 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 Q.t0 a_2227_47.t2 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.09805 ps=0.98 w=0.65 l=0.15
X2 a_1597_329.t2 SET_B.t0 VPWR.t8 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0966 ps=0.88 w=0.42 l=0.15
X3 VPWR.t10 SCD.t0 a_27_369.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_1081_413# a_643_369.t2 a_997_413.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_809_369.t0 a_643_369.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND.t5 a_1597_329.t4 a_2227_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.09805 pd=0.98 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_997_413.t0 a_809_369.t2 a_181_47.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR.t9 SET_B.t1 a_1129_21.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.27 as=0.0714 ps=0.76 w=0.42 l=0.15
X9 a_181_47.t1 SCE.t0 a_109_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_1514_47.t0 a_997_413.t4 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.2384 pd=1.385 as=0.09575 ps=0.965 w=0.64 l=0.15
X11 VGND SET_B a_1347_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09575 pd=0.965 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 a_27_369.t0 a_319_21.t2 a_181_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 VGND.t6 SCE.t1 a_319_21.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_1597_329.t0 a_809_369.t3 a_1514_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1241 pd=1.1 as=0.2384 ps=1.385 w=0.64 l=0.15
X15 a_181_47.t4 D.t0 a_193_369.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X16 VGND SET_B a_1887_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_1597_329.t1 a_643_369.t4 a_1525_329.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.32 as=0.0882 ps=1.05 w=0.84 l=0.15
X18 a_265_47.t0 D.t1 a_181_47.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_997_413.t2 a_643_369.t5 a_181_47.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 a_1781_295.t0 a_1597_329.t5 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_1087_47# a_809_369.t4 a_997_413.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_193_369.t1 SCE.t2 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_809_369.t1 a_643_369.t6 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1525_329.t0 a_997_413.t5 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.1428 ps=1.27 w=0.84 l=0.15
X25 VPWR.t5 SCE.t3 a_319_21.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 Q.t1 a_2227_47.t3 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1506 ps=1.33 w=1 l=0.15
X27 VPWR.t4 CLK.t0 a_643_369.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 VGND.t8 a_319_21.t3 a_265_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0567 ps=0.69 w=0.42 l=0.15
X29 VGND.t7 CLK.t1 a_643_369.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 a_1781_295.t1 a_1597_329.t6 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_109_47.t0 SCD.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1597_329.t1 a_1597_329.n4 778.22
R1 a_1597_329.n4 a_1597_329.t2 648.322
R2 a_1597_329.n0 a_1597_329.t0 473.219
R3 a_1597_329.n1 a_1597_329.t4 356.68
R4 a_1597_329.n2 a_1597_329.n1 291.342
R5 a_1597_329.n4 a_1597_329.n3 186.715
R6 a_1597_329.n2 a_1597_329.t6 144.601
R7 a_1597_329.n1 a_1597_329.t3 133.353
R8 a_1597_329.n0 a_1597_329.t5 132.282
R9 a_1597_329.n3 a_1597_329.n0 111.575
R10 a_1597_329.n3 a_1597_329.n2 32.1338
R11 a_2227_47.t0 a_2227_47.n1 391.599
R12 a_2227_47.n1 a_2227_47.t1 250.895
R13 a_2227_47.n0 a_2227_47.t3 241.536
R14 a_2227_47.n1 a_2227_47.n0 178.183
R15 a_2227_47.n0 a_2227_47.t2 169.237
R16 VPWR.n41 VPWR.t5 734.085
R17 VPWR.n18 VPWR.t8 688.083
R18 VPWR.n16 VPWR.t7 663.062
R19 VPWR.n48 VPWR.n1 602.067
R20 VPWR.n5 VPWR.n4 598.965
R21 VPWR.n10 VPWR.n9 585
R22 VPWR.n15 VPWR.n14 319.486
R23 VPWR.n9 VPWR.t1 87.9469
R24 VPWR.n9 VPWR.t9 84.4291
R25 VPWR.n14 VPWR.t6 60.0239
R26 VPWR.n1 VPWR.t2 41.5552
R27 VPWR.n1 VPWR.t10 41.5552
R28 VPWR.n4 VPWR.t0 41.5552
R29 VPWR.n4 VPWR.t4 41.5552
R30 VPWR.n42 VPWR.n2 34.6358
R31 VPWR.n46 VPWR.n2 34.6358
R32 VPWR.n47 VPWR.n46 34.6358
R33 VPWR.n40 VPWR.n39 34.6358
R34 VPWR.n33 VPWR.n7 34.6358
R35 VPWR.n34 VPWR.n33 34.6358
R36 VPWR.n35 VPWR.n34 34.6358
R37 VPWR.n22 VPWR.n12 34.6358
R38 VPWR.n23 VPWR.n22 34.6358
R39 VPWR.n35 VPWR.n5 33.5064
R40 VPWR.n14 VPWR.t3 31.1381
R41 VPWR.n28 VPWR.n27 30.6829
R42 VPWR.n18 VPWR.n17 30.1181
R43 VPWR.n29 VPWR.n28 28.4986
R44 VPWR.n48 VPWR.n47 27.4829
R45 VPWR.n29 VPWR.n7 21.0829
R46 VPWR.n17 VPWR.n16 19.9534
R47 VPWR.n18 VPWR.n12 14.3064
R48 VPWR.n42 VPWR.n41 12.0476
R49 VPWR.n39 VPWR.n5 10.9181
R50 VPWR.n24 VPWR.n23 10.6358
R51 VPWR.n17 VPWR.n13 9.3005
R52 VPWR.n19 VPWR.n18 9.3005
R53 VPWR.n20 VPWR.n12 9.3005
R54 VPWR.n22 VPWR.n21 9.3005
R55 VPWR.n23 VPWR.n11 9.3005
R56 VPWR.n25 VPWR.n24 9.3005
R57 VPWR.n27 VPWR.n26 9.3005
R58 VPWR.n28 VPWR.n8 9.3005
R59 VPWR.n30 VPWR.n29 9.3005
R60 VPWR.n31 VPWR.n7 9.3005
R61 VPWR.n33 VPWR.n32 9.3005
R62 VPWR.n34 VPWR.n6 9.3005
R63 VPWR.n36 VPWR.n35 9.3005
R64 VPWR.n37 VPWR.n5 9.3005
R65 VPWR.n39 VPWR.n38 9.3005
R66 VPWR.n40 VPWR.n3 9.3005
R67 VPWR.n43 VPWR.n42 9.3005
R68 VPWR.n44 VPWR.n2 9.3005
R69 VPWR.n46 VPWR.n45 9.3005
R70 VPWR.n47 VPWR.n0 9.3005
R71 VPWR.n49 VPWR.n48 7.12063
R72 VPWR.n16 VPWR.n15 7.10319
R73 VPWR.n24 VPWR.n10 6.87109
R74 VPWR.n27 VPWR.n10 1.78874
R75 VPWR.n41 VPWR.n40 0.376971
R76 VPWR.n15 VPWR.n13 0.234117
R77 VPWR.n49 VPWR.n0 0.148519
R78 VPWR.n19 VPWR.n13 0.120292
R79 VPWR.n20 VPWR.n19 0.120292
R80 VPWR.n21 VPWR.n20 0.120292
R81 VPWR.n21 VPWR.n11 0.120292
R82 VPWR.n25 VPWR.n11 0.120292
R83 VPWR.n26 VPWR.n25 0.120292
R84 VPWR.n26 VPWR.n8 0.120292
R85 VPWR.n30 VPWR.n8 0.120292
R86 VPWR.n31 VPWR.n30 0.120292
R87 VPWR.n32 VPWR.n31 0.120292
R88 VPWR.n32 VPWR.n6 0.120292
R89 VPWR.n36 VPWR.n6 0.120292
R90 VPWR.n37 VPWR.n36 0.120292
R91 VPWR.n38 VPWR.n37 0.120292
R92 VPWR.n38 VPWR.n3 0.120292
R93 VPWR.n43 VPWR.n3 0.120292
R94 VPWR.n44 VPWR.n43 0.120292
R95 VPWR.n45 VPWR.n44 0.120292
R96 VPWR.n45 VPWR.n0 0.120292
R97 VPWR VPWR.n49 0.114842
R98 VPB.t1 VPB.t13 994.394
R99 VPB.t4 VPB.t14 970.716
R100 VPB.t10 VPB.t11 556.386
R101 VPB.t13 VPB.t10 556.386
R102 VPB.t2 VPB.t0 556.386
R103 VPB.t9 VPB.t8 556.386
R104 VPB.t6 VPB.t9 556.386
R105 VPB.t14 VPB.t3 343.303
R106 VPB.t11 VPB.t7 284.113
R107 VPB.t0 VPB.t4 248.599
R108 VPB.t8 VPB.t2 248.599
R109 VPB.t12 VPB.t6 248.599
R110 VPB.t15 VPB.t5 248.599
R111 VPB.t3 VPB.t1 213.084
R112 VPB.t5 VPB.t12 213.084
R113 VPB VPB.t15 192.369
R114 VGND.n42 VGND.t8 250.499
R115 VGND.n13 VGND.t4 242.004
R116 VGND.n21 VGND.t2 224.153
R117 VGND.n48 VGND.t0 223.571
R118 VGND.n40 VGND.t6 223.571
R119 VGND.n12 VGND.n11 205.856
R120 VGND.n35 VGND.n34 198.964
R121 VGND.n11 VGND.t5 55.7148
R122 VGND.n34 VGND.t1 38.5719
R123 VGND.n34 VGND.t7 38.5719
R124 VGND.n15 VGND.n14 34.6358
R125 VGND.n15 VGND.n9 34.6358
R126 VGND.n19 VGND.n9 34.6358
R127 VGND.n20 VGND.n19 34.6358
R128 VGND.n27 VGND.n26 34.6358
R129 VGND.n32 VGND.n5 34.6358
R130 VGND.n33 VGND.n32 34.6358
R131 VGND.n46 VGND.n1 34.6358
R132 VGND.n47 VGND.n46 34.0711
R133 VGND.n42 VGND.n41 33.1299
R134 VGND.n35 VGND.n33 31.2476
R135 VGND.n39 VGND.n3 28.5534
R136 VGND.n28 VGND.n5 27.3528
R137 VGND.n22 VGND.n20 27.0218
R138 VGND.n11 VGND.t3 25.9346
R139 VGND.n14 VGND.n13 16.9417
R140 VGND.n28 VGND.n27 16.6884
R141 VGND.n42 VGND.n1 16.1887
R142 VGND.n41 VGND.n40 15.2476
R143 VGND.n35 VGND.n3 13.177
R144 VGND.n49 VGND.n48 9.86521
R145 VGND.n14 VGND.n10 9.3005
R146 VGND.n16 VGND.n15 9.3005
R147 VGND.n17 VGND.n9 9.3005
R148 VGND.n19 VGND.n18 9.3005
R149 VGND.n20 VGND.n8 9.3005
R150 VGND.n23 VGND.n22 9.3005
R151 VGND.n24 VGND.n7 9.3005
R152 VGND.n26 VGND.n25 9.3005
R153 VGND.n27 VGND.n6 9.3005
R154 VGND.n29 VGND.n28 9.3005
R155 VGND.n30 VGND.n5 9.3005
R156 VGND.n32 VGND.n31 9.3005
R157 VGND.n33 VGND.n4 9.3005
R158 VGND.n36 VGND.n35 9.3005
R159 VGND.n37 VGND.n3 9.3005
R160 VGND.n39 VGND.n38 9.3005
R161 VGND.n41 VGND.n2 9.3005
R162 VGND.n43 VGND.n42 9.3005
R163 VGND.n44 VGND.n1 9.3005
R164 VGND.n46 VGND.n45 9.3005
R165 VGND.n47 VGND.n0 9.3005
R166 VGND.n26 VGND.n7 8.74815
R167 VGND.n48 VGND.n47 8.09462
R168 VGND.n13 VGND.n12 7.4962
R169 VGND.n22 VGND.n21 5.03421
R170 VGND.n40 VGND.n39 2.8005
R171 VGND.n21 VGND.n7 1.58252
R172 VGND.n12 VGND.n10 0.213852
R173 VGND.n16 VGND.n10 0.120292
R174 VGND.n17 VGND.n16 0.120292
R175 VGND.n18 VGND.n17 0.120292
R176 VGND.n18 VGND.n8 0.120292
R177 VGND.n23 VGND.n8 0.120292
R178 VGND.n24 VGND.n23 0.120292
R179 VGND.n25 VGND.n24 0.120292
R180 VGND.n25 VGND.n6 0.120292
R181 VGND.n29 VGND.n6 0.120292
R182 VGND.n30 VGND.n29 0.120292
R183 VGND.n31 VGND.n30 0.120292
R184 VGND.n31 VGND.n4 0.120292
R185 VGND.n36 VGND.n4 0.120292
R186 VGND.n37 VGND.n36 0.120292
R187 VGND.n38 VGND.n37 0.120292
R188 VGND.n38 VGND.n2 0.120292
R189 VGND.n43 VGND.n2 0.120292
R190 VGND.n44 VGND.n43 0.120292
R191 VGND.n45 VGND.n44 0.120292
R192 VGND.n45 VGND.n0 0.120292
R193 VGND.n49 VGND.n0 0.120292
R194 VGND VGND.n49 0.0226354
R195 Q.n0 Q 591.024
R196 Q.n1 Q.n0 585
R197 Q.n4 Q.t0 209.923
R198 Q.n0 Q.t1 26.5955
R199 Q.n3 Q 18.8637
R200 Q Q.n4 12.2358
R201 Q.n2 Q 10.9181
R202 Q.n1 Q 6.77697
R203 Q Q.n1 6.02403
R204 Q.n3 Q 4.04261
R205 Q Q.n2 3.36892
R206 Q Q.n3 2.25932
R207 Q.n2 Q 1.88285
R208 Q.n4 Q 0.565206
R209 VNB.t7 VNB.t4 6080.26
R210 VNB.t0 VNB.t9 5752.75
R211 VNB.t9 VNB.t10 3018.77
R212 VNB.t13 VNB.t11 2762.46
R213 VNB.t3 VNB.t1 2677.02
R214 VNB.t11 VNB.t12 2677.02
R215 VNB.t4 VNB.t0 2548.87
R216 VNB.t10 VNB.t5 1366.99
R217 VNB.t1 VNB.t7 1196.12
R218 VNB.t12 VNB.t3 1196.12
R219 VNB.t8 VNB.t13 1196.12
R220 VNB.t6 VNB.t8 1196.12
R221 VNB.t2 VNB.t6 1025.24
R222 VNB VNB.t2 925.567
R223 SET_B.n1 SET_B.n0 360.18
R224 SET_B.n3 SET_B.n2 357.216
R225 SET_B.n4 SET_B.n3 223.113
R226 SET_B.n1 SET_B.t1 166.577
R227 SET_B.n3 SET_B.t0 161.03
R228 SET_B.n4 SET_B.n1 159
R229 SET_B SET_B.n4 3.4005
R230 SCD.n0 SCD.t0 299.433
R231 SCD.n0 SCD.t1 206.245
R232 SCD.n1 SCD.n0 152
R233 SCD.n1 SCD 19.828
R234 SCD SCD.n1 14.3064
R235 a_27_369.t0 a_27_369.t1 1468.74
R236 a_643_369.t0 a_643_369.n6 670.312
R237 a_643_369.n4 a_643_369.t4 419.243
R238 a_643_369.n4 a_643_369.n3 413.587
R239 a_643_369.n0 a_643_369.t5 393.634
R240 a_643_369.n5 a_643_369.t2 317.574
R241 a_643_369.n2 a_643_369.t1 291.962
R242 a_643_369.n1 a_643_369.t6 267.3
R243 a_643_369.n2 a_643_369.n1 152
R244 a_643_369.n1 a_643_369.n0 100.206
R245 a_643_369.n0 a_643_369.t3 91.5805
R246 a_643_369.n5 a_643_369.n4 53.8068
R247 a_643_369.n6 a_643_369.n2 30.2774
R248 a_643_369.n6 a_643_369.n5 10.4313
R249 a_997_413.n7 a_997_413.n6 662.052
R250 a_997_413.n3 a_997_413.n1 312.132
R251 a_997_413.n0 a_997_413.t5 262.64
R252 a_997_413.n3 a_997_413.n2 238.226
R253 a_997_413.n6 a_997_413.n5 234.409
R254 a_997_413.n4 a_997_413.n0 200.561
R255 a_997_413.n0 a_997_413.t4 166.24
R256 a_997_413.n4 a_997_413.n3 152
R257 a_997_413.n7 a_997_413.t3 63.3219
R258 a_997_413.t0 a_997_413.n7 63.3219
R259 a_997_413.n6 a_997_413.n4 53.8358
R260 a_997_413.n5 a_997_413.t1 38.5719
R261 a_997_413.n5 a_997_413.t2 38.5719
R262 a_809_369.t1 a_809_369.n4 672.456
R263 a_809_369.n3 a_809_369.t4 433.509
R264 a_809_369.n1 a_809_369.t3 385.065
R265 a_809_369.n3 a_809_369.t2 321.334
R266 a_809_369.n2 a_809_369.t0 275.591
R267 a_809_369.n2 a_809_369.n1 205.534
R268 a_809_369.n4 a_809_369.n3 182.673
R269 a_809_369.n1 a_809_369.n0 148.35
R270 a_809_369.n4 a_809_369.n2 2.5605
R271 a_181_47.n1 a_181_47.t2 693.452
R272 a_181_47.n3 a_181_47.n2 613.688
R273 a_181_47.n2 a_181_47.n0 574.096
R274 a_181_47.n1 a_181_47.t5 288.805
R275 a_181_47.t0 a_181_47.n3 41.5552
R276 a_181_47.n3 a_181_47.t4 41.5552
R277 a_181_47.n0 a_181_47.t3 38.5719
R278 a_181_47.n0 a_181_47.t1 38.5719
R279 a_181_47.n2 a_181_47.n1 22.6251
R280 a_1129_21.t0 a_1129_21.n2 896.688
R281 a_1129_21.n2 a_1129_21.n1 336.712
R282 a_1129_21.n2 a_1129_21.n0 139.822
R283 SCE.n1 SCE.t3 295.168
R284 SCE.n0 SCE.t2 263.18
R285 SCE.n0 SCE.t0 231.73
R286 SCE.n1 SCE.t1 201.982
R287 SCE.n2 SCE.n1 173.305
R288 SCE.n2 SCE.n0 154.744
R289 SCE SCE.n2 3.88621
R290 a_109_47.t0 a_109_47.t1 60.0005
R291 a_1514_47.t0 a_1514_47.t1 139.689
R292 a_1781_295.n3 a_1781_295.t1 697.798
R293 a_1781_295.n2 a_1781_295.n0 453.616
R294 a_1781_295.t0 a_1781_295.n3 302.202
R295 a_1781_295.n3 a_1781_295.n2 252.554
R296 a_1781_295.n2 a_1781_295.n1 161.202
R297 a_319_21.t1 a_319_21.n1 754.953
R298 a_319_21.n0 a_319_21.t2 283.286
R299 a_319_21.n1 a_319_21.t0 259.202
R300 a_319_21.n0 a_319_21.t3 190.101
R301 a_319_21.n1 a_319_21.n0 152
R302 D.n0 D.t0 373.283
R303 D.n1 D.n0 152
R304 D.n0 D.t1 132.282
R305 D.n1 D 23.1303
R306 D D.n1 7.41103
R307 a_193_369.t0 a_193_369.t1 64.6411
R308 a_1525_329.t0 a_1525_329.t1 49.2505
R309 a_265_47.t0 a_265_47.t1 77.1434
R310 CLK.n0 CLK.t0 255.077
R311 CLK.n0 CLK.t1 218.642
R312 CLK.n1 CLK.n0 152
R313 CLK.n1 CLK 19.0712
R314 CLK CLK.n1 2.90959
C0 Q VPWR 0.103233f
C1 VPB Q 0.012688f
C2 VPB VPWR 0.266622f
C3 a_1723_413# VPWR 8.96e-19
C4 VGND Q 0.090934f
C5 Q SET_B 1.23e-19
C6 VGND VPWR 0.082476f
C7 SET_B VPWR 0.100473f
C8 CLK VPWR 0.03f
C9 SCE VPWR 0.064479f
C10 VPB VGND 0.016405f
C11 VPB SET_B 0.198194f
C12 VPB CLK 0.080439f
C13 a_1887_47# VPWR 2.81e-19
C14 VPB SCE 0.130585f
C15 a_1723_413# SET_B 2.84e-19
C16 a_1081_413# VPWR 9.08e-19
C17 VGND SET_B 0.041467f
C18 VGND CLK 0.040331f
C19 D VPWR 0.007869f
C20 SCE VGND 0.142351f
C21 SCD VPWR 0.017326f
C22 SCE CLK 0.090396f
C23 VPB D 0.043648f
C24 a_1887_47# VGND 0.001665f
C25 a_1815_47# VPWR 1.13e-19
C26 VPB SCD 0.070898f
C27 VGND a_1347_47# 0.004877f
C28 VGND a_1087_47# 0.005211f
C29 VGND D 0.008596f
C30 SCD VGND 0.045223f
C31 SCE D 0.20207f
C32 a_1815_47# VGND 0.001224f
C33 a_1815_47# SET_B 4.89e-19
C34 SCD SCE 0.170177f
C35 Q VNB 0.091182f
C36 VGND VNB 1.37378f
C37 VPWR VNB 1.08748f
C38 SET_B VNB 0.219168f
C39 CLK VNB 0.13687f
C40 D VNB 0.104133f
C41 SCE VNB 0.253779f
C42 SCD VNB 0.205442f
C43 VPB VNB 2.46528f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfstp_2 VPWR VGND VPB VNB SCD SCE D CLK SET_B Q
X0 VPWR.t7 a_1597_329.t3 a_2227_47.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 VPWR.t9 a_2227_47.t2 Q.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 Q.t3 a_2227_47.t3 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.097 ps=0.975 w=0.65 l=0.15
X3 a_1597_329.t2 SET_B.t0 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0966 ps=0.88 w=0.42 l=0.15
X4 VPWR.t3 SCD.t0 a_27_369.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_1081_413.t0 a_643_369.t2 a_997_413.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_809_369.t1 a_643_369.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND.t7 a_1597_329.t4 a_2227_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_997_413.t0 a_809_369.t2 a_181_47.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VPWR.t2 SET_B.t1 a_1129_21# VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.27 as=0.0714 ps=0.76 w=0.42 l=0.15
X10 a_181_47.t2 SCE.t0 a_109_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 a_1514_47.t0 a_997_413.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.2384 pd=1.385 as=0.09575 ps=0.965 w=0.64 l=0.15
X12 VGND SET_B a_1347_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09575 pd=0.965 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 a_27_369.t1 a_319_21.t2 a_181_47.t5 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14 VGND.t4 SCE.t1 a_319_21.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1597_329.t0 a_809_369.t3 a_1514_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1241 pd=1.1 as=0.2384 ps=1.385 w=0.64 l=0.15
X16 a_181_47.t0 D.t0 a_193_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X17 VGND SET_B a_1887_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1597_329.t1 a_643_369.t4 a_1525_329.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.32 as=0.0882 ps=1.05 w=0.84 l=0.15
X19 a_265_47.t0 D.t1 a_181_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_997_413.t2 a_643_369.t5 a_181_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VGND.t8 a_2227_47.t4 Q.t2 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X22 Q.t0 a_2227_47.t5 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.149 ps=1.325 w=1 l=0.15
X23 a_1781_295.t1 a_1597_329.t5 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.0882 ps=0.84 w=0.42 l=0.15
X24 a_1087_47.t0 a_809_369.t4 a_997_413.t3 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X25 a_193_369.t0 SCE.t2 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 a_809_369.t0 a_643_369.t6 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_1525_329.t1 a_997_413.t5 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.1428 ps=1.27 w=0.84 l=0.15
X28 VPWR.t5 SCE.t3 a_319_21.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 VPWR.t11 CLK.t0 a_643_369.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X30 VGND.t5 a_319_21.t3 a_265_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0567 ps=0.69 w=0.42 l=0.15
X31 VGND.t3 CLK.t1 a_643_369.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_1781_295.t0 a_1597_329.t6 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 a_109_47.t1 SCD.t1 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1597_329.t1 a_1597_329.n4 778.22
R1 a_1597_329.n4 a_1597_329.t2 648.322
R2 a_1597_329.n0 a_1597_329.t0 473.219
R3 a_1597_329.n1 a_1597_329.t4 356.68
R4 a_1597_329.n2 a_1597_329.n1 291.342
R5 a_1597_329.n4 a_1597_329.n3 186.715
R6 a_1597_329.n2 a_1597_329.t6 144.601
R7 a_1597_329.n1 a_1597_329.t3 133.353
R8 a_1597_329.n0 a_1597_329.t5 132.282
R9 a_1597_329.n3 a_1597_329.n0 111.575
R10 a_1597_329.n3 a_1597_329.n2 32.1338
R11 a_2227_47.t1 a_2227_47.n2 392.002
R12 a_2227_47.n2 a_2227_47.t0 251.633
R13 a_2227_47.n0 a_2227_47.t2 212.081
R14 a_2227_47.n1 a_2227_47.t5 212.081
R15 a_2227_47.n2 a_2227_47.n1 186.215
R16 a_2227_47.n0 a_2227_47.t4 139.78
R17 a_2227_47.n1 a_2227_47.t3 139.78
R18 a_2227_47.n1 a_2227_47.n0 67.9187
R19 VPWR.n47 VPWR.t5 734.085
R20 VPWR.n24 VPWR.t1 688.083
R21 VPWR.n22 VPWR.t6 663.062
R22 VPWR.n54 VPWR.n1 602.067
R23 VPWR.n5 VPWR.n4 598.965
R24 VPWR.n10 VPWR.n9 585
R25 VPWR.n17 VPWR.n16 318.55
R26 VPWR.n18 VPWR.t9 256.387
R27 VPWR.n9 VPWR.t0 87.9469
R28 VPWR.n9 VPWR.t2 84.4291
R29 VPWR.n16 VPWR.t7 58.4849
R30 VPWR.n1 VPWR.t4 41.5552
R31 VPWR.n1 VPWR.t3 41.5552
R32 VPWR.n4 VPWR.t10 41.5552
R33 VPWR.n4 VPWR.t11 41.5552
R34 VPWR.n48 VPWR.n2 34.6358
R35 VPWR.n52 VPWR.n2 34.6358
R36 VPWR.n53 VPWR.n52 34.6358
R37 VPWR.n46 VPWR.n45 34.6358
R38 VPWR.n39 VPWR.n7 34.6358
R39 VPWR.n40 VPWR.n39 34.6358
R40 VPWR.n41 VPWR.n40 34.6358
R41 VPWR.n28 VPWR.n12 34.6358
R42 VPWR.n29 VPWR.n28 34.6358
R43 VPWR.n21 VPWR.n15 34.6358
R44 VPWR.n41 VPWR.n5 33.5064
R45 VPWR.n16 VPWR.t8 31.1381
R46 VPWR.n34 VPWR.n33 30.6829
R47 VPWR.n24 VPWR.n23 30.1181
R48 VPWR.n35 VPWR.n34 28.4986
R49 VPWR.n54 VPWR.n53 27.4829
R50 VPWR.n22 VPWR.n21 24.4711
R51 VPWR.n17 VPWR.n15 22.5887
R52 VPWR.n35 VPWR.n7 21.0829
R53 VPWR.n23 VPWR.n22 19.9534
R54 VPWR.n24 VPWR.n12 14.3064
R55 VPWR.n48 VPWR.n47 12.0476
R56 VPWR.n45 VPWR.n5 10.9181
R57 VPWR.n30 VPWR.n29 10.6358
R58 VPWR.n19 VPWR.n15 9.3005
R59 VPWR.n21 VPWR.n20 9.3005
R60 VPWR.n22 VPWR.n14 9.3005
R61 VPWR.n23 VPWR.n13 9.3005
R62 VPWR.n25 VPWR.n24 9.3005
R63 VPWR.n26 VPWR.n12 9.3005
R64 VPWR.n28 VPWR.n27 9.3005
R65 VPWR.n29 VPWR.n11 9.3005
R66 VPWR.n31 VPWR.n30 9.3005
R67 VPWR.n33 VPWR.n32 9.3005
R68 VPWR.n34 VPWR.n8 9.3005
R69 VPWR.n36 VPWR.n35 9.3005
R70 VPWR.n37 VPWR.n7 9.3005
R71 VPWR.n39 VPWR.n38 9.3005
R72 VPWR.n40 VPWR.n6 9.3005
R73 VPWR.n42 VPWR.n41 9.3005
R74 VPWR.n43 VPWR.n5 9.3005
R75 VPWR.n45 VPWR.n44 9.3005
R76 VPWR.n46 VPWR.n3 9.3005
R77 VPWR.n49 VPWR.n48 9.3005
R78 VPWR.n50 VPWR.n2 9.3005
R79 VPWR.n52 VPWR.n51 9.3005
R80 VPWR.n53 VPWR.n0 9.3005
R81 VPWR.n55 VPWR.n54 7.12063
R82 VPWR.n18 VPWR.n17 6.93035
R83 VPWR.n30 VPWR.n10 6.87109
R84 VPWR.n33 VPWR.n10 1.78874
R85 VPWR.n19 VPWR.n18 0.554139
R86 VPWR.n47 VPWR.n46 0.376971
R87 VPWR.n55 VPWR.n0 0.148519
R88 VPWR.n20 VPWR.n19 0.120292
R89 VPWR.n20 VPWR.n14 0.120292
R90 VPWR.n14 VPWR.n13 0.120292
R91 VPWR.n25 VPWR.n13 0.120292
R92 VPWR.n26 VPWR.n25 0.120292
R93 VPWR.n27 VPWR.n26 0.120292
R94 VPWR.n27 VPWR.n11 0.120292
R95 VPWR.n31 VPWR.n11 0.120292
R96 VPWR.n32 VPWR.n31 0.120292
R97 VPWR.n32 VPWR.n8 0.120292
R98 VPWR.n36 VPWR.n8 0.120292
R99 VPWR.n37 VPWR.n36 0.120292
R100 VPWR.n38 VPWR.n37 0.120292
R101 VPWR.n38 VPWR.n6 0.120292
R102 VPWR.n42 VPWR.n6 0.120292
R103 VPWR.n43 VPWR.n42 0.120292
R104 VPWR.n44 VPWR.n43 0.120292
R105 VPWR.n44 VPWR.n3 0.120292
R106 VPWR.n49 VPWR.n3 0.120292
R107 VPWR.n50 VPWR.n49 0.120292
R108 VPWR.n51 VPWR.n50 0.120292
R109 VPWR.n51 VPWR.n0 0.120292
R110 VPWR VPWR.n55 0.114842
R111 VPB.t4 VPB.t5 994.394
R112 VPB.t3 VPB.t6 970.716
R113 VPB.t10 VPB.t11 556.386
R114 VPB.t5 VPB.t10 556.386
R115 VPB.t14 VPB.t0 556.386
R116 VPB.t9 VPB.t15 556.386
R117 VPB.t16 VPB.t9 556.386
R118 VPB.t6 VPB.t2 343.303
R119 VPB.t11 VPB.t12 281.154
R120 VPB.t12 VPB.t13 275.235
R121 VPB.t0 VPB.t3 248.599
R122 VPB.t15 VPB.t14 248.599
R123 VPB.t1 VPB.t16 248.599
R124 VPB.t7 VPB.t8 248.599
R125 VPB.t2 VPB.t4 213.084
R126 VPB.t8 VPB.t1 213.084
R127 VPB VPB.t7 192.369
R128 Q.n1 Q 593.34
R129 Q.n1 Q.n0 585
R130 Q.n2 Q.n1 585
R131 Q.n5 Q 187.522
R132 Q.n6 Q.n5 185
R133 Q.n1 Q.t0 35.4605
R134 Q.n5 Q.t3 33.2313
R135 Q.n1 Q.t1 26.5955
R136 Q.n5 Q.t2 24.9236
R137 Q.n4 Q 16.2914
R138 Q.n6 Q 10.6672
R139 Q.n0 Q 8.33989
R140 Q.n3 Q.n2 6.4005
R141 Q.n0 Q 4.84898
R142 Q.n2 Q 4.84898
R143 Q.n4 Q 3.49141
R144 Q Q.n3 2.90959
R145 Q Q.n6 2.52171
R146 Q Q.n4 2.32777
R147 Q.n3 Q 1.93989
R148 VGND.n48 VGND.t5 250.499
R149 VGND.n19 VGND.t6 242.004
R150 VGND.n27 VGND.t0 224.153
R151 VGND.n54 VGND.t2 223.571
R152 VGND.n46 VGND.t4 223.571
R153 VGND.n14 VGND.n13 200.62
R154 VGND.n41 VGND.n40 198.964
R155 VGND.n12 VGND.t8 161.581
R156 VGND.n13 VGND.t7 54.2862
R157 VGND.n40 VGND.t1 38.5719
R158 VGND.n40 VGND.t3 38.5719
R159 VGND.n15 VGND.n11 34.6358
R160 VGND.n21 VGND.n20 34.6358
R161 VGND.n21 VGND.n9 34.6358
R162 VGND.n25 VGND.n9 34.6358
R163 VGND.n26 VGND.n25 34.6358
R164 VGND.n33 VGND.n32 34.6358
R165 VGND.n38 VGND.n5 34.6358
R166 VGND.n39 VGND.n38 34.6358
R167 VGND.n52 VGND.n1 34.6358
R168 VGND.n53 VGND.n52 34.0711
R169 VGND.n19 VGND.n11 33.5064
R170 VGND.n48 VGND.n47 33.1299
R171 VGND.n41 VGND.n39 31.2476
R172 VGND.n45 VGND.n3 28.5534
R173 VGND.n34 VGND.n5 27.3528
R174 VGND.n28 VGND.n26 27.0218
R175 VGND.n13 VGND.t9 25.9346
R176 VGND.n15 VGND.n14 22.5887
R177 VGND.n20 VGND.n19 16.9417
R178 VGND.n34 VGND.n33 16.6884
R179 VGND.n48 VGND.n1 16.1887
R180 VGND.n47 VGND.n46 15.2476
R181 VGND.n41 VGND.n3 13.177
R182 VGND.n55 VGND.n54 9.86521
R183 VGND.n16 VGND.n15 9.3005
R184 VGND.n17 VGND.n11 9.3005
R185 VGND.n19 VGND.n18 9.3005
R186 VGND.n20 VGND.n10 9.3005
R187 VGND.n22 VGND.n21 9.3005
R188 VGND.n23 VGND.n9 9.3005
R189 VGND.n25 VGND.n24 9.3005
R190 VGND.n26 VGND.n8 9.3005
R191 VGND.n29 VGND.n28 9.3005
R192 VGND.n30 VGND.n7 9.3005
R193 VGND.n32 VGND.n31 9.3005
R194 VGND.n33 VGND.n6 9.3005
R195 VGND.n35 VGND.n34 9.3005
R196 VGND.n36 VGND.n5 9.3005
R197 VGND.n38 VGND.n37 9.3005
R198 VGND.n39 VGND.n4 9.3005
R199 VGND.n42 VGND.n41 9.3005
R200 VGND.n43 VGND.n3 9.3005
R201 VGND.n45 VGND.n44 9.3005
R202 VGND.n47 VGND.n2 9.3005
R203 VGND.n49 VGND.n48 9.3005
R204 VGND.n50 VGND.n1 9.3005
R205 VGND.n52 VGND.n51 9.3005
R206 VGND.n53 VGND.n0 9.3005
R207 VGND.n32 VGND.n7 8.74815
R208 VGND.n54 VGND.n53 8.09462
R209 VGND.n14 VGND.n12 6.73566
R210 VGND.n28 VGND.n27 5.03421
R211 VGND.n46 VGND.n45 2.8005
R212 VGND.n27 VGND.n7 1.58252
R213 VGND.n16 VGND.n12 0.589728
R214 VGND.n17 VGND.n16 0.120292
R215 VGND.n18 VGND.n17 0.120292
R216 VGND.n18 VGND.n10 0.120292
R217 VGND.n22 VGND.n10 0.120292
R218 VGND.n23 VGND.n22 0.120292
R219 VGND.n24 VGND.n23 0.120292
R220 VGND.n24 VGND.n8 0.120292
R221 VGND.n29 VGND.n8 0.120292
R222 VGND.n30 VGND.n29 0.120292
R223 VGND.n31 VGND.n30 0.120292
R224 VGND.n31 VGND.n6 0.120292
R225 VGND.n35 VGND.n6 0.120292
R226 VGND.n36 VGND.n35 0.120292
R227 VGND.n37 VGND.n36 0.120292
R228 VGND.n37 VGND.n4 0.120292
R229 VGND.n42 VGND.n4 0.120292
R230 VGND.n43 VGND.n42 0.120292
R231 VGND.n44 VGND.n43 0.120292
R232 VGND.n44 VGND.n2 0.120292
R233 VGND.n49 VGND.n2 0.120292
R234 VGND.n50 VGND.n49 0.120292
R235 VGND.n51 VGND.n50 0.120292
R236 VGND.n51 VGND.n0 0.120292
R237 VGND.n55 VGND.n0 0.120292
R238 VGND VGND.n55 0.0226354
R239 VNB.t14 VNB.t1 6080.26
R240 VNB.t0 VNB.t10 5752.75
R241 VNB.t10 VNB.t11 3018.77
R242 VNB.t9 VNB.t8 2762.46
R243 VNB.t2 VNB.t3 2677.02
R244 VNB.t8 VNB.t5 2677.02
R245 VNB.t1 VNB.t0 2548.87
R246 VNB.t11 VNB.t13 1352.75
R247 VNB.t13 VNB.t12 1324.27
R248 VNB.t3 VNB.t14 1196.12
R249 VNB.t5 VNB.t2 1196.12
R250 VNB.t6 VNB.t9 1196.12
R251 VNB.t7 VNB.t6 1196.12
R252 VNB.t4 VNB.t7 1025.24
R253 VNB VNB.t4 925.567
R254 SET_B.n1 SET_B.n0 360.18
R255 SET_B.n3 SET_B.n2 357.216
R256 SET_B.n4 SET_B.n3 223.113
R257 SET_B.n1 SET_B.t1 166.577
R258 SET_B.n3 SET_B.t0 161.03
R259 SET_B.n4 SET_B.n1 159
R260 SET_B SET_B.n4 3.4005
R261 SCD.n0 SCD.t0 299.433
R262 SCD.n0 SCD.t1 206.245
R263 SCD.n1 SCD.n0 152
R264 SCD.n1 SCD 19.828
R265 SCD SCD.n1 14.3064
R266 a_27_369.t0 a_27_369.t1 1468.74
R267 a_643_369.t1 a_643_369.n6 670.312
R268 a_643_369.n4 a_643_369.t4 419.243
R269 a_643_369.n4 a_643_369.n3 413.587
R270 a_643_369.n0 a_643_369.t5 393.634
R271 a_643_369.n5 a_643_369.t2 317.574
R272 a_643_369.n2 a_643_369.t0 291.962
R273 a_643_369.n1 a_643_369.t6 267.3
R274 a_643_369.n2 a_643_369.n1 152
R275 a_643_369.n1 a_643_369.n0 100.206
R276 a_643_369.n0 a_643_369.t3 91.5805
R277 a_643_369.n5 a_643_369.n4 53.8068
R278 a_643_369.n6 a_643_369.n2 30.2774
R279 a_643_369.n6 a_643_369.n5 10.4313
R280 a_997_413.n7 a_997_413.n6 662.052
R281 a_997_413.n3 a_997_413.n1 312.132
R282 a_997_413.n0 a_997_413.t5 262.64
R283 a_997_413.n3 a_997_413.n2 238.226
R284 a_997_413.n6 a_997_413.n5 234.409
R285 a_997_413.n4 a_997_413.n0 200.561
R286 a_997_413.n0 a_997_413.t4 166.24
R287 a_997_413.n4 a_997_413.n3 152
R288 a_997_413.n7 a_997_413.t1 63.3219
R289 a_997_413.t0 a_997_413.n7 63.3219
R290 a_997_413.n6 a_997_413.n4 53.8358
R291 a_997_413.n5 a_997_413.t3 38.5719
R292 a_997_413.n5 a_997_413.t2 38.5719
R293 a_809_369.t0 a_809_369.n4 672.456
R294 a_809_369.n3 a_809_369.t4 433.509
R295 a_809_369.n1 a_809_369.t3 385.065
R296 a_809_369.n3 a_809_369.t2 321.334
R297 a_809_369.n2 a_809_369.t1 275.591
R298 a_809_369.n2 a_809_369.n1 205.534
R299 a_809_369.n4 a_809_369.n3 182.673
R300 a_809_369.n1 a_809_369.n0 148.35
R301 a_809_369.n4 a_809_369.n2 2.5605
R302 a_181_47.n1 a_181_47.t4 693.452
R303 a_181_47.n3 a_181_47.n2 613.688
R304 a_181_47.n2 a_181_47.n0 574.096
R305 a_181_47.n1 a_181_47.t3 288.805
R306 a_181_47.n3 a_181_47.t5 41.5552
R307 a_181_47.t0 a_181_47.n3 41.5552
R308 a_181_47.n0 a_181_47.t1 38.5719
R309 a_181_47.n0 a_181_47.t2 38.5719
R310 a_181_47.n2 a_181_47.n1 22.6251
R311 SCE.n1 SCE.t3 295.168
R312 SCE.n0 SCE.t2 263.18
R313 SCE.n0 SCE.t0 231.73
R314 SCE.n1 SCE.t1 201.982
R315 SCE.n2 SCE.n1 173.305
R316 SCE.n2 SCE.n0 154.744
R317 SCE SCE.n2 3.88621
R318 a_109_47.t0 a_109_47.t1 60.0005
R319 a_1514_47.t0 a_1514_47.t1 139.689
R320 a_1781_295.t0 a_1781_295.n3 697.798
R321 a_1781_295.n2 a_1781_295.n0 453.616
R322 a_1781_295.n3 a_1781_295.t1 302.202
R323 a_1781_295.n3 a_1781_295.n2 252.554
R324 a_1781_295.n2 a_1781_295.n1 161.202
R325 a_319_21.t0 a_319_21.n1 754.953
R326 a_319_21.n0 a_319_21.t2 283.286
R327 a_319_21.n1 a_319_21.t1 259.202
R328 a_319_21.n0 a_319_21.t3 190.101
R329 a_319_21.n1 a_319_21.n0 152
R330 D.n0 D.t0 373.283
R331 D.n1 D.n0 152
R332 D.n0 D.t1 132.282
R333 D.n1 D 23.1303
R334 D D.n1 7.41103
R335 a_193_369.t0 a_193_369.t1 64.6411
R336 a_1525_329.t0 a_1525_329.t1 49.2505
R337 a_265_47.t0 a_265_47.t1 77.1434
R338 CLK.n0 CLK.t0 255.077
R339 CLK.n0 CLK.t1 218.642
R340 CLK.n1 CLK.n0 152
R341 CLK.n1 CLK 19.0712
R342 CLK CLK.n1 2.90959
C0 Q VPB 0.006405f
C1 VPWR VPB 0.283079f
C2 SET_B a_1723_413# 2.84e-19
C3 a_1129_21# VPB 0.10089f
C4 SCE SCD 0.170177f
C5 D VPB 0.043648f
C6 Q VGND 0.146818f
C7 VPWR VGND 0.104607f
C8 a_1129_21# VGND 0.160635f
C9 D VGND 0.008596f
C10 SCE CLK 0.090396f
C11 a_1815_47# VPWR 1.13e-19
C12 SCE VPB 0.130585f
C13 SET_B VPB 0.19822f
C14 Q VPWR 0.176468f
C15 a_1129_21# VPWR 0.132033f
C16 D VPWR 0.007869f
C17 SCE VGND 0.142351f
C18 SET_B VGND 0.041467f
C19 VPB SCD 0.070898f
C20 SET_B a_1815_47# 4.89e-19
C21 VGND SCD 0.045223f
C22 CLK VPB 0.080439f
C23 SET_B Q 1.32e-19
C24 SCE VPWR 0.064479f
C25 CLK VGND 0.040331f
C26 SET_B VPWR 0.100556f
C27 SET_B a_1129_21# 0.030541f
C28 SCE D 0.20207f
C29 a_1887_47# VGND 0.001665f
C30 a_1723_413# VPWR 8.96e-19
C31 a_1723_413# a_1129_21# 7.11e-20
C32 VPWR SCD 0.017326f
C33 VGND VPB 0.01788f
C34 CLK VPWR 0.03f
C35 a_1347_47# VGND 0.004877f
C36 a_1815_47# VGND 0.001224f
C37 a_1887_47# VPWR 2.81e-19
C38 Q VNB 0.024645f
C39 VGND VNB 1.44867f
C40 VPWR VNB 1.16297f
C41 SET_B VNB 0.21886f
C42 CLK VNB 0.13687f
C43 D VNB 0.104133f
C44 SCE VNB 0.253779f
C45 SCD VNB 0.205442f
C46 VPB VNB 2.55388f
C47 a_1129_21# VNB 0.14521f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfstp_4 VPWR VGND VPB VNB Q SET_B CLK D SCD SCE
X0 VPWR.t11 a_2227_47.t2 Q.t5 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Q.t2 a_2227_47.t3 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X2 a_1597_329.t0 SET_B.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0966 ps=0.88 w=0.42 l=0.15
X3 Q.t4 a_2227_47.t4 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.32 w=1 l=0.15
X4 VPWR.t0 SCD.t0 a_27_369.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_1081_413.t0 a_643_369.t2 a_997_413.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0756 pd=0.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_809_369.t1 a_643_369.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND.t6 a_1597_329.t3 a_2227_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_997_413.t2 a_809_369.t2 a_181_47.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VPWR.t4 SET_B.t1 a_1129_21# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.27 as=0.0714 ps=0.76 w=0.42 l=0.15
X10 a_181_47.t0 SCE.t0 a_109_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 a_1514_47.t0 a_997_413.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.2384 pd=1.385 as=0.09575 ps=0.965 w=0.64 l=0.15
X12 Q.t1 a_2227_47.t5 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.104 ps=0.97 w=0.65 l=0.15
X13 VGND SET_B a_1347_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09575 pd=0.965 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 a_27_369.t1 a_319_21.t2 a_181_47.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 VGND.t3 SCE.t1 a_319_21.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 a_1597_329.t2 a_809_369.t3 a_1514_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1241 pd=1.1 as=0.2384 ps=1.385 w=0.64 l=0.15
X17 a_181_47.t5 D.t0 a_193_369.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X18 VGND SET_B a_1887_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 VGND.t8 a_2227_47.t6 Q.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_1597_329.t1 a_643_369.t4 a_1525_329.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.32 as=0.0882 ps=1.05 w=0.84 l=0.15
X21 a_265_47.t0 D.t1 a_181_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_997_413.t0 a_643_369.t5 a_181_47.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 Q.t3 a_2227_47.t7 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X24 a_1781_295.t1 a_1597_329.t4 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.0882 ps=0.84 w=0.42 l=0.15
X25 a_1087_47# a_809_369.t4 a_997_413.t3 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 a_193_369.t1 SCE.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_809_369.t0 a_643_369.t6 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_1525_329.t0 a_997_413.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.1428 ps=1.27 w=0.84 l=0.15
X29 VPWR.t8 SCE.t3 a_319_21.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.1664 ps=1.8 w=0.64 l=0.15
X30 VPWR.t6 a_1597_329.t5 a_2227_47.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X31 VPWR.t12 CLK.t0 a_643_369.t1 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X32 VGND.t5 a_319_21.t3 a_265_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0567 ps=0.69 w=0.42 l=0.15
X33 VGND a_1129_21# a_1087_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X34 VGND.t4 CLK.t1 a_643_369.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_1781_295.t0 a_1597_329.t6 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X36 a_109_47.t0 SCD.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_2227_47.t1 a_2227_47.n6 354.238
R1 a_2227_47.n6 a_2227_47.t0 237.986
R2 a_2227_47.n2 a_2227_47.t2 212.081
R3 a_2227_47.n3 a_2227_47.t4 212.081
R4 a_2227_47.n4 a_2227_47.n0 212.081
R5 a_2227_47.n5 a_2227_47.t7 212.081
R6 a_2227_47.n6 a_2227_47.n5 186.215
R7 a_2227_47.n2 a_2227_47.t6 139.78
R8 a_2227_47.n3 a_2227_47.t5 139.78
R9 a_2227_47.n4 a_2227_47.n1 139.78
R10 a_2227_47.n5 a_2227_47.t3 139.78
R11 a_2227_47.n4 a_2227_47.n3 68.649
R12 a_2227_47.n3 a_2227_47.n2 61.346
R13 a_2227_47.n5 a_2227_47.n4 61.346
R14 Q Q.t3 810.096
R15 Q.n4 Q.n2 220.989
R16 Q.n0 Q.t2 209.923
R17 Q.n4 Q.n3 114.692
R18 Q.n2 Q.t5 26.5955
R19 Q.n2 Q.t4 26.5955
R20 Q.n3 Q.t0 24.9236
R21 Q.n3 Q.t1 24.9236
R22 Q.n5 Q 19.2005
R23 Q.n5 Q.n1 13.0849
R24 Q Q.n0 12.6066
R25 Q.n6 Q 11.249
R26 Q Q.n4 10.4301
R27 Q Q.n5 6.82717
R28 Q.n1 Q 3.41383
R29 Q.n6 Q 2.84494
R30 Q.n5 Q 2.60791
R31 Q.n1 Q 2.32777
R32 Q Q.n6 1.93989
R33 Q.n0 Q 0.582318
R34 VPWR.n51 VPWR.t8 734.085
R35 VPWR.n28 VPWR.t3 688.083
R36 VPWR.n26 VPWR.t7 663.062
R37 VPWR.n58 VPWR.n1 602.067
R38 VPWR.n5 VPWR.n4 598.965
R39 VPWR.n10 VPWR.n9 585
R40 VPWR.n19 VPWR.t10 257.474
R41 VPWR.n18 VPWR.t11 249.917
R42 VPWR.n21 VPWR.n17 214.662
R43 VPWR.n9 VPWR.t1 87.9469
R44 VPWR.n9 VPWR.t4 84.4291
R45 VPWR.n1 VPWR.t2 41.5552
R46 VPWR.n1 VPWR.t0 41.5552
R47 VPWR.n4 VPWR.t5 41.5552
R48 VPWR.n4 VPWR.t12 41.5552
R49 VPWR.n52 VPWR.n2 34.6358
R50 VPWR.n56 VPWR.n2 34.6358
R51 VPWR.n57 VPWR.n56 34.6358
R52 VPWR.n50 VPWR.n49 34.6358
R53 VPWR.n43 VPWR.n7 34.6358
R54 VPWR.n44 VPWR.n43 34.6358
R55 VPWR.n45 VPWR.n44 34.6358
R56 VPWR.n32 VPWR.n12 34.6358
R57 VPWR.n33 VPWR.n32 34.6358
R58 VPWR.n25 VPWR.n15 34.6358
R59 VPWR.n45 VPWR.n5 33.5064
R60 VPWR.n20 VPWR.n19 32.7534
R61 VPWR.n17 VPWR.t9 32.5055
R62 VPWR.n17 VPWR.t6 31.5205
R63 VPWR.n38 VPWR.n37 30.6829
R64 VPWR.n28 VPWR.n27 30.1181
R65 VPWR.n39 VPWR.n38 28.4986
R66 VPWR.n58 VPWR.n57 27.4829
R67 VPWR.n26 VPWR.n25 24.4711
R68 VPWR.n21 VPWR.n20 24.0946
R69 VPWR.n39 VPWR.n7 21.0829
R70 VPWR.n27 VPWR.n26 19.9534
R71 VPWR.n21 VPWR.n15 18.4476
R72 VPWR.n28 VPWR.n12 14.3064
R73 VPWR.n52 VPWR.n51 12.0476
R74 VPWR.n49 VPWR.n5 10.9181
R75 VPWR.n34 VPWR.n33 10.6358
R76 VPWR.n20 VPWR.n16 9.3005
R77 VPWR.n22 VPWR.n21 9.3005
R78 VPWR.n23 VPWR.n15 9.3005
R79 VPWR.n25 VPWR.n24 9.3005
R80 VPWR.n26 VPWR.n14 9.3005
R81 VPWR.n27 VPWR.n13 9.3005
R82 VPWR.n29 VPWR.n28 9.3005
R83 VPWR.n30 VPWR.n12 9.3005
R84 VPWR.n32 VPWR.n31 9.3005
R85 VPWR.n33 VPWR.n11 9.3005
R86 VPWR.n35 VPWR.n34 9.3005
R87 VPWR.n37 VPWR.n36 9.3005
R88 VPWR.n38 VPWR.n8 9.3005
R89 VPWR.n40 VPWR.n39 9.3005
R90 VPWR.n41 VPWR.n7 9.3005
R91 VPWR.n43 VPWR.n42 9.3005
R92 VPWR.n44 VPWR.n6 9.3005
R93 VPWR.n46 VPWR.n45 9.3005
R94 VPWR.n47 VPWR.n5 9.3005
R95 VPWR.n49 VPWR.n48 9.3005
R96 VPWR.n50 VPWR.n3 9.3005
R97 VPWR.n53 VPWR.n52 9.3005
R98 VPWR.n54 VPWR.n2 9.3005
R99 VPWR.n56 VPWR.n55 9.3005
R100 VPWR.n57 VPWR.n0 9.3005
R101 VPWR.n19 VPWR.n18 9.06231
R102 VPWR.n59 VPWR.n58 7.12063
R103 VPWR.n34 VPWR.n10 6.87109
R104 VPWR.n37 VPWR.n10 1.78874
R105 VPWR.n18 VPWR.n16 0.550633
R106 VPWR.n51 VPWR.n50 0.376971
R107 VPWR.n59 VPWR.n0 0.148519
R108 VPWR.n22 VPWR.n16 0.120292
R109 VPWR.n23 VPWR.n22 0.120292
R110 VPWR.n24 VPWR.n23 0.120292
R111 VPWR.n24 VPWR.n14 0.120292
R112 VPWR.n14 VPWR.n13 0.120292
R113 VPWR.n29 VPWR.n13 0.120292
R114 VPWR.n30 VPWR.n29 0.120292
R115 VPWR.n31 VPWR.n30 0.120292
R116 VPWR.n31 VPWR.n11 0.120292
R117 VPWR.n35 VPWR.n11 0.120292
R118 VPWR.n36 VPWR.n35 0.120292
R119 VPWR.n36 VPWR.n8 0.120292
R120 VPWR.n40 VPWR.n8 0.120292
R121 VPWR.n41 VPWR.n40 0.120292
R122 VPWR.n42 VPWR.n41 0.120292
R123 VPWR.n42 VPWR.n6 0.120292
R124 VPWR.n46 VPWR.n6 0.120292
R125 VPWR.n47 VPWR.n46 0.120292
R126 VPWR.n48 VPWR.n47 0.120292
R127 VPWR.n48 VPWR.n3 0.120292
R128 VPWR.n53 VPWR.n3 0.120292
R129 VPWR.n54 VPWR.n53 0.120292
R130 VPWR.n55 VPWR.n54 0.120292
R131 VPWR.n55 VPWR.n0 0.120292
R132 VPWR VPWR.n59 0.114842
R133 VPB.t6 VPB.t4 994.394
R134 VPB.t2 VPB.t5 970.716
R135 VPB.t9 VPB.t8 556.386
R136 VPB.t4 VPB.t9 556.386
R137 VPB.t7 VPB.t11 556.386
R138 VPB.t10 VPB.t17 556.386
R139 VPB.t12 VPB.t10 556.386
R140 VPB.t14 VPB.t15 526.792
R141 VPB.t5 VPB.t1 343.303
R142 VPB.t8 VPB.t14 281.154
R143 VPB.t15 VPB.t16 248.599
R144 VPB.t11 VPB.t2 248.599
R145 VPB.t17 VPB.t7 248.599
R146 VPB.t13 VPB.t12 248.599
R147 VPB.t0 VPB.t3 248.599
R148 VPB.t1 VPB.t6 213.084
R149 VPB.t3 VPB.t13 213.084
R150 VPB VPB.t0 192.369
R151 VGND.n52 VGND.t5 250.499
R152 VGND.n23 VGND.t7 242.004
R153 VGND.n31 VGND.t1 224.153
R154 VGND.n58 VGND.t0 223.571
R155 VGND.n50 VGND.t3 223.571
R156 VGND.n45 VGND.n44 198.964
R157 VGND.n14 VGND.t8 156.222
R158 VGND.n13 VGND.t9 152.832
R159 VGND.n18 VGND.n17 108.448
R160 VGND.n44 VGND.t2 38.5719
R161 VGND.n44 VGND.t4 38.5719
R162 VGND.n19 VGND.n11 34.6358
R163 VGND.n25 VGND.n24 34.6358
R164 VGND.n25 VGND.n9 34.6358
R165 VGND.n29 VGND.n9 34.6358
R166 VGND.n30 VGND.n29 34.6358
R167 VGND.n37 VGND.n36 34.6358
R168 VGND.n42 VGND.n5 34.6358
R169 VGND.n43 VGND.n42 34.6358
R170 VGND.n56 VGND.n1 34.6358
R171 VGND.n57 VGND.n56 34.0711
R172 VGND.n23 VGND.n11 33.5064
R173 VGND.n52 VGND.n51 33.1299
R174 VGND.n16 VGND.n13 32.7534
R175 VGND.n45 VGND.n43 31.2476
R176 VGND.n17 VGND.t10 30.462
R177 VGND.n17 VGND.t6 29.539
R178 VGND.n49 VGND.n3 28.5534
R179 VGND.n38 VGND.n5 27.3528
R180 VGND.n32 VGND.n30 27.0218
R181 VGND.n18 VGND.n16 24.0946
R182 VGND.n19 VGND.n18 18.4476
R183 VGND.n24 VGND.n23 16.9417
R184 VGND.n38 VGND.n37 16.6884
R185 VGND.n52 VGND.n1 16.1887
R186 VGND.n51 VGND.n50 15.2476
R187 VGND.n45 VGND.n3 13.177
R188 VGND.n59 VGND.n58 9.86521
R189 VGND.n16 VGND.n15 9.3005
R190 VGND.n18 VGND.n12 9.3005
R191 VGND.n20 VGND.n19 9.3005
R192 VGND.n21 VGND.n11 9.3005
R193 VGND.n23 VGND.n22 9.3005
R194 VGND.n24 VGND.n10 9.3005
R195 VGND.n26 VGND.n25 9.3005
R196 VGND.n27 VGND.n9 9.3005
R197 VGND.n29 VGND.n28 9.3005
R198 VGND.n30 VGND.n8 9.3005
R199 VGND.n33 VGND.n32 9.3005
R200 VGND.n34 VGND.n7 9.3005
R201 VGND.n36 VGND.n35 9.3005
R202 VGND.n37 VGND.n6 9.3005
R203 VGND.n39 VGND.n38 9.3005
R204 VGND.n40 VGND.n5 9.3005
R205 VGND.n42 VGND.n41 9.3005
R206 VGND.n43 VGND.n4 9.3005
R207 VGND.n46 VGND.n45 9.3005
R208 VGND.n47 VGND.n3 9.3005
R209 VGND.n49 VGND.n48 9.3005
R210 VGND.n51 VGND.n2 9.3005
R211 VGND.n53 VGND.n52 9.3005
R212 VGND.n54 VGND.n1 9.3005
R213 VGND.n56 VGND.n55 9.3005
R214 VGND.n57 VGND.n0 9.3005
R215 VGND.n14 VGND.n13 9.06231
R216 VGND.n36 VGND.n7 8.74815
R217 VGND.n58 VGND.n57 8.09462
R218 VGND.n32 VGND.n31 5.03421
R219 VGND.n50 VGND.n49 2.8005
R220 VGND.n31 VGND.n7 1.58252
R221 VGND.n15 VGND.n14 0.550633
R222 VGND.n15 VGND.n12 0.120292
R223 VGND.n20 VGND.n12 0.120292
R224 VGND.n21 VGND.n20 0.120292
R225 VGND.n22 VGND.n21 0.120292
R226 VGND.n22 VGND.n10 0.120292
R227 VGND.n26 VGND.n10 0.120292
R228 VGND.n27 VGND.n26 0.120292
R229 VGND.n28 VGND.n27 0.120292
R230 VGND.n28 VGND.n8 0.120292
R231 VGND.n33 VGND.n8 0.120292
R232 VGND.n34 VGND.n33 0.120292
R233 VGND.n35 VGND.n34 0.120292
R234 VGND.n35 VGND.n6 0.120292
R235 VGND.n39 VGND.n6 0.120292
R236 VGND.n40 VGND.n39 0.120292
R237 VGND.n41 VGND.n40 0.120292
R238 VGND.n41 VGND.n4 0.120292
R239 VGND.n46 VGND.n4 0.120292
R240 VGND.n47 VGND.n46 0.120292
R241 VGND.n48 VGND.n47 0.120292
R242 VGND.n48 VGND.n2 0.120292
R243 VGND.n53 VGND.n2 0.120292
R244 VGND.n54 VGND.n53 0.120292
R245 VGND.n55 VGND.n54 0.120292
R246 VGND.n55 VGND.n0 0.120292
R247 VGND.n59 VGND.n0 0.120292
R248 VGND VGND.n59 0.0226354
R249 VNB.t15 VNB.t2 6080.26
R250 VNB.t11 VNB.t10 5752.75
R251 VNB.t10 VNB.t9 3018.77
R252 VNB.t7 VNB.t4 2762.46
R253 VNB.t3 VNB.t8 2677.02
R254 VNB.t4 VNB.t6 2677.02
R255 VNB.t2 VNB.t11 2548.87
R256 VNB.t14 VNB.t13 2534.63
R257 VNB.t9 VNB.t14 1352.75
R258 VNB.t13 VNB.t12 1196.12
R259 VNB.t8 VNB.t15 1196.12
R260 VNB.t6 VNB.t3 1196.12
R261 VNB.t5 VNB.t7 1196.12
R262 VNB.t0 VNB.t5 1196.12
R263 VNB.t1 VNB.t0 1025.24
R264 VNB VNB.t1 925.567
R265 SET_B.n1 SET_B.n0 360.18
R266 SET_B.n3 SET_B.n2 357.216
R267 SET_B.n4 SET_B.n3 223.113
R268 SET_B.n1 SET_B.t1 166.577
R269 SET_B.n3 SET_B.t0 161.03
R270 SET_B.n4 SET_B.n1 159
R271 SET_B SET_B.n4 3.4005
R272 a_1597_329.t1 a_1597_329.n4 778.22
R273 a_1597_329.n4 a_1597_329.t0 648.322
R274 a_1597_329.n1 a_1597_329.t2 473.219
R275 a_1597_329.n2 a_1597_329.n0 277.954
R276 a_1597_329.n0 a_1597_329.t3 207.261
R277 a_1597_329.n0 a_1597_329.t5 202.44
R278 a_1597_329.n4 a_1597_329.n3 181.361
R279 a_1597_329.n3 a_1597_329.t6 161.286
R280 a_1597_329.n1 a_1597_329.t4 132.282
R281 a_1597_329.n2 a_1597_329.n1 58.3623
R282 a_1597_329.n3 a_1597_329.n2 50.6723
R283 SCD.n0 SCD.t0 299.433
R284 SCD.n0 SCD.t1 206.245
R285 SCD.n1 SCD.n0 152
R286 SCD SCD.n1 19.828
R287 SCD.n1 SCD 14.3064
R288 a_27_369.t0 a_27_369.t1 1468.74
R289 a_643_369.t1 a_643_369.n6 670.312
R290 a_643_369.n4 a_643_369.t4 419.243
R291 a_643_369.n4 a_643_369.n3 413.587
R292 a_643_369.n0 a_643_369.t5 393.634
R293 a_643_369.n5 a_643_369.t2 317.574
R294 a_643_369.n2 a_643_369.t0 291.962
R295 a_643_369.n1 a_643_369.t6 267.3
R296 a_643_369.n2 a_643_369.n1 152
R297 a_643_369.n1 a_643_369.n0 100.206
R298 a_643_369.n0 a_643_369.t3 91.5805
R299 a_643_369.n5 a_643_369.n4 53.8068
R300 a_643_369.n6 a_643_369.n2 30.2774
R301 a_643_369.n6 a_643_369.n5 10.4313
R302 a_997_413.n6 a_997_413.n0 662.052
R303 a_997_413.n4 a_997_413.n2 312.132
R304 a_997_413.n1 a_997_413.t5 262.64
R305 a_997_413.n4 a_997_413.n3 238.226
R306 a_997_413.n7 a_997_413.n6 234.409
R307 a_997_413.n5 a_997_413.n1 200.561
R308 a_997_413.n1 a_997_413.t4 166.24
R309 a_997_413.n5 a_997_413.n4 152
R310 a_997_413.n0 a_997_413.t1 63.3219
R311 a_997_413.n0 a_997_413.t2 63.3219
R312 a_997_413.n6 a_997_413.n5 53.8358
R313 a_997_413.n7 a_997_413.t3 38.5719
R314 a_997_413.t0 a_997_413.n7 38.5719
R315 a_809_369.t0 a_809_369.n4 672.456
R316 a_809_369.n3 a_809_369.t4 433.509
R317 a_809_369.n1 a_809_369.t3 385.065
R318 a_809_369.n3 a_809_369.t2 321.334
R319 a_809_369.n2 a_809_369.t1 275.591
R320 a_809_369.n2 a_809_369.n1 205.534
R321 a_809_369.n4 a_809_369.n3 182.673
R322 a_809_369.n1 a_809_369.n0 148.35
R323 a_809_369.n4 a_809_369.n2 2.5605
R324 a_181_47.n1 a_181_47.t3 693.452
R325 a_181_47.n3 a_181_47.n2 613.688
R326 a_181_47.n2 a_181_47.n0 574.096
R327 a_181_47.n1 a_181_47.t2 288.805
R328 a_181_47.t4 a_181_47.n3 41.5552
R329 a_181_47.n3 a_181_47.t5 41.5552
R330 a_181_47.n0 a_181_47.t1 38.5719
R331 a_181_47.n0 a_181_47.t0 38.5719
R332 a_181_47.n2 a_181_47.n1 22.6251
R333 SCE.n1 SCE.t3 295.168
R334 SCE.n0 SCE.t2 263.18
R335 SCE.n0 SCE.t0 231.73
R336 SCE.n1 SCE.t1 201.982
R337 SCE.n2 SCE.n1 173.305
R338 SCE.n2 SCE.n0 154.744
R339 SCE SCE.n2 3.88621
R340 a_109_47.t0 a_109_47.t1 60.0005
R341 a_1514_47.t0 a_1514_47.t1 139.689
R342 a_1781_295.t0 a_1781_295.n3 697.798
R343 a_1781_295.n2 a_1781_295.n0 453.616
R344 a_1781_295.n3 a_1781_295.t1 302.202
R345 a_1781_295.n3 a_1781_295.n2 252.554
R346 a_1781_295.n2 a_1781_295.n1 161.202
R347 a_319_21.t0 a_319_21.n1 754.953
R348 a_319_21.n0 a_319_21.t2 283.286
R349 a_319_21.n1 a_319_21.t1 259.202
R350 a_319_21.n0 a_319_21.t3 190.101
R351 a_319_21.n1 a_319_21.n0 152
R352 D.n0 D.t0 373.283
R353 D.n1 D.n0 152
R354 D.n0 D.t1 132.282
R355 D D.n1 23.1303
R356 D.n1 D 7.41103
R357 a_193_369.t0 a_193_369.t1 64.6411
R358 a_1525_329.t0 a_1525_329.t1 49.2505
R359 a_265_47.t0 a_265_47.t1 77.1434
R360 CLK.n0 CLK.t0 255.077
R361 CLK.n0 CLK.t1 218.642
R362 CLK.n1 CLK.n0 152
R363 CLK.n1 CLK 19.0712
R364 CLK CLK.n1 2.90959
C0 SET_B a_1129_21# 0.030541f
C1 VPWR SCD 0.017326f
C2 VPWR VPB 0.301274f
C3 a_1087_47# a_1129_21# 7.75e-19
C4 VPWR Q 0.440815f
C5 SET_B a_1815_47# 4.89e-19
C6 D VPB 0.043648f
C7 CLK VGND 0.040331f
C8 SCD SCE 0.170177f
C9 a_1129_21# VPB 0.10089f
C10 VPB SCE 0.130585f
C11 SET_B VPB 0.198032f
C12 SET_B Q 2.18e-19
C13 VPWR VGND 0.127528f
C14 VPWR CLK 0.03f
C15 D VGND 0.008596f
C16 a_1887_47# VGND 0.001665f
C17 VPB SCD 0.070898f
C18 a_1129_21# VGND 0.160635f
C19 a_1347_47# VGND 0.004877f
C20 VGND SCE 0.142351f
C21 SET_B VGND 0.041467f
C22 Q VPB 0.011192f
C23 CLK SCE 0.090396f
C24 VPWR D 0.007869f
C25 VPWR a_1887_47# 2.81e-19
C26 VPWR a_1723_413# 8.96e-19
C27 a_1815_47# VGND 0.001224f
C28 a_1087_47# VGND 0.005211f
C29 VPWR a_1129_21# 0.132033f
C30 VPWR SCE 0.064479f
C31 SET_B VPWR 0.100614f
C32 VGND SCD 0.045223f
C33 a_1723_413# a_1129_21# 7.11e-20
C34 VGND VPB 0.018556f
C35 D SCE 0.20207f
C36 VGND Q 0.322044f
C37 VPWR a_1815_47# 1.13e-19
C38 SET_B a_1723_413# 2.84e-19
C39 CLK VPB 0.080439f
C40 Q VNB 0.028198f
C41 VGND VNB 1.5421f
C42 VPWR VNB 1.23728f
C43 SET_B VNB 0.218391f
C44 CLK VNB 0.13687f
C45 D VNB 0.104133f
C46 SCE VNB 0.253779f
C47 SCD VNB 0.205442f
C48 VPB VNB 2.73107f
C49 a_1129_21# VNB 0.14521f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxbp_1 VGND VPWR VNB VPB Q Q_N SCD SCE D CLK
X0 a_640_369.t1 a_299_47.t2 a_556_369.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1008 pd=0.955 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_1346_413.t1 a_193_47.t2 a_1089_183# VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR.t4 SCE.t0 a_299_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_556_369.t4 D.t0 a_465_369.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X4 a_1430_413.t0 a_193_47.t3 a_1346_413.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 Q.t0 a_1517_315.t2 VGND.t6 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Q_N.t0 a_1948_47.t2 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X7 VPWR.t6 CLK.t0 a_27_47.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_1346_413.t0 a_27_47.t2 a_1089_183# VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9 a_657_47.t0 SCE.t1 a_556_369.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND.t9 a_1346_413.t3 a_1517_315.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_930_413.t2 a_27_47.t3 a_556_369.t2 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1008 ps=1.28 w=0.36 l=0.15
X12 VPWR.t2 SCD.t0 a_640_369.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1824 pd=1.85 as=0.1008 ps=0.955 w=0.64 l=0.15
X13 a_193_47.t0 a_27_47.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_483_47.t0 a_299_47.t3 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X15 VGND.t1 a_1089_183# a_1027_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X16 a_930_413.t1 a_193_47.t4 a_556_369.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 Q_N.t1 a_1948_47.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X18 VGND.t4 a_1517_315.t3 a_1475_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X19 Q.t1 a_1517_315.t4 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t8 a_1346_413.t4 a_1517_315.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 a_193_47.t1 a_27_47.t5 VPWR.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1023_413# a_27_47.t6 a_930_413.t3 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X23 VGND.t5 a_1517_315.t5 a_1948_47.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VGND.t7 SCE.t2 a_299_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 VGND.t10 SCD.t1 a_657_47.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0483 ps=0.65 w=0.42 l=0.15
X26 a_1027_47.t1 a_193_47.t5 a_930_413.t0 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 VPWR a_1089_183# a_1023_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 VPWR.t7 a_1517_315.t6 a_1948_47.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 a_465_369.t0 SCE.t3 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 VGND.t3 CLK.t1 a_27_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_556_369.t5 D.t1 a_483_47.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_299_47.t0 a_299_47.n1 635.986
R1 a_299_47.n0 a_299_47.t2 416.856
R2 a_299_47.n0 a_299_47.t3 382.026
R3 a_299_47.n1 a_299_47.t1 331.699
R4 a_299_47.n1 a_299_47.n0 28.5772
R5 a_556_369.n3 a_556_369.n2 704.341
R6 a_556_369.n2 a_556_369.t1 663.176
R7 a_556_369.n1 a_556_369.n0 299.825
R8 a_556_369.n1 a_556_369.t2 257.75
R9 a_556_369.n2 a_556_369.n1 70.777
R10 a_556_369.n0 a_556_369.t5 54.2862
R11 a_556_369.t3 a_556_369.n3 41.5552
R12 a_556_369.n3 a_556_369.t4 41.5552
R13 a_556_369.n0 a_556_369.t0 40.0005
R14 a_640_369.t0 a_640_369.t1 96.9614
R15 VPB.t6 VPB.t0 970.716
R16 VPB.t14 VPB.t3 955.919
R17 VPB.t5 VPB.t7 583.023
R18 VPB.t1 VPB.t13 556.386
R19 VPB.t9 VPB.t4 556.386
R20 VPB.t13 VPB.t2 287.072
R21 VPB.t7 VPB.t14 275.235
R22 VPB.t10 VPB.t5 275.235
R23 VPB.t8 VPB.t11 269.315
R24 VPB.t0 VPB.t1 248.599
R25 VPB.t3 VPB.t6 248.599
R26 VPB.t11 VPB.t10 248.599
R27 VPB.t4 VPB.t8 248.599
R28 VPB.t12 VPB.t9 248.599
R29 VPB VPB.t12 142.056
R30 a_193_47.t1 a_193_47.n3 446.825
R31 a_193_47.n0 a_193_47.t3 348.661
R32 a_193_47.n1 a_193_47.t4 345.803
R33 a_193_47.n1 a_193_47.t5 281.236
R34 a_193_47.n0 a_193_47.t2 271.262
R35 a_193_47.n3 a_193_47.t0 249.172
R36 a_193_47.n2 a_193_47.n0 18.9875
R37 a_193_47.n3 a_193_47.n2 12.5295
R38 a_193_47.n2 a_193_47.n1 9.3005
R39 a_1346_413.n2 a_1346_413.n1 693.449
R40 a_1346_413.n1 a_1346_413.t1 317.325
R41 a_1346_413.n1 a_1346_413.n0 253.677
R42 a_1346_413.n0 a_1346_413.t4 212.081
R43 a_1346_413.n0 a_1346_413.t3 139.78
R44 a_1346_413.n2 a_1346_413.t2 63.3219
R45 a_1346_413.t0 a_1346_413.n2 63.3219
R46 VNB.t1 VNB.t7 3517.15
R47 VNB.t7 VNB.t3 2819.42
R48 VNB.t15 VNB.t10 2819.42
R49 VNB.t2 VNB.t13 2677.02
R50 VNB.t3 VNB.t14 2677.02
R51 VNB.t0 VNB.t9 2677.02
R52 VNB.t9 VNB.t11 1452.43
R53 VNB.t6 VNB.t1 1395.47
R54 VNB.t13 VNB.t4 1381.23
R55 VNB.t10 VNB.t6 1366.99
R56 VNB.t12 VNB.t8 1366.99
R57 VNB.t14 VNB.t2 1196.12
R58 VNB.t5 VNB.t0 1196.12
R59 VNB.t11 VNB.t12 1110.68
R60 VNB.t8 VNB.t15 1082.2
R61 VNB VNB.t5 683.495
R62 SCE.n2 SCE.t1 342.286
R63 SCE.n1 SCE.t2 321.772
R64 SCE.n2 SCE.n1 305.351
R65 SCE.n0 SCE.t3 241
R66 SCE.n0 SCE.t0 174.835
R67 SCE SCE.n2 20.1148
R68 SCE.n1 SCE.n0 8.76414
R69 VPWR.n5 VPWR.t2 722.018
R70 VPWR.n41 VPWR.n1 604.394
R71 VPWR.n3 VPWR.n2 600.128
R72 VPWR.n12 VPWR.n11 333.348
R73 VPWR.n14 VPWR.n13 237.108
R74 VPWR.n13 VPWR.t7 61.9924
R75 VPWR.n1 VPWR.t3 41.5552
R76 VPWR.n1 VPWR.t6 41.5552
R77 VPWR.n2 VPWR.t5 41.5552
R78 VPWR.n2 VPWR.t4 41.5552
R79 VPWR.n40 VPWR.n39 34.6358
R80 VPWR.n18 VPWR.n9 34.6358
R81 VPWR.n22 VPWR.n9 34.6358
R82 VPWR.n23 VPWR.n22 34.6358
R83 VPWR.n24 VPWR.n23 34.6358
R84 VPWR.n24 VPWR.n7 34.6358
R85 VPWR.n28 VPWR.n7 34.6358
R86 VPWR.n29 VPWR.n28 34.6358
R87 VPWR.n30 VPWR.n29 34.6358
R88 VPWR.n34 VPWR.n33 34.6358
R89 VPWR.n35 VPWR.n34 34.6358
R90 VPWR.n17 VPWR.n16 33.1299
R91 VPWR.n16 VPWR.n12 31.2476
R92 VPWR.n13 VPWR.t1 30.164
R93 VPWR.n33 VPWR.n5 28.2358
R94 VPWR.n11 VPWR.t0 26.5955
R95 VPWR.n11 VPWR.t8 26.5955
R96 VPWR.n35 VPWR.n3 24.4711
R97 VPWR.n41 VPWR.n40 22.9652
R98 VPWR.n39 VPWR.n3 19.9534
R99 VPWR.n18 VPWR.n17 13.177
R100 VPWR.n14 VPWR.n12 10.9351
R101 VPWR.n16 VPWR.n15 9.3005
R102 VPWR.n17 VPWR.n10 9.3005
R103 VPWR.n19 VPWR.n18 9.3005
R104 VPWR.n20 VPWR.n9 9.3005
R105 VPWR.n22 VPWR.n21 9.3005
R106 VPWR.n23 VPWR.n8 9.3005
R107 VPWR.n25 VPWR.n24 9.3005
R108 VPWR.n26 VPWR.n7 9.3005
R109 VPWR.n28 VPWR.n27 9.3005
R110 VPWR.n29 VPWR.n6 9.3005
R111 VPWR.n31 VPWR.n30 9.3005
R112 VPWR.n33 VPWR.n32 9.3005
R113 VPWR.n34 VPWR.n4 9.3005
R114 VPWR.n36 VPWR.n35 9.3005
R115 VPWR.n37 VPWR.n3 9.3005
R116 VPWR.n39 VPWR.n38 9.3005
R117 VPWR.n40 VPWR.n0 9.3005
R118 VPWR.n42 VPWR.n41 7.12063
R119 VPWR.n30 VPWR.n5 6.4005
R120 VPWR.n15 VPWR.n14 0.200927
R121 VPWR.n42 VPWR.n0 0.148519
R122 VPWR.n15 VPWR.n10 0.120292
R123 VPWR.n19 VPWR.n10 0.120292
R124 VPWR.n20 VPWR.n19 0.120292
R125 VPWR.n21 VPWR.n20 0.120292
R126 VPWR.n21 VPWR.n8 0.120292
R127 VPWR.n25 VPWR.n8 0.120292
R128 VPWR.n26 VPWR.n25 0.120292
R129 VPWR.n27 VPWR.n26 0.120292
R130 VPWR.n27 VPWR.n6 0.120292
R131 VPWR.n31 VPWR.n6 0.120292
R132 VPWR.n32 VPWR.n31 0.120292
R133 VPWR.n32 VPWR.n4 0.120292
R134 VPWR.n36 VPWR.n4 0.120292
R135 VPWR.n37 VPWR.n36 0.120292
R136 VPWR.n38 VPWR.n37 0.120292
R137 VPWR.n38 VPWR.n0 0.120292
R138 VPWR VPWR.n42 0.114842
R139 D.n0 D.t1 321.87
R140 D.n0 D.t0 183.696
R141 D D.n0 161.504
R142 a_465_369.t0 a_465_369.t1 93.8833
R143 a_930_413.n5 a_930_413.n4 693.048
R144 a_930_413.n4 a_930_413.n3 300.243
R145 a_930_413.n2 a_930_413.n1 226.541
R146 a_930_413.n2 a_930_413.n0 196.013
R147 a_930_413.n4 a_930_413.n2 168.738
R148 a_930_413.t1 a_930_413.n5 75.0481
R149 a_930_413.n5 a_930_413.t3 72.7029
R150 a_930_413.n3 a_930_413.t2 65.0005
R151 a_930_413.n3 a_930_413.t0 45.0005
R152 a_1517_315.n4 a_1517_315.t3 383.5
R153 a_1517_315.t1 a_1517_315.n5 324.786
R154 a_1517_315.n0 a_1517_315.t6 256.988
R155 a_1517_315.n1 a_1517_315.t4 212.081
R156 a_1517_315.n5 a_1517_315.n4 178.571
R157 a_1517_315.n2 a_1517_315.n1 173.721
R158 a_1517_315.n0 a_1517_315.t5 163.803
R159 a_1517_315.n2 a_1517_315.t0 150.524
R160 a_1517_315.n1 a_1517_315.t2 139.78
R161 a_1517_315.n4 a_1517_315.n3 139.286
R162 a_1517_315.n1 a_1517_315.n0 129.264
R163 a_1517_315.n5 a_1517_315.n2 19.2372
R164 VGND.n6 VGND.t1 286.673
R165 VGND.n4 VGND.t10 256.464
R166 VGND.n15 VGND.t4 239.139
R167 VGND.n13 VGND.n10 218.506
R168 VGND.n40 VGND.n39 199.739
R169 VGND.n2 VGND.n1 198.964
R170 VGND.n12 VGND.n11 116.692
R171 VGND.n1 VGND.t7 61.4291
R172 VGND.n11 VGND.t5 57.8264
R173 VGND.n1 VGND.t8 41.4291
R174 VGND.n39 VGND.t0 38.5719
R175 VGND.n39 VGND.t3 38.5719
R176 VGND.n19 VGND.n8 34.6358
R177 VGND.n20 VGND.n19 34.6358
R178 VGND.n21 VGND.n20 34.6358
R179 VGND.n26 VGND.n25 34.6358
R180 VGND.n27 VGND.n26 34.6358
R181 VGND.n32 VGND.n31 34.6358
R182 VGND.n33 VGND.n32 34.6358
R183 VGND.n38 VGND.n37 34.6358
R184 VGND.n15 VGND.n14 33.1299
R185 VGND.n27 VGND.n4 32.0005
R186 VGND.n14 VGND.n13 31.2476
R187 VGND.n25 VGND.n6 28.9887
R188 VGND.n37 VGND.n2 25.977
R189 VGND.n10 VGND.t6 24.9236
R190 VGND.n10 VGND.t9 24.9236
R191 VGND.n11 VGND.t2 24.7418
R192 VGND.n40 VGND.n38 22.9652
R193 VGND.n31 VGND.n4 22.2123
R194 VGND.n33 VGND.n2 18.4476
R195 VGND.n21 VGND.n6 12.424
R196 VGND.n13 VGND.n12 10.9322
R197 VGND.n38 VGND.n0 9.3005
R198 VGND.n37 VGND.n36 9.3005
R199 VGND.n35 VGND.n2 9.3005
R200 VGND.n34 VGND.n33 9.3005
R201 VGND.n32 VGND.n3 9.3005
R202 VGND.n31 VGND.n30 9.3005
R203 VGND.n29 VGND.n4 9.3005
R204 VGND.n28 VGND.n27 9.3005
R205 VGND.n26 VGND.n5 9.3005
R206 VGND.n25 VGND.n24 9.3005
R207 VGND.n23 VGND.n6 9.3005
R208 VGND.n22 VGND.n21 9.3005
R209 VGND.n20 VGND.n7 9.3005
R210 VGND.n19 VGND.n18 9.3005
R211 VGND.n17 VGND.n8 9.3005
R212 VGND.n16 VGND.n15 9.3005
R213 VGND.n14 VGND.n9 9.3005
R214 VGND.n15 VGND.n8 8.28285
R215 VGND.n41 VGND.n40 7.12063
R216 VGND.n12 VGND.n9 0.203707
R217 VGND.n41 VGND.n0 0.148519
R218 VGND.n16 VGND.n9 0.120292
R219 VGND.n17 VGND.n16 0.120292
R220 VGND.n18 VGND.n17 0.120292
R221 VGND.n18 VGND.n7 0.120292
R222 VGND.n22 VGND.n7 0.120292
R223 VGND.n23 VGND.n22 0.120292
R224 VGND.n24 VGND.n23 0.120292
R225 VGND.n24 VGND.n5 0.120292
R226 VGND.n28 VGND.n5 0.120292
R227 VGND.n29 VGND.n28 0.120292
R228 VGND.n30 VGND.n29 0.120292
R229 VGND.n30 VGND.n3 0.120292
R230 VGND.n34 VGND.n3 0.120292
R231 VGND.n35 VGND.n34 0.120292
R232 VGND.n36 VGND.n35 0.120292
R233 VGND.n36 VGND.n0 0.120292
R234 VGND VGND.n41 0.114842
R235 Q.n0 Q.t1 558.89
R236 Q.n0 Q.t0 129.232
R237 Q Q.n0 5.4997
R238 a_1948_47.t1 a_1948_47.n1 390.777
R239 a_1948_47.n1 a_1948_47.t0 258.99
R240 a_1948_47.n0 a_1948_47.t3 239.04
R241 a_1948_47.n1 a_1948_47.n0 174.109
R242 a_1948_47.n0 a_1948_47.t2 166.739
R243 Q_N Q_N.t1 379.89
R244 Q_N Q_N.t0 257.825
R245 CLK.n0 CLK.t0 292.95
R246 CLK.n0 CLK.t1 209.403
R247 CLK CLK.n0 154.069
R248 a_27_47.n4 a_27_47.t3 501.817
R249 a_27_47.n3 a_27_47.n2 448.26
R250 a_27_47.t1 a_27_47.n6 390.443
R251 a_27_47.n1 a_27_47.t0 290.872
R252 a_27_47.n0 a_27_47.t5 263.406
R253 a_27_47.n3 a_27_47.t2 254.389
R254 a_27_47.n0 a_27_47.t4 228.06
R255 a_27_47.n5 a_27_47.n3 193.447
R256 a_27_47.n5 a_27_47.n4 166.708
R257 a_27_47.n1 a_27_47.n0 152
R258 a_27_47.n4 a_27_47.t6 148.35
R259 a_27_47.n6 a_27_47.n1 35.3396
R260 a_27_47.n6 a_27_47.n5 13.2349
R261 a_657_47.t0 a_657_47.t1 65.7148
R262 SCD.n0 SCD.t1 268.849
R263 SCD.n0 SCD.t0 236.716
R264 SCD SCD.n0 158.667
R265 a_483_47.t0 a_483_47.t1 68.5719
R266 a_1027_47.t0 a_1027_47.t1 98.0601
R267 a_1475_47.n0 a_1475_47.t0 11.0774
C0 SCE VPB 0.108963f
C1 Q VPB 0.012184f
C2 SCD SCE 0.044967f
C3 SCE VGND 0.112398f
C4 Q VGND 0.081895f
C5 Q_N VPWR 0.099695f
C6 VPWR a_1089_183# 0.102299f
C7 CLK VPB 0.069635f
C8 D SCE 0.104236f
C9 CLK VGND 0.019296f
C10 SCE VPWR 0.025911f
C11 Q VPWR 0.116712f
C12 SCD VPB 0.06725f
C13 VGND VPB 0.015998f
C14 SCD VGND 0.010122f
C15 VPWR a_1023_413# 0.002662f
C16 CLK VPWR 0.019263f
C17 D VPB 0.054102f
C18 VPWR VPB 0.240795f
C19 D SCD 0.006114f
C20 SCD VPWR 0.010663f
C21 D VGND 0.00928f
C22 VPWR VGND 0.100535f
C23 Q_N VPB 0.010916f
C24 VPB a_1089_183# 0.073615f
C25 Q_N VGND 0.082678f
C26 D VPWR 0.008024f
C27 VGND a_1089_183# 0.124169f
C28 Q_N VNB 0.087247f
C29 Q VNB 0.008531f
C30 VGND VNB 1.20729f
C31 VPWR VNB 0.988242f
C32 SCD VNB 0.121325f
C33 D VNB 0.101787f
C34 SCE VNB 0.241707f
C35 CLK VNB 0.195128f
C36 VPB VNB 2.19949f
C37 a_1089_183# VNB 0.150154f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxbp_2 VGND VPWR VNB VPB Q_N Q SCD SCE D CLK
X0 VPWR.t8 a_1525_315.t2 Q.t2 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 a_466_369.t1 SCE.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1024 pd=0.96 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_938_413.t3 a_27_47.t2 a_560_369.t5 VNB.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1008 ps=1.28 w=0.36 l=0.15
X3 Q.t3 a_1525_315.t3 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X4 VPWR.t4 SCD.t0 a_644_369.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1824 pd=1.85 as=0.1008 ps=0.955 w=0.64 l=0.15
X5 Q.t1 a_1525_315.t4 VPWR.t7 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X6 VPWR.t3 SCE.t1 a_299_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_1354_413.t0 a_193_47.t2 a_1097_183# VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X8 VGND.t8 a_1525_315.t5 a_1483_47.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_1097_183# a_1031_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_487_47.t1 a_299_47.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X12 Q_N.t1 a_2049_47.t2 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X13 a_193_47.t0 a_27_47.t3 VGND.t11 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1031_413# a_27_47.t4 a_938_413.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X15 VGND.t2 a_1354_413.t3 a_1525_315.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VGND.t7 a_1525_315.t6 a_2049_47.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 a_1438_413.t0 a_193_47.t3 a_1354_413.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR.t1 a_1354_413.t4 a_1525_315.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.26 ps=2.52 w=1 l=0.15
X19 a_1354_413.t2 a_27_47.t5 a_1097_183# VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X20 VGND.t6 SCE.t2 a_299_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.1176 ps=1.4 w=0.42 l=0.15
X21 a_644_369.t0 a_299_47.t3 a_560_369.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1008 pd=0.955 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_661_47.t1 SCE.t3 a_560_369.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 VGND.t3 SCD.t1 a_661_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0483 ps=0.65 w=0.42 l=0.15
X24 VGND.t4 a_1097_183# a_1035_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X25 a_560_369.t3 D.t0 a_466_369.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1024 ps=0.96 w=0.64 l=0.15
X26 VPWR.t9 a_1525_315.t7 a_2049_47.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X27 a_560_369.t0 D.t1 a_487_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0504 ps=0.66 w=0.42 l=0.15
X28 Q_N.t0 a_2049_47.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X29 a_193_47.t1 a_27_47.t6 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 a_1035_47.t1 a_193_47.t4 a_938_413.t0 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X31 VGND.t9 a_1525_315.t8 Q.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_938_413.t1 a_193_47.t5 a_560_369.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1113 ps=1.37 w=0.42 l=0.15
X33 VGND.t5 CLK.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1525_315.n5 a_1525_315.t5 383.5
R1 a_1525_315.n0 a_1525_315.t7 256.988
R2 a_1525_315.t1 a_1525_315.n6 224.66
R3 a_1525_315.n1 a_1525_315.t2 212.081
R4 a_1525_315.n2 a_1525_315.t4 212.081
R5 a_1525_315.n6 a_1525_315.n5 178.376
R6 a_1525_315.n3 a_1525_315.n2 176.643
R7 a_1525_315.n0 a_1525_315.t6 163.803
R8 a_1525_315.n3 a_1525_315.t0 149.856
R9 a_1525_315.n1 a_1525_315.t8 139.78
R10 a_1525_315.n2 a_1525_315.t3 139.78
R11 a_1525_315.n5 a_1525_315.n4 139.286
R12 a_1525_315.n1 a_1525_315.n0 130.725
R13 a_1525_315.n2 a_1525_315.n1 61.346
R14 a_1525_315.n6 a_1525_315.n3 20.0129
R15 Q.n1 Q.n0 324.151
R16 Q Q.n2 187.522
R17 Q.n2 Q.n1 185
R18 Q.n0 Q.t2 26.5955
R19 Q.n0 Q.t1 26.5955
R20 Q.n2 Q.t0 24.9236
R21 Q.n2 Q.t3 24.9236
R22 Q Q.n1 10.6672
R23 VPWR.n5 VPWR.t4 722.018
R24 VPWR.n45 VPWR.n1 604.394
R25 VPWR.n3 VPWR.n2 600.128
R26 VPWR.n15 VPWR.t8 426.704
R27 VPWR.n12 VPWR.n11 337.132
R28 VPWR.n14 VPWR.n13 236.686
R29 VPWR.n13 VPWR.t9 61.9924
R30 VPWR.n1 VPWR.t6 41.5552
R31 VPWR.n1 VPWR.t0 41.5552
R32 VPWR.n2 VPWR.t2 41.5552
R33 VPWR.n2 VPWR.t3 41.5552
R34 VPWR.n44 VPWR.n43 34.6358
R35 VPWR.n22 VPWR.n9 34.6358
R36 VPWR.n26 VPWR.n9 34.6358
R37 VPWR.n27 VPWR.n26 34.6358
R38 VPWR.n28 VPWR.n27 34.6358
R39 VPWR.n28 VPWR.n7 34.6358
R40 VPWR.n32 VPWR.n7 34.6358
R41 VPWR.n33 VPWR.n32 34.6358
R42 VPWR.n34 VPWR.n33 34.6358
R43 VPWR.n38 VPWR.n37 34.6358
R44 VPWR.n39 VPWR.n38 34.6358
R45 VPWR.n16 VPWR.n15 31.624
R46 VPWR.n13 VPWR.t5 30.164
R47 VPWR.n21 VPWR.n20 30.1181
R48 VPWR.n37 VPWR.n5 29.7417
R49 VPWR.n20 VPWR.n12 28.9887
R50 VPWR.n11 VPWR.t7 28.5655
R51 VPWR.n11 VPWR.t1 28.5655
R52 VPWR.n16 VPWR.n12 26.7299
R53 VPWR.n39 VPWR.n3 24.0946
R54 VPWR.n45 VPWR.n44 22.5887
R55 VPWR.n43 VPWR.n3 20.3299
R56 VPWR.n22 VPWR.n21 16.1887
R57 VPWR.n15 VPWR.n14 10.3382
R58 VPWR.n17 VPWR.n16 9.3005
R59 VPWR.n18 VPWR.n12 9.3005
R60 VPWR.n20 VPWR.n19 9.3005
R61 VPWR.n21 VPWR.n10 9.3005
R62 VPWR.n23 VPWR.n22 9.3005
R63 VPWR.n24 VPWR.n9 9.3005
R64 VPWR.n26 VPWR.n25 9.3005
R65 VPWR.n27 VPWR.n8 9.3005
R66 VPWR.n29 VPWR.n28 9.3005
R67 VPWR.n30 VPWR.n7 9.3005
R68 VPWR.n32 VPWR.n31 9.3005
R69 VPWR.n33 VPWR.n6 9.3005
R70 VPWR.n35 VPWR.n34 9.3005
R71 VPWR.n37 VPWR.n36 9.3005
R72 VPWR.n38 VPWR.n4 9.3005
R73 VPWR.n40 VPWR.n39 9.3005
R74 VPWR.n41 VPWR.n3 9.3005
R75 VPWR.n43 VPWR.n42 9.3005
R76 VPWR.n44 VPWR.n0 9.3005
R77 VPWR.n46 VPWR.n45 7.14087
R78 VPWR.n34 VPWR.n5 4.89462
R79 VPWR.n17 VPWR.n14 0.412086
R80 VPWR.n46 VPWR.n0 0.148262
R81 VPWR.n18 VPWR.n17 0.120292
R82 VPWR.n19 VPWR.n18 0.120292
R83 VPWR.n19 VPWR.n10 0.120292
R84 VPWR.n23 VPWR.n10 0.120292
R85 VPWR.n24 VPWR.n23 0.120292
R86 VPWR.n25 VPWR.n24 0.120292
R87 VPWR.n25 VPWR.n8 0.120292
R88 VPWR.n29 VPWR.n8 0.120292
R89 VPWR.n30 VPWR.n29 0.120292
R90 VPWR.n31 VPWR.n30 0.120292
R91 VPWR.n31 VPWR.n6 0.120292
R92 VPWR.n35 VPWR.n6 0.120292
R93 VPWR.n36 VPWR.n35 0.120292
R94 VPWR.n36 VPWR.n4 0.120292
R95 VPWR.n40 VPWR.n4 0.120292
R96 VPWR.n41 VPWR.n40 0.120292
R97 VPWR.n42 VPWR.n41 0.120292
R98 VPWR.n42 VPWR.n0 0.120292
R99 VPWR VPWR.n46 0.115103
R100 VPB.t6 VPB.t1 979.596
R101 VPB.t3 VPB.t10 955.919
R102 VPB.t7 VPB.t8 594.861
R103 VPB.t15 VPB.t13 562.306
R104 VPB.t11 VPB.t5 556.386
R105 VPB.t13 VPB.t9 287.072
R106 VPB.t4 VPB.t12 278.193
R107 VPB.t8 VPB.t3 275.235
R108 VPB.t2 VPB.t7 275.235
R109 VPB.t1 VPB.t14 260.437
R110 VPB.t14 VPB.t15 248.599
R111 VPB.t10 VPB.t6 248.599
R112 VPB.t12 VPB.t2 248.599
R113 VPB.t5 VPB.t4 248.599
R114 VPB.t0 VPB.t11 248.599
R115 VPB VPB.t0 145.017
R116 SCE.n2 SCE.t3 342.286
R117 SCE.n1 SCE.t2 321.772
R118 SCE.n2 SCE.n1 253.272
R119 SCE.n0 SCE.t0 236.18
R120 SCE.n0 SCE.t1 174.835
R121 SCE SCE.n2 20.1148
R122 SCE.n1 SCE.n0 8.76414
R123 a_466_369.t0 a_466_369.t1 98.5005
R124 a_27_47.n4 a_27_47.t2 501.817
R125 a_27_47.n3 a_27_47.n2 448.26
R126 a_27_47.t0 a_27_47.n6 390.067
R127 a_27_47.n1 a_27_47.t1 290.872
R128 a_27_47.n0 a_27_47.t6 263.173
R129 a_27_47.n3 a_27_47.t5 254.389
R130 a_27_47.n0 a_27_47.t3 227.826
R131 a_27_47.n5 a_27_47.n3 193.457
R132 a_27_47.n5 a_27_47.n4 166.708
R133 a_27_47.n1 a_27_47.n0 152
R134 a_27_47.n4 a_27_47.t4 148.35
R135 a_27_47.n6 a_27_47.n1 35.3396
R136 a_27_47.n6 a_27_47.n5 13.2706
R137 a_560_369.n3 a_560_369.n2 705.847
R138 a_560_369.n2 a_560_369.t2 665.538
R139 a_560_369.n1 a_560_369.n0 299.825
R140 a_560_369.n1 a_560_369.t5 256.243
R141 a_560_369.n2 a_560_369.n1 72.2828
R142 a_560_369.n0 a_560_369.t0 54.2862
R143 a_560_369.t1 a_560_369.n3 41.5552
R144 a_560_369.n3 a_560_369.t3 41.5552
R145 a_560_369.n0 a_560_369.t4 40.0005
R146 a_938_413.n5 a_938_413.n4 693.048
R147 a_938_413.n4 a_938_413.n3 300.243
R148 a_938_413.n2 a_938_413.n1 226.541
R149 a_938_413.n2 a_938_413.n0 196.013
R150 a_938_413.n4 a_938_413.n2 168.738
R151 a_938_413.t1 a_938_413.n5 75.0481
R152 a_938_413.n5 a_938_413.t2 72.7029
R153 a_938_413.n3 a_938_413.t3 65.0005
R154 a_938_413.n3 a_938_413.t0 45.0005
R155 VNB.t5 VNB.t7 3517.15
R156 VNB.t4 VNB.t16 2876.38
R157 VNB.t7 VNB.t13 2819.42
R158 VNB.t15 VNB.t10 2733.98
R159 VNB.t13 VNB.t3 2719.74
R160 VNB.t11 VNB.t12 2705.5
R161 VNB.t10 VNB.t2 1452.43
R162 VNB.t8 VNB.t5 1395.47
R163 VNB.t12 VNB.t1 1381.23
R164 VNB.t16 VNB.t8 1366.99
R165 VNB.t0 VNB.t9 1366.99
R166 VNB.t3 VNB.t14 1253.07
R167 VNB.t14 VNB.t11 1196.12
R168 VNB.t6 VNB.t15 1196.12
R169 VNB.t2 VNB.t0 1110.68
R170 VNB.t9 VNB.t4 1082.2
R171 VNB VNB.t6 683.495
R172 VGND.n6 VGND.t4 286.673
R173 VGND.n4 VGND.t3 255.184
R174 VGND.n13 VGND.t9 240.988
R175 VGND.n19 VGND.t8 239.139
R176 VGND.n17 VGND.n11 220.706
R177 VGND.n44 VGND.n43 199.739
R178 VGND.n2 VGND.n1 198.964
R179 VGND.n14 VGND.n12 116.216
R180 VGND.n1 VGND.t6 61.4291
R181 VGND.n12 VGND.t7 57.8264
R182 VGND.n1 VGND.t1 41.4291
R183 VGND.n43 VGND.t11 38.5719
R184 VGND.n43 VGND.t5 38.5719
R185 VGND.n23 VGND.n8 34.6358
R186 VGND.n24 VGND.n23 34.6358
R187 VGND.n25 VGND.n24 34.6358
R188 VGND.n30 VGND.n29 34.6358
R189 VGND.n31 VGND.n30 34.6358
R190 VGND.n36 VGND.n35 34.6358
R191 VGND.n37 VGND.n36 34.6358
R192 VGND.n42 VGND.n41 34.6358
R193 VGND.n29 VGND.n6 32.0005
R194 VGND.n31 VGND.n4 30.4946
R195 VGND.n19 VGND.n18 30.1181
R196 VGND.n18 VGND.n17 28.9887
R197 VGND.n41 VGND.n2 27.4829
R198 VGND.n11 VGND.t10 26.7697
R199 VGND.n11 VGND.t2 26.7697
R200 VGND.n17 VGND.n10 25.977
R201 VGND.n12 VGND.t0 24.7418
R202 VGND.n13 VGND.n10 24.4711
R203 VGND.n35 VGND.n4 23.7181
R204 VGND.n44 VGND.n42 22.9652
R205 VGND.n37 VGND.n2 16.9417
R206 VGND.n19 VGND.n8 11.2946
R207 VGND.n25 VGND.n6 9.41227
R208 VGND.n42 VGND.n0 9.3005
R209 VGND.n41 VGND.n40 9.3005
R210 VGND.n39 VGND.n2 9.3005
R211 VGND.n38 VGND.n37 9.3005
R212 VGND.n36 VGND.n3 9.3005
R213 VGND.n35 VGND.n34 9.3005
R214 VGND.n33 VGND.n4 9.3005
R215 VGND.n32 VGND.n31 9.3005
R216 VGND.n30 VGND.n5 9.3005
R217 VGND.n29 VGND.n28 9.3005
R218 VGND.n27 VGND.n6 9.3005
R219 VGND.n26 VGND.n25 9.3005
R220 VGND.n24 VGND.n7 9.3005
R221 VGND.n23 VGND.n22 9.3005
R222 VGND.n21 VGND.n8 9.3005
R223 VGND.n20 VGND.n19 9.3005
R224 VGND.n18 VGND.n9 9.3005
R225 VGND.n17 VGND.n16 9.3005
R226 VGND.n15 VGND.n10 9.3005
R227 VGND.n45 VGND.n44 7.12063
R228 VGND.n14 VGND.n13 6.98836
R229 VGND.n15 VGND.n14 0.473965
R230 VGND.n45 VGND.n0 0.148519
R231 VGND.n16 VGND.n15 0.120292
R232 VGND.n16 VGND.n9 0.120292
R233 VGND.n20 VGND.n9 0.120292
R234 VGND.n21 VGND.n20 0.120292
R235 VGND.n22 VGND.n21 0.120292
R236 VGND.n22 VGND.n7 0.120292
R237 VGND.n26 VGND.n7 0.120292
R238 VGND.n27 VGND.n26 0.120292
R239 VGND.n28 VGND.n27 0.120292
R240 VGND.n28 VGND.n5 0.120292
R241 VGND.n32 VGND.n5 0.120292
R242 VGND.n33 VGND.n32 0.120292
R243 VGND.n34 VGND.n33 0.120292
R244 VGND.n34 VGND.n3 0.120292
R245 VGND.n38 VGND.n3 0.120292
R246 VGND.n39 VGND.n38 0.120292
R247 VGND.n40 VGND.n39 0.120292
R248 VGND.n40 VGND.n0 0.120292
R249 VGND VGND.n45 0.114842
R250 SCD.n0 SCD.t1 268.849
R251 SCD.n0 SCD.t0 236.716
R252 SCD SCD.n0 158.4
R253 a_644_369.t0 a_644_369.t1 96.9614
R254 a_299_47.t1 a_299_47.n1 636.33
R255 a_299_47.n0 a_299_47.t3 416.856
R256 a_299_47.n0 a_299_47.t2 382.026
R257 a_299_47.n1 a_299_47.t0 344.036
R258 a_299_47.n1 a_299_47.n0 29.4703
R259 a_193_47.t1 a_193_47.n3 424.863
R260 a_193_47.n0 a_193_47.t3 348.661
R261 a_193_47.n1 a_193_47.t5 344.252
R262 a_193_47.n1 a_193_47.t4 282.788
R263 a_193_47.n0 a_193_47.t2 271.262
R264 a_193_47.n3 a_193_47.t0 242.661
R265 a_193_47.n2 a_193_47.n0 18.4548
R266 a_193_47.n3 a_193_47.n2 12.4983
R267 a_193_47.n2 a_193_47.n1 9.3005
R268 a_1354_413.n2 a_1354_413.n1 693.449
R269 a_1354_413.n1 a_1354_413.t0 317.325
R270 a_1354_413.n1 a_1354_413.n0 254.258
R271 a_1354_413.n0 a_1354_413.t4 212.081
R272 a_1354_413.n0 a_1354_413.t3 139.78
R273 a_1354_413.t1 a_1354_413.n2 63.3219
R274 a_1354_413.n2 a_1354_413.t2 63.3219
R275 a_1483_47.n0 a_1483_47.t0 11.0774
R276 CLK.n0 CLK.t0 294.557
R277 CLK.n0 CLK.t1 209.403
R278 CLK CLK.n0 153.871
R279 a_2049_47.t1 a_2049_47.n4 386.31
R280 a_2049_47.n4 a_2049_47.t0 249.956
R281 a_2049_47.n2 a_2049_47.n0 212.081
R282 a_2049_47.n3 a_2049_47.t2 212.081
R283 a_2049_47.n4 a_2049_47.n3 188.077
R284 a_2049_47.n2 a_2049_47.n1 139.78
R285 a_2049_47.n3 a_2049_47.t3 139.78
R286 a_2049_47.n3 a_2049_47.n2 61.346
R287 Q_N Q_N.t1 377.966
R288 Q_N Q_N.t0 258.957
R289 a_487_47.t0 a_487_47.t1 68.5719
R290 a_661_47.t0 a_661_47.t1 65.7148
R291 a_1035_47.t0 a_1035_47.t1 98.0601
R292 D.n0 D.t1 321.87
R293 D.n0 D.t0 183.696
R294 D D.n0 161.115
C0 VPB SCD 0.067797f
C1 Q_N VGND 0.139845f
C2 SCE VGND 0.110929f
C3 a_1097_183# VPWR 0.101889f
C4 SCE D 0.102564f
C5 VPB VGND 0.020019f
C6 VPB D 0.054539f
C7 Q VGND 0.122626f
C8 Q_N VPWR 0.177426f
C9 CLK VGND 0.019316f
C10 SCE VPWR 0.025893f
C11 VPB a_1097_183# 0.073615f
C12 VPB VPWR 0.26791f
C13 VGND SCD 0.010136f
C14 Q VPWR 0.17786f
C15 CLK VPWR 0.019412f
C16 Q_N VPB 0.004284f
C17 D SCD 0.006114f
C18 SCE VPB 0.108437f
C19 VGND D 0.00928f
C20 VPWR SCD 0.010908f
C21 a_1031_413# VPWR 0.002659f
C22 Q VPB 0.005546f
C23 CLK VPB 0.070163f
C24 a_1097_183# VGND 0.124022f
C25 VPWR VGND 0.141013f
C26 SCE SCD 0.046103f
C27 VPWR D 0.008006f
C28 Q_N VNB 0.020269f
C29 Q VNB 0.0045f
C30 VGND VNB 1.33047f
C31 VPWR VNB 1.10363f
C32 SCD VNB 0.12227f
C33 D VNB 0.101787f
C34 SCE VNB 0.241924f
C35 CLK VNB 0.195347f
C36 VPB VNB 2.37668f
C37 a_1097_183# VNB 0.150154f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxtp_1 VPWR VGND Q CLK D SCE SCD VPB VNB
X0 a_640_369.t0 a_299_47.t2 a_556_369.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1024 pd=0.96 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_933_413.t2 a_193_47.t2 a_556_369.t5 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.45 w=0.42 l=0.15
X2 a_556_369.t2 D.t0 a_467_369.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0944 ps=0.935 w=0.64 l=0.15
X3 a_1030_47.t0 a_193_47.t3 a_933_413.t3 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X4 a_1092_183.t1 a_933_413.t4 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X5 VPWR.t6 a_1349_413.t3 a_1520_315.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR.t0 SCE.t0 a_299_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.088 pd=0.915 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 Q.t1 a_1520_315.t2 VPWR.t7 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X8 VPWR.t4 CLK.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_467_369.t0 SCE.t1 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0944 pd=0.935 as=0.088 ps=0.915 w=0.64 l=0.15
X10 a_1026_413.t1 a_27_47.t2 a_933_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X11 a_657_47.t1 SCE.t2 a_556_369.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 VPWR.t8 a_1520_315.t3 a_1433_413.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.59 as=0.09135 ps=0.855 w=0.42 l=0.15
X13 Q.t0 a_1520_315.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X14 a_933_413.t0 a_27_47.t3 a_556_369.t1 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.099 ps=1.27 w=0.36 l=0.15
X15 VPWR.t1 a_1092_183.t3 a_1026_413.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 VGND.t7 a_1092_183.t4 a_1030_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X17 VGND.t2 a_1520_315.t5 a_1478_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X18 a_193_47.t1 a_27_47.t4 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_483_47.t0 a_299_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0714 ps=0.76 w=0.42 l=0.15
X20 a_1478_47.t0 a_27_47.t5 a_1349_413.t2 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X21 VPWR.t3 SCD.t0 a_640_369.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.1024 ps=0.96 w=0.64 l=0.15
X22 a_1433_413.t0 a_193_47.t4 a_1349_413.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 VGND.t4 SCE.t3 a_299_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0714 pd=0.76 as=0.1176 ps=1.4 w=0.42 l=0.15
X24 a_1092_183.t2 a_933_413.t5 VPWR.t9 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X25 a_1349_413.t0 a_27_47.t6 a_1092_183.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X26 VGND.t3 a_1349_413.t4 a_1520_315.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X27 VGND.t5 SCD.t1 a_657_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0483 ps=0.65 w=0.42 l=0.15
X28 a_193_47.t0 a_27_47.t7 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X29 VGND.t9 CLK.t1 a_27_47.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 a_556_369.t3 D.t1 a_483_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 a_299_47.t0 a_299_47.n1 635.824
R1 a_299_47.n0 a_299_47.t2 433.969
R2 a_299_47.n0 a_299_47.t3 380.75
R3 a_299_47.n1 a_299_47.t1 345.021
R4 a_299_47.n1 a_299_47.n0 29.1726
R5 a_556_369.n3 a_556_369.n2 705.471
R6 a_556_369.n2 a_556_369.t5 685.899
R7 a_556_369.n1 a_556_369.n0 300.954
R8 a_556_369.n1 a_556_369.t1 250.072
R9 a_556_369.n2 a_556_369.n1 70.777
R10 a_556_369.n0 a_556_369.t3 54.2862
R11 a_556_369.t0 a_556_369.n3 41.5552
R12 a_556_369.n3 a_556_369.t2 41.5552
R13 a_556_369.n0 a_556_369.t4 40.0005
R14 a_640_369.t0 a_640_369.t1 98.5005
R15 VPB.t15 VPB.t8 624.456
R16 VPB.t6 VPB.t11 588.942
R17 VPB.t4 VPB.t2 556.386
R18 VPB.t13 VPB.t1 390.654
R19 VPB.t12 VPB.t15 346.262
R20 VPB.t7 VPB.t13 284.113
R21 VPB.t1 VPB.t3 281.154
R22 VPB.t0 VPB.t6 278.193
R23 VPB.t11 VPB.t7 275.235
R24 VPB.t8 VPB.t14 269.315
R25 VPB.t10 VPB.t5 263.397
R26 VPB.t2 VPB.t10 251.559
R27 VPB.t3 VPB.t12 248.599
R28 VPB.t5 VPB.t0 248.599
R29 VPB.t9 VPB.t4 248.599
R30 VPB VPB.t9 145.017
R31 a_193_47.t0 a_193_47.n4 429.714
R32 a_193_47.n1 a_193_47.t4 348.661
R33 a_193_47.n2 a_193_47.t2 347.389
R34 a_193_47.n2 a_193_47.t3 283.928
R35 a_193_47.n1 a_193_47.n0 271.262
R36 a_193_47.n4 a_193_47.t1 244.006
R37 a_193_47.n3 a_193_47.n1 17.864
R38 a_193_47.n4 a_193_47.n3 12.5072
R39 a_193_47.n3 a_193_47.n2 9.3005
R40 a_933_413.n3 a_933_413.n2 693.048
R41 a_933_413.n2 a_933_413.n1 300.243
R42 a_933_413.n0 a_933_413.t4 226.541
R43 a_933_413.n0 a_933_413.t5 196.013
R44 a_933_413.n2 a_933_413.n0 168.738
R45 a_933_413.n3 a_933_413.t2 75.0481
R46 a_933_413.t1 a_933_413.n3 72.7029
R47 a_933_413.n1 a_933_413.t0 65.0005
R48 a_933_413.n1 a_933_413.t3 45.0005
R49 D.n0 D.t1 321.87
R50 D.n0 D.t0 183.696
R51 D D.n0 159.758
R52 a_467_369.t0 a_467_369.t1 90.8052
R53 a_1030_47.t1 a_1030_47.t0 98.0601
R54 VNB.t12 VNB.t10 2904.85
R55 VNB.t7 VNB.t1 2862.14
R56 VNB.t9 VNB.t6 2733.98
R57 VNB.t3 VNB.t5 2677.02
R58 VNB.t11 VNB.t12 2078.96
R59 VNB.t8 VNB.t11 1395.47
R60 VNB.t6 VNB.t0 1395.47
R61 VNB.t1 VNB.t8 1366.99
R62 VNB.t14 VNB.t4 1366.99
R63 VNB.t10 VNB.t3 1352.75
R64 VNB.t5 VNB.t2 1295.79
R65 VNB.t13 VNB.t9 1196.12
R66 VNB.t0 VNB.t14 1110.68
R67 VNB.t4 VNB.t7 1082.2
R68 VNB VNB.t13 683.495
R69 VGND.n4 VGND.t5 262.178
R70 VGND.n10 VGND.t2 239.139
R71 VGND.n12 VGND.n11 225.395
R72 VGND.n36 VGND.n35 199.739
R73 VGND.n7 VGND.n6 199.53
R74 VGND.n2 VGND.n1 198.357
R75 VGND.n6 VGND.t7 87.1434
R76 VGND.n6 VGND.t8 66.2951
R77 VGND.n1 VGND.t4 57.1434
R78 VGND.n1 VGND.t0 40.0005
R79 VGND.n35 VGND.t6 38.5719
R80 VGND.n35 VGND.t9 38.5719
R81 VGND.n15 VGND.n9 34.6358
R82 VGND.n16 VGND.n15 34.6358
R83 VGND.n17 VGND.n16 34.6358
R84 VGND.n22 VGND.n21 34.6358
R85 VGND.n23 VGND.n22 34.6358
R86 VGND.n28 VGND.n27 34.6358
R87 VGND.n29 VGND.n28 34.6358
R88 VGND.n34 VGND.n33 34.6358
R89 VGND.n23 VGND.n4 30.8711
R90 VGND.n21 VGND.n7 30.1181
R91 VGND.n11 VGND.t3 28.6159
R92 VGND.n11 VGND.t1 27.6928
R93 VGND.n33 VGND.n2 26.3534
R94 VGND.n27 VGND.n4 23.3417
R95 VGND.n36 VGND.n34 22.9652
R96 VGND.n29 VGND.n2 16.9417
R97 VGND.n17 VGND.n7 11.2946
R98 VGND.n10 VGND.n9 9.41227
R99 VGND.n34 VGND.n0 9.3005
R100 VGND.n33 VGND.n32 9.3005
R101 VGND.n31 VGND.n2 9.3005
R102 VGND.n30 VGND.n29 9.3005
R103 VGND.n28 VGND.n3 9.3005
R104 VGND.n27 VGND.n26 9.3005
R105 VGND.n13 VGND.n9 9.3005
R106 VGND.n15 VGND.n14 9.3005
R107 VGND.n16 VGND.n8 9.3005
R108 VGND.n18 VGND.n17 9.3005
R109 VGND.n19 VGND.n7 9.3005
R110 VGND.n21 VGND.n20 9.3005
R111 VGND.n22 VGND.n5 9.3005
R112 VGND.n24 VGND.n23 9.3005
R113 VGND.n25 VGND.n4 9.3005
R114 VGND.n12 VGND.n10 7.22337
R115 VGND.n37 VGND.n36 7.12063
R116 VGND.n13 VGND.n12 0.435082
R117 VGND.n37 VGND.n0 0.148519
R118 VGND.n14 VGND.n13 0.120292
R119 VGND.n14 VGND.n8 0.120292
R120 VGND.n18 VGND.n8 0.120292
R121 VGND.n19 VGND.n18 0.120292
R122 VGND.n20 VGND.n19 0.120292
R123 VGND.n20 VGND.n5 0.120292
R124 VGND.n24 VGND.n5 0.120292
R125 VGND.n25 VGND.n24 0.120292
R126 VGND.n26 VGND.n25 0.120292
R127 VGND.n26 VGND.n3 0.120292
R128 VGND.n30 VGND.n3 0.120292
R129 VGND.n31 VGND.n30 0.120292
R130 VGND.n32 VGND.n31 0.120292
R131 VGND.n32 VGND.n0 0.120292
R132 VGND VGND.n37 0.114842
R133 a_1092_183.n2 a_1092_183.n1 674.014
R134 a_1092_183.n0 a_1092_183.t3 433.8
R135 a_1092_183.n1 a_1092_183.t1 254.9
R136 a_1092_183.n1 a_1092_183.n0 185.308
R137 a_1092_183.n0 a_1092_183.t4 128.1
R138 a_1092_183.n2 a_1092_183.t0 89.1195
R139 a_1092_183.t2 a_1092_183.n2 37.5243
R140 a_1349_413.n2 a_1349_413.n1 693.449
R141 a_1349_413.n1 a_1349_413.t2 292.325
R142 a_1349_413.n1 a_1349_413.n0 249.922
R143 a_1349_413.n0 a_1349_413.t3 212.081
R144 a_1349_413.n0 a_1349_413.t4 139.78
R145 a_1349_413.n2 a_1349_413.t1 63.3219
R146 a_1349_413.t0 a_1349_413.n2 63.3219
R147 a_1520_315.t0 a_1520_315.n2 834.348
R148 a_1520_315.t0 a_1520_315.n4 816.096
R149 a_1520_315.n3 a_1520_315.t5 383.5
R150 a_1520_315.n0 a_1520_315.t2 236.934
R151 a_1520_315.n4 a_1520_315.n3 177.794
R152 a_1520_315.n1 a_1520_315.n0 172.559
R153 a_1520_315.n0 a_1520_315.t4 164.633
R154 a_1520_315.n1 a_1520_315.t1 151.163
R155 a_1520_315.n3 a_1520_315.t3 139.286
R156 a_1520_315.n2 a_1520_315.n1 20.7634
R157 a_1520_315.n4 a_1520_315.n2 1.93989
R158 VPWR.n5 VPWR.t3 730.99
R159 VPWR.n10 VPWR.t8 717.543
R160 VPWR.n37 VPWR.n1 604.394
R161 VPWR.n3 VPWR.n2 600.128
R162 VPWR.n12 VPWR.n11 340.231
R163 VPWR.n18 VPWR.n17 320.976
R164 VPWR.n17 VPWR.t1 113.98
R165 VPWR.n2 VPWR.t5 43.0943
R166 VPWR.n1 VPWR.t2 41.5552
R167 VPWR.n1 VPWR.t4 41.5552
R168 VPWR.n2 VPWR.t0 41.5552
R169 VPWR.n17 VPWR.t9 35.4605
R170 VPWR.n36 VPWR.n35 34.6358
R171 VPWR.n30 VPWR.n29 34.6358
R172 VPWR.n31 VPWR.n30 34.6358
R173 VPWR.n15 VPWR.n9 34.6358
R174 VPWR.n16 VPWR.n15 34.6358
R175 VPWR.n19 VPWR.n16 34.6358
R176 VPWR.n23 VPWR.n7 34.6358
R177 VPWR.n24 VPWR.n23 34.6358
R178 VPWR.n25 VPWR.n24 34.6358
R179 VPWR.n25 VPWR.n5 33.5064
R180 VPWR.n11 VPWR.t6 30.5355
R181 VPWR.n11 VPWR.t7 29.5505
R182 VPWR.n31 VPWR.n3 24.0946
R183 VPWR.n37 VPWR.n36 22.5887
R184 VPWR.n29 VPWR.n5 21.0829
R185 VPWR.n35 VPWR.n3 20.3299
R186 VPWR.n18 VPWR.n7 17.6946
R187 VPWR.n19 VPWR.n18 16.9417
R188 VPWR.n10 VPWR.n9 15.0593
R189 VPWR.n13 VPWR.n9 9.3005
R190 VPWR.n15 VPWR.n14 9.3005
R191 VPWR.n16 VPWR.n8 9.3005
R192 VPWR.n20 VPWR.n19 9.3005
R193 VPWR.n21 VPWR.n7 9.3005
R194 VPWR.n23 VPWR.n22 9.3005
R195 VPWR.n24 VPWR.n6 9.3005
R196 VPWR.n26 VPWR.n25 9.3005
R197 VPWR.n27 VPWR.n5 9.3005
R198 VPWR.n29 VPWR.n28 9.3005
R199 VPWR.n30 VPWR.n4 9.3005
R200 VPWR.n32 VPWR.n31 9.3005
R201 VPWR.n33 VPWR.n3 9.3005
R202 VPWR.n35 VPWR.n34 9.3005
R203 VPWR.n36 VPWR.n0 9.3005
R204 VPWR.n12 VPWR.n10 7.19098
R205 VPWR.n38 VPWR.n37 7.14087
R206 VPWR.n13 VPWR.n12 0.439982
R207 VPWR.n38 VPWR.n0 0.148262
R208 VPWR.n14 VPWR.n13 0.120292
R209 VPWR.n14 VPWR.n8 0.120292
R210 VPWR.n20 VPWR.n8 0.120292
R211 VPWR.n21 VPWR.n20 0.120292
R212 VPWR.n22 VPWR.n21 0.120292
R213 VPWR.n22 VPWR.n6 0.120292
R214 VPWR.n26 VPWR.n6 0.120292
R215 VPWR.n27 VPWR.n26 0.120292
R216 VPWR.n28 VPWR.n27 0.120292
R217 VPWR.n28 VPWR.n4 0.120292
R218 VPWR.n32 VPWR.n4 0.120292
R219 VPWR.n33 VPWR.n32 0.120292
R220 VPWR.n34 VPWR.n33 0.120292
R221 VPWR.n34 VPWR.n0 0.120292
R222 VPWR VPWR.n38 0.115103
R223 SCE.n2 SCE.t2 331.443
R224 SCE.n1 SCE.t3 319.83
R225 SCE.n2 SCE.n1 260.62
R226 SCE.n0 SCE.t1 244.214
R227 SCE.n0 SCE.t0 175.542
R228 SCE SCE.n2 20.1148
R229 SCE.n1 SCE.n0 9.32953
R230 Q Q.n0 591.865
R231 Q.n3 Q.n0 585
R232 Q.n2 Q.n0 585
R233 Q.n1 Q.t0 129.19
R234 Q.n2 Q.n1 65.0342
R235 Q.n0 Q.t1 26.5955
R236 Q.n3 Q 6.86427
R237 Q Q.n3 5.75122
R238 Q Q.n2 5.75122
R239 Q.n1 Q 5.5918
R240 CLK.n0 CLK.t0 294.557
R241 CLK.n0 CLK.t1 209.403
R242 CLK CLK.n0 154.069
R243 a_27_47.n3 a_27_47.t3 501.817
R244 a_27_47.n2 a_27_47.t5 448.26
R245 a_27_47.t1 a_27_47.n5 390.067
R246 a_27_47.n1 a_27_47.t0 290.872
R247 a_27_47.n0 a_27_47.t7 263.173
R248 a_27_47.n2 a_27_47.t6 254.389
R249 a_27_47.n0 a_27_47.t4 227.826
R250 a_27_47.n4 a_27_47.n2 193.425
R251 a_27_47.n4 a_27_47.n3 167.611
R252 a_27_47.n1 a_27_47.n0 152
R253 a_27_47.n3 a_27_47.t2 148.35
R254 a_27_47.n5 a_27_47.n1 35.3396
R255 a_27_47.n5 a_27_47.n4 13.2751
R256 a_1026_413.t0 a_1026_413.t1 154.786
R257 a_657_47.t0 a_657_47.t1 65.7148
R258 a_1433_413.t0 a_1433_413.t1 204.036
R259 a_1478_47.t1 a_1478_47.t0 93.0601
R260 a_483_47.t0 a_483_47.t1 68.5719
R261 SCD.n0 SCD.t1 255.15
R262 SCD.n0 SCD.t0 236.115
R263 SCD SCD.n0 158.958
C0 VPWR VGND 0.070564f
C1 VGND SCE 0.112116f
C2 VPB VGND 0.012232f
C3 SCD D 0.00528f
C4 VPWR SCE 0.026023f
C5 VPB VPWR 0.208187f
C6 VPB SCE 0.108049f
C7 SCD VGND 0.010424f
C8 SCD VPWR 0.011404f
C9 SCD SCE 0.043305f
C10 VPB SCD 0.067042f
C11 VGND Q 0.075059f
C12 VPWR Q 0.10335f
C13 VGND D 0.009413f
C14 VPB Q 0.011076f
C15 CLK VGND 0.019316f
C16 VPWR D 0.008393f
C17 CLK VPWR 0.019412f
C18 SCE D 0.103105f
C19 VPB D 0.053104f
C20 VPB CLK 0.070163f
C21 Q VNB 0.088175f
C22 VGND VNB 1.06298f
C23 VPWR VNB 0.871436f
C24 SCD VNB 0.123851f
C25 D VNB 0.101763f
C26 SCE VNB 0.240657f
C27 CLK VNB 0.195347f
C28 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxtp_2 VGND VPWR VNB VPB SCD SCE D CLK Q
X0 VPWR.t8 SCD.t0 a_643_369.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1824 pd=1.85 as=0.1008 ps=0.955 w=0.64 l=0.15
X1 Q.t1 a_1526_315# VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X2 a_939_413.t3 a_193_47.t2 a_559_369.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1302 ps=1.46 w=0.42 l=0.15
X3 VGND a_1526_315# a_1484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4 VPWR.t9 SCE.t0 a_299_47.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.088 pd=0.915 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR a_1355_413# a_1526_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X6 a_1355_413# a_193_47.t3 a_1098_183.t2 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X7 VPWR.t4 a_1526_315# Q.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t7 CLK.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_467_369.t0 SCE.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0992 pd=0.95 as=0.088 ps=0.915 w=0.64 l=0.15
X10 VPWR.t5 a_1526_315# a_1439_413.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.59 as=0.09135 ps=0.855 w=0.42 l=0.15
X11 Q.t2 a_1526_315# VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X12 a_486_47.t1 a_299_47.t2 VGND.t6 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.07455 ps=0.775 w=0.42 l=0.15
X13 VPWR.t1 a_1098_183.t3 a_1032_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_193_47.t1 a_27_47.t2 VGND.t8 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1098_183.t0 a_939_413.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X16 a_643_369.t1 a_299_47.t3 a_559_369.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1008 pd=0.955 as=0.0864 ps=0.91 w=0.64 l=0.15
X17 VGND a_1355_413# a_1526_315# VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X18 a_559_369.t1 D.t0 a_467_369.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0992 ps=0.95 w=0.64 l=0.15
X19 a_939_413.t0 a_27_47.t3 a_559_369.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1008 ps=1.28 w=0.36 l=0.15
X20 a_1032_413.t0 a_27_47.t4 a_939_413.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X21 VGND.t1 SCE.t2 a_299_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.07455 pd=0.775 as=0.1176 ps=1.4 w=0.42 l=0.15
X22 VGND.t4 a_1098_183.t4 a_1036_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X23 a_1098_183.t1 a_939_413.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X24 a_660_47.t0 SCE.t3 a_559_369.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 VGND.t5 SCD.t1 a_660_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0483 ps=0.65 w=0.42 l=0.15
X26 a_1484_47# a_27_47.t5 a_1355_413# VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X27 a_193_47.t0 a_27_47.t6 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_559_369.t0 D.t1 a_486_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0504 ps=0.66 w=0.42 l=0.15
X29 a_1036_47.t1 a_193_47.t4 a_939_413.t2 VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X30 VGND.t2 a_1526_315# Q.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VGND.t7 CLK.t1 a_27_47.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 SCD.n0 SCD.t1 268.849
R1 SCD.n0 SCD.t0 236.716
R2 SCD SCD.n0 158.531
R3 a_643_369.t0 a_643_369.t1 96.9614
R4 VPWR.n5 VPWR.t8 722.018
R5 VPWR.n16 VPWR.t5 717.543
R6 VPWR.n41 VPWR.n1 604.394
R7 VPWR.n3 VPWR.n2 600.128
R8 VPWR.n12 VPWR.t3 403.082
R9 VPWR.n23 VPWR.n9 320.976
R10 VPWR.n13 VPWR.t4 271.363
R11 VPWR.n9 VPWR.t1 113.98
R12 VPWR.n2 VPWR.t0 43.0943
R13 VPWR.n1 VPWR.t6 41.5552
R14 VPWR.n1 VPWR.t7 41.5552
R15 VPWR.n2 VPWR.t9 41.5552
R16 VPWR.n9 VPWR.t2 35.4605
R17 VPWR.n40 VPWR.n39 34.6358
R18 VPWR.n17 VPWR.n10 34.6358
R19 VPWR.n21 VPWR.n10 34.6358
R20 VPWR.n22 VPWR.n21 34.6358
R21 VPWR.n24 VPWR.n7 34.6358
R22 VPWR.n28 VPWR.n7 34.6358
R23 VPWR.n29 VPWR.n28 34.6358
R24 VPWR.n30 VPWR.n29 34.6358
R25 VPWR.n34 VPWR.n33 34.6358
R26 VPWR.n35 VPWR.n34 34.6358
R27 VPWR.n15 VPWR.n12 29.7417
R28 VPWR.n16 VPWR.n15 29.7417
R29 VPWR.n33 VPWR.n5 29.3652
R30 VPWR.n35 VPWR.n3 24.0946
R31 VPWR.n41 VPWR.n40 22.5887
R32 VPWR.n39 VPWR.n3 20.3299
R33 VPWR.n24 VPWR.n23 19.9534
R34 VPWR.n17 VPWR.n16 16.5652
R35 VPWR.n23 VPWR.n22 14.6829
R36 VPWR.n15 VPWR.n14 9.3005
R37 VPWR.n16 VPWR.n11 9.3005
R38 VPWR.n18 VPWR.n17 9.3005
R39 VPWR.n19 VPWR.n10 9.3005
R40 VPWR.n21 VPWR.n20 9.3005
R41 VPWR.n22 VPWR.n8 9.3005
R42 VPWR.n25 VPWR.n24 9.3005
R43 VPWR.n26 VPWR.n7 9.3005
R44 VPWR.n28 VPWR.n27 9.3005
R45 VPWR.n29 VPWR.n6 9.3005
R46 VPWR.n31 VPWR.n30 9.3005
R47 VPWR.n33 VPWR.n32 9.3005
R48 VPWR.n34 VPWR.n4 9.3005
R49 VPWR.n36 VPWR.n35 9.3005
R50 VPWR.n37 VPWR.n3 9.3005
R51 VPWR.n39 VPWR.n38 9.3005
R52 VPWR.n40 VPWR.n0 9.3005
R53 VPWR.n42 VPWR.n41 7.14087
R54 VPWR.n13 VPWR.n12 6.84914
R55 VPWR.n30 VPWR.n5 5.27109
R56 VPWR.n14 VPWR.n13 0.582214
R57 VPWR.n42 VPWR.n0 0.148262
R58 VPWR.n14 VPWR.n11 0.120292
R59 VPWR.n18 VPWR.n11 0.120292
R60 VPWR.n19 VPWR.n18 0.120292
R61 VPWR.n20 VPWR.n19 0.120292
R62 VPWR.n20 VPWR.n8 0.120292
R63 VPWR.n25 VPWR.n8 0.120292
R64 VPWR.n26 VPWR.n25 0.120292
R65 VPWR.n27 VPWR.n26 0.120292
R66 VPWR.n27 VPWR.n6 0.120292
R67 VPWR.n31 VPWR.n6 0.120292
R68 VPWR.n32 VPWR.n31 0.120292
R69 VPWR.n32 VPWR.n4 0.120292
R70 VPWR.n36 VPWR.n4 0.120292
R71 VPWR.n37 VPWR.n36 0.120292
R72 VPWR.n38 VPWR.n37 0.120292
R73 VPWR.n38 VPWR.n0 0.120292
R74 VPWR VPWR.n42 0.115103
R75 VPB.t5 VPB.t4 893.769
R76 VPB.t2 VPB.t5 876.013
R77 VPB.t10 VPB.t3 600.779
R78 VPB.t7 VPB.t11 556.386
R79 VPB.t1 VPB.t2 390.654
R80 VPB.t12 VPB.t1 284.113
R81 VPB.t3 VPB.t12 275.235
R82 VPB.t13 VPB.t10 275.235
R83 VPB.t0 VPB.t8 272.274
R84 VPB.t11 VPB.t0 251.559
R85 VPB.t4 VPB.t6 248.599
R86 VPB.t8 VPB.t13 248.599
R87 VPB.t9 VPB.t7 248.599
R88 VPB VPB.t9 145.017
R89 VGND.n4 VGND.t5 255.184
R90 VGND.n11 VGND.t3 246.198
R91 VGND.n41 VGND.n40 199.739
R92 VGND.n7 VGND.n6 199.53
R93 VGND.n2 VGND.n1 198.964
R94 VGND.n12 VGND.t2 166.008
R95 VGND.n6 VGND.t4 87.1434
R96 VGND.n6 VGND.t0 66.2951
R97 VGND.n1 VGND.t1 61.4291
R98 VGND.n1 VGND.t6 40.0005
R99 VGND.n12 VGND.n11 38.7738
R100 VGND.n40 VGND.t8 38.5719
R101 VGND.n40 VGND.t7 38.5719
R102 VGND.n15 VGND.n14 34.6358
R103 VGND.n20 VGND.n9 34.6358
R104 VGND.n21 VGND.n20 34.6358
R105 VGND.n22 VGND.n21 34.6358
R106 VGND.n27 VGND.n26 34.6358
R107 VGND.n28 VGND.n27 34.6358
R108 VGND.n33 VGND.n32 34.6358
R109 VGND.n34 VGND.n33 34.6358
R110 VGND.n39 VGND.n38 34.6358
R111 VGND.n26 VGND.n7 32.377
R112 VGND.n28 VGND.n4 30.8711
R113 VGND.n16 VGND.n15 29.7417
R114 VGND.n38 VGND.n2 27.4829
R115 VGND.n32 VGND.n4 23.3417
R116 VGND.n41 VGND.n39 22.9652
R117 VGND.n34 VGND.n2 16.9417
R118 VGND.n16 VGND.n9 11.6711
R119 VGND.n14 VGND.n13 9.3005
R120 VGND.n15 VGND.n10 9.3005
R121 VGND.n17 VGND.n16 9.3005
R122 VGND.n18 VGND.n9 9.3005
R123 VGND.n20 VGND.n19 9.3005
R124 VGND.n21 VGND.n8 9.3005
R125 VGND.n23 VGND.n22 9.3005
R126 VGND.n24 VGND.n7 9.3005
R127 VGND.n26 VGND.n25 9.3005
R128 VGND.n27 VGND.n5 9.3005
R129 VGND.n29 VGND.n28 9.3005
R130 VGND.n30 VGND.n4 9.3005
R131 VGND.n32 VGND.n31 9.3005
R132 VGND.n33 VGND.n3 9.3005
R133 VGND.n35 VGND.n34 9.3005
R134 VGND.n36 VGND.n2 9.3005
R135 VGND.n38 VGND.n37 9.3005
R136 VGND.n39 VGND.n0 9.3005
R137 VGND.n22 VGND.n7 9.03579
R138 VGND.n42 VGND.n41 7.12063
R139 VGND.n13 VGND.n12 2.15642
R140 VGND.n14 VGND.n11 1.50638
R141 VGND.n42 VGND.n0 0.148519
R142 VGND.n13 VGND.n10 0.120292
R143 VGND.n17 VGND.n10 0.120292
R144 VGND.n18 VGND.n17 0.120292
R145 VGND.n19 VGND.n18 0.120292
R146 VGND.n19 VGND.n8 0.120292
R147 VGND.n23 VGND.n8 0.120292
R148 VGND.n24 VGND.n23 0.120292
R149 VGND.n25 VGND.n24 0.120292
R150 VGND.n25 VGND.n5 0.120292
R151 VGND.n29 VGND.n5 0.120292
R152 VGND.n30 VGND.n29 0.120292
R153 VGND.n31 VGND.n30 0.120292
R154 VGND.n31 VGND.n3 0.120292
R155 VGND.n35 VGND.n3 0.120292
R156 VGND.n36 VGND.n35 0.120292
R157 VGND.n37 VGND.n36 0.120292
R158 VGND.n37 VGND.n0 0.120292
R159 VGND VGND.n42 0.114842
R160 Q Q.n0 591.865
R161 Q.n4 Q.n0 585
R162 Q.n3 Q.n0 585
R163 Q.n1 Q 186.113
R164 Q.n2 Q.n1 185
R165 Q.n3 Q.n2 59.3683
R166 Q.n0 Q.t3 26.5955
R167 Q.n0 Q.t2 26.5955
R168 Q.n1 Q.t0 24.9236
R169 Q.n1 Q.t1 24.9236
R170 Q.n2 Q 11.5019
R171 Q.n4 Q 6.86427
R172 Q Q.n4 5.75122
R173 Q Q.n3 5.75122
R174 VNB.t7 VNB.t6 5325.57
R175 VNB.t10 VNB.t11 2904.85
R176 VNB.t14 VNB.t4 2733.98
R177 VNB.t8 VNB.t1 2078.96
R178 VNB.t2 VNB.t7 1466.67
R179 VNB.t1 VNB.t2 1438.19
R180 VNB.t4 VNB.t12 1438.19
R181 VNB.t3 VNB.t8 1395.47
R182 VNB.t11 VNB.t3 1366.99
R183 VNB.t0 VNB.t9 1366.99
R184 VNB.t6 VNB.t5 1196.12
R185 VNB.t13 VNB.t14 1196.12
R186 VNB.t12 VNB.t0 1110.68
R187 VNB.t9 VNB.t10 1082.2
R188 VNB VNB.t13 683.495
R189 a_193_47.t0 a_193_47.n4 424.863
R190 a_193_47.n1 a_193_47.n0 348.661
R191 a_193_47.n2 a_193_47.t2 344.058
R192 a_193_47.n2 a_193_47.t4 282.983
R193 a_193_47.n1 a_193_47.t3 271.262
R194 a_193_47.n4 a_193_47.t1 242.661
R195 a_193_47.n3 a_193_47.n1 19.0277
R196 a_193_47.n4 a_193_47.n3 12.4983
R197 a_193_47.n3 a_193_47.n2 9.3005
R198 a_559_369.n3 a_559_369.n2 706.601
R199 a_559_369.n2 a_559_369.t4 688.484
R200 a_559_369.n1 a_559_369.n0 300.577
R201 a_559_369.n1 a_559_369.t3 256.243
R202 a_559_369.n2 a_559_369.n1 72.2828
R203 a_559_369.n0 a_559_369.t0 54.2862
R204 a_559_369.n3 a_559_369.t5 41.5552
R205 a_559_369.t1 a_559_369.n3 41.5552
R206 a_559_369.n0 a_559_369.t2 40.0005
R207 a_939_413.n3 a_939_413.n2 693.048
R208 a_939_413.n2 a_939_413.n1 300.243
R209 a_939_413.n0 a_939_413.t4 226.541
R210 a_939_413.n0 a_939_413.t5 196.013
R211 a_939_413.n2 a_939_413.n0 168.738
R212 a_939_413.n3 a_939_413.t3 75.0481
R213 a_939_413.t1 a_939_413.n3 72.7029
R214 a_939_413.n1 a_939_413.t0 65.0005
R215 a_939_413.n1 a_939_413.t2 45.0005
R216 SCE.n2 SCE.t3 341.909
R217 SCE.n1 SCE.t2 321.305
R218 SCE.n2 SCE.n1 253.272
R219 SCE.n0 SCE.t1 237.787
R220 SCE.n0 SCE.t0 174.835
R221 SCE SCE.n2 20.1148
R222 SCE.n1 SCE.n0 8.76414
R223 a_299_47.t1 a_299_47.n1 636.33
R224 a_299_47.n0 a_299_47.t3 416.56
R225 a_299_47.n0 a_299_47.t2 381.649
R226 a_299_47.n1 a_299_47.t0 344.036
R227 a_299_47.n1 a_299_47.n0 29.4703
R228 a_1098_183.n3 a_1098_183.n2 689.168
R229 a_1098_183.n1 a_1098_183.t3 433.8
R230 a_1098_183.n2 a_1098_183.n0 218.13
R231 a_1098_183.n2 a_1098_183.n1 185.308
R232 a_1098_183.n1 a_1098_183.t4 128.1
R233 a_1098_183.n3 a_1098_183.t1 100.016
R234 a_1098_183.n0 a_1098_183.t2 63.3338
R235 a_1098_183.n0 a_1098_183.t0 36.7713
R236 CLK.n0 CLK.t0 294.557
R237 CLK.n0 CLK.t1 209.403
R238 CLK CLK.n0 154.069
R239 a_27_47.n4 a_27_47.t3 501.817
R240 a_27_47.n3 a_27_47.t5 448.26
R241 a_27_47.t1 a_27_47.n6 390.067
R242 a_27_47.n1 a_27_47.t0 290.872
R243 a_27_47.n0 a_27_47.t6 263.173
R244 a_27_47.n3 a_27_47.n2 254.389
R245 a_27_47.n0 a_27_47.t2 227.826
R246 a_27_47.n5 a_27_47.n3 193.452
R247 a_27_47.n5 a_27_47.n4 166.529
R248 a_27_47.n1 a_27_47.n0 152
R249 a_27_47.n4 a_27_47.t4 148.35
R250 a_27_47.n6 a_27_47.n1 35.3396
R251 a_27_47.n6 a_27_47.n5 13.2751
R252 a_467_369.t0 a_467_369.t1 95.4224
R253 a_486_47.t0 a_486_47.t1 68.5719
R254 a_1032_413.t0 a_1032_413.t1 154.786
R255 D.n0 D.t1 321.87
R256 D.n0 D.t0 183.696
R257 D D.n0 159.758
R258 a_1036_47.t0 a_1036_47.t1 98.0601
R259 a_660_47.t0 a_660_47.t1 65.7148
C0 VGND Q 0.128185f
C1 VGND SCD 0.010095f
C2 VGND D 0.00939f
C3 SCD SCE 0.046103f
C4 VPB VGND 0.013929f
C5 SCE D 0.103738f
C6 VPB SCE 0.108717f
C7 VGND a_1484_47# 0.006699f
C8 VGND a_1355_413# 0.12177f
C9 Q a_1526_315# 0.111382f
C10 VPB a_1526_315# 0.184682f
C11 a_1526_315# a_1484_47# 1.79e-19
C12 a_1526_315# a_1355_413# 0.290659f
C13 VGND SCE 0.110817f
C14 VGND a_1526_315# 0.174119f
C15 CLK VPWR 0.019412f
C16 Q VPWR 0.188144f
C17 SCD VPWR 0.010859f
C18 VPWR D 0.008006f
C19 VPB VPWR 0.222304f
C20 VPWR a_1484_47# 7.15e-19
C21 VPB CLK 0.070163f
C22 VPWR a_1355_413# 0.114791f
C23 VGND VPWR 0.091311f
C24 SCD D 0.006114f
C25 VPWR SCE 0.026019f
C26 CLK VGND 0.019316f
C27 VPB Q 0.004049f
C28 VPB SCD 0.067873f
C29 VPB D 0.054165f
C30 Q a_1355_413# 0.001732f
C31 VPWR a_1526_315# 0.246438f
C32 VPB a_1355_413# 0.071437f
C33 a_1355_413# a_1484_47# 0.005862f
C34 Q VNB 0.021869f
C35 VGND VNB 1.14122f
C36 VPWR VNB 0.950572f
C37 SCD VNB 0.122371f
C38 D VNB 0.101775f
C39 SCE VNB 0.242046f
C40 CLK VNB 0.195347f
C41 VPB VNB 2.0223f
C42 a_1355_413# VNB 0.159814f
C43 a_1526_315# VNB 0.33821f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxtp_4 VGND VPWR VNB VPB Q CLK D SCE SCD
X0 Q.t1 a_1527_315.t2 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1 a_466_369.t1 SCE.t0 VPWR.t9 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1024 pd=0.96 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_1356_413.t2 a_193_47.t2 a_1099_183.t1 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X3 VPWR.t7 SCD.t0 a_644_369.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1824 pd=1.85 as=0.1008 ps=0.955 w=0.64 l=0.15
X4 VPWR.t10 SCE.t1 a_299_47.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_940_413.t1 a_193_47.t3 a_560_369.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1302 ps=1.46 w=0.42 l=0.15
X6 VPWR.t5 CLK.t0 a_27_47.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_487_47.t1 a_299_47.t2 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X8 VPWR.t8 a_1356_413.t4 a_1527_315.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X9 a_1099_183.t3 a_940_413.t4 VGND.t8 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X10 a_193_47.t0 a_27_47.t2 VGND.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VPWR.t1 a_1527_315.t3 a_1440_413.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.59 as=0.09135 ps=0.855 w=0.42 l=0.15
X12 VGND.t1 a_1356_413.t5 a_1527_315.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VPWR.t0 a_1099_183.t4 a_1033_413.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_940_413.t3 a_27_47.t3 a_560_369.t5 VNB.t14 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1008 ps=1.28 w=0.36 l=0.15
X15 VGND.t2 SCE.t2 a_299_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.1176 ps=1.4 w=0.42 l=0.15
X16 VGND.t5 a_1527_315.t4 a_1485_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X17 Q.t3 a_1527_315.t5 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_644_369.t1 a_299_47.t3 a_560_369.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1008 pd=0.955 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 a_661_47.t0 SCE.t3 a_560_369.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 VGND.t6 SCD.t1 a_661_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_560_369.t1 D.t0 a_466_369.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1024 ps=0.96 w=0.64 l=0.15
X22 a_560_369.t0 D.t1 a_487_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0504 ps=0.66 w=0.42 l=0.15
X23 VPWR.t3 a_1527_315.t6 Q.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1485_47.t0 a_27_47.t4 a_1356_413.t1 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X25 a_1033_413.t0 a_27_47.t5 a_940_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X26 a_193_47.t1 a_27_47.t6 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 a_1099_183.t2 a_940_413.t5 VPWR.t6 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X28 a_1440_413.t1 a_193_47.t4 a_1356_413.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X29 a_1037_47# a_193_47.t5 a_940_413.t2 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X30 VGND.t9 CLK.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_1356_413.t0 a_27_47.t7 a_1099_183.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X32 VGND.t3 a_1527_315.t7 Q.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_1527_315.n16 a_1527_315.t4 383.5
R1 a_1527_315.t0 a_1527_315.n17 324.885
R2 a_1527_315.n4 a_1527_315.t6 212.081
R3 a_1527_315.n3 a_1527_315.t2 212.081
R4 a_1527_315.n8 a_1527_315.n1 212.081
R5 a_1527_315.n12 a_1527_315.n10 212.081
R6 a_1527_315.n17 a_1527_315.n16 179.928
R7 a_1527_315.n6 a_1527_315.n5 169.409
R8 a_1527_315.n15 a_1527_315.t1 155.958
R9 a_1527_315.n14 a_1527_315.n13 152
R10 a_1527_315.n9 a_1527_315.n0 152
R11 a_1527_315.n7 a_1527_315.n6 152
R12 a_1527_315.n4 a_1527_315.t7 139.78
R13 a_1527_315.n3 a_1527_315.t5 139.78
R14 a_1527_315.n8 a_1527_315.n2 139.78
R15 a_1527_315.n12 a_1527_315.n11 139.78
R16 a_1527_315.n16 a_1527_315.t3 139.286
R17 a_1527_315.n13 a_1527_315.n9 49.6611
R18 a_1527_315.n8 a_1527_315.n7 46.7399
R19 a_1527_315.n5 a_1527_315.n3 33.5944
R20 a_1527_315.n15 a_1527_315.n14 32.7685
R21 a_1527_315.n5 a_1527_315.n4 27.752
R22 a_1527_315.n17 a_1527_315.n15 19.2372
R23 a_1527_315.n6 a_1527_315.n0 17.4085
R24 a_1527_315.n14 a_1527_315.n0 17.4085
R25 a_1527_315.n7 a_1527_315.n3 16.0672
R26 a_1527_315.n13 a_1527_315.n12 8.76414
R27 a_1527_315.n9 a_1527_315.n8 2.92171
R28 VPWR.n5 VPWR.t7 722.018
R29 VPWR.n20 VPWR.t1 717.543
R30 VPWR.n45 VPWR.n1 604.394
R31 VPWR.n3 VPWR.n2 600.128
R32 VPWR.n12 VPWR.t8 397.829
R33 VPWR.n13 VPWR.t3 357.522
R34 VPWR.n14 VPWR.t2 346.818
R35 VPWR.n27 VPWR.n9 320.976
R36 VPWR.n9 VPWR.t0 113.98
R37 VPWR.n1 VPWR.t4 41.5552
R38 VPWR.n1 VPWR.t5 41.5552
R39 VPWR.n2 VPWR.t9 41.5552
R40 VPWR.n2 VPWR.t10 41.5552
R41 VPWR.n9 VPWR.t6 35.4605
R42 VPWR.n44 VPWR.n43 34.6358
R43 VPWR.n21 VPWR.n10 34.6358
R44 VPWR.n25 VPWR.n10 34.6358
R45 VPWR.n26 VPWR.n25 34.6358
R46 VPWR.n28 VPWR.n7 34.6358
R47 VPWR.n32 VPWR.n7 34.6358
R48 VPWR.n33 VPWR.n32 34.6358
R49 VPWR.n34 VPWR.n33 34.6358
R50 VPWR.n38 VPWR.n37 34.6358
R51 VPWR.n39 VPWR.n38 34.6358
R52 VPWR.n15 VPWR.n14 33.8829
R53 VPWR.n19 VPWR.n12 31.2476
R54 VPWR.n37 VPWR.n5 29.7417
R55 VPWR.n20 VPWR.n19 29.3652
R56 VPWR.n15 VPWR.n12 24.4711
R57 VPWR.n39 VPWR.n3 24.0946
R58 VPWR.n45 VPWR.n44 22.5887
R59 VPWR.n43 VPWR.n3 20.3299
R60 VPWR.n28 VPWR.n27 20.3299
R61 VPWR.n21 VPWR.n20 16.9417
R62 VPWR.n27 VPWR.n26 14.3064
R63 VPWR.n16 VPWR.n15 9.3005
R64 VPWR.n17 VPWR.n12 9.3005
R65 VPWR.n19 VPWR.n18 9.3005
R66 VPWR.n20 VPWR.n11 9.3005
R67 VPWR.n22 VPWR.n21 9.3005
R68 VPWR.n23 VPWR.n10 9.3005
R69 VPWR.n25 VPWR.n24 9.3005
R70 VPWR.n26 VPWR.n8 9.3005
R71 VPWR.n29 VPWR.n28 9.3005
R72 VPWR.n30 VPWR.n7 9.3005
R73 VPWR.n32 VPWR.n31 9.3005
R74 VPWR.n33 VPWR.n6 9.3005
R75 VPWR.n35 VPWR.n34 9.3005
R76 VPWR.n37 VPWR.n36 9.3005
R77 VPWR.n38 VPWR.n4 9.3005
R78 VPWR.n40 VPWR.n39 9.3005
R79 VPWR.n41 VPWR.n3 9.3005
R80 VPWR.n43 VPWR.n42 9.3005
R81 VPWR.n44 VPWR.n0 9.3005
R82 VPWR.n14 VPWR.n13 7.85305
R83 VPWR.n46 VPWR.n45 7.14087
R84 VPWR.n34 VPWR.n5 4.89462
R85 VPWR.n16 VPWR.n13 0.649897
R86 VPWR.n46 VPWR.n0 0.148262
R87 VPWR.n17 VPWR.n16 0.120292
R88 VPWR.n18 VPWR.n17 0.120292
R89 VPWR.n18 VPWR.n11 0.120292
R90 VPWR.n22 VPWR.n11 0.120292
R91 VPWR.n23 VPWR.n22 0.120292
R92 VPWR.n24 VPWR.n23 0.120292
R93 VPWR.n24 VPWR.n8 0.120292
R94 VPWR.n29 VPWR.n8 0.120292
R95 VPWR.n30 VPWR.n29 0.120292
R96 VPWR.n31 VPWR.n30 0.120292
R97 VPWR.n31 VPWR.n6 0.120292
R98 VPWR.n35 VPWR.n6 0.120292
R99 VPWR.n36 VPWR.n35 0.120292
R100 VPWR.n36 VPWR.n4 0.120292
R101 VPWR.n40 VPWR.n4 0.120292
R102 VPWR.n41 VPWR.n40 0.120292
R103 VPWR.n42 VPWR.n41 0.120292
R104 VPWR.n42 VPWR.n0 0.120292
R105 VPWR VPWR.n46 0.115103
R106 Q Q.n0 238.727
R107 Q Q.n1 125.448
R108 Q.n0 Q.t0 26.5955
R109 Q.n0 Q.t1 26.5955
R110 Q.n1 Q.t2 24.9236
R111 Q.n1 Q.t3 24.9236
R112 VPB.t14 VPB.t8 784.269
R113 VPB.t7 VPB.t14 624.456
R114 VPB.t13 VPB.t2 600.779
R115 VPB.t9 VPB.t16 556.386
R116 VPB.t5 VPB.t12 390.654
R117 VPB.t3 VPB.t7 346.262
R118 VPB.t0 VPB.t5 284.113
R119 VPB.t12 VPB.t4 281.154
R120 VPB.t15 VPB.t1 278.193
R121 VPB.t2 VPB.t0 275.235
R122 VPB.t11 VPB.t13 275.235
R123 VPB.t8 VPB.t6 248.599
R124 VPB.t4 VPB.t3 248.599
R125 VPB.t1 VPB.t11 248.599
R126 VPB.t16 VPB.t15 248.599
R127 VPB.t10 VPB.t9 248.599
R128 VPB VPB.t10 145.017
R129 SCE.n2 SCE.t3 342.286
R130 SCE.n1 SCE.t2 321.772
R131 SCE.n2 SCE.n1 253.272
R132 SCE.n0 SCE.t0 236.18
R133 SCE.n0 SCE.t1 174.835
R134 SCE SCE.n2 20.1148
R135 SCE.n1 SCE.n0 8.76414
R136 a_466_369.t0 a_466_369.t1 98.5005
R137 a_193_47.t1 a_193_47.n3 424.863
R138 a_193_47.n0 a_193_47.t4 348.661
R139 a_193_47.n1 a_193_47.t3 344.252
R140 a_193_47.n1 a_193_47.t5 282.788
R141 a_193_47.n0 a_193_47.t2 271.262
R142 a_193_47.n3 a_193_47.t0 242.661
R143 a_193_47.n2 a_193_47.n0 19.4022
R144 a_193_47.n3 a_193_47.n2 12.5028
R145 a_193_47.n2 a_193_47.n1 9.3005
R146 a_1099_183.n4 a_1099_183.n3 674.014
R147 a_1099_183.n2 a_1099_183.t4 433.8
R148 a_1099_183.n3 a_1099_183.n0 218.13
R149 a_1099_183.n3 a_1099_183.n2 185.308
R150 a_1099_183.n2 a_1099_183.n1 128.1
R151 a_1099_183.n4 a_1099_183.t0 89.1195
R152 a_1099_183.n0 a_1099_183.t1 63.3338
R153 a_1099_183.t2 a_1099_183.n4 37.5243
R154 a_1099_183.n0 a_1099_183.t3 36.7713
R155 a_1356_413.n3 a_1356_413.n2 693.449
R156 a_1356_413.n2 a_1356_413.n0 249.922
R157 a_1356_413.n2 a_1356_413.n1 243.993
R158 a_1356_413.n0 a_1356_413.t4 212.081
R159 a_1356_413.n0 a_1356_413.t5 139.78
R160 a_1356_413.n1 a_1356_413.t2 73.3338
R161 a_1356_413.n3 a_1356_413.t3 63.3219
R162 a_1356_413.t0 a_1356_413.n3 63.3219
R163 a_1356_413.n1 a_1356_413.t1 48.3338
R164 VNB.t2 VNB.t6 3773.46
R165 VNB.t10 VNB.t15 3474.43
R166 VNB.t9 VNB.t14 2904.85
R167 VNB.t12 VNB.t4 2733.98
R168 VNB.t7 VNB.t2 2677.02
R169 VNB.t11 VNB.t8 1466.67
R170 VNB.t4 VNB.t13 1452.43
R171 VNB.t15 VNB.t11 1438.19
R172 VNB.t14 VNB.t10 1366.99
R173 VNB.t0 VNB.t3 1366.99
R174 VNB.t8 VNB.t7 1352.75
R175 VNB.t6 VNB.t5 1196.12
R176 VNB.t1 VNB.t12 1196.12
R177 VNB.t13 VNB.t0 1110.68
R178 VNB.t3 VNB.t9 1082.2
R179 VNB VNB.t1 683.495
R180 SCD.n0 SCD.t1 268.849
R181 SCD.n0 SCD.t0 236.716
R182 SCD SCD.n0 158.531
R183 a_644_369.t0 a_644_369.t1 96.9614
R184 a_299_47.t0 a_299_47.n1 636.33
R185 a_299_47.n0 a_299_47.t3 416.856
R186 a_299_47.n0 a_299_47.t2 382.026
R187 a_299_47.n1 a_299_47.t1 344.036
R188 a_299_47.n1 a_299_47.n0 29.4703
R189 a_560_369.n3 a_560_369.n2 706.601
R190 a_560_369.n2 a_560_369.t4 688.484
R191 a_560_369.n1 a_560_369.n0 300.577
R192 a_560_369.n1 a_560_369.t5 256.243
R193 a_560_369.n2 a_560_369.n1 72.2828
R194 a_560_369.n0 a_560_369.t0 54.2862
R195 a_560_369.n3 a_560_369.t3 41.5552
R196 a_560_369.t1 a_560_369.n3 41.5552
R197 a_560_369.n0 a_560_369.t2 40.0005
R198 a_940_413.n3 a_940_413.n2 693.048
R199 a_940_413.n2 a_940_413.n1 300.243
R200 a_940_413.n0 a_940_413.t4 226.541
R201 a_940_413.n0 a_940_413.t5 196.013
R202 a_940_413.n2 a_940_413.n0 168.738
R203 a_940_413.n3 a_940_413.t1 75.0481
R204 a_940_413.t0 a_940_413.n3 72.7029
R205 a_940_413.n1 a_940_413.t3 65.0005
R206 a_940_413.n1 a_940_413.t2 45.0005
R207 CLK.n0 CLK.t0 294.557
R208 CLK.n0 CLK.t1 209.403
R209 CLK CLK.n0 154.069
R210 a_27_47.n3 a_27_47.t3 501.817
R211 a_27_47.n2 a_27_47.t4 448.26
R212 a_27_47.t0 a_27_47.n5 390.067
R213 a_27_47.n1 a_27_47.t1 290.872
R214 a_27_47.n0 a_27_47.t6 263.173
R215 a_27_47.n2 a_27_47.t7 254.389
R216 a_27_47.n0 a_27_47.t2 227.826
R217 a_27_47.n4 a_27_47.n2 193.447
R218 a_27_47.n4 a_27_47.n3 166.708
R219 a_27_47.n1 a_27_47.n0 152
R220 a_27_47.n3 a_27_47.t5 148.35
R221 a_27_47.n5 a_27_47.n1 35.3396
R222 a_27_47.n5 a_27_47.n4 13.3063
R223 VGND.n11 VGND.t3 293.764
R224 VGND.n12 VGND.t4 279.055
R225 VGND.n6 VGND.t8 265.825
R226 VGND.n4 VGND.t6 255.184
R227 VGND.n10 VGND.t1 249.891
R228 VGND.n18 VGND.t5 239.139
R229 VGND.n43 VGND.n42 199.739
R230 VGND.n2 VGND.n1 198.964
R231 VGND.n1 VGND.t2 61.4291
R232 VGND.n1 VGND.t7 41.4291
R233 VGND.n42 VGND.t0 38.5719
R234 VGND.n42 VGND.t9 38.5719
R235 VGND.n17 VGND.n16 34.6358
R236 VGND.n22 VGND.n8 34.6358
R237 VGND.n23 VGND.n22 34.6358
R238 VGND.n24 VGND.n23 34.6358
R239 VGND.n29 VGND.n28 34.6358
R240 VGND.n30 VGND.n29 34.6358
R241 VGND.n35 VGND.n34 34.6358
R242 VGND.n36 VGND.n35 34.6358
R243 VGND.n41 VGND.n40 34.6358
R244 VGND.n13 VGND.n12 33.8829
R245 VGND.n28 VGND.n6 32.7534
R246 VGND.n13 VGND.n10 31.624
R247 VGND.n30 VGND.n4 30.4946
R248 VGND.n18 VGND.n17 29.3652
R249 VGND.n40 VGND.n2 27.4829
R250 VGND.n34 VGND.n4 23.7181
R251 VGND.n43 VGND.n41 22.9652
R252 VGND.n36 VGND.n2 16.9417
R253 VGND.n18 VGND.n8 12.0476
R254 VGND.n14 VGND.n13 9.3005
R255 VGND.n16 VGND.n15 9.3005
R256 VGND.n17 VGND.n9 9.3005
R257 VGND.n19 VGND.n18 9.3005
R258 VGND.n20 VGND.n8 9.3005
R259 VGND.n22 VGND.n21 9.3005
R260 VGND.n23 VGND.n7 9.3005
R261 VGND.n25 VGND.n24 9.3005
R262 VGND.n26 VGND.n6 9.3005
R263 VGND.n28 VGND.n27 9.3005
R264 VGND.n29 VGND.n5 9.3005
R265 VGND.n31 VGND.n30 9.3005
R266 VGND.n32 VGND.n4 9.3005
R267 VGND.n34 VGND.n33 9.3005
R268 VGND.n35 VGND.n3 9.3005
R269 VGND.n37 VGND.n36 9.3005
R270 VGND.n38 VGND.n2 9.3005
R271 VGND.n40 VGND.n39 9.3005
R272 VGND.n41 VGND.n0 9.3005
R273 VGND.n24 VGND.n6 8.65932
R274 VGND.n12 VGND.n11 7.85305
R275 VGND.n44 VGND.n43 7.12063
R276 VGND.n16 VGND.n10 3.01226
R277 VGND.n14 VGND.n11 0.649897
R278 VGND.n44 VGND.n0 0.148519
R279 VGND.n15 VGND.n14 0.120292
R280 VGND.n15 VGND.n9 0.120292
R281 VGND.n19 VGND.n9 0.120292
R282 VGND.n20 VGND.n19 0.120292
R283 VGND.n21 VGND.n20 0.120292
R284 VGND.n21 VGND.n7 0.120292
R285 VGND.n25 VGND.n7 0.120292
R286 VGND.n26 VGND.n25 0.120292
R287 VGND.n27 VGND.n26 0.120292
R288 VGND.n27 VGND.n5 0.120292
R289 VGND.n31 VGND.n5 0.120292
R290 VGND.n32 VGND.n31 0.120292
R291 VGND.n33 VGND.n32 0.120292
R292 VGND.n33 VGND.n3 0.120292
R293 VGND.n37 VGND.n3 0.120292
R294 VGND.n38 VGND.n37 0.120292
R295 VGND.n39 VGND.n38 0.120292
R296 VGND.n39 VGND.n0 0.120292
R297 VGND VGND.n44 0.114842
R298 a_487_47.t0 a_487_47.t1 68.5719
R299 a_1440_413.t0 a_1440_413.t1 204.036
R300 a_1033_413.t0 a_1033_413.t1 154.786
R301 a_1485_47.t1 a_1485_47.t0 93.0601
R302 a_661_47.t0 a_661_47.t1 65.7148
R303 D.n0 D.t1 321.87
R304 D.n0 D.t0 183.696
R305 D D.n0 158.207
C0 Q VGND 0.251251f
C1 SCD VPWR 0.010916f
C2 D VGND 0.00928f
C3 VPB Q 0.013373f
C4 VGND SCE 0.110929f
C5 VPB VGND 0.013912f
C6 D SCE 0.102564f
C7 VPB D 0.054539f
C8 VPB SCE 0.108437f
C9 a_1037_47# VGND 0.004185f
C10 Q VPWR 0.343459f
C11 VPWR VGND 0.098533f
C12 D VPWR 0.008006f
C13 VGND CLK 0.019316f
C14 VPWR SCE 0.025893f
C15 VPB VPWR 0.235851f
C16 VPB CLK 0.070163f
C17 VPWR CLK 0.019412f
C18 SCD VGND 0.010144f
C19 D SCD 0.006114f
C20 SCD SCE 0.046103f
C21 VPB SCD 0.067875f
C22 Q VNB 0.062104f
C23 VGND VNB 1.21529f
C24 VPWR VNB 1.00901f
C25 SCD VNB 0.122377f
C26 D VNB 0.101787f
C27 SCE VNB 0.241946f
C28 CLK VNB 0.195347f
C29 VPB VNB 2.19949f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdlclkp_1 VGND VPWR VPB VNB GCLK CLK GATE SCE
X0 a_1094_47.t0 a_464_315.t2 a_1012_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0861 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_464_315.t1 a_286_413.t4 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2533 pd=2.52 as=0.1838 ps=1.53 w=1 l=0.15
X2 a_464_315.t0 a_286_413.t5 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134375 ps=1.09 w=0.65 l=0.15
X3 VPWR.t6 CLK.t0 a_1012_47.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 a_1012_47.t0 a_464_315.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_109_369.t1 SCE.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 VPWR.t2 a_464_315.t4 a_382_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1838 pd=1.53 as=0.0924 ps=0.86 w=0.42 l=0.15
X7 a_382_413.t1 a_256_147.t2 a_286_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_286_413.t3 a_256_243.t2 a_27_47.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.11175 ps=1.015 w=0.42 l=0.15
X9 a_27_47.t2 GATE.t0 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.06705 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_256_147.t1 CLK.t1 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.16925 ps=1.37 w=0.64 l=0.15
X11 VGND.t5 a_256_147.t3 a_256_243.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 GCLK.t1 a_1012_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X13 a_27_47.t1 GATE.t1 a_109_369.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.11175 pd=1.015 as=0.0672 ps=0.85 w=0.64 l=0.15
X14 a_256_147.t0 CLK.t2 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 GCLK.t0 a_1012_47.t4 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X16 VPWR.t3 a_256_147.t4 a_256_243.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.16925 pd=1.37 as=0.1629 ps=1.8 w=0.64 l=0.15
X17 a_286_413.t2 a_256_147.t5 a_27_47.t0 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0675 pd=0.735 as=0.06705 ps=0.75 w=0.36 l=0.15
X18 VGND.t6 CLK.t3 a_1094_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0861 ps=0.83 w=0.42 l=0.15
X19 a_394_47.t1 a_256_243.t3 a_286_413.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0903 pd=0.88 as=0.0675 ps=0.735 w=0.36 l=0.15
X20 VGND.t2 a_464_315.t5 a_394_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.134375 pd=1.09 as=0.0903 ps=0.88 w=0.42 l=0.15
X21 VGND.t1 SCE.t1 a_27_47.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_464_315.n4 a_464_315.n3 602.456
R1 a_464_315.n1 a_464_315.t5 392.562
R2 a_464_315.n0 a_464_315.t2 321.772
R3 a_464_315.n2 a_464_315.t0 320.307
R4 a_464_315.n3 a_464_315.n0 302.832
R5 a_464_315.n2 a_464_315.n1 191.585
R6 a_464_315.n0 a_464_315.t3 183.599
R7 a_464_315.n4 a_464_315.t1 175.532
R8 a_464_315.n1 a_464_315.t4 148.35
R9 a_464_315.n5 a_464_315.n4 15.1543
R10 a_464_315.n3 a_464_315.n2 5.52777
R11 a_1012_47.n2 a_1012_47.n1 625.039
R12 a_1012_47.n1 a_1012_47.t1 334.692
R13 a_1012_47.n0 a_1012_47.t3 241.536
R14 a_1012_47.n0 a_1012_47.t4 169.237
R15 a_1012_47.n1 a_1012_47.n0 152
R16 a_1012_47.n2 a_1012_47.t2 41.5552
R17 a_1012_47.t0 a_1012_47.n2 41.5552
R18 a_1094_47.t0 a_1094_47.t1 117.144
R19 VNB.t10 VNB.t5 2677.02
R20 VNB.t3 VNB.t7 2677.02
R21 VNB.t0 VNB.t4 1737.22
R22 VNB.t4 VNB.t3 1680.26
R23 VNB.t5 VNB.t9 1594.82
R24 VNB.t8 VNB.t0 1495.15
R25 VNB.t6 VNB.t8 1366.99
R26 VNB.t9 VNB.t1 1352.75
R27 VNB.t7 VNB.t10 1196.12
R28 VNB.t2 VNB.t6 1196.12
R29 VNB VNB.t2 925.567
R30 a_286_413.n3 a_286_413.n2 679.722
R31 a_286_413.n2 a_286_413.n0 255.292
R32 a_286_413.n1 a_286_413.t4 232.472
R33 a_286_413.n2 a_286_413.n1 169.347
R34 a_286_413.n1 a_286_413.t5 160.173
R35 a_286_413.t1 a_286_413.n3 77.3934
R36 a_286_413.n3 a_286_413.t3 77.3934
R37 a_286_413.n0 a_286_413.t0 63.3338
R38 a_286_413.n0 a_286_413.t2 61.6672
R39 VPWR.n14 VPWR.n13 730.78
R40 VPWR.n6 VPWR.t1 717.596
R41 VPWR.n8 VPWR.n7 603.077
R42 VPWR.n21 VPWR.n20 585
R43 VPWR.n29 VPWR.t5 379.784
R44 VPWR.n20 VPWR.t2 136.024
R45 VPWR.n20 VPWR.t4 78.566
R46 VPWR.n13 VPWR.t7 61.563
R47 VPWR.n13 VPWR.t3 61.563
R48 VPWR.n7 VPWR.t6 50.7896
R49 VPWR.n7 VPWR.t0 39.301
R50 VPWR.n23 VPWR.n1 34.6358
R51 VPWR.n27 VPWR.n1 34.6358
R52 VPWR.n28 VPWR.n27 34.6358
R53 VPWR.n19 VPWR.n3 33.4806
R54 VPWR.n8 VPWR.n6 28.6118
R55 VPWR.n29 VPWR.n28 25.977
R56 VPWR.n23 VPWR.n22 25.3942
R57 VPWR.n15 VPWR.n3 17.4687
R58 VPWR.n11 VPWR.n5 10.706
R59 VPWR.n12 VPWR.n11 10.706
R60 VPWR.n15 VPWR.n14 9.30959
R61 VPWR.n9 VPWR.n5 9.3005
R62 VPWR.n11 VPWR.n10 9.3005
R63 VPWR.n12 VPWR.n4 9.3005
R64 VPWR.n16 VPWR.n15 9.3005
R65 VPWR.n17 VPWR.n3 9.3005
R66 VPWR.n19 VPWR.n18 9.3005
R67 VPWR.n22 VPWR.n2 9.3005
R68 VPWR.n24 VPWR.n23 9.3005
R69 VPWR.n25 VPWR.n1 9.3005
R70 VPWR.n27 VPWR.n26 9.3005
R71 VPWR.n28 VPWR.n0 9.3005
R72 VPWR.n30 VPWR.n29 9.3005
R73 VPWR.n22 VPWR.n21 4.5594
R74 VPWR.n21 VPWR.n19 3.50735
R75 VPWR.n9 VPWR.n8 1.93504
R76 VPWR.n14 VPWR.n12 1.39686
R77 VPWR.n6 VPWR.n5 0.815045
R78 VPWR.n10 VPWR.n9 0.120292
R79 VPWR.n10 VPWR.n4 0.120292
R80 VPWR.n16 VPWR.n4 0.120292
R81 VPWR.n17 VPWR.n16 0.120292
R82 VPWR.n18 VPWR.n17 0.120292
R83 VPWR.n18 VPWR.n2 0.120292
R84 VPWR.n24 VPWR.n2 0.120292
R85 VPWR.n25 VPWR.n24 0.120292
R86 VPWR.n26 VPWR.n25 0.120292
R87 VPWR.n26 VPWR.n0 0.120292
R88 VPWR.n30 VPWR.n0 0.120292
R89 VPWR VPWR.n30 0.0226354
R90 VPB.t10 VPB.t2 562.306
R91 VPB.t5 VPB.t3 550.467
R92 VPB.t1 VPB.t5 402.493
R93 VPB.t7 VPB.t1 349.221
R94 VPB.t3 VPB.t10 325.546
R95 VPB.t4 VPB.t9 310.748
R96 VPB.t9 VPB.t7 284.113
R97 VPB.t8 VPB.t0 281.154
R98 VPB.t2 VPB.t8 248.599
R99 VPB.t6 VPB.t4 213.084
R100 VPB VPB.t6 192.369
R101 VGND.n12 VGND.n11 203.923
R102 VGND.n5 VGND.n4 198.964
R103 VGND.n20 VGND.n19 198.964
R104 VGND.n7 VGND.n6 191.016
R105 VGND.n11 VGND.t2 65.7148
R106 VGND.n6 VGND.t0 41.6488
R107 VGND.n11 VGND.t4 41.2972
R108 VGND.n6 VGND.t6 38.5719
R109 VGND.n4 VGND.t7 38.5719
R110 VGND.n4 VGND.t5 38.5719
R111 VGND.n19 VGND.t3 38.5719
R112 VGND.n19 VGND.t1 38.5719
R113 VGND.n10 VGND.n3 34.6358
R114 VGND.n13 VGND.n1 34.6358
R115 VGND.n17 VGND.n1 34.6358
R116 VGND.n18 VGND.n17 34.6358
R117 VGND.n12 VGND.n10 33.1299
R118 VGND.n20 VGND.n18 22.9652
R119 VGND.n5 VGND.n3 12.8005
R120 VGND.n13 VGND.n12 10.1652
R121 VGND.n18 VGND.n0 9.3005
R122 VGND.n17 VGND.n16 9.3005
R123 VGND.n15 VGND.n1 9.3005
R124 VGND.n14 VGND.n13 9.3005
R125 VGND.n8 VGND.n3 9.3005
R126 VGND.n10 VGND.n9 9.3005
R127 VGND.n12 VGND.n2 9.3005
R128 VGND.n7 VGND.n5 7.4704
R129 VGND.n21 VGND.n20 7.12063
R130 VGND.n8 VGND.n7 0.173613
R131 VGND.n21 VGND.n0 0.148519
R132 VGND.n9 VGND.n8 0.120292
R133 VGND.n9 VGND.n2 0.120292
R134 VGND.n14 VGND.n2 0.120292
R135 VGND.n15 VGND.n14 0.120292
R136 VGND.n16 VGND.n15 0.120292
R137 VGND.n16 VGND.n0 0.120292
R138 VGND VGND.n21 0.114842
R139 CLK.n0 CLK.t0 333.498
R140 CLK.n3 CLK.n0 194.323
R141 CLK.n1 CLK.t1 182.816
R142 CLK.n0 CLK.t3 169.619
R143 CLK.n2 CLK.n1 152
R144 CLK.n1 CLK.t2 149.792
R145 CLK CLK.n3 9.30959
R146 CLK.n2 CLK 1.65211
R147 CLK.n3 CLK.n2 1.03276
R148 SCE.n0 SCE.t0 287.995
R149 SCE.n0 SCE.t1 194.809
R150 SCE.n1 SCE.n0 152
R151 SCE.n1 SCE 14.3064
R152 SCE SCE.n1 2.76128
R153 a_109_369.t0 a_109_369.t1 64.6411
R154 a_382_413.t0 a_382_413.t1 206.381
R155 a_256_147.t1 a_256_147.n3 738.269
R156 a_256_147.n2 a_256_147.t2 306.257
R157 a_256_147.n2 a_256_147.t5 295.997
R158 a_256_147.n1 a_256_147.t0 265.705
R159 a_256_147.n0 a_256_147.t3 215.732
R160 a_256_147.n0 a_256_147.t4 183.599
R161 a_256_147.n1 a_256_147.n0 157.648
R162 a_256_147.n3 a_256_147.n2 20.9724
R163 a_256_147.n3 a_256_147.n1 14.2694
R164 a_256_243.n2 a_256_243.n1 648.533
R165 a_256_243.n0 a_256_243.t2 553.23
R166 a_256_243.n1 a_256_243.t0 238.506
R167 a_256_243.n1 a_256_243.n0 177.364
R168 a_256_243.n2 a_256_243.t1 127.046
R169 a_256_243.n0 a_256_243.t3 122.642
R170 a_27_47.n2 a_27_47.n1 700.068
R171 a_27_47.n1 a_27_47.t3 255.688
R172 a_27_47.n1 a_27_47.n0 237.105
R173 a_27_47.n2 a_27_47.t4 89.1195
R174 a_27_47.n0 a_27_47.t0 65.0005
R175 a_27_47.t1 a_27_47.n2 62.589
R176 a_27_47.n0 a_27_47.t2 29.5347
R177 GATE.n0 GATE.t1 295.168
R178 GATE.n0 GATE.t0 201.982
R179 GATE GATE.n0 163.167
R180 GCLK.n0 GCLK.t1 353.795
R181 GCLK GCLK.t0 249.84
R182 GCLK.n0 GCLK 8.2361
R183 GCLK GCLK.n0 6.90173
R184 a_394_47.t0 a_394_47.t1 138.06
C0 GCLK VGND 0.057449f
C1 GATE VGND 0.018562f
C2 GCLK VPB 0.011021f
C3 VGND VPB 0.008877f
C4 GATE VPB 0.054737f
C5 CLK GCLK 0.003607f
C6 CLK VGND 0.041261f
C7 GCLK VPWR 0.0598f
C8 VPWR VGND 0.075584f
C9 GATE VPWR 0.01333f
C10 SCE VGND 0.017084f
C11 SCE GATE 0.102519f
C12 CLK VPB 0.133548f
C13 VPWR VPB 0.154292f
C14 SCE VPB 0.06429f
C15 CLK VPWR 0.039562f
C16 SCE VPWR 0.042528f
C17 GCLK VNB 0.09138f
C18 CLK VNB 0.285077f
C19 VGND VNB 0.769211f
C20 VPWR VNB 0.646415f
C21 GATE VNB 0.112247f
C22 SCE VNB 0.188734f
C23 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdlclkp_2 VGND VPWR VPB VNB SCE GATE CLK GCLK
X0 GCLK.t1 a_1020_47.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1 a_109_369.t1 SCE.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 a_465_315.t1 a_287_413.t4 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1838 ps=1.53 w=1 l=0.15
X3 a_257_147.t1 CLK.t0 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.16925 ps=1.37 w=0.64 l=0.15
X4 a_1102_47.t1 a_465_315.t2 a_1020_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t5 a_1020_47.t4 GCLK.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_287_413.t2 a_257_147.t2 a_27_47.t3 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0675 pd=0.735 as=0.0681 ps=0.755 w=0.36 l=0.15
X7 VGND.t6 a_257_147.t3 a_257_243.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR.t3 a_465_315.t3 a_383_413.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1838 pd=1.53 as=0.0924 ps=0.86 w=0.42 l=0.15
X9 VGND.t2 CLK.t1 a_1102_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.175 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_27_47.t1 GATE.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0681 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VPWR.t7 CLK.t2 a_1020_47.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 GCLK.t2 a_1020_47.t5 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.139 ps=1.175 w=0.65 l=0.15
X13 a_287_413.t1 a_257_243.t2 a_27_47.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.11335 ps=1.02 w=0.42 l=0.15
X14 a_383_413.t0 a_257_147.t4 a_287_413.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_257_147.t0 CLK.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_27_47.t0 GATE.t1 a_109_369.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.11335 pd=1.02 as=0.0672 ps=0.85 w=0.64 l=0.15
X17 VPWR.t8 a_257_147.t5 a_257_243.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.16925 pd=1.37 as=0.1664 ps=1.8 w=0.64 l=0.15
X18 a_1020_47.t1 a_465_315.t4 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X19 a_395_47.t0 a_257_243.t3 a_287_413.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0903 pd=0.88 as=0.0675 ps=0.735 w=0.36 l=0.15
X20 VGND.t7 a_465_315.t5 a_395_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.137625 pd=1.1 as=0.0903 ps=0.88 w=0.42 l=0.15
X21 VPWR.t1 a_1020_47.t6 GCLK.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND.t8 SCE.t1 a_27_47.t4 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 a_465_315.t0 a_287_413.t5 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.137625 ps=1.1 w=0.65 l=0.15
R0 a_1020_47.n3 a_1020_47.n2 625.039
R1 a_1020_47.n2 a_1020_47.t0 337.505
R2 a_1020_47.n0 a_1020_47.t6 212.081
R3 a_1020_47.n1 a_1020_47.t3 212.081
R4 a_1020_47.n2 a_1020_47.n1 160.034
R5 a_1020_47.n0 a_1020_47.t4 139.78
R6 a_1020_47.n1 a_1020_47.t5 139.78
R7 a_1020_47.n1 a_1020_47.n0 61.346
R8 a_1020_47.n3 a_1020_47.t2 41.5552
R9 a_1020_47.t1 a_1020_47.n3 41.5552
R10 VPWR.n17 VPWR.n16 730.78
R11 VPWR.n9 VPWR.t4 717.596
R12 VPWR.n8 VPWR.n7 598.965
R13 VPWR.n24 VPWR.n23 585
R14 VPWR.n32 VPWR.t0 379.784
R15 VPWR.n6 VPWR.t1 255.738
R16 VPWR.n23 VPWR.t3 136.024
R17 VPWR.n23 VPWR.t5 78.566
R18 VPWR.n16 VPWR.t6 61.563
R19 VPWR.n16 VPWR.t8 61.563
R20 VPWR.n7 VPWR.t7 50.7896
R21 VPWR.n7 VPWR.t2 39.301
R22 VPWR.n26 VPWR.n1 34.6358
R23 VPWR.n30 VPWR.n1 34.6358
R24 VPWR.n31 VPWR.n30 34.6358
R25 VPWR.n22 VPWR.n3 33.1918
R26 VPWR.n32 VPWR.n31 25.977
R27 VPWR.n26 VPWR.n25 25.683
R28 VPWR.n10 VPWR.n8 24.0946
R29 VPWR.n10 VPWR.n9 20.4052
R30 VPWR.n18 VPWR.n3 17.2086
R31 VPWR.n14 VPWR.n5 10.706
R32 VPWR.n15 VPWR.n14 10.706
R33 VPWR.n18 VPWR.n17 10.4732
R34 VPWR.n11 VPWR.n10 9.3005
R35 VPWR.n12 VPWR.n5 9.3005
R36 VPWR.n14 VPWR.n13 9.3005
R37 VPWR.n15 VPWR.n4 9.3005
R38 VPWR.n19 VPWR.n18 9.3005
R39 VPWR.n20 VPWR.n3 9.3005
R40 VPWR.n22 VPWR.n21 9.3005
R41 VPWR.n25 VPWR.n2 9.3005
R42 VPWR.n27 VPWR.n26 9.3005
R43 VPWR.n28 VPWR.n1 9.3005
R44 VPWR.n30 VPWR.n29 9.3005
R45 VPWR.n31 VPWR.n0 9.3005
R46 VPWR.n33 VPWR.n32 9.3005
R47 VPWR.n8 VPWR.n6 6.44399
R48 VPWR.n25 VPWR.n24 4.64707
R49 VPWR.n24 VPWR.n22 3.41968
R50 VPWR.n9 VPWR.n5 1.74595
R51 VPWR.n11 VPWR.n6 0.646455
R52 VPWR.n17 VPWR.n15 0.233227
R53 VPWR.n12 VPWR.n11 0.120292
R54 VPWR.n13 VPWR.n12 0.120292
R55 VPWR.n13 VPWR.n4 0.120292
R56 VPWR.n19 VPWR.n4 0.120292
R57 VPWR.n20 VPWR.n19 0.120292
R58 VPWR.n21 VPWR.n20 0.120292
R59 VPWR.n21 VPWR.n2 0.120292
R60 VPWR.n27 VPWR.n2 0.120292
R61 VPWR.n28 VPWR.n27 0.120292
R62 VPWR.n29 VPWR.n28 0.120292
R63 VPWR.n29 VPWR.n0 0.120292
R64 VPWR.n33 VPWR.n0 0.120292
R65 VPWR VPWR.n33 0.0213333
R66 GCLK.n0 GCLK 586.423
R67 GCLK.n1 GCLK.n0 585
R68 GCLK GCLK.n2 185.238
R69 GCLK.n3 GCLK 36.2811
R70 GCLK.n3 GCLK 27.3016
R71 GCLK.n0 GCLK.t0 26.5955
R72 GCLK.n0 GCLK.t1 26.5955
R73 GCLK.n2 GCLK.t3 24.9236
R74 GCLK.n2 GCLK.t2 24.9236
R75 GCLK GCLK.n3 17.2313
R76 GCLK.n1 GCLK 14.6968
R77 GCLK GCLK.n1 1.42272
R78 VPB.t7 VPB.t11 577.104
R79 VPB.t8 VPB.t5 556.386
R80 VPB.t4 VPB.t7 402.493
R81 VPB.t10 VPB.t4 349.221
R82 VPB.t11 VPB.t8 325.546
R83 VPB.t1 VPB.t6 313.707
R84 VPB.t6 VPB.t10 284.113
R85 VPB.t9 VPB.t3 281.154
R86 VPB.t3 VPB.t2 248.599
R87 VPB.t5 VPB.t9 248.599
R88 VPB.t0 VPB.t1 213.084
R89 VPB VPB.t0 189.409
R90 SCE.n0 SCE.t0 287.995
R91 SCE.n0 SCE.t1 194.809
R92 SCE.n1 SCE.n0 152
R93 SCE.n1 SCE 14.3064
R94 SCE SCE.n1 2.76128
R95 a_109_369.t0 a_109_369.t1 64.6411
R96 a_287_413.n3 a_287_413.n2 679.722
R97 a_287_413.n2 a_287_413.n0 255.292
R98 a_287_413.n1 a_287_413.t4 232.472
R99 a_287_413.n2 a_287_413.n1 169.347
R100 a_287_413.n1 a_287_413.t5 160.173
R101 a_287_413.n3 a_287_413.t3 77.3934
R102 a_287_413.t1 a_287_413.n3 77.3934
R103 a_287_413.n0 a_287_413.t0 63.3338
R104 a_287_413.n0 a_287_413.t2 61.6672
R105 a_465_315.t1 a_465_315.n3 763.62
R106 a_465_315.n1 a_465_315.t5 392.562
R107 a_465_315.n0 a_465_315.t2 321.772
R108 a_465_315.n2 a_465_315.t0 320.307
R109 a_465_315.n3 a_465_315.n0 305.466
R110 a_465_315.n2 a_465_315.n1 191.585
R111 a_465_315.n0 a_465_315.t4 183.599
R112 a_465_315.n1 a_465_315.t3 148.35
R113 a_465_315.n3 a_465_315.n2 5.52777
R114 CLK.n0 CLK.t2 333.498
R115 CLK.n3 CLK.n0 196.181
R116 CLK.n1 CLK.t0 182.816
R117 CLK.n0 CLK.t1 169.619
R118 CLK.n2 CLK.n1 152
R119 CLK.n1 CLK.t3 146.172
R120 CLK CLK.n3 9.30959
R121 CLK.n2 CLK 1.65211
R122 CLK.n3 CLK.n2 1.03276
R123 a_257_147.t1 a_257_147.n3 741.66
R124 a_257_147.n2 a_257_147.t4 306.257
R125 a_257_147.n2 a_257_147.t2 295.997
R126 a_257_147.n1 a_257_147.t0 268.442
R127 a_257_147.n0 a_257_147.t3 215.732
R128 a_257_147.n0 a_257_147.t5 183.599
R129 a_257_147.n1 a_257_147.n0 158.776
R130 a_257_147.n3 a_257_147.n2 20.9635
R131 a_257_147.n3 a_257_147.n1 17.0642
R132 a_1102_47.t0 a_1102_47.t1 60.0005
R133 VNB.t2 VNB.t10 2748.22
R134 VNB.t1 VNB.t7 2677.02
R135 VNB.t3 VNB.t5 1922.33
R136 VNB.t0 VNB.t9 1737.22
R137 VNB.t9 VNB.t1 1708.74
R138 VNB.t8 VNB.t0 1495.15
R139 VNB.t4 VNB.t8 1381.23
R140 VNB.t5 VNB.t6 1196.12
R141 VNB.t7 VNB.t2 1196.12
R142 VNB.t11 VNB.t4 1196.12
R143 VNB.t10 VNB.t3 1025.24
R144 VNB VNB.t11 911.327
R145 VGND.n20 VGND.n19 203.923
R146 VGND.n14 VGND.n13 198.964
R147 VGND.n28 VGND.n27 198.964
R148 VGND.n7 VGND.n6 185
R149 VGND.n8 VGND.t5 161.135
R150 VGND.n6 VGND.t2 78.5719
R151 VGND.n19 VGND.t7 65.7148
R152 VGND.n6 VGND.t4 58.7917
R153 VGND.n19 VGND.t0 43.6488
R154 VGND.n13 VGND.t1 38.5719
R155 VGND.n13 VGND.t6 38.5719
R156 VGND.n27 VGND.t3 38.5719
R157 VGND.n27 VGND.t8 38.5719
R158 VGND.n12 VGND.n11 34.6358
R159 VGND.n18 VGND.n3 34.6358
R160 VGND.n21 VGND.n1 34.6358
R161 VGND.n25 VGND.n1 34.6358
R162 VGND.n26 VGND.n25 34.6358
R163 VGND.n20 VGND.n18 32.7534
R164 VGND.n14 VGND.n12 30.4946
R165 VGND.n28 VGND.n26 22.9652
R166 VGND.n11 VGND.n5 21.3386
R167 VGND.n14 VGND.n3 13.9299
R168 VGND.n21 VGND.n20 10.5417
R169 VGND.n7 VGND.n5 9.54012
R170 VGND.n26 VGND.n0 9.3005
R171 VGND.n25 VGND.n24 9.3005
R172 VGND.n23 VGND.n1 9.3005
R173 VGND.n22 VGND.n21 9.3005
R174 VGND.n9 VGND.n5 9.3005
R175 VGND.n11 VGND.n10 9.3005
R176 VGND.n12 VGND.n4 9.3005
R177 VGND.n15 VGND.n14 9.3005
R178 VGND.n16 VGND.n3 9.3005
R179 VGND.n18 VGND.n17 9.3005
R180 VGND.n20 VGND.n2 9.3005
R181 VGND.n8 VGND.n7 8.32828
R182 VGND.n29 VGND.n28 7.12063
R183 VGND.n9 VGND.n8 0.588593
R184 VGND.n29 VGND.n0 0.148519
R185 VGND.n10 VGND.n9 0.120292
R186 VGND.n10 VGND.n4 0.120292
R187 VGND.n15 VGND.n4 0.120292
R188 VGND.n16 VGND.n15 0.120292
R189 VGND.n17 VGND.n16 0.120292
R190 VGND.n17 VGND.n2 0.120292
R191 VGND.n22 VGND.n2 0.120292
R192 VGND.n23 VGND.n22 0.120292
R193 VGND.n24 VGND.n23 0.120292
R194 VGND.n24 VGND.n0 0.120292
R195 VGND VGND.n29 0.11354
R196 a_27_47.n2 a_27_47.n1 704.529
R197 a_27_47.n1 a_27_47.t4 256.065
R198 a_27_47.n1 a_27_47.n0 236.159
R199 a_27_47.n2 a_27_47.t2 89.1195
R200 a_27_47.n0 a_27_47.t3 66.6672
R201 a_27_47.t0 a_27_47.n2 64.9343
R202 a_27_47.n0 a_27_47.t1 28.3186
R203 a_257_243.t1 a_257_243.n1 785.082
R204 a_257_243.n0 a_257_243.t2 553.23
R205 a_257_243.n1 a_257_243.t0 237.651
R206 a_257_243.n1 a_257_243.n0 176.602
R207 a_257_243.n0 a_257_243.t3 122.642
R208 a_383_413.t0 a_383_413.t1 206.381
R209 GATE.n0 GATE.t1 294.774
R210 GATE.n0 GATE.t0 201.587
R211 GATE GATE.n0 162.73
R212 a_395_47.t1 a_395_47.t0 138.06
C0 CLK VPB 0.134874f
C1 SCE VPB 0.06429f
C2 SCE GATE 0.102519f
C3 VPWR VGND 0.08704f
C4 GCLK VGND 0.137495f
C5 VGND VPB 0.009443f
C6 GATE VGND 0.018598f
C7 CLK VGND 0.044657f
C8 GCLK VPWR 0.166738f
C9 VPWR VPB 0.17067f
C10 GATE VPWR 0.013473f
C11 SCE VGND 0.017029f
C12 GCLK VPB 0.005504f
C13 GATE VPB 0.055386f
C14 CLK VPWR 0.040381f
C15 CLK GCLK 0.003098f
C16 SCE VPWR 0.041218f
C17 GCLK VNB 0.027777f
C18 CLK VNB 0.281327f
C19 VGND VNB 0.841702f
C20 VPWR VNB 0.717826f
C21 GATE VNB 0.112864f
C22 SCE VNB 0.188734f
C23 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdlclkp_4 VGND VPWR VPB VNB GCLK CLK GATE SCE
X0 a_257_147.t1 CLK.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.16925 ps=1.37 w=0.64 l=0.15
X1 a_109_369.t1 SCE.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 a_465_315.t1 a_287_413.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1838 ps=1.53 w=1 l=0.15
X3 VPWR.t8 a_1045_47# GCLK.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t0 a_257_147.t2 a_257_243.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.16925 pd=1.37 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 GCLK.t2 a_1045_47# VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_287_413.t2 a_257_147.t3 a_27_47.t1 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0675 pd=0.735 as=0.0681 ps=0.755 w=0.36 l=0.15
X7 VGND.t1 a_257_147.t4 a_257_243.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND.t6 a_1045_47# GCLK.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t1 a_465_315.t2 a_383_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1838 pd=1.53 as=0.0924 ps=0.86 w=0.42 l=0.15
X10 VPWR.t6 a_1045_47# GCLK.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47.t2 GATE.t0 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0681 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 GCLK.t0 a_1045_47# VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X13 a_287_413.t3 a_257_243.t2 a_27_47.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.11335 ps=1.02 w=0.42 l=0.15
X14 a_383_413.t0 a_257_147.t5 a_287_413.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 VGND CLK a_1127_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.06825 ps=0.86 w=0.65 l=0.15
X16 a_257_147.t0 CLK.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 GCLK.t6 a_1045_47# VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X18 GCLK.t5 a_1045_47# VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_47.t0 GATE.t1 a_109_369.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.11335 pd=1.02 as=0.0672 ps=0.85 w=0.64 l=0.15
X20 VPWR CLK a_1045_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND.t3 a_1045_47# GCLK.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_395_47.t0 a_257_243.t3 a_287_413.t0 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0903 pd=0.88 as=0.0675 ps=0.735 w=0.36 l=0.15
X23 VGND.t9 a_465_315.t3 a_395_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.137625 pd=1.1 as=0.0903 ps=0.88 w=0.42 l=0.15
X24 VGND.t8 SCE.t1 a_27_47.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_465_315.t0 a_287_413.t5 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.137625 ps=1.1 w=0.65 l=0.15
R0 CLK.n2 CLK.n0 241.536
R1 CLK.n3 CLK.t0 182.816
R2 CLK.n4 CLK.n2 180.26
R3 CLK.n2 CLK.n1 169.237
R4 CLK.n4 CLK.n3 152
R5 CLK.n3 CLK.t1 149.792
R6 CLK CLK.n4 1.55202
R7 VPWR.n12 VPWR.t5 826.271
R8 VPWR.n20 VPWR.n19 730.78
R9 VPWR.n27 VPWR.n26 585
R10 VPWR.n35 VPWR.t2 379.784
R11 VPWR.n8 VPWR.n7 316.245
R12 VPWR.n9 VPWR.t8 261.925
R13 VPWR.n26 VPWR.t1 136.024
R14 VPWR.n26 VPWR.t3 78.566
R15 VPWR.n19 VPWR.t4 61.563
R16 VPWR.n19 VPWR.t0 61.563
R17 VPWR.n29 VPWR.n1 34.6358
R18 VPWR.n33 VPWR.n1 34.6358
R19 VPWR.n34 VPWR.n33 34.6358
R20 VPWR.n25 VPWR.n3 33.1918
R21 VPWR.n7 VPWR.t7 26.5955
R22 VPWR.n7 VPWR.t6 26.5955
R23 VPWR.n35 VPWR.n34 25.977
R24 VPWR.n29 VPWR.n28 25.683
R25 VPWR.n11 VPWR.n8 24.8476
R26 VPWR.n13 VPWR.n12 22.9652
R27 VPWR.n13 VPWR.n5 22.931
R28 VPWR.n12 VPWR.n11 21.4593
R29 VPWR.n21 VPWR.n3 18.2491
R30 VPWR.n17 VPWR.n5 10.706
R31 VPWR.n18 VPWR.n17 10.706
R32 VPWR.n21 VPWR.n20 9.65868
R33 VPWR.n11 VPWR.n10 9.3005
R34 VPWR.n12 VPWR.n6 9.3005
R35 VPWR.n14 VPWR.n13 9.3005
R36 VPWR.n15 VPWR.n5 9.3005
R37 VPWR.n17 VPWR.n16 9.3005
R38 VPWR.n18 VPWR.n4 9.3005
R39 VPWR.n22 VPWR.n21 9.3005
R40 VPWR.n23 VPWR.n3 9.3005
R41 VPWR.n25 VPWR.n24 9.3005
R42 VPWR.n28 VPWR.n2 9.3005
R43 VPWR.n30 VPWR.n29 9.3005
R44 VPWR.n31 VPWR.n1 9.3005
R45 VPWR.n33 VPWR.n32 9.3005
R46 VPWR.n34 VPWR.n0 9.3005
R47 VPWR.n36 VPWR.n35 9.3005
R48 VPWR.n9 VPWR.n8 6.75922
R49 VPWR.n28 VPWR.n27 4.64707
R50 VPWR.n27 VPWR.n25 3.41968
R51 VPWR.n20 VPWR.n18 1.04777
R52 VPWR.n10 VPWR.n9 0.614355
R53 VPWR.n10 VPWR.n6 0.120292
R54 VPWR.n14 VPWR.n6 0.120292
R55 VPWR.n15 VPWR.n14 0.120292
R56 VPWR.n16 VPWR.n15 0.120292
R57 VPWR.n16 VPWR.n4 0.120292
R58 VPWR.n22 VPWR.n4 0.120292
R59 VPWR.n23 VPWR.n22 0.120292
R60 VPWR.n24 VPWR.n23 0.120292
R61 VPWR.n24 VPWR.n2 0.120292
R62 VPWR.n30 VPWR.n2 0.120292
R63 VPWR.n31 VPWR.n30 0.120292
R64 VPWR.n32 VPWR.n31 0.120292
R65 VPWR.n32 VPWR.n0 0.120292
R66 VPWR.n36 VPWR.n0 0.120292
R67 VPWR VPWR.n36 0.0213333
R68 a_257_147.t1 a_257_147.n3 738.269
R69 a_257_147.n2 a_257_147.t5 306.257
R70 a_257_147.n2 a_257_147.t3 295.997
R71 a_257_147.n1 a_257_147.t0 265.705
R72 a_257_147.n0 a_257_147.t4 215.732
R73 a_257_147.n0 a_257_147.t2 183.599
R74 a_257_147.n1 a_257_147.n0 157.648
R75 a_257_147.n3 a_257_147.n2 20.9813
R76 a_257_147.n3 a_257_147.n1 14.2694
R77 VPB.t4 VPB.t7 1097.97
R78 VPB.t3 VPB.t6 556.386
R79 VPB.t1 VPB.t3 402.493
R80 VPB.t5 VPB.t1 349.221
R81 VPB.t6 VPB.t4 325.546
R82 VPB.t0 VPB.t11 313.707
R83 VPB.t11 VPB.t5 284.113
R84 VPB.t9 VPB.t10 248.599
R85 VPB.t8 VPB.t9 248.599
R86 VPB.t7 VPB.t8 248.599
R87 VPB.t2 VPB.t0 213.084
R88 VPB VPB.t2 189.409
R89 SCE.n0 SCE.t0 288.204
R90 SCE.n0 SCE.t1 195.017
R91 SCE.n1 SCE.n0 152
R92 SCE.n1 SCE 14.0313
R93 SCE SCE.n1 2.70819
R94 a_109_369.t0 a_109_369.t1 64.6411
R95 a_287_413.n3 a_287_413.n2 679.722
R96 a_287_413.n2 a_287_413.n0 255.292
R97 a_287_413.n1 a_287_413.t4 232.472
R98 a_287_413.n2 a_287_413.n1 169.347
R99 a_287_413.n1 a_287_413.t5 160.173
R100 a_287_413.t1 a_287_413.n3 77.3934
R101 a_287_413.n3 a_287_413.t3 77.3934
R102 a_287_413.n0 a_287_413.t0 63.3338
R103 a_287_413.n0 a_287_413.t2 61.6672
R104 a_465_315.t1 a_465_315.n5 763.62
R105 a_465_315.n3 a_465_315.t3 392.562
R106 a_465_315.n4 a_465_315.t0 320.307
R107 a_465_315.n5 a_465_315.n2 315.238
R108 a_465_315.n2 a_465_315.n0 233.01
R109 a_465_315.n4 a_465_315.n3 191.585
R110 a_465_315.n2 a_465_315.n1 160.709
R111 a_465_315.n3 a_465_315.t2 148.35
R112 a_465_315.n5 a_465_315.n4 5.52777
R113 GCLK.n0 GCLK 586.537
R114 GCLK.n1 GCLK.n0 585
R115 GCLK.n5 GCLK.n4 289.55
R116 GCLK GCLK.n7 199.72
R117 GCLK GCLK.n2 188.328
R118 GCLK.n3 GCLK 54.9652
R119 GCLK.n3 GCLK 46.7732
R120 GCLK.n0 GCLK.t1 26.5955
R121 GCLK.n0 GCLK.t0 26.5955
R122 GCLK.n4 GCLK.t3 26.5955
R123 GCLK.n4 GCLK.t2 26.5955
R124 GCLK.n2 GCLK.t7 24.9236
R125 GCLK.n2 GCLK.t6 24.9236
R126 GCLK.n7 GCLK.t4 24.9236
R127 GCLK.n7 GCLK.t5 24.9236
R128 GCLK.n1 GCLK 15.8725
R129 GCLK.n6 GCLK 14.2774
R130 GCLK.n6 GCLK.n3 14.0313
R131 GCLK.n6 GCLK 11.0938
R132 GCLK GCLK.n5 7.81334
R133 GCLK.n5 GCLK 6.54763
R134 GCLK GCLK.n6 3.41383
R135 GCLK.n3 GCLK 2.21588
R136 GCLK GCLK.n1 1.5365
R137 a_257_243.t1 a_257_243.n1 781.129
R138 a_257_243.n0 a_257_243.t2 553.23
R139 a_257_243.n1 a_257_243.t0 238.506
R140 a_257_243.n1 a_257_243.n0 177.374
R141 a_257_243.n0 a_257_243.t3 122.642
R142 a_27_47.n2 a_27_47.n1 704.529
R143 a_27_47.n1 a_27_47.t3 256.065
R144 a_27_47.n1 a_27_47.n0 236.159
R145 a_27_47.n2 a_27_47.t4 89.1195
R146 a_27_47.n0 a_27_47.t1 66.6672
R147 a_27_47.t0 a_27_47.n2 64.9343
R148 a_27_47.n0 a_27_47.t2 28.3186
R149 VNB.t0 VNB.t6 5653.07
R150 VNB.t3 VNB.t1 2677.02
R151 VNB.t10 VNB.t11 1737.22
R152 VNB.t11 VNB.t3 1708.74
R153 VNB.t2 VNB.t10 1495.15
R154 VNB.t8 VNB.t2 1381.23
R155 VNB.t5 VNB.t4 1196.12
R156 VNB.t7 VNB.t5 1196.12
R157 VNB.t6 VNB.t7 1196.12
R158 VNB.t1 VNB.t0 1196.12
R159 VNB.t9 VNB.t8 1196.12
R160 VNB VNB.t9 911.327
R161 VGND.n11 VGND.t5 224.692
R162 VGND.n9 VGND.n8 204.457
R163 VGND.n25 VGND.n24 203.923
R164 VGND.n19 VGND.n18 198.964
R165 VGND.n33 VGND.n32 198.964
R166 VGND.n7 VGND.t3 152.817
R167 VGND.n24 VGND.t9 65.7148
R168 VGND.n24 VGND.t2 43.6488
R169 VGND.n18 VGND.t0 38.5719
R170 VGND.n18 VGND.t1 38.5719
R171 VGND.n32 VGND.t7 38.5719
R172 VGND.n32 VGND.t8 38.5719
R173 VGND.n17 VGND.n16 34.6358
R174 VGND.n23 VGND.n3 34.6358
R175 VGND.n26 VGND.n1 34.6358
R176 VGND.n30 VGND.n1 34.6358
R177 VGND.n31 VGND.n30 34.6358
R178 VGND.n25 VGND.n23 32.7534
R179 VGND.n19 VGND.n17 30.4946
R180 VGND.n12 VGND.n10 28.4986
R181 VGND.n16 VGND.n5 27.22
R182 VGND.n8 VGND.t4 24.9236
R183 VGND.n8 VGND.t6 24.9236
R184 VGND.n10 VGND.n9 24.8476
R185 VGND.n33 VGND.n31 22.9652
R186 VGND.n19 VGND.n3 13.9299
R187 VGND.n26 VGND.n25 10.5417
R188 VGND.n11 VGND.n5 10.0231
R189 VGND.n31 VGND.n0 9.3005
R190 VGND.n30 VGND.n29 9.3005
R191 VGND.n28 VGND.n1 9.3005
R192 VGND.n27 VGND.n26 9.3005
R193 VGND.n10 VGND.n6 9.3005
R194 VGND.n13 VGND.n12 9.3005
R195 VGND.n14 VGND.n5 9.3005
R196 VGND.n16 VGND.n15 9.3005
R197 VGND.n17 VGND.n4 9.3005
R198 VGND.n20 VGND.n19 9.3005
R199 VGND.n21 VGND.n3 9.3005
R200 VGND.n23 VGND.n22 9.3005
R201 VGND.n25 VGND.n2 9.3005
R202 VGND.n34 VGND.n33 7.12063
R203 VGND.n9 VGND.n7 6.75922
R204 VGND.n12 VGND.n11 1.08729
R205 VGND.n7 VGND.n6 0.614355
R206 VGND.n34 VGND.n0 0.148519
R207 VGND.n13 VGND.n6 0.120292
R208 VGND.n14 VGND.n13 0.120292
R209 VGND.n15 VGND.n14 0.120292
R210 VGND.n15 VGND.n4 0.120292
R211 VGND.n20 VGND.n4 0.120292
R212 VGND.n21 VGND.n20 0.120292
R213 VGND.n22 VGND.n21 0.120292
R214 VGND.n22 VGND.n2 0.120292
R215 VGND.n27 VGND.n2 0.120292
R216 VGND.n28 VGND.n27 0.120292
R217 VGND.n29 VGND.n28 0.120292
R218 VGND.n29 VGND.n0 0.120292
R219 VGND VGND.n34 0.11354
R220 a_383_413.t0 a_383_413.t1 206.381
R221 GATE.n0 GATE.t1 294.774
R222 GATE.n0 GATE.t0 201.587
R223 GATE GATE.n0 162.73
R224 a_395_47.t1 a_395_47.t0 138.06
C0 SCE CLK 1.15e-19
C1 GATE VGND 0.018598f
C2 GATE VPB 0.055386f
C3 GCLK CLK 0.002897f
C4 VGND CLK 0.083363f
C5 SCE VGND 0.017037f
C6 VPB CLK 0.105897f
C7 a_1127_47# CLK 0.001439f
C8 VPB SCE 0.064109f
C9 a_1045_47# CLK 0.191018f
C10 GCLK VGND 0.281161f
C11 GCLK VPB 0.010832f
C12 GCLK a_1127_47# 5.98e-19
C13 VPB VGND 0.007288f
C14 a_1045_47# GCLK 0.326708f
C15 a_1127_47# VGND 0.004506f
C16 a_1045_47# VGND 0.222214f
C17 a_1045_47# VPB 0.127717f
C18 a_1045_47# a_1127_47# 0.004638f
C19 GATE VPWR 0.013473f
C20 VPWR CLK 0.075636f
C21 VPWR SCE 0.041572f
C22 GCLK VPWR 0.355598f
C23 VPWR VGND 0.082222f
C24 GATE CLK 1.41e-19
C25 GATE SCE 0.102519f
C26 VPWR VPB 0.187575f
C27 a_1127_47# VPWR 1.88e-20
C28 a_1045_47# VPWR 0.193241f
C29 GCLK VNB 0.038644f
C30 CLK VNB 0.256336f
C31 VGND VNB 0.934457f
C32 VPWR VNB 0.789477f
C33 GATE VNB 0.112864f
C34 SCE VNB 0.188314f
C35 VPB VNB 1.66792f
C36 a_1045_47# VNB 0.404271f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxbp_1 VPWR VGND CLK SCD DE Q D Q_N SCE VPB VNB
X0 a_381_369.t1 D.t0 a_299_47.t5 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_2177_47# a_27_47.t2 a_2051_413.t1 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2 a_1537_413.t1 a_27_47.t3 a_1446_413.t3 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 VPWR.t6 DE.t0 a_423_343.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VPWR.t9 CLK.t0 a_27_47.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t3 SCE.t0 a_885_21.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1264 pd=1.035 as=0.1696 ps=1.81 w=0.64 l=0.15
X6 Q.t1 a_2051_413.t2 VGND.t11 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10025 ps=0.985 w=0.65 l=0.15
X7 VGND.t6 SCE.t1 a_885_21.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 Q_N.t1 a_791_264.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9 VPWR.t1 a_1610_159.t2 a_1537_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_1610_159.t0 a_1446_413.t4 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X11 VGND.t8 DE.t1 a_423_343.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_1561_47# a_193_47.t2 a_1446_413.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X13 a_1974_47.t0 a_1610_159.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_193_47.t1 a_27_47.t4 VGND.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_729_47.t0 a_423_343.t2 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X16 Q_N.t0 a_791_264.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14575 ps=1.335 w=1 l=0.15
X17 a_729_369.t1 DE.t2 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X18 Q.t0 a_2051_413.t3 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.154 ps=1.335 w=1 l=0.15
X19 a_299_47.t0 a_791_264.t4 a_729_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0756 ps=0.78 w=0.42 l=0.15
X20 a_2135_413.t0 a_193_47.t3 a_2051_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 a_1446_413.t2 a_27_47.t5 a_915_47# VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.22515 ps=1.505 w=0.36 l=0.15
X22 a_193_47.t0 a_27_47.t6 VPWR.t4 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_1231_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1056 pd=0.97 as=0.1264 ps=1.035 w=0.64 l=0.15
X24 a_915_47# SCE.t2 a_1226_119.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.22515 pd=1.505 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 VPWR.t10 a_2051_413.t4 a_791_264.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1728 ps=1.82 w=0.64 l=0.15
X26 a_299_47.t1 a_791_264.t5 a_729_369.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0992 pd=0.95 as=0.1152 ps=1 w=0.64 l=0.15
X27 a_381_47.t1 D.t1 a_299_47.t4 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 VPWR.t12 a_791_264.t6 a_2135_413.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0882 ps=0.84 w=0.42 l=0.15
X29 VPWR.t0 a_423_343.t3 a_381_369.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X30 a_915_47# SCE.t3 a_299_47.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1984 pd=1.9 as=0.0992 ps=0.95 w=0.64 l=0.15
X31 a_1960_413.t0 a_1610_159.t4 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 VGND.t10 a_2051_413.t5 a_791_264.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 a_1226_119.t1 SCD.t0 VGND.t7 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X34 a_1446_413.t1 a_193_47.t4 a_915_47# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.13415 ps=1.085 w=0.42 l=0.15
X35 a_915_47# a_885_21.t2 a_299_47.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X36 VGND.t4 CLK.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 VGND.t9 DE.t3 a_381_47.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X38 a_1610_159.t1 a_1446_413.t5 VGND.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
R0 D.n0 D.t1 220.367
R1 D.n0 D.t0 216.796
R2 D D.n0 71.33
R3 a_299_47.n1 a_299_47.t5 467.892
R4 a_299_47.n3 a_299_47.n2 380.248
R5 a_299_47.n1 a_299_47.t4 232.434
R6 a_299_47.n2 a_299_47.n0 188.082
R7 a_299_47.n3 a_299_47.t2 53.8677
R8 a_299_47.t1 a_299_47.n3 41.5552
R9 a_299_47.n0 a_299_47.t3 38.5719
R10 a_299_47.n0 a_299_47.t0 38.5719
R11 a_299_47.n2 a_299_47.n1 20.4743
R12 a_381_369.t0 a_381_369.t1 64.6411
R13 VPB.t6 VPB.t1 1043.39
R14 VPB.t3 VPB.t14 787.227
R15 VPB.t5 VPB.t6 622.851
R16 VPB.t7 VPB.t9 556.386
R17 VPB.t11 VPB.t12 556.386
R18 VPB.t18 VPB.t15 556.386
R19 VPB.t9 VPB.t0 517.913
R20 VPB.t2 VPB.t7 390.654
R21 VPB.t0 VPB.t16 337.384
R22 VPB.t17 VPB.t2 304.829
R23 VPB.t8 VPB.t4 301.87
R24 VPB.t14 VPB.t13 287.072
R25 VPB.t16 VPB.t3 287.072
R26 VPB.t4 VPB.t5 272.274
R27 VPB.t12 VPB.t8 260.437
R28 VPB.t1 VPB.t17 256.56
R29 VPB.t10 VPB.t18 248.599
R30 VPB.t15 VPB.t11 213.084
R31 VPB VPB.t10 142.056
R32 a_27_47.n3 a_27_47.t2 443.44
R33 a_27_47.t1 a_27_47.n6 390.443
R34 a_27_47.n4 a_27_47.t5 344.428
R35 a_27_47.n4 a_27_47.t3 296.969
R36 a_27_47.n1 a_27_47.t0 288.373
R37 a_27_47.n0 a_27_47.t6 263.406
R38 a_27_47.n3 a_27_47.n2 254.389
R39 a_27_47.n0 a_27_47.t4 228.06
R40 a_27_47.n5 a_27_47.n3 194.501
R41 a_27_47.n1 a_27_47.n0 152
R42 a_27_47.n6 a_27_47.n1 35.3396
R43 a_27_47.n6 a_27_47.n5 15.3376
R44 a_27_47.n5 a_27_47.n4 12.879
R45 a_2051_413.t0 a_2051_413.n3 705.342
R46 a_2051_413.n3 a_2051_413.t1 362.557
R47 a_2051_413.n3 a_2051_413.n2 329.163
R48 a_2051_413.n0 a_2051_413.t3 212.081
R49 a_2051_413.n1 a_2051_413.t5 176.733
R50 a_2051_413.n2 a_2051_413.t4 163.881
R51 a_2051_413.n0 a_2051_413.t2 139.78
R52 a_2051_413.n1 a_2051_413.n0 70.8399
R53 a_2051_413.n2 a_2051_413.n1 33.7405
R54 VNB.t3 VNB.t16 3460.19
R55 VNB.t0 VNB.t12 3203.88
R56 VNB.t8 VNB.t5 3066.59
R57 VNB.t1 VNB.t11 2890.61
R58 VNB.t11 VNB.t3 2733.98
R59 VNB.t12 VNB.t1 2677.02
R60 VNB.t14 VNB.t13 2677.02
R61 VNB.t10 VNB.t18 2677.02
R62 VNB.t6 VNB.t9 2318.4
R63 VNB.t2 VNB.t4 1452.43
R64 VNB.t16 VNB.t17 1381.23
R65 VNB.t9 VNB.t0 1253.07
R66 VNB.t13 VNB.t2 1253.07
R67 VNB.t4 VNB.t8 1196.12
R68 VNB.t7 VNB.t10 1196.12
R69 VNB.t5 VNB.t15 1103.28
R70 VNB.t18 VNB.t14 1025.24
R71 VNB.t15 VNB.t6 945.673
R72 VNB VNB.t7 683.495
R73 a_1446_413.n3 a_1446_413.n2 680.737
R74 a_1446_413.n2 a_1446_413.n1 276.272
R75 a_1446_413.n0 a_1446_413.t5 230.484
R76 a_1446_413.n0 a_1446_413.t4 196.013
R77 a_1446_413.n2 a_1446_413.n0 171.939
R78 a_1446_413.n3 a_1446_413.t3 72.7029
R79 a_1446_413.t1 a_1446_413.n3 70.3576
R80 a_1446_413.n1 a_1446_413.t0 51.6672
R81 a_1446_413.n1 a_1446_413.t2 45.0005
R82 a_1537_413.t0 a_1537_413.t1 171.202
R83 DE.n0 DE.t2 319.728
R84 DE.n2 DE.n1 238.69
R85 DE.n0 DE.t0 178.34
R86 DE DE.n2 158.893
R87 DE.n1 DE.n0 147.814
R88 DE.n2 DE.t3 130.387
R89 DE.n1 DE.t1 130.141
R90 a_423_343.t1 a_423_343.n1 376.974
R91 a_423_343.n1 a_423_343.t3 375.568
R92 a_423_343.n0 a_423_343.t2 334.038
R93 a_423_343.n0 a_423_343.t0 244.181
R94 a_423_343.n1 a_423_343.n0 11.1343
R95 VPWR.n26 VPWR.t8 667.963
R96 VPWR.n38 VPWR.t3 659.122
R97 VPWR.n53 VPWR.n1 604.394
R98 VPWR.n47 VPWR.t0 374.937
R99 VPWR.n45 VPWR.n5 323.079
R100 VPWR.n12 VPWR.n11 317.757
R101 VPWR.n18 VPWR.n17 245.905
R102 VPWR.n19 VPWR.n16 231.042
R103 VPWR.n11 VPWR.t1 106.1
R104 VPWR.n16 VPWR.t12 95.3126
R105 VPWR.n17 VPWR.t10 61.9802
R106 VPWR.n5 VPWR.t7 44.6333
R107 VPWR.n5 VPWR.t6 44.6333
R108 VPWR.n11 VPWR.t5 43.3405
R109 VPWR.n1 VPWR.t4 41.5552
R110 VPWR.n1 VPWR.t9 41.5552
R111 VPWR.n51 VPWR.n2 34.6358
R112 VPWR.n52 VPWR.n51 34.6358
R113 VPWR.n40 VPWR.n39 34.6358
R114 VPWR.n40 VPWR.n6 34.6358
R115 VPWR.n44 VPWR.n6 34.6358
R116 VPWR.n32 VPWR.n31 34.6358
R117 VPWR.n33 VPWR.n32 34.6358
R118 VPWR.n33 VPWR.n9 34.6358
R119 VPWR.n37 VPWR.n9 34.6358
R120 VPWR.n21 VPWR.n20 34.6358
R121 VPWR.n21 VPWR.n14 34.6358
R122 VPWR.n25 VPWR.n14 34.6358
R123 VPWR.n45 VPWR.n44 33.8829
R124 VPWR.n47 VPWR.n46 32.0005
R125 VPWR.n17 VPWR.t11 30.1762
R126 VPWR.n27 VPWR.n26 30.1181
R127 VPWR.n19 VPWR.n18 29.0203
R128 VPWR.n39 VPWR.n38 28.2358
R129 VPWR.n31 VPWR.n12 28.2358
R130 VPWR.n16 VPWR.t2 26.4482
R131 VPWR.n27 VPWR.n12 23.3417
R132 VPWR.n53 VPWR.n52 22.9652
R133 VPWR.n46 VPWR.n45 20.7064
R134 VPWR.n26 VPWR.n25 17.3181
R135 VPWR.n38 VPWR.n37 15.0593
R136 VPWR.n20 VPWR.n19 13.177
R137 VPWR.n47 VPWR.n2 12.424
R138 VPWR.n20 VPWR.n15 9.3005
R139 VPWR.n22 VPWR.n21 9.3005
R140 VPWR.n23 VPWR.n14 9.3005
R141 VPWR.n25 VPWR.n24 9.3005
R142 VPWR.n26 VPWR.n13 9.3005
R143 VPWR.n28 VPWR.n27 9.3005
R144 VPWR.n29 VPWR.n12 9.3005
R145 VPWR.n31 VPWR.n30 9.3005
R146 VPWR.n32 VPWR.n10 9.3005
R147 VPWR.n34 VPWR.n33 9.3005
R148 VPWR.n35 VPWR.n9 9.3005
R149 VPWR.n37 VPWR.n36 9.3005
R150 VPWR.n38 VPWR.n8 9.3005
R151 VPWR.n39 VPWR.n7 9.3005
R152 VPWR.n41 VPWR.n40 9.3005
R153 VPWR.n42 VPWR.n6 9.3005
R154 VPWR.n44 VPWR.n43 9.3005
R155 VPWR.n45 VPWR.n4 9.3005
R156 VPWR.n46 VPWR.n3 9.3005
R157 VPWR.n48 VPWR.n47 9.3005
R158 VPWR.n49 VPWR.n2 9.3005
R159 VPWR.n51 VPWR.n50 9.3005
R160 VPWR.n52 VPWR.n0 9.3005
R161 VPWR.n54 VPWR.n53 7.12063
R162 VPWR.n18 VPWR.n15 0.186831
R163 VPWR.n54 VPWR.n0 0.148519
R164 VPWR.n22 VPWR.n15 0.120292
R165 VPWR.n23 VPWR.n22 0.120292
R166 VPWR.n24 VPWR.n23 0.120292
R167 VPWR.n24 VPWR.n13 0.120292
R168 VPWR.n28 VPWR.n13 0.120292
R169 VPWR.n29 VPWR.n28 0.120292
R170 VPWR.n30 VPWR.n29 0.120292
R171 VPWR.n30 VPWR.n10 0.120292
R172 VPWR.n34 VPWR.n10 0.120292
R173 VPWR.n35 VPWR.n34 0.120292
R174 VPWR.n36 VPWR.n35 0.120292
R175 VPWR.n36 VPWR.n8 0.120292
R176 VPWR.n8 VPWR.n7 0.120292
R177 VPWR.n41 VPWR.n7 0.120292
R178 VPWR.n42 VPWR.n41 0.120292
R179 VPWR.n43 VPWR.n42 0.120292
R180 VPWR.n43 VPWR.n4 0.120292
R181 VPWR.n4 VPWR.n3 0.120292
R182 VPWR.n48 VPWR.n3 0.120292
R183 VPWR.n49 VPWR.n48 0.120292
R184 VPWR.n50 VPWR.n49 0.120292
R185 VPWR.n50 VPWR.n0 0.120292
R186 VPWR VPWR.n54 0.114842
R187 CLK.n0 CLK.t0 292.95
R188 CLK.n0 CLK.t1 209.403
R189 CLK CLK.n0 154.069
R190 SCE.t1 SCE.t2 604.107
R191 SCE.n1 SCE.t3 352.397
R192 SCE.n0 SCE.t0 189.588
R193 SCE SCE.n1 153.631
R194 SCE.n0 SCE.t1 142.03
R195 SCE.n1 SCE.n0 74.0857
R196 a_885_21.n0 a_885_21.t2 571.547
R197 a_885_21.n2 a_885_21.n1 427.555
R198 a_885_21.t0 a_885_21.n2 372.423
R199 a_885_21.n0 a_885_21.t1 223.571
R200 a_885_21.n2 a_885_21.n0 74.941
R201 VGND.n26 VGND.t5 273.476
R202 VGND.n20 VGND.t1 244.518
R203 VGND.n47 VGND.t9 238.311
R204 VGND.n34 VGND.n33 222.888
R205 VGND.n45 VGND.n4 202.262
R206 VGND.n54 VGND.n53 199.739
R207 VGND.n14 VGND.t2 141.867
R208 VGND.n15 VGND.n13 123.651
R209 VGND.n13 VGND.t10 57.8184
R210 VGND.n4 VGND.t0 41.4291
R211 VGND.n4 VGND.t8 41.4291
R212 VGND.n33 VGND.t7 38.5719
R213 VGND.n33 VGND.t6 38.5719
R214 VGND.n53 VGND.t3 38.5719
R215 VGND.n53 VGND.t4 38.5719
R216 VGND.n18 VGND.n12 34.6358
R217 VGND.n19 VGND.n18 34.6358
R218 VGND.n21 VGND.n19 34.6358
R219 VGND.n25 VGND.n10 34.6358
R220 VGND.n27 VGND.n8 34.6358
R221 VGND.n31 VGND.n8 34.6358
R222 VGND.n32 VGND.n31 34.6358
R223 VGND.n35 VGND.n32 34.6358
R224 VGND.n39 VGND.n6 34.6358
R225 VGND.n40 VGND.n39 34.6358
R226 VGND.n41 VGND.n40 34.6358
R227 VGND.n41 VGND.n3 34.6358
R228 VGND.n51 VGND.n1 34.6358
R229 VGND.n52 VGND.n51 34.6358
R230 VGND.n47 VGND.n46 32.0005
R231 VGND.n45 VGND.n3 29.7417
R232 VGND.n26 VGND.n25 24.8476
R233 VGND.n13 VGND.t11 24.7498
R234 VGND.n54 VGND.n52 22.9652
R235 VGND.n35 VGND.n34 15.0593
R236 VGND.n27 VGND.n26 14.6829
R237 VGND.n46 VGND.n45 14.6829
R238 VGND.n15 VGND.n14 13.9614
R239 VGND.n47 VGND.n1 12.424
R240 VGND.n21 VGND.n20 11.2946
R241 VGND.n14 VGND.n12 9.41227
R242 VGND.n52 VGND.n0 9.3005
R243 VGND.n51 VGND.n50 9.3005
R244 VGND.n49 VGND.n1 9.3005
R245 VGND.n48 VGND.n47 9.3005
R246 VGND.n46 VGND.n2 9.3005
R247 VGND.n45 VGND.n44 9.3005
R248 VGND.n43 VGND.n3 9.3005
R249 VGND.n42 VGND.n41 9.3005
R250 VGND.n40 VGND.n5 9.3005
R251 VGND.n39 VGND.n38 9.3005
R252 VGND.n37 VGND.n6 9.3005
R253 VGND.n16 VGND.n12 9.3005
R254 VGND.n18 VGND.n17 9.3005
R255 VGND.n19 VGND.n11 9.3005
R256 VGND.n22 VGND.n21 9.3005
R257 VGND.n23 VGND.n10 9.3005
R258 VGND.n25 VGND.n24 9.3005
R259 VGND.n26 VGND.n9 9.3005
R260 VGND.n28 VGND.n27 9.3005
R261 VGND.n29 VGND.n8 9.3005
R262 VGND.n31 VGND.n30 9.3005
R263 VGND.n32 VGND.n7 9.3005
R264 VGND.n36 VGND.n35 9.3005
R265 VGND.n55 VGND.n54 7.12063
R266 VGND.n20 VGND.n10 2.63579
R267 VGND.n34 VGND.n6 0.753441
R268 VGND.n16 VGND.n15 0.186831
R269 VGND.n55 VGND.n0 0.148519
R270 VGND.n17 VGND.n16 0.120292
R271 VGND.n17 VGND.n11 0.120292
R272 VGND.n22 VGND.n11 0.120292
R273 VGND.n23 VGND.n22 0.120292
R274 VGND.n24 VGND.n23 0.120292
R275 VGND.n24 VGND.n9 0.120292
R276 VGND.n28 VGND.n9 0.120292
R277 VGND.n29 VGND.n28 0.120292
R278 VGND.n30 VGND.n29 0.120292
R279 VGND.n30 VGND.n7 0.120292
R280 VGND.n36 VGND.n7 0.120292
R281 VGND.n37 VGND.n36 0.120292
R282 VGND.n38 VGND.n37 0.120292
R283 VGND.n38 VGND.n5 0.120292
R284 VGND.n42 VGND.n5 0.120292
R285 VGND.n43 VGND.n42 0.120292
R286 VGND.n44 VGND.n43 0.120292
R287 VGND.n44 VGND.n2 0.120292
R288 VGND.n48 VGND.n2 0.120292
R289 VGND.n49 VGND.n48 0.120292
R290 VGND.n50 VGND.n49 0.120292
R291 VGND.n50 VGND.n0 0.120292
R292 VGND VGND.n55 0.114842
R293 Q Q.t0 251.107
R294 Q Q.t1 146.542
R295 a_791_264.t0 a_791_264.n6 394.808
R296 a_791_264.n1 a_791_264.t6 368.969
R297 a_791_264.n4 a_791_264.t4 310.623
R298 a_791_264.n6 a_791_264.n3 308.443
R299 a_791_264.n2 a_791_264.t3 245.821
R300 a_791_264.n5 a_791_264.t1 241.077
R301 a_791_264.n5 a_791_264.n4 221.578
R302 a_791_264.n4 a_791_264.t5 194.942
R303 a_791_264.n1 a_791_264.n0 189.588
R304 a_791_264.n3 a_791_264.t2 152.633
R305 a_791_264.n2 a_791_264.n1 96.4005
R306 a_791_264.n3 a_791_264.n2 29.9627
R307 a_791_264.n6 a_791_264.n5 7.71815
R308 Q_N Q_N.t0 246.079
R309 Q_N Q_N.t1 148.946
R310 a_1610_159.t0 a_1610_159.n4 408.848
R311 a_1610_159.n2 a_1610_159.t2 406.401
R312 a_1610_159.n0 a_1610_159.t4 318.12
R313 a_1610_159.n0 a_1610_159.t3 194.477
R314 a_1610_159.n3 a_1610_159.n2 176.534
R315 a_1610_159.n4 a_1610_159.n0 168.486
R316 a_1610_159.n3 a_1610_159.t1 140.249
R317 a_1610_159.n2 a_1610_159.n1 130.054
R318 a_1610_159.n4 a_1610_159.n3 9.32396
R319 a_193_47.t0 a_193_47.n4 395.625
R320 a_193_47.n2 a_193_47.t2 389.545
R321 a_193_47.n1 a_193_47.t3 308.651
R322 a_193_47.n4 a_193_47.t1 300.372
R323 a_193_47.n1 a_193_47.n0 298.373
R324 a_193_47.n2 a_193_47.t4 273.572
R325 a_193_47.n3 a_193_47.n2 173.755
R326 a_193_47.n4 a_193_47.n3 14.6322
R327 a_193_47.n3 a_193_47.n1 12.2528
R328 a_1974_47.n0 a_1974_47.t0 45.1697
R329 a_729_47.t0 a_729_47.t1 102.858
R330 a_729_369.t0 a_729_369.t1 110.812
R331 a_2135_413.t0 a_2135_413.t1 197
R332 SCD.n1 SCD.t0 206.19
R333 SCD.n1 SCD.n0 183.696
R334 SCD SCD.n1 163.675
R335 a_1226_119.t0 a_1226_119.t1 60.0005
R336 a_381_47.t0 a_381_47.t1 60.0005
C0 SCE Q 1.83e-20
C1 VPWR VGND 0.07604f
C2 VPB Q 0.016876f
C3 a_915_47# VGND 0.383404f
C4 a_1561_47# a_915_47# 4.9e-19
C5 VPWR CLK 0.019263f
C6 VPB DE 0.114449f
C7 VGND Q 0.100622f
C8 DE VGND 0.057232f
C9 SCE SCD 0.095395f
C10 SCD VPB 0.045339f
C11 SCD VGND 0.032521f
C12 SCE Q_N 3.14e-20
C13 VPB Q_N 0.015582f
C14 VPB D 0.068631f
C15 VGND Q_N 0.097568f
C16 VPWR a_1231_369# 0.0081f
C17 a_915_47# a_1231_369# 0.003336f
C18 D VGND 0.014495f
C19 SCE VPB 0.1417f
C20 a_915_47# a_2177_47# 1.55e-20
C21 a_915_47# VPWR 0.097411f
C22 SCE VGND 0.047506f
C23 VPB VGND 0.014939f
C24 VPWR Q 0.122443f
C25 VPB CLK 0.069635f
C26 a_915_47# Q 2.61e-20
C27 VPWR DE 0.04692f
C28 a_1561_47# VGND 0.004442f
C29 CLK VGND 0.019296f
C30 SCD VPWR 0.013425f
C31 a_915_47# SCD 0.018533f
C32 VPWR Q_N 0.124307f
C33 a_915_47# Q_N 4.59e-20
C34 VPWR D 0.01674f
C35 D DE 0.099354f
C36 SCE VPWR 0.028732f
C37 VPWR VPB 0.316481f
C38 a_915_47# SCE 0.086615f
C39 a_915_47# VPB 0.021894f
C40 a_2177_47# VGND 0.002966f
C41 Q VNB 0.083148f
C42 Q_N VNB 0.012608f
C43 VGND VNB 1.56683f
C44 VPWR VNB 1.26744f
C45 SCD VNB 0.08884f
C46 SCE VNB 0.334233f
C47 DE VNB 0.282831f
C48 D VNB 0.122269f
C49 CLK VNB 0.195128f
C50 VPB VNB 2.78355f
C51 a_915_47# VNB 0.038144f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxbp_2 VPWR VGND CLK SCD DE Q D Q_N SCE VPB VNB
X0 VGND.t4 a_791_264# Q_N.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_381_369.t1 D.t0 a_299_47.t5 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 a_2177_47# a_27_47.t2 a_2051_413.t1 VNB.t19 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3 a_1537_413.t1 a_27_47.t3 a_1446_413.t2 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 VPWR.t3 DE.t0 a_423_343.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t9 CLK.t0 a_27_47.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 VPWR.t0 SCE.t0 a_885_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1264 pd=1.035 as=0.1696 ps=1.81 w=0.64 l=0.15
X7 VGND.t8 SCE.t1 a_885_21.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND.t5 a_2051_413.t2 Q.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Q_N.t0 a_791_264# VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X10 VPWR.t1 a_1610_159.t2 a_1537_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11 a_1610_159.t0 a_1446_413.t4 VPWR.t2 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 VGND.t1 DE.t1 a_423_343.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_1561_47# a_193_47.t2 a_1446_413.t1 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X14 a_1974_47.t0 a_1610_159.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VPWR.t7 a_791_264# Q_N.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR.t10 a_2051_413.t3 Q.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_193_47.t1 a_27_47.t4 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_729_47.t0 a_423_343.t2 VGND.t12 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X19 Q.t0 a_2051_413.t4 VPWR.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X20 Q_N.t2 a_791_264# VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X21 a_729_369.t0 DE.t2 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X22 a_299_47.t0 a_791_264# a_729_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0756 ps=0.78 w=0.42 l=0.15
X23 a_2135_413.t0 a_193_47.t3 a_2051_413.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 a_1446_413.t3 a_27_47.t5 a_915_47# VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.22515 ps=1.505 w=0.36 l=0.15
X25 a_193_47.t0 a_27_47.t6 VPWR.t12 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 a_1231_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1056 pd=0.97 as=0.1264 ps=1.035 w=0.64 l=0.15
X27 a_915_47# SCE.t2 a_1226_119.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.22515 pd=1.505 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_299_47.t1 a_791_264# a_729_369.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0992 pd=0.95 as=0.1152 ps=1 w=0.64 l=0.15
X29 a_381_47.t1 D.t1 a_299_47.t4 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 VPWR.t8 a_791_264# a_2135_413.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0882 ps=0.84 w=0.42 l=0.15
X31 VPWR.t5 a_423_343.t3 a_381_369.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X32 a_915_47# SCE.t3 a_299_47.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1984 pd=1.9 as=0.0992 ps=0.95 w=0.64 l=0.15
X33 a_1960_413.t0 a_1610_159.t4 VPWR.t13 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X34 a_1226_119.t0 SCD.t0 VGND.t11 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X35 VGND a_791_264# a_2177_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.066 ps=0.745 w=0.42 l=0.15
X36 a_1446_413.t0 a_193_47.t4 a_915_47# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.13415 ps=1.085 w=0.42 l=0.15
X37 a_915_47# a_885_21.t2 a_299_47.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X38 VGND.t7 CLK.t1 a_27_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X39 VGND.t2 DE.t3 a_381_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X40 a_1610_159.t1 a_1446_413.t5 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
X41 Q.t2 a_2051_413.t5 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
R0 Q_N Q_N.n0 220.587
R1 Q_N Q_N.n1 109.635
R2 Q_N.n0 Q_N.t3 26.5955
R3 Q_N.n0 Q_N.t2 26.5955
R4 Q_N.n1 Q_N.t1 24.9236
R5 Q_N.n1 Q_N.t0 24.9236
R6 VGND.n35 VGND.t9 273.476
R7 VGND.n29 VGND.t0 244.518
R8 VGND.n56 VGND.t2 238.311
R9 VGND.n43 VGND.n42 222.888
R10 VGND.n54 VGND.n4 202.262
R11 VGND.n63 VGND.n62 199.739
R12 VGND.n16 VGND.t5 158.077
R13 VGND.n20 VGND.t4 156.085
R14 VGND.n15 VGND.t10 143.409
R15 VGND.n22 VGND.t3 141.867
R16 VGND.n4 VGND.t12 41.4291
R17 VGND.n4 VGND.t1 41.4291
R18 VGND.n42 VGND.t11 38.5719
R19 VGND.n42 VGND.t8 38.5719
R20 VGND.n62 VGND.t6 38.5719
R21 VGND.n62 VGND.t7 38.5719
R22 VGND.n19 VGND.n14 34.6358
R23 VGND.n23 VGND.n21 34.6358
R24 VGND.n27 VGND.n12 34.6358
R25 VGND.n28 VGND.n27 34.6358
R26 VGND.n30 VGND.n28 34.6358
R27 VGND.n34 VGND.n10 34.6358
R28 VGND.n36 VGND.n8 34.6358
R29 VGND.n40 VGND.n8 34.6358
R30 VGND.n41 VGND.n40 34.6358
R31 VGND.n44 VGND.n41 34.6358
R32 VGND.n48 VGND.n6 34.6358
R33 VGND.n49 VGND.n48 34.6358
R34 VGND.n50 VGND.n49 34.6358
R35 VGND.n50 VGND.n3 34.6358
R36 VGND.n60 VGND.n1 34.6358
R37 VGND.n61 VGND.n60 34.6358
R38 VGND.n56 VGND.n55 32.0005
R39 VGND.n15 VGND.n14 31.624
R40 VGND.n54 VGND.n3 29.7417
R41 VGND.n35 VGND.n34 24.8476
R42 VGND.n63 VGND.n61 22.9652
R43 VGND.n44 VGND.n43 15.0593
R44 VGND.n36 VGND.n35 14.6829
R45 VGND.n55 VGND.n54 14.6829
R46 VGND.n56 VGND.n1 12.424
R47 VGND.n30 VGND.n29 11.2946
R48 VGND.n21 VGND.n20 9.41227
R49 VGND.n22 VGND.n12 9.41227
R50 VGND.n61 VGND.n0 9.3005
R51 VGND.n60 VGND.n59 9.3005
R52 VGND.n58 VGND.n1 9.3005
R53 VGND.n57 VGND.n56 9.3005
R54 VGND.n55 VGND.n2 9.3005
R55 VGND.n54 VGND.n53 9.3005
R56 VGND.n52 VGND.n3 9.3005
R57 VGND.n51 VGND.n50 9.3005
R58 VGND.n49 VGND.n5 9.3005
R59 VGND.n48 VGND.n47 9.3005
R60 VGND.n46 VGND.n6 9.3005
R61 VGND.n17 VGND.n14 9.3005
R62 VGND.n19 VGND.n18 9.3005
R63 VGND.n21 VGND.n13 9.3005
R64 VGND.n24 VGND.n23 9.3005
R65 VGND.n25 VGND.n12 9.3005
R66 VGND.n27 VGND.n26 9.3005
R67 VGND.n28 VGND.n11 9.3005
R68 VGND.n31 VGND.n30 9.3005
R69 VGND.n32 VGND.n10 9.3005
R70 VGND.n34 VGND.n33 9.3005
R71 VGND.n35 VGND.n9 9.3005
R72 VGND.n37 VGND.n36 9.3005
R73 VGND.n38 VGND.n8 9.3005
R74 VGND.n40 VGND.n39 9.3005
R75 VGND.n41 VGND.n7 9.3005
R76 VGND.n45 VGND.n44 9.3005
R77 VGND.n64 VGND.n63 7.12063
R78 VGND.n16 VGND.n15 6.56513
R79 VGND.n20 VGND.n19 6.4005
R80 VGND.n23 VGND.n22 6.4005
R81 VGND.n29 VGND.n10 2.63579
R82 VGND.n43 VGND.n6 0.753441
R83 VGND.n17 VGND.n16 0.508363
R84 VGND.n64 VGND.n0 0.148519
R85 VGND.n18 VGND.n17 0.120292
R86 VGND.n18 VGND.n13 0.120292
R87 VGND.n24 VGND.n13 0.120292
R88 VGND.n25 VGND.n24 0.120292
R89 VGND.n26 VGND.n25 0.120292
R90 VGND.n26 VGND.n11 0.120292
R91 VGND.n31 VGND.n11 0.120292
R92 VGND.n32 VGND.n31 0.120292
R93 VGND.n33 VGND.n32 0.120292
R94 VGND.n33 VGND.n9 0.120292
R95 VGND.n37 VGND.n9 0.120292
R96 VGND.n38 VGND.n37 0.120292
R97 VGND.n39 VGND.n38 0.120292
R98 VGND.n39 VGND.n7 0.120292
R99 VGND.n45 VGND.n7 0.120292
R100 VGND.n46 VGND.n45 0.120292
R101 VGND.n47 VGND.n46 0.120292
R102 VGND.n47 VGND.n5 0.120292
R103 VGND.n51 VGND.n5 0.120292
R104 VGND.n52 VGND.n51 0.120292
R105 VGND.n53 VGND.n52 0.120292
R106 VGND.n53 VGND.n2 0.120292
R107 VGND.n57 VGND.n2 0.120292
R108 VGND.n58 VGND.n57 0.120292
R109 VGND.n59 VGND.n58 0.120292
R110 VGND.n59 VGND.n0 0.120292
R111 VGND VGND.n64 0.114842
R112 VNB.t5 VNB.t14 4841.42
R113 VNB.t11 VNB.t13 3203.88
R114 VNB.t12 VNB.t10 3066.59
R115 VNB.t0 VNB.t19 2890.61
R116 VNB.t19 VNB.t4 2733.98
R117 VNB.t13 VNB.t0 2677.02
R118 VNB.t2 VNB.t1 2677.02
R119 VNB.t7 VNB.t18 2677.02
R120 VNB.t16 VNB.t8 2318.4
R121 VNB.t17 VNB.t3 1452.43
R122 VNB.t8 VNB.t11 1253.07
R123 VNB.t1 VNB.t17 1253.07
R124 VNB.t14 VNB.t6 1196.12
R125 VNB.t4 VNB.t5 1196.12
R126 VNB.t3 VNB.t12 1196.12
R127 VNB.t9 VNB.t7 1196.12
R128 VNB.t10 VNB.t15 1103.28
R129 VNB.t18 VNB.t2 1025.24
R130 VNB.t15 VNB.t16 945.673
R131 VNB VNB.t9 683.495
R132 D.n0 D.t1 220.367
R133 D.n0 D.t0 216.796
R134 D D.n0 71.33
R135 a_299_47.n1 a_299_47.t5 467.892
R136 a_299_47.n3 a_299_47.n2 380.248
R137 a_299_47.n1 a_299_47.t4 232.434
R138 a_299_47.n2 a_299_47.n0 188.082
R139 a_299_47.n3 a_299_47.t2 53.8677
R140 a_299_47.t1 a_299_47.n3 41.5552
R141 a_299_47.n0 a_299_47.t3 38.5719
R142 a_299_47.n0 a_299_47.t0 38.5719
R143 a_299_47.n2 a_299_47.n1 20.4743
R144 a_381_369.t0 a_381_369.t1 64.6411
R145 VPB.t7 VPB.t9 1074.3
R146 VPB.t0 VPB.t1 1043.39
R147 VPB.t10 VPB.t0 622.851
R148 VPB.t15 VPB.t19 556.386
R149 VPB.t12 VPB.t14 556.386
R150 VPB.t11 VPB.t17 556.386
R151 VPB.t19 VPB.t16 517.913
R152 VPB.t2 VPB.t15 390.654
R153 VPB.t16 VPB.t4 337.384
R154 VPB.t18 VPB.t2 304.829
R155 VPB.t3 VPB.t5 301.87
R156 VPB.t4 VPB.t6 287.072
R157 VPB.t5 VPB.t10 272.274
R158 VPB.t14 VPB.t3 260.437
R159 VPB.t1 VPB.t18 256.56
R160 VPB.t9 VPB.t8 248.599
R161 VPB.t6 VPB.t7 248.599
R162 VPB.t13 VPB.t11 248.599
R163 VPB.t17 VPB.t12 213.084
R164 VPB VPB.t13 142.056
R165 a_27_47.n3 a_27_47.t2 443.44
R166 a_27_47.t0 a_27_47.n6 390.443
R167 a_27_47.n4 a_27_47.t5 344.428
R168 a_27_47.n4 a_27_47.t3 296.969
R169 a_27_47.n1 a_27_47.t1 288.373
R170 a_27_47.n0 a_27_47.t6 263.406
R171 a_27_47.n3 a_27_47.n2 254.389
R172 a_27_47.n0 a_27_47.t4 228.06
R173 a_27_47.n5 a_27_47.n3 194.501
R174 a_27_47.n1 a_27_47.n0 152
R175 a_27_47.n6 a_27_47.n1 35.3396
R176 a_27_47.n6 a_27_47.n5 15.3376
R177 a_27_47.n5 a_27_47.n4 12.879
R178 a_2051_413.t0 a_2051_413.n6 705.342
R179 a_2051_413.n6 a_2051_413.t1 362.557
R180 a_2051_413.n6 a_2051_413.n5 329.538
R181 a_2051_413.n2 a_2051_413.t3 212.081
R182 a_2051_413.n3 a_2051_413.t4 212.081
R183 a_2051_413.n4 a_2051_413.n1 176.733
R184 a_2051_413.n5 a_2051_413.n0 163.881
R185 a_2051_413.n2 a_2051_413.t2 139.78
R186 a_2051_413.n3 a_2051_413.t5 139.78
R187 a_2051_413.n4 a_2051_413.n3 70.8399
R188 a_2051_413.n3 a_2051_413.n2 61.346
R189 a_2051_413.n5 a_2051_413.n4 33.7405
R190 a_1446_413.n3 a_1446_413.n2 680.737
R191 a_1446_413.n2 a_1446_413.n1 276.272
R192 a_1446_413.n0 a_1446_413.t5 230.484
R193 a_1446_413.n0 a_1446_413.t4 196.013
R194 a_1446_413.n2 a_1446_413.n0 171.939
R195 a_1446_413.n3 a_1446_413.t2 72.7029
R196 a_1446_413.t0 a_1446_413.n3 70.3576
R197 a_1446_413.n1 a_1446_413.t1 51.6672
R198 a_1446_413.n1 a_1446_413.t3 45.0005
R199 a_1537_413.t0 a_1537_413.t1 171.202
R200 DE.n0 DE.t2 319.728
R201 DE.n2 DE.n1 238.69
R202 DE.n0 DE.t0 178.34
R203 DE DE.n2 158.893
R204 DE.n1 DE.n0 147.814
R205 DE.n2 DE.t3 130.387
R206 DE.n1 DE.t1 130.141
R207 a_423_343.t1 a_423_343.n1 376.974
R208 a_423_343.n1 a_423_343.t3 375.568
R209 a_423_343.n0 a_423_343.t2 334.038
R210 a_423_343.n0 a_423_343.t0 244.181
R211 a_423_343.n1 a_423_343.n0 11.1343
R212 VPWR.n35 VPWR.t13 667.963
R213 VPWR.n47 VPWR.t0 659.122
R214 VPWR.n62 VPWR.n1 604.394
R215 VPWR.n56 VPWR.t5 374.937
R216 VPWR.n54 VPWR.n5 323.079
R217 VPWR.n12 VPWR.n11 317.757
R218 VPWR.n20 VPWR.t11 271.303
R219 VPWR.n19 VPWR.t10 258.531
R220 VPWR.n22 VPWR.t7 252
R221 VPWR.n28 VPWR.n16 231.042
R222 VPWR.n11 VPWR.t1 106.1
R223 VPWR.n16 VPWR.t8 95.3126
R224 VPWR.n5 VPWR.t4 44.6333
R225 VPWR.n5 VPWR.t3 44.6333
R226 VPWR.n11 VPWR.t2 43.3405
R227 VPWR.n1 VPWR.t12 41.5552
R228 VPWR.n1 VPWR.t9 41.5552
R229 VPWR.n60 VPWR.n2 34.6358
R230 VPWR.n61 VPWR.n60 34.6358
R231 VPWR.n49 VPWR.n48 34.6358
R232 VPWR.n49 VPWR.n6 34.6358
R233 VPWR.n53 VPWR.n6 34.6358
R234 VPWR.n41 VPWR.n40 34.6358
R235 VPWR.n42 VPWR.n41 34.6358
R236 VPWR.n42 VPWR.n9 34.6358
R237 VPWR.n46 VPWR.n9 34.6358
R238 VPWR.n27 VPWR.n17 34.6358
R239 VPWR.n30 VPWR.n29 34.6358
R240 VPWR.n30 VPWR.n14 34.6358
R241 VPWR.n34 VPWR.n14 34.6358
R242 VPWR.n23 VPWR.n21 34.6358
R243 VPWR.n54 VPWR.n53 33.8829
R244 VPWR.n56 VPWR.n55 32.0005
R245 VPWR.n21 VPWR.n20 31.624
R246 VPWR.n36 VPWR.n35 30.1181
R247 VPWR.n48 VPWR.n47 28.2358
R248 VPWR.n40 VPWR.n12 28.2358
R249 VPWR.n16 VPWR.t6 26.4482
R250 VPWR.n36 VPWR.n12 23.3417
R251 VPWR.n62 VPWR.n61 22.9652
R252 VPWR.n28 VPWR.n27 21.4593
R253 VPWR.n55 VPWR.n54 20.7064
R254 VPWR.n35 VPWR.n34 17.3181
R255 VPWR.n47 VPWR.n46 15.0593
R256 VPWR.n23 VPWR.n22 15.0593
R257 VPWR.n29 VPWR.n28 13.177
R258 VPWR.n56 VPWR.n2 12.424
R259 VPWR.n21 VPWR.n18 9.3005
R260 VPWR.n24 VPWR.n23 9.3005
R261 VPWR.n25 VPWR.n17 9.3005
R262 VPWR.n27 VPWR.n26 9.3005
R263 VPWR.n29 VPWR.n15 9.3005
R264 VPWR.n31 VPWR.n30 9.3005
R265 VPWR.n32 VPWR.n14 9.3005
R266 VPWR.n34 VPWR.n33 9.3005
R267 VPWR.n35 VPWR.n13 9.3005
R268 VPWR.n37 VPWR.n36 9.3005
R269 VPWR.n38 VPWR.n12 9.3005
R270 VPWR.n40 VPWR.n39 9.3005
R271 VPWR.n41 VPWR.n10 9.3005
R272 VPWR.n43 VPWR.n42 9.3005
R273 VPWR.n44 VPWR.n9 9.3005
R274 VPWR.n46 VPWR.n45 9.3005
R275 VPWR.n47 VPWR.n8 9.3005
R276 VPWR.n48 VPWR.n7 9.3005
R277 VPWR.n50 VPWR.n49 9.3005
R278 VPWR.n51 VPWR.n6 9.3005
R279 VPWR.n53 VPWR.n52 9.3005
R280 VPWR.n54 VPWR.n4 9.3005
R281 VPWR.n55 VPWR.n3 9.3005
R282 VPWR.n57 VPWR.n56 9.3005
R283 VPWR.n58 VPWR.n2 9.3005
R284 VPWR.n60 VPWR.n59 9.3005
R285 VPWR.n61 VPWR.n0 9.3005
R286 VPWR.n63 VPWR.n62 7.12063
R287 VPWR.n20 VPWR.n19 6.56513
R288 VPWR.n22 VPWR.n17 0.753441
R289 VPWR.n19 VPWR.n18 0.508363
R290 VPWR.n63 VPWR.n0 0.148519
R291 VPWR.n24 VPWR.n18 0.120292
R292 VPWR.n25 VPWR.n24 0.120292
R293 VPWR.n26 VPWR.n25 0.120292
R294 VPWR.n26 VPWR.n15 0.120292
R295 VPWR.n31 VPWR.n15 0.120292
R296 VPWR.n32 VPWR.n31 0.120292
R297 VPWR.n33 VPWR.n32 0.120292
R298 VPWR.n33 VPWR.n13 0.120292
R299 VPWR.n37 VPWR.n13 0.120292
R300 VPWR.n38 VPWR.n37 0.120292
R301 VPWR.n39 VPWR.n38 0.120292
R302 VPWR.n39 VPWR.n10 0.120292
R303 VPWR.n43 VPWR.n10 0.120292
R304 VPWR.n44 VPWR.n43 0.120292
R305 VPWR.n45 VPWR.n44 0.120292
R306 VPWR.n45 VPWR.n8 0.120292
R307 VPWR.n8 VPWR.n7 0.120292
R308 VPWR.n50 VPWR.n7 0.120292
R309 VPWR.n51 VPWR.n50 0.120292
R310 VPWR.n52 VPWR.n51 0.120292
R311 VPWR.n52 VPWR.n4 0.120292
R312 VPWR.n4 VPWR.n3 0.120292
R313 VPWR.n57 VPWR.n3 0.120292
R314 VPWR.n58 VPWR.n57 0.120292
R315 VPWR.n59 VPWR.n58 0.120292
R316 VPWR.n59 VPWR.n0 0.120292
R317 VPWR VPWR.n63 0.114842
R318 CLK.n0 CLK.t0 292.95
R319 CLK.n0 CLK.t1 209.403
R320 CLK CLK.n0 154.069
R321 SCE.t1 SCE.t2 604.107
R322 SCE.n1 SCE.t3 352.397
R323 SCE.n0 SCE.t0 189.588
R324 SCE SCE.n1 153.631
R325 SCE.n0 SCE.t1 142.03
R326 SCE.n1 SCE.n0 74.0857
R327 a_885_21.n0 a_885_21.t2 571.547
R328 a_885_21.n2 a_885_21.n1 427.555
R329 a_885_21.t0 a_885_21.n2 372.423
R330 a_885_21.n0 a_885_21.t1 223.571
R331 a_885_21.n2 a_885_21.n0 74.941
R332 Q Q.n0 222.542
R333 Q Q.n1 110.037
R334 Q.n0 Q.t1 26.5955
R335 Q.n0 Q.t0 26.5955
R336 Q.n1 Q.t3 24.9236
R337 Q.n1 Q.t2 24.9236
R338 a_1610_159.t0 a_1610_159.n4 408.848
R339 a_1610_159.n2 a_1610_159.t2 406.401
R340 a_1610_159.n0 a_1610_159.t4 318.12
R341 a_1610_159.n0 a_1610_159.t3 194.477
R342 a_1610_159.n3 a_1610_159.n2 176.534
R343 a_1610_159.n4 a_1610_159.n0 168.486
R344 a_1610_159.n3 a_1610_159.t1 140.249
R345 a_1610_159.n2 a_1610_159.n1 130.054
R346 a_1610_159.n4 a_1610_159.n3 9.32396
R347 a_193_47.t0 a_193_47.n4 395.625
R348 a_193_47.n2 a_193_47.t2 389.545
R349 a_193_47.n1 a_193_47.t3 308.651
R350 a_193_47.n4 a_193_47.t1 300.372
R351 a_193_47.n1 a_193_47.n0 298.373
R352 a_193_47.n2 a_193_47.t4 273.572
R353 a_193_47.n3 a_193_47.n2 173.755
R354 a_193_47.n4 a_193_47.n3 14.6322
R355 a_193_47.n3 a_193_47.n1 12.2528
R356 a_1974_47.n0 a_1974_47.t0 45.1697
R357 a_729_47.t0 a_729_47.t1 102.858
R358 a_729_369.t0 a_729_369.t1 110.812
R359 a_2135_413.t0 a_2135_413.t1 197
R360 SCD.n1 SCD.t0 206.19
R361 SCD.n1 SCD.n0 183.696
R362 SCD SCD.n1 163.675
R363 a_1226_119.t0 a_1226_119.t1 60.0005
R364 a_381_47.t0 a_381_47.t1 60.0005
C0 VPB SCD 0.045339f
C1 a_915_47# a_1231_369# 0.003336f
C2 a_791_264# VPB 0.24965f
C3 a_1561_47# a_915_47# 4.9e-19
C4 SCE SCD 0.095395f
C5 DE VPWR 0.04692f
C6 D VGND 0.014495f
C7 SCE a_791_264# 0.050297f
C8 a_915_47# VGND 0.383468f
C9 a_1231_369# VPWR 0.0081f
C10 VPB Q 0.005756f
C11 VPWR VGND 0.109199f
C12 SCE Q 1.64e-20
C13 a_791_264# Q_N 0.141342f
C14 SCE VPB 0.1417f
C15 D VPWR 0.01674f
C16 DE a_791_264# 0.037542f
C17 CLK VGND 0.019296f
C18 a_915_47# VPWR 0.097411f
C19 a_791_264# a_1561_47# 0.001532f
C20 VPB Q_N 0.00579f
C21 a_2177_47# VGND 0.002966f
C22 SCD VGND 0.032521f
C23 a_791_264# VGND 0.642531f
C24 SCE Q_N 3.14e-20
C25 VGND Q 0.154932f
C26 DE VPB 0.114449f
C27 D a_791_264# 2.15e-19
C28 VPB VGND 0.019902f
C29 CLK VPWR 0.019263f
C30 a_2177_47# a_915_47# 1.55e-20
C31 a_915_47# SCD 0.018533f
C32 a_791_264# a_915_47# 0.276458f
C33 SCE VGND 0.047528f
C34 SCD VPWR 0.013425f
C35 a_791_264# VPWR 0.243886f
C36 a_915_47# Q 2.33e-20
C37 VGND Q_N 0.151675f
C38 VPWR Q 0.203055f
C39 D VPB 0.068631f
C40 VPB a_915_47# 0.021894f
C41 SCE a_915_47# 0.086615f
C42 VPB VPWR 0.358858f
C43 a_791_264# CLK 9.43e-20
C44 SCE VPWR 0.028732f
C45 DE VGND 0.057232f
C46 a_1561_47# VGND 0.004442f
C47 a_791_264# a_2177_47# 6.6e-19
C48 a_791_264# SCD 0.011942f
C49 a_915_47# Q_N 4.59e-20
C50 VPWR Q_N 0.207984f
C51 a_791_264# Q 0.021899f
C52 VPB CLK 0.069635f
C53 D DE 0.099354f
C54 Q VNB 0.021728f
C55 Q_N VNB 0.006861f
C56 VGND VNB 1.69966f
C57 VPWR VNB 1.37565f
C58 SCD VNB 0.08884f
C59 SCE VNB 0.334233f
C60 DE VNB 0.282831f
C61 D VNB 0.122269f
C62 CLK VNB 0.195128f
C63 VPB VNB 2.96074f
C64 a_915_47# VNB 0.037965f
C65 a_791_264# VNB 0.563279f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxtp_1 VPWR VGND CLK SCD DE Q D SCE VPB VNB
X0 a_381_369.t0 D.t0 a_299_47.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_2177_47# a_27_47.t2 a_2051_413# VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2 a_1537_413.t0 a_27_47.t3 a_1446_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 VPWR.t8 DE.t0 a_423_343.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VPWR.t9 CLK.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t5 SCE.t0 a_885_21.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1264 pd=1.035 as=0.1696 ps=1.81 w=0.64 l=0.15
X6 VGND.t0 SCE.t1 a_885_21.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR.t4 a_1610_159.t2 a_1537_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8 a_1610_159.t0 a_1446_413.t4 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X9 VGND.t8 a_2051_413# a_791_264.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND.t6 DE.t1 a_423_343.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_1561_47# a_193_47.t2 a_1446_413.t2 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X12 a_1974_47.t0 a_1610_159.t3 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_193_47.t1 a_27_47.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_729_47.t1 a_423_343.t2 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X15 a_729_369.t1 DE.t2 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X16 Q.t1 a_2051_413# VGND.t9 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10025 ps=0.985 w=0.65 l=0.15
X17 a_299_47.t5 a_791_264.t2 a_729_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0756 ps=0.78 w=0.42 l=0.15
X18 a_2135_413.t1 a_193_47.t3 a_2051_413# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1446_413.t0 a_27_47.t5 a_915_47# VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.22515 ps=1.505 w=0.36 l=0.15
X20 a_193_47.t0 a_27_47.t6 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 a_1231_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1056 pd=0.97 as=0.1264 ps=1.035 w=0.64 l=0.15
X22 a_915_47# SCE.t2 a_1226_119.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.22515 pd=1.505 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 a_299_47.t4 a_791_264.t3 a_729_369.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0992 pd=0.95 as=0.1152 ps=1 w=0.64 l=0.15
X24 a_381_47.t0 D.t1 a_299_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 VPWR.t1 a_791_264.t4 a_2135_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X26 Q.t0 a_2051_413# VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.154 ps=1.335 w=1 l=0.15
X27 VPWR.t6 a_423_343.t3 a_381_369.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X28 a_915_47# SCE.t3 a_299_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1984 pd=1.9 as=0.0992 ps=0.95 w=0.64 l=0.15
X29 a_1960_413# a_1610_159.t4 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 a_1226_119.t1 SCD.t0 VGND.t4 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X31 a_1446_413.t3 a_193_47.t4 a_915_47# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.13415 ps=1.085 w=0.42 l=0.15
X32 a_915_47# a_885_21.t2 a_299_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X33 VPWR.t11 a_2051_413# a_791_264.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1728 ps=1.82 w=0.64 l=0.15
X34 VGND.t10 CLK.t1 a_27_47.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 VGND.t7 DE.t3 a_381_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 a_1610_159.t1 a_1446_413.t5 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
R0 D.n0 D.t1 220.367
R1 D.n0 D.t0 216.796
R2 D D.n0 71.33
R3 a_299_47.n1 a_299_47.t2 467.892
R4 a_299_47.n3 a_299_47.n2 380.248
R5 a_299_47.n1 a_299_47.t1 232.434
R6 a_299_47.n2 a_299_47.n0 188.082
R7 a_299_47.t0 a_299_47.n3 53.8677
R8 a_299_47.n3 a_299_47.t4 41.5552
R9 a_299_47.n0 a_299_47.t3 38.5719
R10 a_299_47.n0 a_299_47.t5 38.5719
R11 a_299_47.n2 a_299_47.n1 20.4743
R12 a_381_369.t0 a_381_369.t1 64.6411
R13 VPB.t5 VPB.t1 1043.39
R14 VPB.t0 VPB.t5 622.851
R15 VPB.t6 VPB.t11 556.386
R16 VPB.t4 VPB.t2 556.386
R17 VPB.t12 VPB.t7 301.87
R18 VPB.t7 VPB.t0 272.274
R19 VPB.t11 VPB.t12 260.437
R20 VPB.t8 VPB.t4 248.599
R21 VPB.t2 VPB.t6 213.084
R22 VPB VPB.t8 142.056
R23 VPB.t3 VPB.t10 18.7604
R24 VPB.t1 VPB.t9 10.959
R25 VPB.t9 VPB.t3 8.25484
R26 a_27_47.n3 a_27_47.t2 443.44
R27 a_27_47.t0 a_27_47.n6 390.443
R28 a_27_47.n4 a_27_47.t5 344.428
R29 a_27_47.n4 a_27_47.t3 296.969
R30 a_27_47.n1 a_27_47.t1 288.373
R31 a_27_47.n0 a_27_47.t6 263.406
R32 a_27_47.n3 a_27_47.n2 254.389
R33 a_27_47.n0 a_27_47.t4 228.06
R34 a_27_47.n5 a_27_47.n3 194.501
R35 a_27_47.n1 a_27_47.n0 152
R36 a_27_47.n6 a_27_47.n1 35.3396
R37 a_27_47.n6 a_27_47.n5 15.3376
R38 a_27_47.n5 a_27_47.n4 12.879
R39 VNB.t3 VNB.t15 4029.77
R40 VNB.t12 VNB.t6 3203.88
R41 VNB.t5 VNB.t8 3066.59
R42 VNB.t7 VNB.t3 2890.61
R43 VNB.t6 VNB.t7 2677.02
R44 VNB.t13 VNB.t16 2677.02
R45 VNB.t2 VNB.t4 2677.02
R46 VNB.t0 VNB.t1 2318.4
R47 VNB.t9 VNB.t11 1452.43
R48 VNB.t15 VNB.t14 1381.23
R49 VNB.t1 VNB.t12 1253.07
R50 VNB.t16 VNB.t9 1253.07
R51 VNB.t11 VNB.t5 1196.12
R52 VNB.t17 VNB.t2 1196.12
R53 VNB.t8 VNB.t10 1103.28
R54 VNB.t4 VNB.t13 1025.24
R55 VNB.t10 VNB.t0 945.673
R56 VNB VNB.t17 683.495
R57 a_1446_413.n3 a_1446_413.n2 680.737
R58 a_1446_413.n2 a_1446_413.n1 276.272
R59 a_1446_413.n0 a_1446_413.t5 230.484
R60 a_1446_413.n0 a_1446_413.t4 196.013
R61 a_1446_413.n2 a_1446_413.n0 171.939
R62 a_1446_413.t1 a_1446_413.n3 72.7029
R63 a_1446_413.n3 a_1446_413.t3 70.3576
R64 a_1446_413.n1 a_1446_413.t2 51.6672
R65 a_1446_413.n1 a_1446_413.t0 45.0005
R66 a_1537_413.t0 a_1537_413.t1 171.202
R67 DE.n0 DE.t2 319.728
R68 DE.n2 DE.n1 238.69
R69 DE.n0 DE.t0 178.34
R70 DE DE.n2 158.893
R71 DE.n1 DE.n0 147.814
R72 DE.n2 DE.t3 130.387
R73 DE.n1 DE.t1 130.141
R74 a_423_343.t0 a_423_343.n1 376.974
R75 a_423_343.n1 a_423_343.t3 375.568
R76 a_423_343.n0 a_423_343.t2 334.038
R77 a_423_343.n0 a_423_343.t1 244.181
R78 a_423_343.n1 a_423_343.n0 11.1343
R79 VPWR.n18 VPWR.t1 671.345
R80 VPWR.n25 VPWR.t2 667.963
R81 VPWR.n37 VPWR.t5 659.122
R82 VPWR.n52 VPWR.n1 604.394
R83 VPWR.n46 VPWR.t6 374.937
R84 VPWR.n44 VPWR.n5 323.079
R85 VPWR.n12 VPWR.n11 317.757
R86 VPWR.n17 VPWR.n16 246.773
R87 VPWR.n11 VPWR.t4 106.1
R88 VPWR.n16 VPWR.t11 61.9802
R89 VPWR.n5 VPWR.t7 44.6333
R90 VPWR.n5 VPWR.t8 44.6333
R91 VPWR.n11 VPWR.t3 43.3405
R92 VPWR.n1 VPWR.t0 41.5552
R93 VPWR.n1 VPWR.t9 41.5552
R94 VPWR.n50 VPWR.n2 34.6358
R95 VPWR.n51 VPWR.n50 34.6358
R96 VPWR.n39 VPWR.n38 34.6358
R97 VPWR.n39 VPWR.n6 34.6358
R98 VPWR.n43 VPWR.n6 34.6358
R99 VPWR.n31 VPWR.n30 34.6358
R100 VPWR.n32 VPWR.n31 34.6358
R101 VPWR.n32 VPWR.n9 34.6358
R102 VPWR.n36 VPWR.n9 34.6358
R103 VPWR.n20 VPWR.n19 34.6358
R104 VPWR.n20 VPWR.n14 34.6358
R105 VPWR.n24 VPWR.n14 34.6358
R106 VPWR.n44 VPWR.n43 33.8829
R107 VPWR.n46 VPWR.n45 32.0005
R108 VPWR.n16 VPWR.t10 30.1762
R109 VPWR.n26 VPWR.n25 30.1181
R110 VPWR.n38 VPWR.n37 28.2358
R111 VPWR.n30 VPWR.n12 28.2358
R112 VPWR.n26 VPWR.n12 23.3417
R113 VPWR.n52 VPWR.n51 22.9652
R114 VPWR.n18 VPWR.n17 21.2697
R115 VPWR.n45 VPWR.n44 20.7064
R116 VPWR.n25 VPWR.n24 17.3181
R117 VPWR.n37 VPWR.n36 15.0593
R118 VPWR.n46 VPWR.n2 12.424
R119 VPWR.n19 VPWR.n15 9.3005
R120 VPWR.n21 VPWR.n20 9.3005
R121 VPWR.n22 VPWR.n14 9.3005
R122 VPWR.n24 VPWR.n23 9.3005
R123 VPWR.n25 VPWR.n13 9.3005
R124 VPWR.n27 VPWR.n26 9.3005
R125 VPWR.n28 VPWR.n12 9.3005
R126 VPWR.n30 VPWR.n29 9.3005
R127 VPWR.n31 VPWR.n10 9.3005
R128 VPWR.n33 VPWR.n32 9.3005
R129 VPWR.n34 VPWR.n9 9.3005
R130 VPWR.n36 VPWR.n35 9.3005
R131 VPWR.n37 VPWR.n8 9.3005
R132 VPWR.n38 VPWR.n7 9.3005
R133 VPWR.n40 VPWR.n39 9.3005
R134 VPWR.n41 VPWR.n6 9.3005
R135 VPWR.n43 VPWR.n42 9.3005
R136 VPWR.n44 VPWR.n4 9.3005
R137 VPWR.n45 VPWR.n3 9.3005
R138 VPWR.n47 VPWR.n46 9.3005
R139 VPWR.n48 VPWR.n2 9.3005
R140 VPWR.n50 VPWR.n49 9.3005
R141 VPWR.n51 VPWR.n0 9.3005
R142 VPWR.n53 VPWR.n52 7.12063
R143 VPWR.n17 VPWR.n15 0.754043
R144 VPWR.n19 VPWR.n18 0.753441
R145 VPWR.n53 VPWR.n0 0.148519
R146 VPWR.n21 VPWR.n15 0.120292
R147 VPWR.n22 VPWR.n21 0.120292
R148 VPWR.n23 VPWR.n22 0.120292
R149 VPWR.n23 VPWR.n13 0.120292
R150 VPWR.n27 VPWR.n13 0.120292
R151 VPWR.n28 VPWR.n27 0.120292
R152 VPWR.n29 VPWR.n28 0.120292
R153 VPWR.n29 VPWR.n10 0.120292
R154 VPWR.n33 VPWR.n10 0.120292
R155 VPWR.n34 VPWR.n33 0.120292
R156 VPWR.n35 VPWR.n34 0.120292
R157 VPWR.n35 VPWR.n8 0.120292
R158 VPWR.n8 VPWR.n7 0.120292
R159 VPWR.n40 VPWR.n7 0.120292
R160 VPWR.n41 VPWR.n40 0.120292
R161 VPWR.n42 VPWR.n41 0.120292
R162 VPWR.n42 VPWR.n4 0.120292
R163 VPWR.n4 VPWR.n3 0.120292
R164 VPWR.n47 VPWR.n3 0.120292
R165 VPWR.n48 VPWR.n47 0.120292
R166 VPWR.n49 VPWR.n48 0.120292
R167 VPWR.n49 VPWR.n0 0.120292
R168 VPWR VPWR.n53 0.114842
R169 CLK.n0 CLK.t0 292.95
R170 CLK.n0 CLK.t1 209.403
R171 CLK CLK.n0 154.069
R172 SCE.t1 SCE.t2 604.107
R173 SCE.n1 SCE.t3 352.397
R174 SCE.n0 SCE.t0 189.588
R175 SCE SCE.n1 153.631
R176 SCE.n0 SCE.t1 142.03
R177 SCE.n1 SCE.n0 74.0857
R178 a_885_21.n0 a_885_21.t2 571.547
R179 a_885_21.n2 a_885_21.n1 427.555
R180 a_885_21.t0 a_885_21.n2 372.423
R181 a_885_21.n0 a_885_21.t1 223.571
R182 a_885_21.n2 a_885_21.n0 74.941
R183 VGND.n17 VGND.t2 273.476
R184 VGND.n11 VGND.t3 244.518
R185 VGND.n38 VGND.t7 238.311
R186 VGND.n25 VGND.n24 222.888
R187 VGND.n36 VGND.n4 202.262
R188 VGND.n45 VGND.n44 199.739
R189 VGND.n13 VGND.n12 125.585
R190 VGND.n12 VGND.t8 57.8184
R191 VGND.n4 VGND.t5 41.4291
R192 VGND.n4 VGND.t6 41.4291
R193 VGND.n24 VGND.t4 38.5719
R194 VGND.n24 VGND.t0 38.5719
R195 VGND.n44 VGND.t1 38.5719
R196 VGND.n44 VGND.t10 38.5719
R197 VGND.n16 VGND.n10 34.6358
R198 VGND.n18 VGND.n8 34.6358
R199 VGND.n22 VGND.n8 34.6358
R200 VGND.n23 VGND.n22 34.6358
R201 VGND.n26 VGND.n23 34.6358
R202 VGND.n30 VGND.n6 34.6358
R203 VGND.n31 VGND.n30 34.6358
R204 VGND.n32 VGND.n31 34.6358
R205 VGND.n32 VGND.n3 34.6358
R206 VGND.n42 VGND.n1 34.6358
R207 VGND.n43 VGND.n42 34.6358
R208 VGND.n38 VGND.n37 32.0005
R209 VGND.n36 VGND.n3 29.7417
R210 VGND.n17 VGND.n16 24.8476
R211 VGND.n12 VGND.t9 24.7498
R212 VGND.n45 VGND.n43 22.9652
R213 VGND.n13 VGND.n11 18.8938
R214 VGND.n26 VGND.n25 15.0593
R215 VGND.n18 VGND.n17 14.6829
R216 VGND.n37 VGND.n36 14.6829
R217 VGND.n38 VGND.n1 12.424
R218 VGND.n43 VGND.n0 9.3005
R219 VGND.n42 VGND.n41 9.3005
R220 VGND.n40 VGND.n1 9.3005
R221 VGND.n39 VGND.n38 9.3005
R222 VGND.n37 VGND.n2 9.3005
R223 VGND.n36 VGND.n35 9.3005
R224 VGND.n34 VGND.n3 9.3005
R225 VGND.n33 VGND.n32 9.3005
R226 VGND.n31 VGND.n5 9.3005
R227 VGND.n30 VGND.n29 9.3005
R228 VGND.n28 VGND.n6 9.3005
R229 VGND.n14 VGND.n10 9.3005
R230 VGND.n16 VGND.n15 9.3005
R231 VGND.n17 VGND.n9 9.3005
R232 VGND.n19 VGND.n18 9.3005
R233 VGND.n20 VGND.n8 9.3005
R234 VGND.n22 VGND.n21 9.3005
R235 VGND.n23 VGND.n7 9.3005
R236 VGND.n27 VGND.n26 9.3005
R237 VGND.n46 VGND.n45 7.12063
R238 VGND.n11 VGND.n10 2.63579
R239 VGND.n25 VGND.n6 0.753441
R240 VGND.n14 VGND.n13 0.148563
R241 VGND.n46 VGND.n0 0.148519
R242 VGND.n15 VGND.n14 0.120292
R243 VGND.n15 VGND.n9 0.120292
R244 VGND.n19 VGND.n9 0.120292
R245 VGND.n20 VGND.n19 0.120292
R246 VGND.n21 VGND.n20 0.120292
R247 VGND.n21 VGND.n7 0.120292
R248 VGND.n27 VGND.n7 0.120292
R249 VGND.n28 VGND.n27 0.120292
R250 VGND.n29 VGND.n28 0.120292
R251 VGND.n29 VGND.n5 0.120292
R252 VGND.n33 VGND.n5 0.120292
R253 VGND.n34 VGND.n33 0.120292
R254 VGND.n35 VGND.n34 0.120292
R255 VGND.n35 VGND.n2 0.120292
R256 VGND.n39 VGND.n2 0.120292
R257 VGND.n40 VGND.n39 0.120292
R258 VGND.n41 VGND.n40 0.120292
R259 VGND.n41 VGND.n0 0.120292
R260 VGND VGND.n46 0.114842
R261 a_1610_159.t0 a_1610_159.n4 408.848
R262 a_1610_159.n2 a_1610_159.t2 406.401
R263 a_1610_159.n0 a_1610_159.t4 318.12
R264 a_1610_159.n0 a_1610_159.t3 194.477
R265 a_1610_159.n3 a_1610_159.n2 176.534
R266 a_1610_159.n4 a_1610_159.n0 168.486
R267 a_1610_159.n3 a_1610_159.t1 140.249
R268 a_1610_159.n2 a_1610_159.n1 130.054
R269 a_1610_159.n4 a_1610_159.n3 9.32396
R270 a_791_264.n3 a_791_264.n2 382.745
R271 a_791_264.t0 a_791_264.n4 362.808
R272 a_791_264.n0 a_791_264.t2 310.623
R273 a_791_264.n1 a_791_264.t1 242.322
R274 a_791_264.n1 a_791_264.n0 220.962
R275 a_791_264.n0 a_791_264.t3 194.942
R276 a_791_264.n4 a_791_264.n3 174.017
R277 a_791_264.n3 a_791_264.t4 138.53
R278 a_791_264.n4 a_791_264.n1 48.371
R279 a_193_47.t0 a_193_47.n4 395.625
R280 a_193_47.n2 a_193_47.t2 389.545
R281 a_193_47.n1 a_193_47.t3 308.651
R282 a_193_47.n4 a_193_47.t1 300.372
R283 a_193_47.n1 a_193_47.n0 298.373
R284 a_193_47.n2 a_193_47.t4 273.572
R285 a_193_47.n3 a_193_47.n2 173.755
R286 a_193_47.n4 a_193_47.n3 14.6322
R287 a_193_47.n3 a_193_47.n1 12.2528
R288 a_1974_47.n0 a_1974_47.t0 45.1697
R289 a_729_47.t0 a_729_47.t1 102.858
R290 a_729_369.t0 a_729_369.t1 110.812
R291 Q Q.t0 251.107
R292 Q Q.t1 146.542
R293 a_2135_413.t0 a_2135_413.t1 197
R294 SCD.n1 SCD.t0 206.19
R295 SCD.n1 SCD.n0 183.696
R296 SCD SCD.n1 163.675
R297 a_1226_119.t0 a_1226_119.t1 60.0005
R298 a_381_47.t0 a_381_47.t1 60.0005
C0 VPWR DE 0.04692f
C1 VPWR VPB 0.295394f
C2 VPWR a_1960_413# 0.007488f
C3 VPB DE 0.114449f
C4 VPWR a_915_47# 0.097411f
C5 VPB a_915_47# 0.021894f
C6 Q a_2051_413# 0.036123f
C7 VGND Q 0.092175f
C8 Q SCE 1.95e-20
C9 VGND SCD 0.032521f
C10 VGND D 0.014495f
C11 VGND a_1561_47# 0.004442f
C12 SCE SCD 0.095395f
C13 VGND a_2051_413# 0.173214f
C14 SCE a_2051_413# 8.01e-20
C15 a_2177_47# a_2051_413# 0.006472f
C16 VPWR Q 0.122606f
C17 VPWR SCD 0.013425f
C18 VGND SCE 0.047517f
C19 Q VPB 0.013891f
C20 VPWR D 0.01674f
C21 VGND CLK 0.019296f
C22 VGND a_2177_47# 0.004743f
C23 D DE 0.099354f
C24 VPB SCD 0.045339f
C25 VPB D 0.068631f
C26 Q a_915_47# 3.29e-20
C27 VPWR a_2051_413# 0.160369f
C28 SCD a_915_47# 0.018533f
C29 VPB a_2051_413# 0.147526f
C30 a_1561_47# a_915_47# 4.9e-19
C31 a_1960_413# a_2051_413# 0.002082f
C32 a_2051_413# a_915_47# 2.43e-19
C33 VPWR VGND 0.05975f
C34 VPWR SCE 0.028732f
C35 VGND DE 0.057232f
C36 VPWR CLK 0.019263f
C37 VGND VPB 0.012131f
C38 VGND a_1960_413# 2.3e-19
C39 VPB SCE 0.1417f
C40 VPB CLK 0.069635f
C41 VGND a_915_47# 0.383397f
C42 VPWR a_1231_369# 0.0081f
C43 SCE a_915_47# 0.086615f
C44 a_2177_47# a_915_47# 5.05e-20
C45 a_915_47# a_1231_369# 0.003336f
C46 Q VNB 0.084065f
C47 VGND VNB 1.46617f
C48 VPWR VNB 1.18094f
C49 SCD VNB 0.08884f
C50 SCE VNB 0.334233f
C51 DE VNB 0.282831f
C52 D VNB 0.122269f
C53 CLK VNB 0.195128f
C54 VPB VNB 2.60636f
C55 a_915_47# VNB 0.03825f
C56 a_2051_413# VNB 0.312829f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxtp_2 VPWR VGND CLK SCD DE Q D SCE VPB VNB
X0 a_381_369.t1 D.t0 a_299_47.t5 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_2177_47# a_27_47.t2 a_2051_413# VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2 a_1537_413.t0 a_27_47.t3 a_1446_413.t1 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 VPWR.t2 DE.t0 a_423_343.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VPWR.t7 CLK.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t0 SCE.t0 a_885_21.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1264 pd=1.035 as=0.1696 ps=1.81 w=0.64 l=0.15
X6 VGND.t7 SCE.t1 a_885_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR.t8 a_1610_159.t2 a_1537_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8 a_1610_159.t1 a_1446_413.t4 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X9 VGND.t6 a_2051_413# a_791_264.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND.t3 DE.t1 a_423_343.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_1561_47# a_193_47.t2 a_1446_413.t2 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X12 a_1974_47.t0 a_1610_159.t3 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 VGND.t4 a_2051_413# Q.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_193_47.t0 a_27_47.t4 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_729_47.t1 a_423_343.t2 VGND.t10 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X16 a_729_369.t0 DE.t2 VPWR.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X17 Q.t0 a_2051_413# VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X18 a_299_47.t1 a_791_264.t2 a_729_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0756 ps=0.78 w=0.42 l=0.15
X19 a_2135_413.t0 a_193_47.t3 a_2051_413# VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1446_413.t0 a_27_47.t5 a_915_47.t0 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.22515 ps=1.505 w=0.36 l=0.15
X21 a_193_47.t1 a_27_47.t6 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1231_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1056 pd=0.97 as=0.1264 ps=1.035 w=0.64 l=0.15
X23 a_915_47.t2 SCE.t2 a_1226_119.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.22515 pd=1.505 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 VPWR.t4 a_2051_413# Q.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X25 a_299_47.t2 a_791_264.t3 a_729_369.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0992 pd=0.95 as=0.1152 ps=1 w=0.64 l=0.15
X26 a_381_47.t1 D.t1 a_299_47.t4 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR.t12 a_791_264.t4 a_2135_413.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X28 Q.t2 a_2051_413# VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X29 VPWR.t10 a_423_343.t3 a_381_369.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X30 a_915_47.t3 SCE.t3 a_299_47.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1984 pd=1.9 as=0.0992 ps=0.95 w=0.64 l=0.15
X31 a_1960_413# a_1610_159.t4 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_1226_119.t0 SCD.t0 VGND.t8 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X33 a_1446_413.t3 a_193_47.t4 a_915_47.t1 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.13415 ps=1.085 w=0.42 l=0.15
X34 a_915_47.t4 a_885_21.t2 a_299_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X35 VPWR.t5 a_2051_413# a_791_264.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1728 ps=1.82 w=0.64 l=0.15
X36 VGND.t1 CLK.t1 a_27_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 VGND.t2 DE.t3 a_381_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X38 a_1610_159.t0 a_1446_413.t5 VGND.t11 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
R0 D.n0 D.t1 220.367
R1 D.n0 D.t0 216.796
R2 D D.n0 71.33
R3 a_299_47.n1 a_299_47.t5 467.892
R4 a_299_47.n3 a_299_47.n2 380.248
R5 a_299_47.n1 a_299_47.t4 232.434
R6 a_299_47.n2 a_299_47.n0 188.082
R7 a_299_47.n3 a_299_47.t3 53.8677
R8 a_299_47.t2 a_299_47.n3 41.5552
R9 a_299_47.n0 a_299_47.t0 38.5719
R10 a_299_47.n0 a_299_47.t1 38.5719
R11 a_299_47.n2 a_299_47.n1 20.4743
R12 a_381_369.t0 a_381_369.t1 64.6411
R13 VPB.t0 VPB.t18 1043.39
R14 VPB.t16 VPB.t6 624.456
R15 VPB.t13 VPB.t0 622.851
R16 VPB.t14 VPB.t12 556.386
R17 VPB.t10 VPB.t5 556.386
R18 VPB.t4 VPB.t15 556.386
R19 VPB.t12 VPB.t2 517.913
R20 VPB.t11 VPB.t14 390.654
R21 VPB.t2 VPB.t16 337.384
R22 VPB.t17 VPB.t11 304.829
R23 VPB.t1 VPB.t3 301.87
R24 VPB.t6 VPB.t7 287.072
R25 VPB.t3 VPB.t13 272.274
R26 VPB.t5 VPB.t1 260.437
R27 VPB.t18 VPB.t17 256.56
R28 VPB.t7 VPB.t8 248.599
R29 VPB.t9 VPB.t4 248.599
R30 VPB.t15 VPB.t10 213.084
R31 VPB VPB.t9 142.056
R32 a_27_47.n3 a_27_47.t2 443.44
R33 a_27_47.t1 a_27_47.n6 390.443
R34 a_27_47.n4 a_27_47.t5 344.428
R35 a_27_47.n4 a_27_47.t3 296.969
R36 a_27_47.n1 a_27_47.t0 288.373
R37 a_27_47.n0 a_27_47.t6 263.406
R38 a_27_47.n3 a_27_47.n2 254.389
R39 a_27_47.n0 a_27_47.t4 228.06
R40 a_27_47.n5 a_27_47.n3 194.501
R41 a_27_47.n1 a_27_47.n0 152
R42 a_27_47.n6 a_27_47.n1 35.3396
R43 a_27_47.n6 a_27_47.n5 15.3376
R44 a_27_47.n5 a_27_47.n4 12.879
R45 VNB.t4 VNB.t12 4029.77
R46 VNB.t8 VNB.t17 3203.88
R47 VNB.t0 VNB.t1 3066.59
R48 VNB.t15 VNB.t4 2890.61
R49 VNB.t17 VNB.t15 2677.02
R50 VNB.t7 VNB.t6 2677.02
R51 VNB.t3 VNB.t18 2677.02
R52 VNB.t16 VNB.t2 2318.4
R53 VNB.t13 VNB.t9 1452.43
R54 VNB.t12 VNB.t10 1381.23
R55 VNB.t2 VNB.t8 1253.07
R56 VNB.t6 VNB.t13 1253.07
R57 VNB.t10 VNB.t11 1196.12
R58 VNB.t9 VNB.t0 1196.12
R59 VNB.t5 VNB.t3 1196.12
R60 VNB.t1 VNB.t14 1103.28
R61 VNB.t18 VNB.t7 1025.24
R62 VNB.t14 VNB.t16 945.673
R63 VNB VNB.t5 683.495
R64 a_1446_413.n3 a_1446_413.n2 680.737
R65 a_1446_413.n2 a_1446_413.n1 276.272
R66 a_1446_413.n0 a_1446_413.t5 230.484
R67 a_1446_413.n0 a_1446_413.t4 196.013
R68 a_1446_413.n2 a_1446_413.n0 171.939
R69 a_1446_413.t1 a_1446_413.n3 72.7029
R70 a_1446_413.n3 a_1446_413.t3 70.3576
R71 a_1446_413.n1 a_1446_413.t2 51.6672
R72 a_1446_413.n1 a_1446_413.t0 45.0005
R73 a_1537_413.t0 a_1537_413.t1 171.202
R74 DE.n0 DE.t2 319.728
R75 DE.n2 DE.n1 238.69
R76 DE.n0 DE.t0 178.34
R77 DE DE.n2 158.893
R78 DE.n1 DE.n0 147.814
R79 DE.n2 DE.t3 130.387
R80 DE.n1 DE.t1 130.141
R81 a_423_343.t0 a_423_343.n1 376.974
R82 a_423_343.n1 a_423_343.t3 375.568
R83 a_423_343.n0 a_423_343.t2 334.038
R84 a_423_343.n0 a_423_343.t1 244.181
R85 a_423_343.n1 a_423_343.n0 11.1343
R86 VPWR.n23 VPWR.t12 671.345
R87 VPWR.n30 VPWR.t9 667.963
R88 VPWR.n42 VPWR.t0 659.122
R89 VPWR.n57 VPWR.n1 604.394
R90 VPWR.n51 VPWR.t10 374.937
R91 VPWR.n49 VPWR.n5 323.079
R92 VPWR.n12 VPWR.n11 317.757
R93 VPWR.n19 VPWR.t4 260.05
R94 VPWR.n18 VPWR.n17 241.126
R95 VPWR.n11 VPWR.t8 106.1
R96 VPWR.n17 VPWR.t5 61.9796
R97 VPWR.n5 VPWR.t3 44.6333
R98 VPWR.n5 VPWR.t2 44.6333
R99 VPWR.n11 VPWR.t11 43.3405
R100 VPWR.n1 VPWR.t1 41.5552
R101 VPWR.n1 VPWR.t7 41.5552
R102 VPWR.n55 VPWR.n2 34.6358
R103 VPWR.n56 VPWR.n55 34.6358
R104 VPWR.n44 VPWR.n43 34.6358
R105 VPWR.n44 VPWR.n6 34.6358
R106 VPWR.n48 VPWR.n6 34.6358
R107 VPWR.n36 VPWR.n35 34.6358
R108 VPWR.n37 VPWR.n36 34.6358
R109 VPWR.n37 VPWR.n9 34.6358
R110 VPWR.n41 VPWR.n9 34.6358
R111 VPWR.n25 VPWR.n24 34.6358
R112 VPWR.n25 VPWR.n14 34.6358
R113 VPWR.n29 VPWR.n14 34.6358
R114 VPWR.n22 VPWR.n16 34.6358
R115 VPWR.n49 VPWR.n48 33.8829
R116 VPWR.n51 VPWR.n50 32.0005
R117 VPWR.n17 VPWR.t6 30.1768
R118 VPWR.n31 VPWR.n30 30.1181
R119 VPWR.n43 VPWR.n42 28.2358
R120 VPWR.n35 VPWR.n12 28.2358
R121 VPWR.n31 VPWR.n12 23.3417
R122 VPWR.n57 VPWR.n56 22.9652
R123 VPWR.n50 VPWR.n49 20.7064
R124 VPWR.n30 VPWR.n29 17.3181
R125 VPWR.n42 VPWR.n41 15.0593
R126 VPWR.n23 VPWR.n22 14.3064
R127 VPWR.n51 VPWR.n2 12.424
R128 VPWR.n18 VPWR.n16 12.0476
R129 VPWR.n19 VPWR.n18 11.7868
R130 VPWR.n20 VPWR.n16 9.3005
R131 VPWR.n22 VPWR.n21 9.3005
R132 VPWR.n24 VPWR.n15 9.3005
R133 VPWR.n26 VPWR.n25 9.3005
R134 VPWR.n27 VPWR.n14 9.3005
R135 VPWR.n29 VPWR.n28 9.3005
R136 VPWR.n30 VPWR.n13 9.3005
R137 VPWR.n32 VPWR.n31 9.3005
R138 VPWR.n33 VPWR.n12 9.3005
R139 VPWR.n35 VPWR.n34 9.3005
R140 VPWR.n36 VPWR.n10 9.3005
R141 VPWR.n38 VPWR.n37 9.3005
R142 VPWR.n39 VPWR.n9 9.3005
R143 VPWR.n41 VPWR.n40 9.3005
R144 VPWR.n42 VPWR.n8 9.3005
R145 VPWR.n43 VPWR.n7 9.3005
R146 VPWR.n45 VPWR.n44 9.3005
R147 VPWR.n46 VPWR.n6 9.3005
R148 VPWR.n48 VPWR.n47 9.3005
R149 VPWR.n49 VPWR.n4 9.3005
R150 VPWR.n50 VPWR.n3 9.3005
R151 VPWR.n52 VPWR.n51 9.3005
R152 VPWR.n53 VPWR.n2 9.3005
R153 VPWR.n55 VPWR.n54 9.3005
R154 VPWR.n56 VPWR.n0 9.3005
R155 VPWR.n58 VPWR.n57 7.12063
R156 VPWR.n20 VPWR.n19 0.826395
R157 VPWR.n24 VPWR.n23 0.753441
R158 VPWR.n58 VPWR.n0 0.148519
R159 VPWR.n21 VPWR.n20 0.120292
R160 VPWR.n21 VPWR.n15 0.120292
R161 VPWR.n26 VPWR.n15 0.120292
R162 VPWR.n27 VPWR.n26 0.120292
R163 VPWR.n28 VPWR.n27 0.120292
R164 VPWR.n28 VPWR.n13 0.120292
R165 VPWR.n32 VPWR.n13 0.120292
R166 VPWR.n33 VPWR.n32 0.120292
R167 VPWR.n34 VPWR.n33 0.120292
R168 VPWR.n34 VPWR.n10 0.120292
R169 VPWR.n38 VPWR.n10 0.120292
R170 VPWR.n39 VPWR.n38 0.120292
R171 VPWR.n40 VPWR.n39 0.120292
R172 VPWR.n40 VPWR.n8 0.120292
R173 VPWR.n8 VPWR.n7 0.120292
R174 VPWR.n45 VPWR.n7 0.120292
R175 VPWR.n46 VPWR.n45 0.120292
R176 VPWR.n47 VPWR.n46 0.120292
R177 VPWR.n47 VPWR.n4 0.120292
R178 VPWR.n4 VPWR.n3 0.120292
R179 VPWR.n52 VPWR.n3 0.120292
R180 VPWR.n53 VPWR.n52 0.120292
R181 VPWR.n54 VPWR.n53 0.120292
R182 VPWR.n54 VPWR.n0 0.120292
R183 VPWR VPWR.n58 0.114842
R184 CLK.n0 CLK.t0 292.95
R185 CLK.n0 CLK.t1 209.403
R186 CLK CLK.n0 154.069
R187 SCE.t1 SCE.t2 604.107
R188 SCE.n1 SCE.t3 352.397
R189 SCE.n0 SCE.t0 189.588
R190 SCE SCE.n1 153.631
R191 SCE.n0 SCE.t1 142.03
R192 SCE.n1 SCE.n0 74.0857
R193 a_885_21.n0 a_885_21.t2 571.547
R194 a_885_21.n2 a_885_21.n1 427.555
R195 a_885_21.t1 a_885_21.n2 372.423
R196 a_885_21.n0 a_885_21.t0 223.571
R197 a_885_21.n2 a_885_21.n0 74.941
R198 VGND.n30 VGND.t11 273.476
R199 VGND.n24 VGND.t9 244.518
R200 VGND.n51 VGND.t2 238.311
R201 VGND.n38 VGND.n37 222.888
R202 VGND.n49 VGND.n4 202.262
R203 VGND.n58 VGND.n57 199.739
R204 VGND.n14 VGND.t4 158.339
R205 VGND.n16 VGND.n15 118.657
R206 VGND.n15 VGND.t6 57.8171
R207 VGND.n4 VGND.t10 41.4291
R208 VGND.n4 VGND.t3 41.4291
R209 VGND.n37 VGND.t8 38.5719
R210 VGND.n37 VGND.t7 38.5719
R211 VGND.n57 VGND.t0 38.5719
R212 VGND.n57 VGND.t1 38.5719
R213 VGND.n18 VGND.n17 34.6358
R214 VGND.n22 VGND.n12 34.6358
R215 VGND.n23 VGND.n22 34.6358
R216 VGND.n25 VGND.n23 34.6358
R217 VGND.n29 VGND.n10 34.6358
R218 VGND.n31 VGND.n8 34.6358
R219 VGND.n35 VGND.n8 34.6358
R220 VGND.n36 VGND.n35 34.6358
R221 VGND.n39 VGND.n36 34.6358
R222 VGND.n43 VGND.n6 34.6358
R223 VGND.n44 VGND.n43 34.6358
R224 VGND.n45 VGND.n44 34.6358
R225 VGND.n45 VGND.n3 34.6358
R226 VGND.n55 VGND.n1 34.6358
R227 VGND.n56 VGND.n55 34.6358
R228 VGND.n51 VGND.n50 32.0005
R229 VGND.n49 VGND.n3 29.7417
R230 VGND.n30 VGND.n29 24.8476
R231 VGND.n15 VGND.t5 24.7511
R232 VGND.n58 VGND.n56 22.9652
R233 VGND.n39 VGND.n38 15.0593
R234 VGND.n31 VGND.n30 14.6829
R235 VGND.n50 VGND.n49 14.6829
R236 VGND.n51 VGND.n1 12.424
R237 VGND.n17 VGND.n16 12.0476
R238 VGND.n16 VGND.n14 11.7868
R239 VGND.n25 VGND.n24 11.2946
R240 VGND.n18 VGND.n12 10.9181
R241 VGND.n56 VGND.n0 9.3005
R242 VGND.n55 VGND.n54 9.3005
R243 VGND.n53 VGND.n1 9.3005
R244 VGND.n52 VGND.n51 9.3005
R245 VGND.n50 VGND.n2 9.3005
R246 VGND.n49 VGND.n48 9.3005
R247 VGND.n47 VGND.n3 9.3005
R248 VGND.n46 VGND.n45 9.3005
R249 VGND.n44 VGND.n5 9.3005
R250 VGND.n43 VGND.n42 9.3005
R251 VGND.n41 VGND.n6 9.3005
R252 VGND.n17 VGND.n13 9.3005
R253 VGND.n19 VGND.n18 9.3005
R254 VGND.n20 VGND.n12 9.3005
R255 VGND.n22 VGND.n21 9.3005
R256 VGND.n23 VGND.n11 9.3005
R257 VGND.n26 VGND.n25 9.3005
R258 VGND.n27 VGND.n10 9.3005
R259 VGND.n29 VGND.n28 9.3005
R260 VGND.n30 VGND.n9 9.3005
R261 VGND.n32 VGND.n31 9.3005
R262 VGND.n33 VGND.n8 9.3005
R263 VGND.n35 VGND.n34 9.3005
R264 VGND.n36 VGND.n7 9.3005
R265 VGND.n40 VGND.n39 9.3005
R266 VGND.n59 VGND.n58 7.12063
R267 VGND.n24 VGND.n10 2.63579
R268 VGND.n14 VGND.n13 0.826395
R269 VGND.n38 VGND.n6 0.753441
R270 VGND.n59 VGND.n0 0.148519
R271 VGND.n19 VGND.n13 0.120292
R272 VGND.n20 VGND.n19 0.120292
R273 VGND.n21 VGND.n20 0.120292
R274 VGND.n21 VGND.n11 0.120292
R275 VGND.n26 VGND.n11 0.120292
R276 VGND.n27 VGND.n26 0.120292
R277 VGND.n28 VGND.n27 0.120292
R278 VGND.n28 VGND.n9 0.120292
R279 VGND.n32 VGND.n9 0.120292
R280 VGND.n33 VGND.n32 0.120292
R281 VGND.n34 VGND.n33 0.120292
R282 VGND.n34 VGND.n7 0.120292
R283 VGND.n40 VGND.n7 0.120292
R284 VGND.n41 VGND.n40 0.120292
R285 VGND.n42 VGND.n41 0.120292
R286 VGND.n42 VGND.n5 0.120292
R287 VGND.n46 VGND.n5 0.120292
R288 VGND.n47 VGND.n46 0.120292
R289 VGND.n48 VGND.n47 0.120292
R290 VGND.n48 VGND.n2 0.120292
R291 VGND.n52 VGND.n2 0.120292
R292 VGND.n53 VGND.n52 0.120292
R293 VGND.n54 VGND.n53 0.120292
R294 VGND.n54 VGND.n0 0.120292
R295 VGND VGND.n59 0.114842
R296 a_1610_159.t1 a_1610_159.n4 408.848
R297 a_1610_159.n2 a_1610_159.t2 406.401
R298 a_1610_159.n0 a_1610_159.t4 318.12
R299 a_1610_159.n0 a_1610_159.t3 194.477
R300 a_1610_159.n3 a_1610_159.n2 176.534
R301 a_1610_159.n4 a_1610_159.n0 168.486
R302 a_1610_159.n3 a_1610_159.t0 140.249
R303 a_1610_159.n2 a_1610_159.n1 130.054
R304 a_1610_159.n4 a_1610_159.n3 9.32396
R305 a_791_264.n3 a_791_264.n2 382.745
R306 a_791_264.t1 a_791_264.n4 362.808
R307 a_791_264.n0 a_791_264.t2 310.623
R308 a_791_264.n1 a_791_264.t0 242.322
R309 a_791_264.n1 a_791_264.n0 220.962
R310 a_791_264.n0 a_791_264.t3 194.942
R311 a_791_264.n4 a_791_264.n3 174.017
R312 a_791_264.n3 a_791_264.t4 138.53
R313 a_791_264.n4 a_791_264.n1 48.371
R314 a_193_47.t1 a_193_47.n4 395.625
R315 a_193_47.n2 a_193_47.t2 389.545
R316 a_193_47.n1 a_193_47.t3 308.651
R317 a_193_47.n4 a_193_47.t0 300.372
R318 a_193_47.n1 a_193_47.n0 298.373
R319 a_193_47.n2 a_193_47.t4 273.572
R320 a_193_47.n3 a_193_47.n2 173.755
R321 a_193_47.n4 a_193_47.n3 14.6322
R322 a_193_47.n3 a_193_47.n1 12.2528
R323 a_1974_47.n0 a_1974_47.t0 45.1697
R324 Q Q.n0 222.542
R325 Q Q.n1 110.037
R326 Q.n0 Q.t3 26.5955
R327 Q.n0 Q.t2 26.5955
R328 Q.n1 Q.t1 24.9236
R329 Q.n1 Q.t0 24.9236
R330 a_915_47.n0 a_915_47.t1 489.325
R331 a_915_47.t3 a_915_47.n4 452.894
R332 a_915_47.n4 a_915_47.t4 227.732
R333 a_915_47.n3 a_915_47.n2 189.981
R334 a_915_47.n1 a_915_47.n0 185
R335 a_915_47.n2 a_915_47.t0 75.3851
R336 a_915_47.n2 a_915_47.n1 51.539
R337 a_915_47.n1 a_915_47.t2 32.1983
R338 a_915_47.n4 a_915_47.n3 19.8561
R339 a_915_47.n3 a_915_47.n0 9.52245
R340 a_729_47.t0 a_729_47.t1 102.858
R341 a_729_369.t0 a_729_369.t1 110.812
R342 a_2135_413.t0 a_2135_413.t1 197
R343 SCD.n1 SCD.t0 206.19
R344 SCD.n1 SCD.n0 183.696
R345 SCD SCD.n1 163.675
R346 a_1226_119.t0 a_1226_119.t1 60.0005
R347 a_381_47.t0 a_381_47.t1 60.0005
C0 VPWR Q 0.203312f
C1 DE VGND 0.057232f
C2 D VPWR 0.01674f
C3 Q VPB 0.005361f
C4 VPWR VPB 0.314821f
C5 D VPB 0.068631f
C6 VPWR a_1960_413# 0.007488f
C7 VGND Q 0.142656f
C8 VPWR VGND 0.0823f
C9 D VGND 0.014495f
C10 SCD VPWR 0.013425f
C11 CLK VPWR 0.019263f
C12 VGND VPB 0.013793f
C13 a_1561_47# VGND 0.004442f
C14 a_1960_413# VGND 2.3e-19
C15 SCD VPB 0.045339f
C16 CLK VPB 0.069635f
C17 a_1231_369# VPWR 0.0081f
C18 Q a_2051_413# 0.075634f
C19 VPWR a_2051_413# 0.174159f
C20 a_2051_413# VPB 0.180229f
C21 a_1960_413# a_2051_413# 0.002082f
C22 SCE Q 1.96e-20
C23 SCD VGND 0.032521f
C24 CLK VGND 0.019296f
C25 SCE VPWR 0.028732f
C26 SCE VPB 0.1417f
C27 VGND a_2051_413# 0.186035f
C28 SCE VGND 0.047533f
C29 SCE SCD 0.095395f
C30 VGND a_2177_47# 0.004743f
C31 SCE a_2051_413# 8.01e-20
C32 DE VPWR 0.04692f
C33 D DE 0.099354f
C34 a_2051_413# a_2177_47# 0.006472f
C35 DE VPB 0.114449f
C36 Q VNB 0.022118f
C37 VGND VNB 1.54525f
C38 VPWR VNB 1.25646f
C39 SCD VNB 0.08884f
C40 SCE VNB 0.334233f
C41 DE VNB 0.282831f
C42 D VNB 0.122269f
C43 CLK VNB 0.195128f
C44 VPB VNB 2.69495f
C45 a_2051_413# VNB 0.402271f
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxtp_4 VPWR VGND CLK SCD DE Q D SCE VPB VNB
X0 a_381_369.t1 D.t0 a_299_47.t5 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_2177_47# a_27_47.t2 a_2051_413.t1 VNB.t19 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2 a_1537_413.t1 a_27_47.t3 a_1446_413.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 VPWR.t1 DE.t0 a_423_343.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t9 SCE.t0 a_885_21.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1264 pd=1.035 as=0.1696 ps=1.81 w=0.64 l=0.15
X6 VGND.t10 SCE.t1 a_885_21.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR.t11 a_1610_159.t2 a_1537_413.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8 a_1610_159.t0 a_1446_413.t4 VPWR.t10 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X9 VPWR.t5 a_2051_413.t2 Q.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t4 a_2051_413.t3 a_791_264.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND.t1 DE.t1 a_423_343.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_1561_47# a_193_47.t2 a_1446_413.t0 VNB.t14 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X13 a_1974_47.t0 a_1610_159.t3 VGND.t12 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 Q.t2 a_2051_413.t4 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t8 a_2051_413.t5 Q.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_193_47.t1 a_27_47.t4 VGND.t13 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_729_47.t0 a_423_343.t2 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X18 a_729_369.t0 DE.t2 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X19 Q.t6 a_2051_413.t6 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X20 a_299_47.t1 a_791_264.t2 a_729_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0756 ps=0.78 w=0.42 l=0.15
X21 a_2135_413.t1 a_193_47.t3 a_2051_413.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1446_413.t2 a_27_47.t5 a_915_47# VNB.t17 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.22515 ps=1.505 w=0.36 l=0.15
X23 Q.t5 a_2051_413.t7 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_193_47.t0 a_27_47.t6 VPWR.t13 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1231_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1056 pd=0.97 as=0.1264 ps=1.035 w=0.64 l=0.15
X26 a_915_47# SCE.t2 a_1226_119.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.22515 pd=1.505 as=0.0441 ps=0.63 w=0.42 l=0.15
X27 VPWR.t8 a_2051_413.t8 Q.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_299_47.t3 a_791_264.t3 a_729_369.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0992 pd=0.95 as=0.1152 ps=1 w=0.64 l=0.15
X29 a_381_47.t1 D.t1 a_299_47.t4 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 VPWR.t12 a_791_264.t4 a_2135_413.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X31 Q.t0 a_2051_413.t9 VPWR.t7 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X32 VPWR.t0 a_423_343.t3 a_381_369.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X33 a_915_47# SCE.t3 a_299_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1984 pd=1.9 as=0.0992 ps=0.95 w=0.64 l=0.15
X34 a_1960_413.t0 a_1610_159.t4 VPWR.t14 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_1226_119.t1 SCD.t0 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X36 a_1446_413.t1 a_193_47.t4 a_915_47# VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.13415 ps=1.085 w=0.42 l=0.15
X37 a_915_47# a_885_21.t2 a_299_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X38 VPWR.t6 a_2051_413.t10 a_791_264.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1728 ps=1.82 w=0.64 l=0.15
X39 VGND.t5 a_2051_413.t11 Q.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 VGND.t9 CLK.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X41 VGND.t2 DE.t3 a_381_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X42 a_1610_159.t1 a_1446_413.t5 VGND.t11 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
R0 D.n0 D.t1 220.367
R1 D.n0 D.t0 216.796
R2 D D.n0 71.33
R3 a_299_47.n1 a_299_47.t5 467.892
R4 a_299_47.n3 a_299_47.n2 380.248
R5 a_299_47.n1 a_299_47.t4 232.434
R6 a_299_47.n2 a_299_47.n0 188.082
R7 a_299_47.t0 a_299_47.n3 53.8677
R8 a_299_47.n3 a_299_47.t3 41.5552
R9 a_299_47.n0 a_299_47.t2 38.5719
R10 a_299_47.n0 a_299_47.t1 38.5719
R11 a_299_47.n2 a_299_47.n1 20.4743
R12 a_381_369.t0 a_381_369.t1 64.6411
R13 VPB.t10 VPB.t18 1043.39
R14 VPB.t15 VPB.t9 624.456
R15 VPB.t0 VPB.t10 622.851
R16 VPB.t8 VPB.t19 556.386
R17 VPB.t2 VPB.t7 556.386
R18 VPB.t12 VPB.t20 556.386
R19 VPB.t19 VPB.t5 517.913
R20 VPB.t13 VPB.t8 390.654
R21 VPB.t5 VPB.t15 337.384
R22 VPB.t11 VPB.t13 304.829
R23 VPB.t1 VPB.t14 301.87
R24 VPB.t9 VPB.t17 287.072
R25 VPB.t14 VPB.t0 272.274
R26 VPB.t7 VPB.t1 260.437
R27 VPB.t18 VPB.t11 256.56
R28 VPB.t4 VPB.t3 248.599
R29 VPB.t16 VPB.t4 248.599
R30 VPB.t17 VPB.t16 248.599
R31 VPB.t6 VPB.t12 248.599
R32 VPB.t20 VPB.t2 213.084
R33 VPB VPB.t6 142.056
R34 a_27_47.n3 a_27_47.t2 443.44
R35 a_27_47.t0 a_27_47.n6 390.443
R36 a_27_47.n4 a_27_47.t5 344.428
R37 a_27_47.n4 a_27_47.t3 296.969
R38 a_27_47.n1 a_27_47.t1 288.373
R39 a_27_47.n0 a_27_47.t6 263.406
R40 a_27_47.n3 a_27_47.n2 254.389
R41 a_27_47.n0 a_27_47.t4 228.06
R42 a_27_47.n5 a_27_47.n3 194.501
R43 a_27_47.n1 a_27_47.n0 152
R44 a_27_47.n6 a_27_47.n1 35.3396
R45 a_27_47.n6 a_27_47.n5 15.3376
R46 a_27_47.n5 a_27_47.n4 12.879
R47 a_2051_413.t0 a_2051_413.n5 754.347
R48 a_2051_413.n5 a_2051_413.t1 328.771
R49 a_2051_413.n4 a_2051_413.t10 269.921
R50 a_2051_413.n5 a_2051_413.n4 252.183
R51 a_2051_413.n0 a_2051_413.t2 212.081
R52 a_2051_413.n1 a_2051_413.t4 212.081
R53 a_2051_413.n2 a_2051_413.t8 212.081
R54 a_2051_413.n3 a_2051_413.t9 212.081
R55 a_2051_413.n4 a_2051_413.t3 176.733
R56 a_2051_413.n0 a_2051_413.t11 139.78
R57 a_2051_413.n1 a_2051_413.t7 139.78
R58 a_2051_413.n2 a_2051_413.t5 139.78
R59 a_2051_413.n3 a_2051_413.t6 139.78
R60 a_2051_413.n4 a_2051_413.n3 70.8399
R61 a_2051_413.n1 a_2051_413.n0 61.346
R62 a_2051_413.n2 a_2051_413.n1 61.346
R63 a_2051_413.n3 a_2051_413.n2 61.346
R64 VNB.t19 VNB.t11 4029.77
R65 VNB.t14 VNB.t13 3203.88
R66 VNB.t5 VNB.t15 3066.59
R67 VNB.t16 VNB.t19 2890.61
R68 VNB.t13 VNB.t16 2677.02
R69 VNB.t3 VNB.t12 2677.02
R70 VNB.t18 VNB.t20 2677.02
R71 VNB.t0 VNB.t17 2318.4
R72 VNB.t4 VNB.t1 1452.43
R73 VNB.t11 VNB.t9 1381.23
R74 VNB.t17 VNB.t14 1253.07
R75 VNB.t12 VNB.t4 1253.07
R76 VNB.t8 VNB.t7 1196.12
R77 VNB.t10 VNB.t8 1196.12
R78 VNB.t9 VNB.t10 1196.12
R79 VNB.t1 VNB.t5 1196.12
R80 VNB.t6 VNB.t18 1196.12
R81 VNB.t15 VNB.t2 1103.28
R82 VNB.t20 VNB.t3 1025.24
R83 VNB.t2 VNB.t0 945.673
R84 VNB VNB.t6 683.495
R85 a_1446_413.n3 a_1446_413.n2 680.737
R86 a_1446_413.n2 a_1446_413.n1 276.272
R87 a_1446_413.n0 a_1446_413.t5 230.484
R88 a_1446_413.n0 a_1446_413.t4 196.013
R89 a_1446_413.n2 a_1446_413.n0 171.939
R90 a_1446_413.n3 a_1446_413.t3 72.7029
R91 a_1446_413.t1 a_1446_413.n3 70.3576
R92 a_1446_413.n1 a_1446_413.t0 51.6672
R93 a_1446_413.n1 a_1446_413.t2 45.0005
R94 a_1537_413.t0 a_1537_413.t1 171.202
R95 DE.n0 DE.t2 319.728
R96 DE.n2 DE.n1 238.69
R97 DE.n0 DE.t0 178.34
R98 DE DE.n2 158.893
R99 DE.n1 DE.n0 147.814
R100 DE.n2 DE.t3 130.387
R101 DE.n1 DE.t1 130.141
R102 a_423_343.t0 a_423_343.n1 376.974
R103 a_423_343.n1 a_423_343.t3 375.568
R104 a_423_343.n0 a_423_343.t2 334.038
R105 a_423_343.n0 a_423_343.t1 244.181
R106 a_423_343.n1 a_423_343.n0 11.1343
R107 VPWR.n29 VPWR.t12 671.345
R108 VPWR.n36 VPWR.t14 667.963
R109 VPWR.n48 VPWR.t9 659.122
R110 VPWR.n63 VPWR.n1 604.394
R111 VPWR.n57 VPWR.t0 374.937
R112 VPWR.n55 VPWR.n5 323.079
R113 VPWR.n12 VPWR.n11 317.757
R114 VPWR.n19 VPWR.t5 259.553
R115 VPWR.n23 VPWR.n22 241.126
R116 VPWR.n20 VPWR.n18 233.137
R117 VPWR.n11 VPWR.t11 106.1
R118 VPWR.n22 VPWR.t6 61.9796
R119 VPWR.n5 VPWR.t2 44.6333
R120 VPWR.n5 VPWR.t1 44.6333
R121 VPWR.n11 VPWR.t10 43.3405
R122 VPWR.n1 VPWR.t13 41.5552
R123 VPWR.n1 VPWR.t3 41.5552
R124 VPWR.n61 VPWR.n2 34.6358
R125 VPWR.n62 VPWR.n61 34.6358
R126 VPWR.n50 VPWR.n49 34.6358
R127 VPWR.n50 VPWR.n6 34.6358
R128 VPWR.n54 VPWR.n6 34.6358
R129 VPWR.n42 VPWR.n41 34.6358
R130 VPWR.n43 VPWR.n42 34.6358
R131 VPWR.n43 VPWR.n9 34.6358
R132 VPWR.n47 VPWR.n9 34.6358
R133 VPWR.n31 VPWR.n30 34.6358
R134 VPWR.n31 VPWR.n14 34.6358
R135 VPWR.n35 VPWR.n14 34.6358
R136 VPWR.n28 VPWR.n16 34.6358
R137 VPWR.n24 VPWR.n21 34.6358
R138 VPWR.n55 VPWR.n54 33.8829
R139 VPWR.n57 VPWR.n56 32.0005
R140 VPWR.n22 VPWR.t7 30.1768
R141 VPWR.n37 VPWR.n36 30.1181
R142 VPWR.n49 VPWR.n48 28.2358
R143 VPWR.n41 VPWR.n12 28.2358
R144 VPWR.n18 VPWR.t4 26.5955
R145 VPWR.n18 VPWR.t8 26.5955
R146 VPWR.n20 VPWR.n19 23.9067
R147 VPWR.n37 VPWR.n12 23.3417
R148 VPWR.n63 VPWR.n62 22.9652
R149 VPWR.n56 VPWR.n55 20.7064
R150 VPWR.n36 VPWR.n35 17.3181
R151 VPWR.n21 VPWR.n20 17.3181
R152 VPWR.n48 VPWR.n47 15.0593
R153 VPWR.n29 VPWR.n28 14.3064
R154 VPWR.n57 VPWR.n2 12.424
R155 VPWR.n23 VPWR.n16 12.0476
R156 VPWR.n21 VPWR.n17 9.3005
R157 VPWR.n25 VPWR.n24 9.3005
R158 VPWR.n26 VPWR.n16 9.3005
R159 VPWR.n28 VPWR.n27 9.3005
R160 VPWR.n30 VPWR.n15 9.3005
R161 VPWR.n32 VPWR.n31 9.3005
R162 VPWR.n33 VPWR.n14 9.3005
R163 VPWR.n35 VPWR.n34 9.3005
R164 VPWR.n36 VPWR.n13 9.3005
R165 VPWR.n38 VPWR.n37 9.3005
R166 VPWR.n39 VPWR.n12 9.3005
R167 VPWR.n41 VPWR.n40 9.3005
R168 VPWR.n42 VPWR.n10 9.3005
R169 VPWR.n44 VPWR.n43 9.3005
R170 VPWR.n45 VPWR.n9 9.3005
R171 VPWR.n47 VPWR.n46 9.3005
R172 VPWR.n48 VPWR.n8 9.3005
R173 VPWR.n49 VPWR.n7 9.3005
R174 VPWR.n51 VPWR.n50 9.3005
R175 VPWR.n52 VPWR.n6 9.3005
R176 VPWR.n54 VPWR.n53 9.3005
R177 VPWR.n55 VPWR.n4 9.3005
R178 VPWR.n56 VPWR.n3 9.3005
R179 VPWR.n58 VPWR.n57 9.3005
R180 VPWR.n59 VPWR.n2 9.3005
R181 VPWR.n61 VPWR.n60 9.3005
R182 VPWR.n62 VPWR.n0 9.3005
R183 VPWR.n64 VPWR.n63 7.12063
R184 VPWR.n24 VPWR.n23 4.89462
R185 VPWR.n19 VPWR.n17 1.13003
R186 VPWR.n30 VPWR.n29 0.753441
R187 VPWR.n64 VPWR.n0 0.148519
R188 VPWR.n25 VPWR.n17 0.120292
R189 VPWR.n26 VPWR.n25 0.120292
R190 VPWR.n27 VPWR.n26 0.120292
R191 VPWR.n27 VPWR.n15 0.120292
R192 VPWR.n32 VPWR.n15 0.120292
R193 VPWR.n33 VPWR.n32 0.120292
R194 VPWR.n34 VPWR.n33 0.120292
R195 VPWR.n34 VPWR.n13 0.120292
R196 VPWR.n38 VPWR.n13 0.120292
R197 VPWR.n39 VPWR.n38 0.120292
R198 VPWR.n40 VPWR.n39 0.120292
R199 VPWR.n40 VPWR.n10 0.120292
R200 VPWR.n44 VPWR.n10 0.120292
R201 VPWR.n45 VPWR.n44 0.120292
R202 VPWR.n46 VPWR.n45 0.120292
R203 VPWR.n46 VPWR.n8 0.120292
R204 VPWR.n8 VPWR.n7 0.120292
R205 VPWR.n51 VPWR.n7 0.120292
R206 VPWR.n52 VPWR.n51 0.120292
R207 VPWR.n53 VPWR.n52 0.120292
R208 VPWR.n53 VPWR.n4 0.120292
R209 VPWR.n4 VPWR.n3 0.120292
R210 VPWR.n58 VPWR.n3 0.120292
R211 VPWR.n59 VPWR.n58 0.120292
R212 VPWR.n60 VPWR.n59 0.120292
R213 VPWR.n60 VPWR.n0 0.120292
R214 VPWR VPWR.n64 0.114842
R215 CLK.n0 CLK.t0 292.95
R216 CLK.n0 CLK.t1 209.403
R217 CLK CLK.n0 154.069
R218 SCE.t1 SCE.t2 604.107
R219 SCE.n1 SCE.t3 352.397
R220 SCE.n0 SCE.t0 189.588
R221 SCE SCE.n1 153.631
R222 SCE.n0 SCE.t1 142.03
R223 SCE.n1 SCE.n0 74.0857
R224 a_885_21.n0 a_885_21.t2 571.547
R225 a_885_21.n2 a_885_21.n1 427.555
R226 a_885_21.t0 a_885_21.n2 372.423
R227 a_885_21.n0 a_885_21.t1 223.571
R228 a_885_21.n2 a_885_21.n0 74.941
R229 VGND.n36 VGND.t11 273.476
R230 VGND.n30 VGND.t12 244.518
R231 VGND.n57 VGND.t2 238.311
R232 VGND.n44 VGND.n43 222.888
R233 VGND.n55 VGND.n4 202.262
R234 VGND.n64 VGND.n63 199.739
R235 VGND.n17 VGND.t5 157.841
R236 VGND.n16 VGND.n15 121.828
R237 VGND.n22 VGND.n21 118.657
R238 VGND.n21 VGND.t4 57.8171
R239 VGND.n4 VGND.t0 41.4291
R240 VGND.n4 VGND.t1 41.4291
R241 VGND.n43 VGND.t3 38.5719
R242 VGND.n43 VGND.t10 38.5719
R243 VGND.n63 VGND.t13 38.5719
R244 VGND.n63 VGND.t9 38.5719
R245 VGND.n20 VGND.n14 34.6358
R246 VGND.n24 VGND.n23 34.6358
R247 VGND.n28 VGND.n12 34.6358
R248 VGND.n29 VGND.n28 34.6358
R249 VGND.n31 VGND.n29 34.6358
R250 VGND.n35 VGND.n10 34.6358
R251 VGND.n37 VGND.n8 34.6358
R252 VGND.n41 VGND.n8 34.6358
R253 VGND.n42 VGND.n41 34.6358
R254 VGND.n45 VGND.n42 34.6358
R255 VGND.n49 VGND.n6 34.6358
R256 VGND.n50 VGND.n49 34.6358
R257 VGND.n51 VGND.n50 34.6358
R258 VGND.n51 VGND.n3 34.6358
R259 VGND.n61 VGND.n1 34.6358
R260 VGND.n62 VGND.n61 34.6358
R261 VGND.n57 VGND.n56 32.0005
R262 VGND.n55 VGND.n3 29.7417
R263 VGND.n15 VGND.t6 24.9236
R264 VGND.n15 VGND.t8 24.9236
R265 VGND.n36 VGND.n35 24.8476
R266 VGND.n21 VGND.t7 24.7511
R267 VGND.n17 VGND.n16 23.9067
R268 VGND.n64 VGND.n62 22.9652
R269 VGND.n16 VGND.n14 17.3181
R270 VGND.n45 VGND.n44 15.0593
R271 VGND.n37 VGND.n36 14.6829
R272 VGND.n56 VGND.n55 14.6829
R273 VGND.n57 VGND.n1 12.424
R274 VGND.n23 VGND.n22 12.0476
R275 VGND.n31 VGND.n30 11.2946
R276 VGND.n24 VGND.n12 10.9181
R277 VGND.n62 VGND.n0 9.3005
R278 VGND.n61 VGND.n60 9.3005
R279 VGND.n59 VGND.n1 9.3005
R280 VGND.n58 VGND.n57 9.3005
R281 VGND.n56 VGND.n2 9.3005
R282 VGND.n55 VGND.n54 9.3005
R283 VGND.n53 VGND.n3 9.3005
R284 VGND.n52 VGND.n51 9.3005
R285 VGND.n50 VGND.n5 9.3005
R286 VGND.n49 VGND.n48 9.3005
R287 VGND.n47 VGND.n6 9.3005
R288 VGND.n18 VGND.n14 9.3005
R289 VGND.n20 VGND.n19 9.3005
R290 VGND.n23 VGND.n13 9.3005
R291 VGND.n25 VGND.n24 9.3005
R292 VGND.n26 VGND.n12 9.3005
R293 VGND.n28 VGND.n27 9.3005
R294 VGND.n29 VGND.n11 9.3005
R295 VGND.n32 VGND.n31 9.3005
R296 VGND.n33 VGND.n10 9.3005
R297 VGND.n35 VGND.n34 9.3005
R298 VGND.n36 VGND.n9 9.3005
R299 VGND.n38 VGND.n37 9.3005
R300 VGND.n39 VGND.n8 9.3005
R301 VGND.n41 VGND.n40 9.3005
R302 VGND.n42 VGND.n7 9.3005
R303 VGND.n46 VGND.n45 9.3005
R304 VGND.n65 VGND.n64 7.12063
R305 VGND.n22 VGND.n20 4.89462
R306 VGND.n30 VGND.n10 2.63579
R307 VGND.n18 VGND.n17 1.13003
R308 VGND.n44 VGND.n6 0.753441
R309 VGND.n65 VGND.n0 0.148519
R310 VGND.n19 VGND.n18 0.120292
R311 VGND.n19 VGND.n13 0.120292
R312 VGND.n25 VGND.n13 0.120292
R313 VGND.n26 VGND.n25 0.120292
R314 VGND.n27 VGND.n26 0.120292
R315 VGND.n27 VGND.n11 0.120292
R316 VGND.n32 VGND.n11 0.120292
R317 VGND.n33 VGND.n32 0.120292
R318 VGND.n34 VGND.n33 0.120292
R319 VGND.n34 VGND.n9 0.120292
R320 VGND.n38 VGND.n9 0.120292
R321 VGND.n39 VGND.n38 0.120292
R322 VGND.n40 VGND.n39 0.120292
R323 VGND.n40 VGND.n7 0.120292
R324 VGND.n46 VGND.n7 0.120292
R325 VGND.n47 VGND.n46 0.120292
R326 VGND.n48 VGND.n47 0.120292
R327 VGND.n48 VGND.n5 0.120292
R328 VGND.n52 VGND.n5 0.120292
R329 VGND.n53 VGND.n52 0.120292
R330 VGND.n54 VGND.n53 0.120292
R331 VGND.n54 VGND.n2 0.120292
R332 VGND.n58 VGND.n2 0.120292
R333 VGND.n59 VGND.n58 0.120292
R334 VGND.n60 VGND.n59 0.120292
R335 VGND.n60 VGND.n0 0.120292
R336 VGND VGND.n65 0.114842
R337 a_1610_159.t0 a_1610_159.n4 408.848
R338 a_1610_159.n2 a_1610_159.t2 406.401
R339 a_1610_159.n0 a_1610_159.t4 318.12
R340 a_1610_159.n0 a_1610_159.t3 194.477
R341 a_1610_159.n3 a_1610_159.n2 176.534
R342 a_1610_159.n4 a_1610_159.n0 168.486
R343 a_1610_159.n3 a_1610_159.t1 140.249
R344 a_1610_159.n2 a_1610_159.n1 130.054
R345 a_1610_159.n4 a_1610_159.n3 9.32396
R346 Q.n4 Q.n3 219.632
R347 Q.n2 Q.n0 219.631
R348 Q.n2 Q.n1 112.945
R349 Q Q.n5 110.037
R350 Q.n4 Q.n2 29.0138
R351 Q.n3 Q.t1 26.5955
R352 Q.n3 Q.t0 26.5955
R353 Q.n0 Q.t3 26.5955
R354 Q.n0 Q.t2 26.5955
R355 Q.n5 Q.t7 24.9236
R356 Q.n5 Q.t6 24.9236
R357 Q.n1 Q.t4 24.9236
R358 Q.n1 Q.t5 24.9236
R359 Q Q.n4 2.90959
R360 a_791_264.n3 a_791_264.n2 382.745
R361 a_791_264.t0 a_791_264.n4 362.808
R362 a_791_264.n0 a_791_264.t2 310.623
R363 a_791_264.n1 a_791_264.t1 242.322
R364 a_791_264.n1 a_791_264.n0 220.962
R365 a_791_264.n0 a_791_264.t3 194.942
R366 a_791_264.n4 a_791_264.n3 174.017
R367 a_791_264.n3 a_791_264.t4 138.53
R368 a_791_264.n4 a_791_264.n1 48.371
R369 a_193_47.t0 a_193_47.n4 395.625
R370 a_193_47.n2 a_193_47.t2 389.545
R371 a_193_47.n1 a_193_47.t3 308.651
R372 a_193_47.n4 a_193_47.t1 300.372
R373 a_193_47.n1 a_193_47.n0 298.373
R374 a_193_47.n2 a_193_47.t4 273.572
R375 a_193_47.n3 a_193_47.n2 173.755
R376 a_193_47.n4 a_193_47.n3 14.6322
R377 a_193_47.n3 a_193_47.n1 12.2528
R378 a_1974_47.n0 a_1974_47.t0 45.1697
R379 a_729_47.t0 a_729_47.t1 102.858
R380 a_729_369.t0 a_729_369.t1 110.812
R381 a_2135_413.t0 a_2135_413.t1 197
R382 SCD.n1 SCD.t0 206.19
R383 SCD.n1 SCD.n0 183.696
R384 SCD SCD.n1 163.675
R385 a_1226_119.t0 a_1226_119.t1 60.0005
R386 a_381_47.t0 a_381_47.t1 60.0005
C0 VPB DE 0.114449f
C1 a_915_47# VPB 0.021894f
C2 VPWR DE 0.04692f
C3 a_915_47# VPWR 0.097411f
C4 a_915_47# a_1561_47# 4.9e-19
C5 D VGND 0.014495f
C6 VGND Q 0.342075f
C7 Q SCE 3.49e-20
C8 VGND SCD 0.032521f
C9 SCE SCD 0.095395f
C10 VPB D 0.068631f
C11 CLK VGND 0.019296f
C12 D VPWR 0.01674f
C13 VPB Q 0.010305f
C14 D DE 0.099354f
C15 VPB SCD 0.045339f
C16 VPWR Q 0.429786f
C17 VPWR SCD 0.013425f
C18 VGND SCE 0.047542f
C19 a_915_47# Q 5.86e-20
C20 a_915_47# SCD 0.018533f
C21 a_2177_47# VGND 0.004743f
C22 VPB CLK 0.069635f
C23 CLK VPWR 0.019263f
C24 VPB VGND 0.015334f
C25 VPB SCE 0.1417f
C26 VPWR VGND 0.113339f
C27 VPWR SCE 0.028732f
C28 VGND DE 0.057232f
C29 a_915_47# VGND 0.38346f
C30 a_1231_369# VPWR 0.0081f
C31 a_915_47# SCE 0.086615f
C32 a_915_47# a_1231_369# 0.003336f
C33 VGND a_1561_47# 0.004442f
C34 a_915_47# a_2177_47# 5.05e-20
C35 VPB VPWR 0.334953f
C36 Q VNB 0.011356f
C37 VGND VNB 1.6599f
C38 VPWR VNB 1.33466f
C39 SCD VNB 0.08884f
C40 SCE VNB 0.334233f
C41 DE VNB 0.282831f
C42 D VNB 0.122269f
C43 CLK VNB 0.195128f
C44 VPB VNB 2.87215f
C45 a_915_47# VNB 0.03797f
.ends

* NGSPICE file created from sky130_fd_sc_hd__tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tap_1 VGND VPWR VNB VPB
C0 VPWR VPB 0.054142f
C1 VPWR VGND 0.009821f
C2 VPB VGND 0.005223f
C3 VGND VNB 0.139414f
C4 VPWR VNB 0.091891f
C5 VPB VNB 0.244246f
.ends

* NGSPICE file created from sky130_fd_sc_hd__tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tap_2 VGND VPWR VPB VNB
C0 VPB VGND 0.008596f
C1 VPWR VGND 0.017949f
C2 VPB VPWR 0.121904f
C3 VGND VNB 0.242529f
C4 VPWR VNB 0.13283f
C5 VPB VNB 0.352722f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X.t1 a_35_297.t3 a_285_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X.t0 B.t0 a_285_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297.t1 B.t2 a_35_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR.t1 B.t3 a_285_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t3 A.t0 a_35_297.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND.t2 a_35_297.t4 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297.t0 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t0 A.t2 a_117_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47.t1 A.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_35_297.t1 a_35_297.n2 442.868
R1 a_35_297.n2 a_35_297.n1 343.923
R2 a_35_297.n1 a_35_297.t3 215.482
R3 a_35_297.n2 a_35_297.n0 196.672
R4 a_35_297.n1 a_35_297.t4 139.78
R5 a_35_297.n0 a_35_297.t2 24.9236
R6 a_35_297.n0 a_35_297.t0 24.9236
R7 a_285_297.n0 a_285_297.t2 661.615
R8 a_285_297.n0 a_285_297.t1 26.5955
R9 a_285_297.t0 a_285_297.n0 26.5955
R10 X.n1 X.t1 235.792
R11 X.n1 X.n0 173.87
R12 X.n0 X.t0 66.0319
R13 X.n0 X.t2 59.081
R14 X X.n1 0.2005
R15 VPB.t3 VPB.t4 556.386
R16 VPB.t2 VPB.t3 248.599
R17 VPB.t0 VPB.t2 248.599
R18 VPB.t1 VPB.t0 248.599
R19 VPB VPB.t1 216.044
R20 B.n2 B.n0 249.882
R21 B.n1 B.t2 241.536
R22 B.n0 B.t3 241.536
R23 B.n1 B.t1 169.237
R24 B.n0 B.t0 169.237
R25 B B.n1 166.891
R26 B B.n2 4.89462
R27 B.n2 B 4.44132
R28 a_285_47.t0 a_285_47.t1 49.8467
R29 VNB.t1 VNB.t3 2620.06
R30 VNB.t2 VNB.t1 1196.12
R31 VNB.t4 VNB.t2 1196.12
R32 VNB.t0 VNB.t4 1196.12
R33 VNB VNB.t0 1039.48
R34 VGND.n5 VGND.t0 278.589
R35 VGND.n3 VGND.n2 200.127
R36 VGND.n1 VGND.t2 152.428
R37 VGND.n2 VGND.t1 24.9236
R38 VGND.n2 VGND.t3 24.9236
R39 VGND.n4 VGND.n3 21.4593
R40 VGND.n5 VGND.n4 16.9417
R41 VGND.n6 VGND.n5 9.3005
R42 VGND.n4 VGND.n0 9.3005
R43 VGND.n3 VGND.n1 7.08982
R44 VGND.n1 VGND.n0 0.170346
R45 VGND.n6 VGND.n0 0.120292
R46 VGND VGND.n6 0.0226354
R47 a_117_297.t0 a_117_297.t1 53.1905
R48 VPWR.n1 VPWR.t1 852.101
R49 VPWR.n1 VPWR.n0 331.286
R50 VPWR.n0 VPWR.t2 26.5955
R51 VPWR.n0 VPWR.t0 26.5955
R52 VPWR VPWR.n1 0.648038
R53 A.n0 A.t1 212.081
R54 A.n1 A.t2 212.081
R55 A A.n2 153.28
R56 A.n0 A.t3 139.78
R57 A.n1 A.t0 139.78
R58 A.n2 A.n0 37.246
R59 A.n2 A.n1 24.1005
C0 B VPWR 0.070314f
C1 VPB X 0.015415f
C2 VPB B 0.069694f
C3 VPB VPWR 0.068915f
C4 A VGND 0.032545f
C5 X VGND 0.172898f
C6 B VGND 0.030447f
C7 A X 0.001658f
C8 B A 0.221335f
C9 VPWR VGND 0.064265f
C10 A VPWR 0.034845f
C11 B X 0.014878f
C12 VPB VGND 0.006962f
C13 VPB A 0.051013f
C14 VPWR X 0.053654f
C15 VGND VNB 0.434883f
C16 X VNB 0.064909f
C17 VPWR VNB 0.332777f
C18 A VNB 0.166719f
C19 B VNB 0.213371f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor3_4 VNB VPB VGND VPWR X C B A
X0 a_1382_49.t5 a_1011_297.t2 a_631_49# VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.246 pd=1.525 as=0.2431 ps=1.445 w=0.64 l=0.15
X1 a_1382_49.t3 a_1117_297.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1824 pd=1.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_1117_297.t3 a_1011_297.t3 a_631_49# VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.11 pd=0.99 as=0.140825 ps=1.1 w=0.6 l=0.15
X3 a_1011_297.t0 B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.16515 pd=1.82 as=0.1885 ps=1.88 w=0.65 l=0.15
X4 a_1382_49.t2 a_1117_297.t5 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X5 a_101_21.t2 C.t0 a_631_49# VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0928 pd=0.93 as=0.1728 ps=1.82 w=0.64 l=0.15
X6 VPWR.t2 A.t0 a_1117_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1715 ps=1.355 w=1 l=0.15
X7 VPWR.t4 a_101_21.t4 X.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1011_297.t1 B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.25655 ps=2.52 w=1 l=0.15
X9 X.t2 a_101_21.t5 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X10 VPWR.t6 a_101_21.t6 X.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X11 a_492_93.t0 C.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1792 pd=1.84 as=0.169 ps=1.365 w=0.64 l=0.15
X12 X.t7 a_101_21.t7 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X.t6 a_101_21.t8 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_607_325.t0 B.t2 a_1382_49.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1458 pd=1.205 as=0.246 ps=1.525 w=0.64 l=0.15
X15 X.t0 a_101_21.t9 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 a_631_49# B.t3 a_1382_49.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.140825 pd=1.1 as=0.19265 ps=1.285 w=0.64 l=0.15
X17 a_101_21.t3 C.t2 a_607_325.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.15295 pd=1.315 as=0.273 ps=2.33 w=0.84 l=0.15
X18 VGND.t6 a_101_21.t10 X.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1165 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_631_49# a_492_93.t2 a_101_21.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.32235 pd=2.45 as=0.15295 ps=1.315 w=0.84 l=0.15
X20 VGND.t7 a_101_21.t11 X.t4 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_607_325.t1 a_492_93.t3 a_101_21.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.224 pd=1.98 as=0.0928 ps=0.93 w=0.64 l=0.15
X22 VGND.t2 A.t1 a_1117_297.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.11 ps=0.99 w=0.64 l=0.15
X23 a_1117_297.t2 a_1011_297.t4 a_607_325.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1715 pd=1.355 as=0.1458 ps=1.205 w=0.84 l=0.15
X24 a_1382_49.t4 a_1011_297.t5 a_607_325.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.19265 pd=1.285 as=0.18205 ps=1.245 w=0.42 l=0.15
X25 a_492_93.t1 C.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1785 pd=1.69 as=0.1165 ps=1.035 w=0.42 l=0.15
R0 a_1011_297.t1 a_1011_297.n3 891.352
R1 a_1011_297.n0 a_1011_297.t4 283.257
R2 a_1011_297.n2 a_1011_297.n1 224.038
R3 a_1011_297.n3 a_1011_297.t0 218.472
R4 a_1011_297.n2 a_1011_297.n0 175.175
R5 a_1011_297.n1 a_1011_297.t5 173.52
R6 a_1011_297.n0 a_1011_297.t3 161.202
R7 a_1011_297.n1 a_1011_297.t2 154.24
R8 a_1011_297.n3 a_1011_297.n2 10.4313
R9 a_1382_49.n2 a_1382_49.n1 590.155
R10 a_1382_49.t2 a_1382_49.n3 323.08
R11 a_1382_49.n3 a_1382_49.t3 318.813
R12 a_1382_49.n2 a_1382_49.n0 284.765
R13 a_1382_49.n1 a_1382_49.t5 209.827
R14 a_1382_49.n3 a_1382_49.n2 130.951
R15 a_1382_49.n0 a_1382_49.t4 94.7773
R16 a_1382_49.n1 a_1382_49.t0 41.5557
R17 a_1382_49.n0 a_1382_49.t1 38.438
R18 VPB.t1 VPB.t7 1097.97
R19 VPB.t8 VPB.t1 627.414
R20 VPB.t3 VPB.t4 621.495
R21 VPB.t7 VPB.t2 517.913
R22 VPB.t2 VPB.t6 304.829
R23 VPB.t9 VPB.t3 304.829
R24 VPB.t6 VPB.t0 298.911
R25 VPB.t4 VPB.t8 287.072
R26 VPB.t11 VPB.t10 266.356
R27 VPB VPB.t12 257.478
R28 VPB.t0 VPB.t5 248.599
R29 VPB.t10 VPB.t9 248.599
R30 VPB.t12 VPB.t11 248.599
R31 a_1117_297.n4 a_1117_297.n3 641.726
R32 a_1117_297.n2 a_1117_297.t5 241.536
R33 a_1117_297.n3 a_1117_297.n1 241.438
R34 a_1117_297.n2 a_1117_297.t4 170.843
R35 a_1117_297.n3 a_1117_297.n2 152
R36 a_1117_297.n0 a_1117_297.t2 50.4231
R37 a_1117_297.n1 a_1117_297.t3 43.0005
R38 a_1117_297.n5 a_1117_297.n4 38.6969
R39 a_1117_297.n0 a_1117_297.t0 28.8712
R40 a_1117_297.n1 a_1117_297.t1 23.0795
R41 a_1117_297.n4 a_1117_297.n0 17.5898
R42 VGND.n26 VGND.t5 245.689
R43 VGND.n20 VGND.n19 244.077
R44 VGND.n2 VGND.n1 220.766
R45 VGND.n9 VGND.n8 217.561
R46 VGND.n7 VGND.t1 154.78
R47 VGND.n19 VGND.t3 65.7148
R48 VGND.n12 VGND.n6 34.6358
R49 VGND.n13 VGND.n12 34.6358
R50 VGND.n14 VGND.n13 34.6358
R51 VGND.n14 VGND.n4 34.6358
R52 VGND.n18 VGND.n4 34.6358
R53 VGND.n25 VGND.n24 34.6358
R54 VGND.n9 VGND.n7 33.9541
R55 VGND.n21 VGND.n2 30.1181
R56 VGND.n20 VGND.n18 28.9887
R57 VGND.n1 VGND.t4 26.7697
R58 VGND.n8 VGND.t0 25.313
R59 VGND.n8 VGND.t2 25.313
R60 VGND.n1 VGND.t7 24.9236
R61 VGND.n26 VGND.n25 24.0946
R62 VGND.n21 VGND.n20 21.4593
R63 VGND.n19 VGND.t6 20.0915
R64 VGND.n27 VGND.n26 19.8417
R65 VGND.n10 VGND.n6 9.3005
R66 VGND.n12 VGND.n11 9.3005
R67 VGND.n13 VGND.n5 9.3005
R68 VGND.n15 VGND.n14 9.3005
R69 VGND.n16 VGND.n4 9.3005
R70 VGND.n18 VGND.n17 9.3005
R71 VGND.n20 VGND.n3 9.3005
R72 VGND.n22 VGND.n21 9.3005
R73 VGND.n24 VGND.n23 9.3005
R74 VGND.n25 VGND.n0 9.3005
R75 VGND.n7 VGND.n6 8.28285
R76 VGND.n24 VGND.n2 4.51815
R77 VGND.n10 VGND.n9 0.147198
R78 VGND.n11 VGND.n10 0.120292
R79 VGND.n11 VGND.n5 0.120292
R80 VGND.n15 VGND.n5 0.120292
R81 VGND.n16 VGND.n15 0.120292
R82 VGND.n17 VGND.n16 0.120292
R83 VGND.n17 VGND.n3 0.120292
R84 VGND.n22 VGND.n3 0.120292
R85 VGND.n23 VGND.n22 0.120292
R86 VGND.n23 VGND.n0 0.120292
R87 VGND.n27 VGND.n0 0.120292
R88 VGND VGND.n27 0.0226354
R89 VNB.t1 VNB.t6 4798.71
R90 VNB.t5 VNB.t1 3445.95
R91 VNB.t4 VNB.t8 3175.4
R92 VNB.t6 VNB.t2 2264.08
R93 VNB.t2 VNB.t7 1708.74
R94 VNB.t11 VNB.t4 1523.62
R95 VNB.t7 VNB.t3 1423.95
R96 VNB.t8 VNB.t5 1253.07
R97 VNB VNB.t10 1238.83
R98 VNB.t12 VNB.t9 1224.6
R99 VNB.t3 VNB.t0 1196.12
R100 VNB.t9 VNB.t11 1196.12
R101 VNB.t10 VNB.t12 1196.12
R102 B.t2 B.n3 864.388
R103 B.n2 B.n1 298.841
R104 B.n1 B.t1 295.627
R105 B.n4 B.t2 235.109
R106 B.n3 B.n2 215.293
R107 B B.n4 194.166
R108 B.n1 B.t0 168.701
R109 B.n4 B.t3 167.63
R110 B.n2 B.n0 167.094
R111 VPWR.n7 VPWR.t1 783.061
R112 VPWR.n18 VPWR.n4 719.928
R113 VPWR.n9 VPWR.n8 605.511
R114 VPWR.n24 VPWR.t7 257.474
R115 VPWR.n2 VPWR.n1 230.879
R116 VPWR.n4 VPWR.t3 67.7193
R117 VPWR.n23 VPWR.n22 34.6358
R118 VPWR.n12 VPWR.n11 34.6358
R119 VPWR.n13 VPWR.n12 34.6358
R120 VPWR.n13 VPWR.n5 34.6358
R121 VPWR.n17 VPWR.n5 34.6358
R122 VPWR.n1 VPWR.t5 32.5055
R123 VPWR.n4 VPWR.t4 30.3773
R124 VPWR.n19 VPWR.n2 30.1181
R125 VPWR.n1 VPWR.t6 26.5955
R126 VPWR.n8 VPWR.t0 26.5955
R127 VPWR.n8 VPWR.t2 26.5955
R128 VPWR.n24 VPWR.n23 24.0946
R129 VPWR.n19 VPWR.n18 22.9652
R130 VPWR.n18 VPWR.n17 21.0829
R131 VPWR.n25 VPWR.n24 19.8417
R132 VPWR.n11 VPWR.n7 17.6946
R133 VPWR.n11 VPWR.n10 9.3005
R134 VPWR.n12 VPWR.n6 9.3005
R135 VPWR.n14 VPWR.n13 9.3005
R136 VPWR.n15 VPWR.n5 9.3005
R137 VPWR.n17 VPWR.n16 9.3005
R138 VPWR.n18 VPWR.n3 9.3005
R139 VPWR.n20 VPWR.n19 9.3005
R140 VPWR.n22 VPWR.n21 9.3005
R141 VPWR.n23 VPWR.n0 9.3005
R142 VPWR.n9 VPWR.n7 7.29413
R143 VPWR.n22 VPWR.n2 4.51815
R144 VPWR.n10 VPWR.n9 0.151957
R145 VPWR.n10 VPWR.n6 0.120292
R146 VPWR.n14 VPWR.n6 0.120292
R147 VPWR.n15 VPWR.n14 0.120292
R148 VPWR.n16 VPWR.n15 0.120292
R149 VPWR.n16 VPWR.n3 0.120292
R150 VPWR.n20 VPWR.n3 0.120292
R151 VPWR.n21 VPWR.n20 0.120292
R152 VPWR.n21 VPWR.n0 0.120292
R153 VPWR.n25 VPWR.n0 0.120292
R154 VPWR VPWR.n25 0.0226354
R155 C.n0 C.t2 269.921
R156 C C.n2 155.584
R157 C.n1 C.t1 154.24
R158 C.n0 C.t0 143.286
R159 C.n2 C.n1 132.916
R160 C.n1 C.t3 102.828
R161 C.n2 C.n0 24.8308
R162 a_101_21.n8 a_101_21.n7 774.88
R163 a_101_21.n7 a_101_21.n0 351.414
R164 a_101_21.n6 a_101_21.t4 212.081
R165 a_101_21.n4 a_101_21.t5 212.081
R166 a_101_21.n2 a_101_21.t6 212.081
R167 a_101_21.n1 a_101_21.t9 212.081
R168 a_101_21.n7 a_101_21.n6 165.876
R169 a_101_21.n2 a_101_21.t11 139.78
R170 a_101_21.n1 a_101_21.t8 139.78
R171 a_101_21.n3 a_101_21.t7 139.78
R172 a_101_21.n5 a_101_21.t10 139.78
R173 a_101_21.n3 a_101_21.n2 62.8066
R174 a_101_21.n2 a_101_21.n1 61.346
R175 a_101_21.n5 a_101_21.n4 58.4247
R176 a_101_21.n10 a_101_21.n9 55.1605
R177 a_101_21.n8 a_101_21.t3 32.6122
R178 a_101_21.n9 a_101_21.t1 30.3415
R179 a_101_21.n0 a_101_21.t0 27.188
R180 a_101_21.n0 a_101_21.t2 27.188
R181 a_101_21.n9 a_101_21.n8 21.1076
R182 a_101_21.n6 a_101_21.n5 2.92171
R183 a_101_21.n4 a_101_21.n3 2.92171
R184 A.n0 A.t0 239.505
R185 A.n0 A.t1 168.811
R186 A A.n0 163.52
R187 X.n3 X.n1 215.172
R188 X.n3 X.n2 208.825
R189 X.n4 X.n0 206.626
R190 X.n6 X.n5 198.507
R191 X.n4 X.n3 30.8369
R192 X.n5 X.t3 26.5955
R193 X.n5 X.t2 26.5955
R194 X.n1 X.t1 26.5955
R195 X.n1 X.t0 26.5955
R196 X.n0 X.t5 24.9236
R197 X.n0 X.t7 24.9236
R198 X.n2 X.t4 24.9236
R199 X.n2 X.t6 24.9236
R200 X.n6 X.n4 19.1577
R201 X X.n6 2.5605
R202 a_607_325.n2 a_607_325.n1 783.149
R203 a_607_325.n0 a_607_325.t4 728.472
R204 a_607_325.n1 a_607_325.t3 411.976
R205 a_607_325.n0 a_607_325.t1 355.445
R206 a_607_325.n1 a_607_325.n0 116.707
R207 a_607_325.n2 a_607_325.t0 67.7193
R208 a_607_325.t2 a_607_325.n2 34.3691
R209 a_492_93.t0 a_492_93.n1 726.078
R210 a_492_93.n1 a_492_93.t1 323.353
R211 a_492_93.n1 a_492_93.n0 256.433
R212 a_492_93.n0 a_492_93.t2 215.829
R213 a_492_93.n0 a_492_93.t3 167.63
C0 C a_631_49# 0.047636f
C1 VPWR A 0.014124f
C2 X B 2.49e-21
C3 a_631_49# VGND 0.176954f
C4 VPB a_631_49# 0.024916f
C5 VPWR X 0.369604f
C6 A VGND 0.01316f
C7 X C 0.002305f
C8 VPWR B 0.058719f
C9 VPB A 0.028102f
C10 X VGND 0.198412f
C11 VPB X 0.009243f
C12 C B 0.001529f
C13 B VGND 0.034452f
C14 VPB B 0.295971f
C15 VPWR C 0.020838f
C16 A a_631_49# 2.28e-19
C17 VPWR VGND 0.115211f
C18 VPB VPWR 0.202178f
C19 X a_631_49# 2.94e-19
C20 C VGND 0.018132f
C21 VPB C 0.142646f
C22 B a_631_49# 0.042426f
C23 VPB VGND 0.014343f
C24 VPWR a_631_49# 0.124351f
C25 B A 0.002172f
C26 VGND VNB 1.08407f
C27 A VNB 0.092322f
C28 B VNB 0.422926f
C29 C VNB 0.256456f
C30 X VNB 0.036337f
C31 VPWR VNB 0.90573f
C32 VPB VNB 1.9337f
C33 a_631_49# VNB 0.039097f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor3_2 VNB VPB VGND VPWR X C B A
X0 X.t1 a_87_21.t4 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_1198_49.t2 a_933_297.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1824 pd=1.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_87_21.t0 C.t0 a_423_325.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.15295 pd=1.315 as=0.273 ps=2.33 w=0.84 l=0.15
X3 a_447_49.t3 a_308_93.t2 a_87_21.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.32235 pd=2.45 as=0.15295 ps=1.315 w=0.84 l=0.15
X4 a_447_49.t2 B.t0 a_1198_49.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.140825 pd=1.1 as=0.19265 ps=1.285 w=0.64 l=0.15
X5 a_87_21.t1 C.t1 a_447_49.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0928 pd=0.93 as=0.1728 ps=1.82 w=0.64 l=0.15
X6 a_827_297.t1 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.16515 pd=1.82 as=0.1885 ps=1.88 w=0.65 l=0.15
X7 a_933_297.t0 a_827_297.t2 a_423_325.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1715 pd=1.355 as=0.1458 ps=1.205 w=0.84 l=0.15
X8 X.t3 a_87_21.t5 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.195 ps=1.9 w=0.65 l=0.15
X9 a_423_325.t3 a_308_93.t3 a_87_21.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.224 pd=1.98 as=0.0928 ps=0.93 w=0.64 l=0.15
X10 a_1198_49.t4 a_827_297.t3 a_423_325.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.19265 pd=1.285 as=0.18205 ps=1.245 w=0.42 l=0.15
X11 VGND.t5 A.t0 a_933_297.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.11 ps=0.99 w=0.64 l=0.15
X12 a_308_93.t1 C.t2 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1785 pd=1.69 as=0.1165 ps=1.035 w=0.42 l=0.15
X13 a_1198_49.t5 a_827_297.t4 a_447_49.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.246 pd=1.525 as=0.2431 ps=1.445 w=0.64 l=0.15
X14 a_1198_49.t1 a_933_297.t7 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X15 a_933_297.t1 a_827_297.t5 a_447_49.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.11 pd=0.99 as=0.140825 ps=1.1 w=0.6 l=0.15
X16 VPWR.t1 a_87_21.t6 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR.t3 A.t1 a_933_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1715 ps=1.355 w=1 l=0.15
X18 a_827_297.t0 B.t2 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.25655 ps=2.52 w=1 l=0.15
X19 a_423_325.t5 B.t3 a_933_297.t4 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.18205 pd=1.245 as=0.16275 ps=1.8 w=0.64 l=0.15
X20 VGND.t2 a_87_21.t7 X.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1165 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_308_93.t0 C.t3 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1792 pd=1.84 as=0.169 ps=1.365 w=0.64 l=0.15
X22 a_447_49.t5 B.t4 a_933_297.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.2431 pd=1.445 as=0.3528 ps=2.52 w=0.84 l=0.15
X23 a_423_325.t2 B.t5 a_1198_49.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1458 pd=1.205 as=0.246 ps=1.525 w=0.64 l=0.15
R0 a_87_21.n0 a_87_21.n5 774.88
R1 a_87_21.n5 a_87_21.n1 351.414
R2 a_87_21.n4 a_87_21.t6 212.081
R3 a_87_21.n2 a_87_21.t4 212.081
R4 a_87_21.n5 a_87_21.n4 165.876
R5 a_87_21.n2 a_87_21.t5 142.702
R6 a_87_21.n3 a_87_21.t7 139.78
R7 a_87_21.n3 a_87_21.n2 58.4247
R8 a_87_21.n6 a_87_21.n0 53.039
R9 a_87_21.n0 a_87_21.t3 51.4487
R10 a_87_21.n0 a_87_21.t0 32.6122
R11 a_87_21.n1 a_87_21.t2 27.188
R12 a_87_21.n1 a_87_21.t1 27.188
R13 a_87_21.n4 a_87_21.n3 2.92171
R14 VPWR.n5 VPWR.t5 783.061
R15 VPWR.n16 VPWR.n2 719.928
R16 VPWR.n7 VPWR.n6 605.511
R17 VPWR.n18 VPWR.t2 258.332
R18 VPWR.n2 VPWR.t4 67.7193
R19 VPWR.n10 VPWR.n9 34.6358
R20 VPWR.n11 VPWR.n10 34.6358
R21 VPWR.n11 VPWR.n3 34.6358
R22 VPWR.n15 VPWR.n3 34.6358
R23 VPWR.n2 VPWR.t1 30.3773
R24 VPWR.n6 VPWR.t0 26.5955
R25 VPWR.n6 VPWR.t3 26.5955
R26 VPWR.n18 VPWR.n17 23.7181
R27 VPWR.n17 VPWR.n16 22.9652
R28 VPWR.n16 VPWR.n15 21.0829
R29 VPWR.n9 VPWR.n5 17.6946
R30 VPWR.n9 VPWR.n8 9.3005
R31 VPWR.n10 VPWR.n4 9.3005
R32 VPWR.n12 VPWR.n11 9.3005
R33 VPWR.n13 VPWR.n3 9.3005
R34 VPWR.n15 VPWR.n14 9.3005
R35 VPWR.n16 VPWR.n1 9.3005
R36 VPWR.n17 VPWR.n0 9.3005
R37 VPWR.n19 VPWR.n18 9.3005
R38 VPWR.n7 VPWR.n5 7.29413
R39 VPWR.n8 VPWR.n7 0.151957
R40 VPWR.n8 VPWR.n4 0.120292
R41 VPWR.n12 VPWR.n4 0.120292
R42 VPWR.n13 VPWR.n12 0.120292
R43 VPWR.n14 VPWR.n13 0.120292
R44 VPWR.n14 VPWR.n1 0.120292
R45 VPWR.n1 VPWR.n0 0.120292
R46 VPWR.n19 VPWR.n0 0.120292
R47 VPWR VPWR.n19 0.0226354
R48 X.n2 X.n0 585
R49 X X.n0 304.337
R50 X.n2 X.n1 238.105
R51 X.n0 X.t0 26.5955
R52 X.n0 X.t1 26.5955
R53 X.n1 X.t2 24.9236
R54 X.n1 X.t3 24.9236
R55 X X.n2 7.54336
R56 VPB.t8 VPB.t10 651.091
R57 VPB.t11 VPB.t8 627.414
R58 VPB.t7 VPB.t0 621.495
R59 VPB.t9 VPB.t3 517.913
R60 VPB.t10 VPB.t9 446.885
R61 VPB.t3 VPB.t1 304.829
R62 VPB.t4 VPB.t7 304.829
R63 VPB.t1 VPB.t6 298.911
R64 VPB.t0 VPB.t11 287.072
R65 VPB.t6 VPB.t2 248.599
R66 VPB.t5 VPB.t4 248.599
R67 VPB VPB.t5 227.882
R68 a_933_297.n1 a_933_297.t3 760.636
R69 a_933_297.n6 a_933_297.n5 641.726
R70 a_933_297.n4 a_933_297.t7 241.536
R71 a_933_297.n1 a_933_297.t4 222.47
R72 a_933_297.n3 a_933_297.n2 185
R73 a_933_297.n4 a_933_297.t6 170.843
R74 a_933_297.n5 a_933_297.n4 152
R75 a_933_297.n5 a_933_297.n3 56.4377
R76 a_933_297.n0 a_933_297.t0 50.4231
R77 a_933_297.n2 a_933_297.t1 43.0005
R78 a_933_297.n7 a_933_297.n6 38.6969
R79 a_933_297.n0 a_933_297.t2 28.8712
R80 a_933_297.n3 a_933_297.n1 26.8515
R81 a_933_297.n2 a_933_297.t5 23.0795
R82 a_933_297.n6 a_933_297.n0 17.5898
R83 VGND.n18 VGND.n2 244.077
R84 VGND.n20 VGND.t3 242.025
R85 VGND.n6 VGND.n5 217.561
R86 VGND.n7 VGND.t0 154.78
R87 VGND.n2 VGND.t4 65.7148
R88 VGND.n8 VGND.n4 34.6358
R89 VGND.n12 VGND.n4 34.6358
R90 VGND.n13 VGND.n12 34.6358
R91 VGND.n14 VGND.n13 34.6358
R92 VGND.n14 VGND.n1 34.6358
R93 VGND.n7 VGND.n6 33.9541
R94 VGND.n18 VGND.n1 28.9887
R95 VGND.n5 VGND.t1 25.313
R96 VGND.n5 VGND.t5 25.313
R97 VGND.n20 VGND.n19 23.7181
R98 VGND.n19 VGND.n18 21.4593
R99 VGND.n2 VGND.t2 20.0915
R100 VGND.n21 VGND.n20 9.3005
R101 VGND.n9 VGND.n8 9.3005
R102 VGND.n10 VGND.n4 9.3005
R103 VGND.n12 VGND.n11 9.3005
R104 VGND.n13 VGND.n3 9.3005
R105 VGND.n15 VGND.n14 9.3005
R106 VGND.n16 VGND.n1 9.3005
R107 VGND.n18 VGND.n17 9.3005
R108 VGND.n19 VGND.n0 9.3005
R109 VGND.n8 VGND.n7 8.28285
R110 VGND.n9 VGND.n6 0.147198
R111 VGND.n10 VGND.n9 0.120292
R112 VGND.n11 VGND.n10 0.120292
R113 VGND.n11 VGND.n3 0.120292
R114 VGND.n15 VGND.n3 0.120292
R115 VGND.n16 VGND.n15 0.120292
R116 VGND.n17 VGND.n16 0.120292
R117 VGND.n17 VGND.n0 0.120292
R118 VGND.n21 VGND.n0 0.120292
R119 VGND VGND.n21 0.0213333
R120 a_1198_49.n2 a_1198_49.n1 590.155
R121 a_1198_49.t1 a_1198_49.n3 323.08
R122 a_1198_49.n3 a_1198_49.t2 318.813
R123 a_1198_49.n2 a_1198_49.n0 284.765
R124 a_1198_49.n1 a_1198_49.t5 209.827
R125 a_1198_49.n3 a_1198_49.n2 130.951
R126 a_1198_49.n0 a_1198_49.t4 94.7773
R127 a_1198_49.n1 a_1198_49.t0 41.5557
R128 a_1198_49.n0 a_1198_49.t3 38.438
R129 VNB.t6 VNB.t0 3445.95
R130 VNB.t8 VNB.t5 3175.4
R131 VNB.t0 VNB.t10 2648.54
R132 VNB.t9 VNB.t7 2264.08
R133 VNB.t10 VNB.t9 2150.16
R134 VNB.t7 VNB.t4 1708.74
R135 VNB.t2 VNB.t8 1523.62
R136 VNB.t4 VNB.t11 1423.95
R137 VNB.t5 VNB.t6 1253.07
R138 VNB.t11 VNB.t1 1196.12
R139 VNB.t3 VNB.t2 1196.12
R140 VNB VNB.t3 1025.24
R141 C.n0 C.t0 269.921
R142 C C.n2 155.584
R143 C.n1 C.t3 154.24
R144 C.n0 C.t1 143.286
R145 C.n2 C.n1 132.916
R146 C.n1 C.t2 102.828
R147 C.n2 C.n0 24.8308
R148 a_423_325.n3 a_423_325.n2 783.149
R149 a_423_325.n1 a_423_325.t1 728.472
R150 a_423_325.n1 a_423_325.t3 355.445
R151 a_423_325.n2 a_423_325.n0 313.538
R152 a_423_325.n2 a_423_325.n1 116.707
R153 a_423_325.n0 a_423_325.t4 98.438
R154 a_423_325.n3 a_423_325.t2 67.7193
R155 a_423_325.t0 a_423_325.n3 34.3691
R156 a_423_325.n0 a_423_325.t5 25.313
R157 a_308_93.t0 a_308_93.n1 726.078
R158 a_308_93.n1 a_308_93.t1 323.353
R159 a_308_93.n1 a_308_93.n0 256.433
R160 a_308_93.n0 a_308_93.t2 215.829
R161 a_308_93.n0 a_308_93.t3 167.63
R162 a_447_49.t3 a_447_49.n3 739.606
R163 a_447_49.n3 a_447_49.t0 380.211
R164 a_447_49.n2 a_447_49.n0 342.616
R165 a_447_49.n2 a_447_49.n1 297.875
R166 a_447_49.n4 a_447_49.t3 108.513
R167 a_447_49.n1 a_447_49.t5 85.162
R168 a_447_49.n1 a_447_49.t4 83.1099
R169 a_447_49.n0 a_447_49.t1 51.3868
R170 a_447_49.n0 a_447_49.t2 25.3226
R171 a_447_49.n3 a_447_49.n2 20.5528
R172 B.t5 B.t4 864.388
R173 B.n1 B.n0 298.841
R174 B.n0 B.t2 295.627
R175 B.n2 B.t5 235.109
R176 B.t4 B.n1 215.293
R177 B B.n2 194.166
R178 B.n0 B.t1 168.701
R179 B.n2 B.t0 167.63
R180 B.n1 B.t3 167.094
R181 a_827_297.t0 a_827_297.n3 891.352
R182 a_827_297.n0 a_827_297.t2 283.257
R183 a_827_297.n2 a_827_297.n1 224.038
R184 a_827_297.n3 a_827_297.t1 218.472
R185 a_827_297.n2 a_827_297.n0 175.175
R186 a_827_297.n1 a_827_297.t3 173.52
R187 a_827_297.n0 a_827_297.t5 161.202
R188 a_827_297.n1 a_827_297.t4 154.24
R189 a_827_297.n3 a_827_297.n2 10.4313
R190 A.n0 A.t1 239.505
R191 A.n0 A.t0 168.811
R192 A A.n0 163.52
C0 VPB X 0.004285f
C1 VPB A 0.028102f
C2 C B 0.001529f
C3 B VGND 0.034452f
C4 VPWR B 0.058719f
C5 X B 1.3e-21
C6 B A 0.002172f
C7 C VGND 0.018153f
C8 VPB B 0.295965f
C9 VPWR C 0.020896f
C10 VPWR VGND 0.098649f
C11 X C 0.001861f
C12 X VGND 0.082848f
C13 A VGND 0.01316f
C14 VPB C 0.141335f
C15 VPWR X 0.14684f
C16 VPWR A 0.014124f
C17 VPB VGND 0.012462f
C18 VPB VPWR 0.185896f
C19 VGND VNB 0.986574f
C20 A VNB 0.092322f
C21 B VNB 0.422932f
C22 C VNB 0.257768f
C23 X VNB 0.03113f
C24 VPWR VNB 0.820976f
C25 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor3_1 VNB VPB VGND VPWR X C B A
X0 a_841_297.t3 a_735_297.t2 a_355_49.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.11 pd=0.99 as=0.140825 ps=1.1 w=0.6 l=0.15
X1 a_1106_49.t2 a_841_297.t6 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1824 pd=1.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_78_199.t3 C.t0 a_355_49.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0928 pd=0.93 as=0.1728 ps=1.82 w=0.64 l=0.15
X3 a_1106_49.t1 a_735_297.t3 a_355_49.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.246 pd=1.525 as=0.2431 ps=1.445 w=0.64 l=0.15
X4 a_735_297.t0 B.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.16515 pd=1.82 as=0.1885 ps=1.88 w=0.65 l=0.15
X5 a_1106_49.t3 a_841_297.t7 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t4 A.t0 a_841_297.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1715 ps=1.355 w=1 l=0.15
X7 a_331_325.t2 B.t1 a_841_297.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.18205 pd=1.245 as=0.16275 ps=1.8 w=0.64 l=0.15
X8 a_355_49.t5 B.t2 a_841_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2431 pd=1.445 as=0.3528 ps=2.52 w=0.84 l=0.15
X9 a_216_93.t0 C.t1 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1792 pd=1.84 as=0.169 ps=1.365 w=0.64 l=0.15
X10 a_735_297.t1 B.t3 VPWR.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.25655 ps=2.52 w=1 l=0.15
X11 VPWR.t2 a_78_199.t4 X.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.365 as=0.28 ps=2.56 w=1 l=0.15
X12 a_355_49.t4 B.t4 a_1106_49.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.140825 pd=1.1 as=0.19265 ps=1.285 w=0.64 l=0.15
X13 a_331_325.t1 B.t5 a_1106_49.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1458 pd=1.205 as=0.246 ps=1.525 w=0.64 l=0.15
X14 a_331_325.t0 a_216_93.t2 a_78_199.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.224 pd=1.98 as=0.0928 ps=0.93 w=0.64 l=0.15
X15 a_78_199.t2 C.t2 a_331_325.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.15295 pd=1.315 as=0.273 ps=2.33 w=0.84 l=0.15
X16 a_355_49.t1 a_216_93.t3 a_78_199.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.32235 pd=2.45 as=0.15295 ps=1.315 w=0.84 l=0.15
X17 VGND.t1 A.t1 a_841_297.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.11 ps=0.99 w=0.64 l=0.15
X18 a_216_93.t1 C.t3 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1785 pd=1.69 as=0.1165 ps=1.035 w=0.42 l=0.15
X19 a_1106_49.t0 a_735_297.t4 a_331_325.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.19265 pd=1.285 as=0.18205 ps=1.245 w=0.42 l=0.15
X20 a_841_297.t2 a_735_297.t5 a_331_325.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1715 pd=1.355 as=0.1458 ps=1.205 w=0.84 l=0.15
X21 VGND.t4 a_78_199.t5 X.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1165 pd=1.035 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_735_297.t1 a_735_297.n3 891.352
R1 a_735_297.n0 a_735_297.t5 283.257
R2 a_735_297.n2 a_735_297.n1 224.038
R3 a_735_297.n3 a_735_297.t0 218.472
R4 a_735_297.n2 a_735_297.n0 175.175
R5 a_735_297.n1 a_735_297.t4 173.52
R6 a_735_297.n0 a_735_297.t2 161.202
R7 a_735_297.n1 a_735_297.t3 154.24
R8 a_735_297.n3 a_735_297.n2 10.4313
R9 a_355_49.t1 a_355_49.n3 739.606
R10 a_355_49.n3 a_355_49.t0 380.211
R11 a_355_49.n2 a_355_49.n0 342.616
R12 a_355_49.n2 a_355_49.n1 297.875
R13 a_355_49.n4 a_355_49.t1 108.513
R14 a_355_49.n1 a_355_49.t5 85.162
R15 a_355_49.n1 a_355_49.t2 83.1099
R16 a_355_49.n0 a_355_49.t3 51.3868
R17 a_355_49.n0 a_355_49.t4 25.3226
R18 a_355_49.n3 a_355_49.n2 20.5528
R19 a_841_297.n1 a_841_297.t5 760.636
R20 a_841_297.n6 a_841_297.n5 641.726
R21 a_841_297.n4 a_841_297.t7 241.536
R22 a_841_297.n1 a_841_297.t0 222.47
R23 a_841_297.n3 a_841_297.n2 185
R24 a_841_297.n4 a_841_297.t6 170.843
R25 a_841_297.n5 a_841_297.n4 152
R26 a_841_297.n5 a_841_297.n3 56.4377
R27 a_841_297.n0 a_841_297.t2 50.4231
R28 a_841_297.n2 a_841_297.t3 43.0005
R29 a_841_297.n7 a_841_297.n6 38.6969
R30 a_841_297.n0 a_841_297.t4 28.8712
R31 a_841_297.n3 a_841_297.n1 26.8515
R32 a_841_297.n2 a_841_297.t1 23.0795
R33 a_841_297.n6 a_841_297.n0 17.5898
R34 VNB.t3 VNB.t1 3445.95
R35 VNB.t9 VNB.t0 3175.4
R36 VNB.t1 VNB.t2 2648.54
R37 VNB.t5 VNB.t8 2264.08
R38 VNB.t2 VNB.t5 2150.16
R39 VNB.t8 VNB.t6 1708.74
R40 VNB.t10 VNB.t9 1523.62
R41 VNB.t6 VNB.t4 1423.95
R42 VNB.t0 VNB.t3 1253.07
R43 VNB.t4 VNB.t7 1196.12
R44 VNB VNB.t10 925.567
R45 VGND.n16 VGND.n15 244.077
R46 VGND.n5 VGND.n4 217.561
R47 VGND.n3 VGND.t0 154.78
R48 VGND.n15 VGND.t3 65.7148
R49 VGND.n8 VGND.n7 34.6358
R50 VGND.n9 VGND.n8 34.6358
R51 VGND.n9 VGND.n1 34.6358
R52 VGND.n13 VGND.n1 34.6358
R53 VGND.n14 VGND.n13 34.6358
R54 VGND.n5 VGND.n3 33.9541
R55 VGND.n16 VGND.n14 28.9887
R56 VGND.n4 VGND.t2 25.313
R57 VGND.n4 VGND.t1 25.313
R58 VGND.n15 VGND.t4 20.0915
R59 VGND.n7 VGND.n6 9.3005
R60 VGND.n8 VGND.n2 9.3005
R61 VGND.n10 VGND.n9 9.3005
R62 VGND.n11 VGND.n1 9.3005
R63 VGND.n13 VGND.n12 9.3005
R64 VGND.n14 VGND.n0 9.3005
R65 VGND.n7 VGND.n3 8.28285
R66 VGND.n17 VGND.n16 7.12063
R67 VGND.n17 VGND.n0 0.148519
R68 VGND.n6 VGND.n5 0.147198
R69 VGND.n6 VGND.n2 0.120292
R70 VGND.n10 VGND.n2 0.120292
R71 VGND.n11 VGND.n10 0.120292
R72 VGND.n12 VGND.n11 0.120292
R73 VGND.n12 VGND.n0 0.120292
R74 VGND VGND.n17 0.114842
R75 a_1106_49.n2 a_1106_49.n1 590.155
R76 a_1106_49.t3 a_1106_49.n3 323.08
R77 a_1106_49.n3 a_1106_49.t2 318.813
R78 a_1106_49.n2 a_1106_49.n0 284.765
R79 a_1106_49.n1 a_1106_49.t1 209.827
R80 a_1106_49.n3 a_1106_49.n2 130.951
R81 a_1106_49.n0 a_1106_49.t0 94.7773
R82 a_1106_49.n1 a_1106_49.t5 41.5557
R83 a_1106_49.n0 a_1106_49.t4 38.438
R84 C.n0 C.t2 269.921
R85 C C.n2 155.584
R86 C.n1 C.t1 154.24
R87 C.n0 C.t0 143.286
R88 C.n2 C.n1 132.916
R89 C.n1 C.t3 102.828
R90 C.n2 C.n0 24.8308
R91 a_78_199.n3 a_78_199.n2 774.88
R92 a_78_199.n2 a_78_199.n0 351.414
R93 a_78_199.n1 a_78_199.t4 236.18
R94 a_78_199.n1 a_78_199.t5 163.881
R95 a_78_199.n2 a_78_199.n1 152
R96 a_78_199.n5 a_78_199.n4 55.1605
R97 a_78_199.n3 a_78_199.t2 32.6122
R98 a_78_199.n4 a_78_199.t0 30.3415
R99 a_78_199.n0 a_78_199.t1 27.188
R100 a_78_199.n0 a_78_199.t3 27.188
R101 a_78_199.n4 a_78_199.n3 21.1076
R102 VPB.t10 VPB.t9 651.091
R103 VPB.t0 VPB.t10 627.414
R104 VPB.t6 VPB.t5 621.495
R105 VPB.t2 VPB.t8 517.913
R106 VPB.t9 VPB.t2 446.885
R107 VPB.t8 VPB.t1 304.829
R108 VPB.t4 VPB.t6 304.829
R109 VPB.t1 VPB.t7 298.911
R110 VPB.t5 VPB.t0 287.072
R111 VPB.t7 VPB.t3 248.599
R112 VPB VPB.t4 204.207
R113 B.t5 B.t2 864.388
R114 B.n1 B.n0 298.841
R115 B.n0 B.t3 295.627
R116 B.n2 B.t5 235.109
R117 B.t2 B.n1 215.293
R118 B B.n2 194.166
R119 B.n0 B.t0 168.701
R120 B.n2 B.t4 167.63
R121 B.n1 B.t1 167.094
R122 VPWR.n6 VPWR.t0 783.061
R123 VPWR.n14 VPWR.n1 719.928
R124 VPWR.n5 VPWR.n4 605.511
R125 VPWR.n1 VPWR.t3 67.7193
R126 VPWR.n8 VPWR.n7 34.6358
R127 VPWR.n8 VPWR.n2 34.6358
R128 VPWR.n12 VPWR.n2 34.6358
R129 VPWR.n13 VPWR.n12 34.6358
R130 VPWR.n1 VPWR.t2 30.3773
R131 VPWR.n4 VPWR.t1 26.5955
R132 VPWR.n4 VPWR.t4 26.5955
R133 VPWR.n14 VPWR.n13 21.0829
R134 VPWR.n7 VPWR.n6 17.6946
R135 VPWR.n7 VPWR.n3 9.3005
R136 VPWR.n9 VPWR.n8 9.3005
R137 VPWR.n10 VPWR.n2 9.3005
R138 VPWR.n12 VPWR.n11 9.3005
R139 VPWR.n13 VPWR.n0 9.3005
R140 VPWR.n6 VPWR.n5 7.29413
R141 VPWR.n15 VPWR.n14 7.1994
R142 VPWR.n5 VPWR.n3 0.151957
R143 VPWR.n15 VPWR.n0 0.147518
R144 VPWR.n9 VPWR.n3 0.120292
R145 VPWR.n10 VPWR.n9 0.120292
R146 VPWR.n11 VPWR.n10 0.120292
R147 VPWR.n11 VPWR.n0 0.120292
R148 VPWR VPWR.n15 0.115857
R149 A.n0 A.t0 239.505
R150 A.n0 A.t1 168.811
R151 A A.n0 163.52
R152 a_331_325.n3 a_331_325.n2 783.149
R153 a_331_325.n1 a_331_325.t5 728.472
R154 a_331_325.n1 a_331_325.t0 355.445
R155 a_331_325.n2 a_331_325.n0 313.538
R156 a_331_325.n2 a_331_325.n1 116.707
R157 a_331_325.n0 a_331_325.t3 98.438
R158 a_331_325.n3 a_331_325.t1 67.7193
R159 a_331_325.t4 a_331_325.n3 34.3691
R160 a_331_325.n0 a_331_325.t2 25.313
R161 a_216_93.t0 a_216_93.n1 726.078
R162 a_216_93.n1 a_216_93.t1 323.353
R163 a_216_93.n1 a_216_93.n0 256.433
R164 a_216_93.n0 a_216_93.t3 215.829
R165 a_216_93.n0 a_216_93.t2 167.63
R166 X.n1 X.n0 585
R167 X X.n0 304.337
R168 X.n1 X.t1 263.027
R169 X.n0 X.t0 26.5955
R170 X X.n1 7.54336
C0 X VGND 0.048261f
C1 VGND B 0.034452f
C2 VPB X 0.010844f
C3 X C 0.001861f
C4 VPB B 0.295962f
C5 C B 0.001529f
C6 VPB VGND 0.010825f
C7 A B 0.002172f
C8 VGND C 0.017948f
C9 VPB C 0.140023f
C10 X VPWR 0.064077f
C11 A VGND 0.01316f
C12 VPWR B 0.058718f
C13 VPB A 0.028102f
C14 VGND VPWR 0.075779f
C15 VPB VPWR 0.16937f
C16 VPWR C 0.020376f
C17 A VPWR 0.014124f
C18 X B 1.3e-21
C19 VGND VNB 0.920637f
C20 A VNB 0.092322f
C21 B VNB 0.422935f
C22 C VNB 0.259079f
C23 VPWR VNB 0.747009f
C24 X VNB 0.089675f
C25 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_4 VNB VPB VGND VPWR Y B A
X0 VGND.t7 A.t0 a_902_47.t7 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y.t7 a_38_297.t12 VPWR.t15 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297.t11 B.t0 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297.t7 B.t1 Y.t2 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t14 a_38_297.t13 Y.t6 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND.t6 A.t1 a_902_47.t6 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND.t10 B.t2 a_902_47.t10 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t11 B.t3 a_902_47.t11 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t3 B.t4 a_820_297.t6 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297.t5 A.t2 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297.t9 B.t5 a_38_47.t7 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t2 A.t3 a_38_47.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_902_47.t8 B.t6 VGND.t8 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_820_297.t5 B.t7 Y.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47.t9 B.t8 VGND.t9 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR.t9 A.t4 a_38_297.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y.t11 a_38_297.t14 a_902_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y.t10 a_38_297.t15 a_902_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_38_47.t6 B.t9 a_38_297.t10 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_38_47.t5 B.t10 a_38_297.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_38_297.t1 B.t11 a_38_47.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47.t2 A.t5 VGND.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t0 B.t12 a_38_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47.t1 A.t6 VGND.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_902_47.t1 a_38_297.t16 Y.t9 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_902_47.t2 a_38_297.t17 Y.t8 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y.t0 B.t13 a_820_297.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297.t7 A.t7 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297.t3 A.t8 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR.t7 A.t9 a_38_297.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND.t0 A.t10 a_38_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR.t5 A.t11 a_820_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47.t5 A.t12 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 a_820_297.t1 A.t13 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y.t5 a_38_297.t18 VPWR.t13 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47.t4 A.t14 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297.t3 B.t14 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR.t3 A.t15 a_820_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR.t12 a_38_297.t19 Y.t4 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR.t2 B.t15 a_38_297.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n8 A.t2 212.081
R1 A.n15 A.t4 212.081
R2 A.n9 A.t7 212.081
R3 A.n10 A.t9 212.081
R4 A.n0 A.t8 212.081
R5 A.n1 A.t11 212.081
R6 A.n3 A.t13 212.081
R7 A.n4 A.t15 212.081
R8 A.n12 A.n11 173.761
R9 A.n6 A.n5 152
R10 A.n17 A.n16 152
R11 A.n14 A.n7 152
R12 A.n13 A.n12 152
R13 A.n8 A.t6 139.78
R14 A.n15 A.t10 139.78
R15 A.n9 A.t5 139.78
R16 A.n10 A.t3 139.78
R17 A.n0 A.t0 139.78
R18 A.n1 A.t12 139.78
R19 A.n3 A.t1 139.78
R20 A.n4 A.t14 139.78
R21 A.n6 A.n2 92.1128
R22 A.n1 A.n0 61.346
R23 A.n14 A.n13 49.6611
R24 A A.n6 46.0805
R25 A.n5 A.n3 45.2793
R26 A.n16 A.n15 44.549
R27 A.n11 A.n9 43.0884
R28 A.n2 A.n1 30.289
R29 A A.n17 29.1205
R30 A.n3 A.n2 24.4894
R31 A.n17 A.n7 21.7605
R32 A.n12 A.n7 21.7605
R33 A.n11 A.n10 18.2581
R34 A.n16 A.n8 16.7975
R35 A.n5 A.n4 16.0672
R36 A.n13 A.n9 6.57323
R37 A.n15 A.n14 5.11262
R38 a_902_47.n8 a_902_47.t2 321.104
R39 a_902_47.n9 a_902_47.n8 185
R40 a_902_47.n2 a_902_47.n0 135.248
R41 a_902_47.n7 a_902_47.t3 127.519
R42 a_902_47.n2 a_902_47.n1 98.982
R43 a_902_47.n4 a_902_47.n3 98.982
R44 a_902_47.n6 a_902_47.n5 98.982
R45 a_902_47.n8 a_902_47.n7 65.2737
R46 a_902_47.n7 a_902_47.n6 60.0516
R47 a_902_47.n4 a_902_47.n2 36.2672
R48 a_902_47.n6 a_902_47.n4 36.2672
R49 a_902_47.n0 a_902_47.t6 24.9236
R50 a_902_47.n0 a_902_47.t4 24.9236
R51 a_902_47.n1 a_902_47.t7 24.9236
R52 a_902_47.n1 a_902_47.t5 24.9236
R53 a_902_47.n3 a_902_47.t10 24.9236
R54 a_902_47.n3 a_902_47.t8 24.9236
R55 a_902_47.n5 a_902_47.t11 24.9236
R56 a_902_47.n5 a_902_47.t9 24.9236
R57 a_902_47.t0 a_902_47.n9 24.9236
R58 a_902_47.n9 a_902_47.t1 24.9236
R59 VGND.n10 VGND.t11 286.447
R60 VGND.n11 VGND.n9 207.965
R61 VGND.n14 VGND.n13 207.965
R62 VGND.n20 VGND.n6 207.965
R63 VGND.n28 VGND.n3 207.965
R64 VGND.n1 VGND.n0 207.965
R65 VGND.n22 VGND.t4 153.726
R66 VGND.n32 VGND.n1 35.0835
R67 VGND.n11 VGND.n10 34.8363
R68 VGND.n15 VGND.n12 34.6358
R69 VGND.n19 VGND.n7 34.6358
R70 VGND.n23 VGND.n21 34.6358
R71 VGND.n27 VGND.n4 34.6358
R72 VGND.n30 VGND.n29 34.6358
R73 VGND.n9 VGND.t9 24.9236
R74 VGND.n9 VGND.t10 24.9236
R75 VGND.n13 VGND.t8 24.9236
R76 VGND.n13 VGND.t7 24.9236
R77 VGND.n6 VGND.t5 24.9236
R78 VGND.n6 VGND.t6 24.9236
R79 VGND.n3 VGND.t1 24.9236
R80 VGND.n3 VGND.t0 24.9236
R81 VGND.n0 VGND.t3 24.9236
R82 VGND.n0 VGND.t2 24.9236
R83 VGND.n15 VGND.n14 22.9652
R84 VGND.n29 VGND.n28 21.4593
R85 VGND.n21 VGND.n20 17.6946
R86 VGND.n20 VGND.n19 16.9417
R87 VGND.n28 VGND.n27 13.177
R88 VGND.n14 VGND.n7 11.6711
R89 VGND.n22 VGND.n4 9.41227
R90 VGND.n31 VGND.n30 9.3005
R91 VGND.n29 VGND.n2 9.3005
R92 VGND.n27 VGND.n26 9.3005
R93 VGND.n25 VGND.n4 9.3005
R94 VGND.n12 VGND.n8 9.3005
R95 VGND.n16 VGND.n15 9.3005
R96 VGND.n17 VGND.n7 9.3005
R97 VGND.n19 VGND.n18 9.3005
R98 VGND.n21 VGND.n5 9.3005
R99 VGND.n24 VGND.n23 9.3005
R100 VGND.n30 VGND.n1 7.15344
R101 VGND.n12 VGND.n11 5.64756
R102 VGND.n23 VGND.n22 4.51815
R103 VGND.n10 VGND.n8 1.62176
R104 VGND VGND.n32 0.47746
R105 VGND.n32 VGND.n31 0.147154
R106 VGND.n16 VGND.n8 0.120292
R107 VGND.n17 VGND.n16 0.120292
R108 VGND.n18 VGND.n17 0.120292
R109 VGND.n18 VGND.n5 0.120292
R110 VGND.n24 VGND.n5 0.120292
R111 VGND.n25 VGND.n24 0.120292
R112 VGND.n26 VGND.n25 0.120292
R113 VGND.n26 VGND.n2 0.120292
R114 VGND.n31 VGND.n2 0.120292
R115 VNB.t19 VNB.t5 2733.98
R116 VNB.t9 VNB.t6 2705.5
R117 VNB.t2 VNB.t4 1196.12
R118 VNB.t3 VNB.t2 1196.12
R119 VNB.t5 VNB.t3 1196.12
R120 VNB.t16 VNB.t19 1196.12
R121 VNB.t18 VNB.t16 1196.12
R122 VNB.t15 VNB.t18 1196.12
R123 VNB.t13 VNB.t15 1196.12
R124 VNB.t7 VNB.t13 1196.12
R125 VNB.t12 VNB.t7 1196.12
R126 VNB.t6 VNB.t12 1196.12
R127 VNB.t8 VNB.t9 1196.12
R128 VNB.t10 VNB.t8 1196.12
R129 VNB.t11 VNB.t10 1196.12
R130 VNB.t0 VNB.t11 1196.12
R131 VNB.t14 VNB.t0 1196.12
R132 VNB.t17 VNB.t14 1196.12
R133 VNB.t1 VNB.t17 1196.12
R134 VNB VNB.t1 1139.16
R135 a_38_297.n1 a_38_297.t5 361.038
R136 a_38_297.n1 a_38_297.n0 300.116
R137 a_38_297.n3 a_38_297.n2 300.116
R138 a_38_297.t2 a_38_297.n21 231
R139 a_38_297.n20 a_38_297.n18 226.355
R140 a_38_297.n8 a_38_297.t18 212.081
R141 a_38_297.n7 a_38_297.t19 212.081
R142 a_38_297.n13 a_38_297.t12 212.081
R143 a_38_297.n14 a_38_297.t13 212.081
R144 a_38_297.n17 a_38_297.n16 195.516
R145 a_38_297.n5 a_38_297.n4 195.25
R146 a_38_297.n20 a_38_297.n19 185
R147 a_38_297.n10 a_38_297.n9 173.761
R148 a_38_297.n16 a_38_297.n15 152
R149 a_38_297.n12 a_38_297.n6 152
R150 a_38_297.n11 a_38_297.n10 152
R151 a_38_297.n8 a_38_297.t17 139.78
R152 a_38_297.n7 a_38_297.t15 139.78
R153 a_38_297.n13 a_38_297.t16 139.78
R154 a_38_297.n14 a_38_297.t14 139.78
R155 a_38_297.n21 a_38_297.n20 59.6377
R156 a_38_297.n12 a_38_297.n11 49.6611
R157 a_38_297.n15 a_38_297.n13 45.2793
R158 a_38_297.n21 a_38_297.n17 44.424
R159 a_38_297.n9 a_38_297.n7 42.3581
R160 a_38_297.n5 a_38_297.n3 39.0276
R161 a_38_297.n3 a_38_297.n1 34.3278
R162 a_38_297.n4 a_38_297.t4 26.5955
R163 a_38_297.n4 a_38_297.t11 26.5955
R164 a_38_297.n0 a_38_297.t8 26.5955
R165 a_38_297.n0 a_38_297.t7 26.5955
R166 a_38_297.n2 a_38_297.t6 26.5955
R167 a_38_297.n2 a_38_297.t3 26.5955
R168 a_38_297.n19 a_38_297.t10 24.9236
R169 a_38_297.n19 a_38_297.t1 24.9236
R170 a_38_297.n18 a_38_297.t0 24.9236
R171 a_38_297.n18 a_38_297.t9 24.9236
R172 a_38_297.n10 a_38_297.n6 21.7605
R173 a_38_297.n16 a_38_297.n6 21.7605
R174 a_38_297.n9 a_38_297.n8 18.9884
R175 a_38_297.n15 a_38_297.n14 16.0672
R176 a_38_297.n17 a_38_297.n5 13.7692
R177 a_38_297.n11 a_38_297.n7 7.30353
R178 a_38_297.n13 a_38_297.n12 4.38232
R179 VPWR.n43 VPWR.n3 604.457
R180 VPWR.n5 VPWR.n4 604.457
R181 VPWR.n37 VPWR.n7 604.457
R182 VPWR.n30 VPWR.n29 604.457
R183 VPWR.n27 VPWR.n10 604.457
R184 VPWR.n17 VPWR.n14 321.911
R185 VPWR.n16 VPWR.n15 316.245
R186 VPWR.n45 VPWR.n1 316.245
R187 VPWR.n35 VPWR.n8 34.6358
R188 VPWR.n36 VPWR.n35 34.6358
R189 VPWR.n31 VPWR.n28 34.6358
R190 VPWR.n20 VPWR.n13 34.6358
R191 VPWR.n21 VPWR.n20 34.6358
R192 VPWR.n22 VPWR.n21 34.6358
R193 VPWR.n22 VPWR.n11 34.6358
R194 VPWR.n26 VPWR.n11 34.6358
R195 VPWR.n38 VPWR.n5 32.377
R196 VPWR.n16 VPWR.n13 27.8593
R197 VPWR.n1 VPWR.t11 26.5955
R198 VPWR.n1 VPWR.t0 26.5955
R199 VPWR.n3 VPWR.t1 26.5955
R200 VPWR.n3 VPWR.t2 26.5955
R201 VPWR.n4 VPWR.t8 26.5955
R202 VPWR.n4 VPWR.t7 26.5955
R203 VPWR.n7 VPWR.t10 26.5955
R204 VPWR.n7 VPWR.t9 26.5955
R205 VPWR.n29 VPWR.t4 26.5955
R206 VPWR.n29 VPWR.t3 26.5955
R207 VPWR.n10 VPWR.t6 26.5955
R208 VPWR.n10 VPWR.t5 26.5955
R209 VPWR.n15 VPWR.t15 26.5955
R210 VPWR.n15 VPWR.t14 26.5955
R211 VPWR.n14 VPWR.t13 26.5955
R212 VPWR.n14 VPWR.t12 26.5955
R213 VPWR.n43 VPWR.n42 26.3534
R214 VPWR.n44 VPWR.n43 24.0946
R215 VPWR.n45 VPWR.n44 20.3299
R216 VPWR.n42 VPWR.n5 18.0711
R217 VPWR.n38 VPWR.n37 12.0476
R218 VPWR.n30 VPWR.n8 11.2946
R219 VPWR.n27 VPWR.n26 10.5417
R220 VPWR.n18 VPWR.n13 9.3005
R221 VPWR.n20 VPWR.n19 9.3005
R222 VPWR.n21 VPWR.n12 9.3005
R223 VPWR.n23 VPWR.n22 9.3005
R224 VPWR.n24 VPWR.n11 9.3005
R225 VPWR.n26 VPWR.n25 9.3005
R226 VPWR.n28 VPWR.n9 9.3005
R227 VPWR.n32 VPWR.n31 9.3005
R228 VPWR.n33 VPWR.n8 9.3005
R229 VPWR.n35 VPWR.n34 9.3005
R230 VPWR.n36 VPWR.n6 9.3005
R231 VPWR.n39 VPWR.n38 9.3005
R232 VPWR.n40 VPWR.n5 9.3005
R233 VPWR.n42 VPWR.n41 9.3005
R234 VPWR.n43 VPWR.n2 9.3005
R235 VPWR.n44 VPWR.n0 9.3005
R236 VPWR.n46 VPWR.n45 7.50721
R237 VPWR.n17 VPWR.n16 6.62505
R238 VPWR.n28 VPWR.n27 5.27109
R239 VPWR.n31 VPWR.n30 4.51815
R240 VPWR.n37 VPWR.n36 3.76521
R241 VPWR.n18 VPWR.n17 0.583351
R242 VPWR.n46 VPWR.n0 0.143603
R243 VPWR.n19 VPWR.n18 0.120292
R244 VPWR.n19 VPWR.n12 0.120292
R245 VPWR.n23 VPWR.n12 0.120292
R246 VPWR.n24 VPWR.n23 0.120292
R247 VPWR.n25 VPWR.n24 0.120292
R248 VPWR.n25 VPWR.n9 0.120292
R249 VPWR.n32 VPWR.n9 0.120292
R250 VPWR.n33 VPWR.n32 0.120292
R251 VPWR.n34 VPWR.n33 0.120292
R252 VPWR.n34 VPWR.n6 0.120292
R253 VPWR.n39 VPWR.n6 0.120292
R254 VPWR.n40 VPWR.n39 0.120292
R255 VPWR.n41 VPWR.n40 0.120292
R256 VPWR.n41 VPWR.n2 0.120292
R257 VPWR.n2 VPWR.n0 0.120292
R258 VPWR VPWR.n46 0.119822
R259 Y.n2 Y.n0 626.355
R260 Y.n2 Y.n1 585
R261 Y.n8 Y.n6 226.355
R262 Y.n10 Y.t5 224.377
R263 Y.n3 Y.t6 221.239
R264 Y.n5 Y.n4 207.739
R265 Y.n8 Y.n7 185
R266 Y.n9 Y.n8 61.9695
R267 Y.n5 Y.n3 45.6965
R268 Y.n3 Y.n2 43.4717
R269 Y.n9 Y.n5 34.3278
R270 Y.n0 Y.t1 26.5955
R271 Y.n0 Y.t0 26.5955
R272 Y.n1 Y.t2 26.5955
R273 Y.n1 Y.t3 26.5955
R274 Y.n4 Y.t4 26.5955
R275 Y.n4 Y.t7 26.5955
R276 Y.n6 Y.t9 24.9236
R277 Y.n6 Y.t11 24.9236
R278 Y.n7 Y.t8 24.9236
R279 Y.n7 Y.t10 24.9236
R280 Y.n10 Y.n9 6.24292
R281 Y Y.n10 2.01239
R282 VPB.t14 VPB.t18 568.225
R283 VPB.t11 VPB.t4 562.306
R284 VPB.t16 VPB.t17 248.599
R285 VPB.t19 VPB.t16 248.599
R286 VPB.t18 VPB.t19 248.599
R287 VPB.t15 VPB.t14 248.599
R288 VPB.t12 VPB.t15 248.599
R289 VPB.t1 VPB.t12 248.599
R290 VPB.t8 VPB.t1 248.599
R291 VPB.t6 VPB.t8 248.599
R292 VPB.t5 VPB.t6 248.599
R293 VPB.t4 VPB.t5 248.599
R294 VPB.t10 VPB.t11 248.599
R295 VPB.t9 VPB.t10 248.599
R296 VPB.t7 VPB.t9 248.599
R297 VPB.t2 VPB.t7 248.599
R298 VPB.t3 VPB.t2 248.599
R299 VPB.t13 VPB.t3 248.599
R300 VPB.t0 VPB.t13 248.599
R301 VPB VPB.t0 236.761
R302 B.n15 B.n14 361.526
R303 B.n3 B.t14 212.081
R304 B.n17 B.t15 212.081
R305 B.n19 B.t0 212.081
R306 B.n1 B.t12 212.081
R307 B.n6 B.t1 212.081
R308 B.n5 B.t4 212.081
R309 B.n11 B.t7 212.081
R310 B.n12 B.t13 212.081
R311 B.n8 B.n7 173.761
R312 B.n21 B.n2 173.761
R313 B.n14 B.n13 152
R314 B.n10 B.n4 152
R315 B.n9 B.n8 152
R316 B.n16 B.n15 152
R317 B.n18 B.n0 152
R318 B.n21 B.n20 152
R319 B.n3 B.t10 139.78
R320 B.n17 B.t5 139.78
R321 B.n19 B.t9 139.78
R322 B.n1 B.t11 139.78
R323 B.n6 B.t3 139.78
R324 B.n5 B.t8 139.78
R325 B.n11 B.t2 139.78
R326 B.n12 B.t6 139.78
R327 B.n20 B.n18 49.6611
R328 B.n10 B.n9 49.6611
R329 B.n19 B.n2 45.2793
R330 B.n7 B.n5 44.549
R331 B.n13 B.n11 43.0884
R332 B.n17 B.n16 42.3581
R333 B.n8 B.n4 21.7605
R334 B.n14 B.n4 21.7605
R335 B.n15 B.n0 21.7605
R336 B.n16 B.n3 18.9884
R337 B.n13 B.n12 18.2581
R338 B B.n0 17.2805
R339 B.n7 B.n6 16.7975
R340 B.n2 B.n1 16.0672
R341 B.n18 B.n17 7.30353
R342 B.n11 B.n10 6.57323
R343 B.n9 B.n5 5.11262
R344 B B.n21 4.4805
R345 B.n20 B.n19 4.38232
R346 a_820_297.n1 a_820_297.t7 866.682
R347 a_820_297.n1 a_820_297.n0 585
R348 a_820_297.n3 a_820_297.t0 359.478
R349 a_820_297.n3 a_820_297.n2 300.116
R350 a_820_297.n5 a_820_297.n4 289.375
R351 a_820_297.n4 a_820_297.n1 49.8336
R352 a_820_297.n4 a_820_297.n3 47.2755
R353 a_820_297.n0 a_820_297.t6 26.5955
R354 a_820_297.n0 a_820_297.t5 26.5955
R355 a_820_297.n2 a_820_297.t2 26.5955
R356 a_820_297.n2 a_820_297.t1 26.5955
R357 a_820_297.n5 a_820_297.t4 26.5955
R358 a_820_297.t3 a_820_297.n5 26.5955
R359 a_38_47.n1 a_38_47.t4 306.731
R360 a_38_47.n1 a_38_47.n0 185
R361 a_38_47.n3 a_38_47.t1 174.512
R362 a_38_47.n3 a_38_47.n2 98.982
R363 a_38_47.n5 a_38_47.n4 88.3446
R364 a_38_47.n4 a_38_47.n1 53.5212
R365 a_38_47.n4 a_38_47.n3 48.9326
R366 a_38_47.n0 a_38_47.t7 24.9236
R367 a_38_47.n0 a_38_47.t6 24.9236
R368 a_38_47.n2 a_38_47.t0 24.9236
R369 a_38_47.n2 a_38_47.t2 24.9236
R370 a_38_47.t3 a_38_47.n5 24.9236
R371 a_38_47.n5 a_38_47.t5 24.9236
C0 VPB VPWR 0.188569f
C1 B A 0.475495f
C2 VGND VPWR 0.091246f
C3 VPWR Y 0.437564f
C4 VPB A 0.242642f
C5 VPB B 0.266848f
C6 VGND A 0.130724f
C7 A Y 4.84e-19
C8 B VGND 0.092495f
C9 B Y 0.029596f
C10 A VPWR 0.098039f
C11 VPB VGND 0.012173f
C12 VPB Y 0.031635f
C13 B VPWR 0.124194f
C14 VGND Y 0.034169f
C15 VGND VNB 1.09064f
C16 Y VNB 0.084111f
C17 VPWR VNB 0.886221f
C18 A VNB 0.734684f
C19 B VNB 0.748552f
C20 VPB VNB 2.0223f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297.t1 B.t0 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47.t3 A.t0 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND.t5 B.t1 a_560_47.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X3 Y.t5 B.t2 a_474_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t0 A.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t1 a_27_297.t6 a_560_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_474_297.t3 B.t3 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X7 VGND.t2 A.t2 a_560_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47.t3 B.t4 a_27_297.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297.t2 B.t5 a_27_47.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X10 a_27_47.t0 A.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t2 B.t6 a_27_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297.t1 A.t4 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47.t0 a_27_297.t7 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR.t7 A.t5 a_474_297.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y.t3 a_27_297.t8 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR.t1 a_27_297.t9 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47.t4 B.t7 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297.t4 A.t6 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t5 A.t7 a_27_297.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 B B.n2 355.976
R1 B.n3 B.t0 212.081
R2 B.n4 B.t6 212.081
R3 B.n0 B.t3 212.081
R4 B.n1 B.t2 212.081
R5 B B.n5 192.067
R6 B.n3 B.t4 139.78
R7 B.n4 B.t5 139.78
R8 B.n0 B.t1 139.78
R9 B.n1 B.t7 139.78
R10 B.n2 B.n0 38.7066
R11 B.n5 B.n3 37.246
R12 B.n2 B.n1 27.752
R13 B.n5 B.n4 24.1005
R14 VPWR.n8 VPWR.t0 845.178
R15 VPWR.n21 VPWR.n1 606.505
R16 VPWR.n19 VPWR.n3 606.505
R17 VPWR.n14 VPWR.n6 606.505
R18 VPWR.n9 VPWR.t1 340.128
R19 VPWR.n18 VPWR.n4 34.6358
R20 VPWR.n12 VPWR.n7 34.6358
R21 VPWR.n13 VPWR.n12 34.6358
R22 VPWR.n19 VPWR.n18 30.8711
R23 VPWR.n14 VPWR.n13 29.3652
R24 VPWR.n1 VPWR.t3 26.5955
R25 VPWR.n1 VPWR.t2 26.5955
R26 VPWR.n3 VPWR.t4 26.5955
R27 VPWR.n3 VPWR.t5 26.5955
R28 VPWR.n6 VPWR.t6 26.5955
R29 VPWR.n6 VPWR.t7 26.5955
R30 VPWR.n21 VPWR.n20 24.8476
R31 VPWR.n14 VPWR.n4 21.0829
R32 VPWR.n20 VPWR.n19 19.577
R33 VPWR.n8 VPWR.n7 19.2005
R34 VPWR.n10 VPWR.n7 9.3005
R35 VPWR.n12 VPWR.n11 9.3005
R36 VPWR.n13 VPWR.n5 9.3005
R37 VPWR.n15 VPWR.n14 9.3005
R38 VPWR.n16 VPWR.n4 9.3005
R39 VPWR.n18 VPWR.n17 9.3005
R40 VPWR.n19 VPWR.n2 9.3005
R41 VPWR.n20 VPWR.n0 9.3005
R42 VPWR.n22 VPWR.n21 7.32436
R43 VPWR.n9 VPWR.n8 6.90658
R44 VPWR.n10 VPWR.n9 0.684981
R45 VPWR.n22 VPWR.n0 0.145929
R46 VPWR.n11 VPWR.n10 0.120292
R47 VPWR.n11 VPWR.n5 0.120292
R48 VPWR.n15 VPWR.n5 0.120292
R49 VPWR.n16 VPWR.n15 0.120292
R50 VPWR.n17 VPWR.n16 0.120292
R51 VPWR.n17 VPWR.n2 0.120292
R52 VPWR.n2 VPWR.n0 0.120292
R53 VPWR VPWR.n22 0.117466
R54 a_27_297.n5 a_27_297.n4 409.762
R55 a_27_297.n5 a_27_297.t4 327.736
R56 a_27_297.n1 a_27_297.t0 325.964
R57 a_27_297.n7 a_27_297.n6 301.14
R58 a_27_297.n1 a_27_297.n0 263.533
R59 a_27_297.n2 a_27_297.t9 212.081
R60 a_27_297.n3 a_27_297.t8 212.081
R61 a_27_297.n2 a_27_297.t6 139.78
R62 a_27_297.n3 a_27_297.t7 139.78
R63 a_27_297.n6 a_27_297.n1 41.9561
R64 a_27_297.n6 a_27_297.n5 41.9561
R65 a_27_297.n4 a_27_297.n2 36.5157
R66 a_27_297.n7 a_27_297.t5 26.5955
R67 a_27_297.t1 a_27_297.n7 26.5955
R68 a_27_297.n0 a_27_297.t3 24.9236
R69 a_27_297.n0 a_27_297.t2 24.9236
R70 a_27_297.n4 a_27_297.n3 24.8308
R71 VPB.t6 VPB.t9 580.062
R72 VPB.t3 VPB.t1 556.386
R73 VPB.t4 VPB.t3 269.315
R74 VPB.t1 VPB.t0 248.599
R75 VPB.t8 VPB.t4 248.599
R76 VPB.t9 VPB.t8 248.599
R77 VPB.t7 VPB.t6 248.599
R78 VPB.t5 VPB.t7 248.599
R79 VPB.t2 VPB.t5 248.599
R80 VPB VPB.t2 201.246
R81 A.n0 A.t4 212.081
R82 A.n1 A.t5 212.081
R83 A.n5 A.t6 212.081
R84 A.n3 A.t7 212.081
R85 A.n7 A.n4 173.761
R86 A.n7 A.n6 152
R87 A.n0 A.t2 139.78
R88 A.n1 A.t0 139.78
R89 A.n5 A.t3 139.78
R90 A.n3 A.t1 139.78
R91 A A.n2 77.4468
R92 A.n6 A.n2 70.7153
R93 A.n2 A.n1 62.952
R94 A.n1 A.n0 61.346
R95 A.n5 A.n4 47.4702
R96 A A.n7 14.4005
R97 A.n4 A.n3 13.8763
R98 A.n6 A.n5 2.19141
R99 VGND.n6 VGND.t5 297.526
R100 VGND.n5 VGND.n4 207.965
R101 VGND.n1 VGND.n0 207.965
R102 VGND.n10 VGND.t3 157.993
R103 VGND.n14 VGND.n1 36.5921
R104 VGND.n9 VGND.n3 34.6358
R105 VGND.n12 VGND.n11 34.6358
R106 VGND.n11 VGND.n10 33.5064
R107 VGND.n5 VGND.n3 27.4829
R108 VGND.n4 VGND.t4 24.9236
R109 VGND.n4 VGND.t2 24.9236
R110 VGND.n0 VGND.t1 24.9236
R111 VGND.n0 VGND.t0 24.9236
R112 VGND.n6 VGND.n5 14.1666
R113 VGND.n7 VGND.n3 9.3005
R114 VGND.n9 VGND.n8 9.3005
R115 VGND.n11 VGND.n2 9.3005
R116 VGND.n13 VGND.n12 9.3005
R117 VGND.n12 VGND.n1 5.64756
R118 VGND.n10 VGND.n9 1.12991
R119 VGND.n7 VGND.n6 0.734599
R120 VGND VGND.n14 0.237687
R121 VGND.n14 VGND.n13 0.146169
R122 VGND.n8 VGND.n7 0.120292
R123 VGND.n8 VGND.n2 0.120292
R124 VGND.n13 VGND.n2 0.120292
R125 a_560_47.n2 a_560_47.n0 266.368
R126 a_560_47.n3 a_560_47.n2 135.248
R127 a_560_47.n2 a_560_47.n1 98.3701
R128 a_560_47.n1 a_560_47.t4 31.3851
R129 a_560_47.n0 a_560_47.t1 24.9236
R130 a_560_47.n0 a_560_47.t0 24.9236
R131 a_560_47.n1 a_560_47.t5 24.9236
R132 a_560_47.n3 a_560_47.t2 24.9236
R133 a_560_47.t3 a_560_47.n3 24.9236
R134 VNB.t2 VNB.t5 2790.94
R135 VNB.t9 VNB.t0 2677.02
R136 VNB.t6 VNB.t9 1295.79
R137 VNB.t0 VNB.t1 1196.12
R138 VNB.t3 VNB.t6 1196.12
R139 VNB.t5 VNB.t3 1196.12
R140 VNB.t4 VNB.t2 1196.12
R141 VNB.t8 VNB.t4 1196.12
R142 VNB.t7 VNB.t8 1196.12
R143 VNB VNB.t7 968.285
R144 a_474_297.n0 a_474_297.t3 873.134
R145 a_474_297.n0 a_474_297.t0 830.553
R146 a_474_297.n1 a_474_297.n0 589.33
R147 a_474_297.n1 a_474_297.t2 26.5955
R148 a_474_297.t1 a_474_297.n1 26.5955
R149 Y.n2 Y.n0 680.03
R150 Y.n3 Y.t0 325.774
R151 Y.n2 Y.n1 290.231
R152 Y.n3 Y.t1 129
R153 Y.n0 Y.t5 33.4905
R154 Y Y.n3 28.9314
R155 Y Y.n2 26.941
R156 Y.n1 Y.t2 26.5955
R157 Y.n1 Y.t3 26.5955
R158 Y.n0 Y.t4 26.5955
R159 a_27_47.n0 a_27_47.t2 312.702
R160 a_27_47.n0 a_27_47.t0 184.374
R161 a_27_47.n1 a_27_47.n0 88.3446
R162 a_27_47.t1 a_27_47.n1 24.9236
R163 a_27_47.n1 a_27_47.t3 24.9236
C0 A Y 8.81e-19
C1 VPB A 0.152874f
C2 VGND A 0.092836f
C3 A VPWR 0.063973f
C4 B Y 0.011787f
C5 VPB B 0.132775f
C6 VGND B 0.051005f
C7 VPB Y 0.01823f
C8 B VPWR 0.062845f
C9 VGND Y 0.149684f
C10 VGND VPB 0.01037f
C11 VPWR Y 0.158488f
C12 VPB VPWR 0.134233f
C13 B A 0.306814f
C14 VGND VPWR 0.093974f
C15 VGND VNB 0.67976f
C16 Y VNB 0.079956f
C17 VPWR VNB 0.576977f
C18 A VNB 0.420889f
C19 B VNB 0.385871f
C20 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297.t1 A.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47.t1 B.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47.t0 B.t1 a_47_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47.t0 B.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y.t2 a_47_47.t3 a_285_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t2 A.t1 a_129_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR.t2 A.t2 a_47_47.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t0 a_47_47.t4 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y.t0 B.t3 a_377_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47.t2 A.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n0 A.t0 266.853
R1 A.n2 A.t2 212.081
R2 A.n4 A.n0 173.761
R3 A.n4 A.n3 152
R4 A.n2 A.t1 139.78
R5 A.n1 A.t3 139.78
R6 A.n3 A.n1 37.246
R7 A.n3 A.n2 24.1005
R8 A.n1 A.n0 12.4157
R9 A A.n4 1.9205
R10 VPWR.n9 VPWR.t1 834.331
R11 VPWR.n3 VPWR.t0 777.489
R12 VPWR.n7 VPWR.n6 585
R13 VPWR.n5 VPWR.n4 585
R14 VPWR.n6 VPWR.n5 90.6205
R15 VPWR.n8 VPWR.n7 29.0829
R16 VPWR.n5 VPWR.t3 26.5955
R17 VPWR.n6 VPWR.t2 26.5955
R18 VPWR.n9 VPWR.n8 22.9652
R19 VPWR.n2 VPWR.n1 9.3005
R20 VPWR.n8 VPWR.n0 9.3005
R21 VPWR.n10 VPWR.n9 9.3005
R22 VPWR.n4 VPWR.n1 8.47109
R23 VPWR.n4 VPWR.n3 7.56025
R24 VPWR.n3 VPWR.n2 0.226309
R25 VPWR.n7 VPWR.n1 0.188735
R26 VPWR.n2 VPWR.n0 0.120292
R27 VPWR.n10 VPWR.n0 0.120292
R28 VPWR VPWR.n10 0.0226354
R29 a_377_297.t0 a_377_297.t1 41.3705
R30 VPB.t3 VPB.t4 520.872
R31 VPB.t1 VPB.t0 284.113
R32 VPB.t2 VPB.t3 248.599
R33 VPB VPB.t2 216.044
R34 VPB.t4 VPB.t1 213.084
R35 B.n2 B.n0 284.519
R36 B.n1 B.t0 241.536
R37 B.n0 B.t3 241.536
R38 B.n1 B.t1 169.237
R39 B.n0 B.t2 169.237
R40 B B.n1 166.891
R41 B B.n2 4.89462
R42 B.n2 B 4.44132
R43 a_47_47.n1 a_47_47.n0 323.671
R44 a_47_47.n2 a_47_47.n1 299.252
R45 a_47_47.n0 a_47_47.t4 241.536
R46 a_47_47.n1 a_47_47.t0 237.917
R47 a_47_47.n0 a_47_47.t3 169.237
R48 a_47_47.n2 a_47_47.t2 26.5955
R49 a_47_47.t1 a_47_47.n2 26.5955
R50 a_129_47.t0 a_129_47.t1 38.7697
R51 VNB.t3 VNB.t0 2677.02
R52 VNB VNB.t1 1210.36
R53 VNB.t0 VNB.t2 1196.12
R54 VNB.t4 VNB.t3 1196.12
R55 VNB.t1 VNB.t4 1025.24
R56 VGND.n1 VGND.t0 283.332
R57 VGND.n1 VGND.n0 128.108
R58 VGND.n0 VGND.t1 24.9236
R59 VGND.n0 VGND.t2 24.9236
R60 VGND VGND.n1 0.524018
R61 a_285_47.n0 a_285_47.t2 381.592
R62 a_285_47.n0 a_285_47.t1 24.9236
R63 a_285_47.t0 a_285_47.n0 24.9236
R64 Y Y.n0 628.915
R65 Y Y.t2 307.411
R66 Y.n0 Y.t0 38.4155
R67 Y.n0 Y.t1 26.5955
C0 B VGND 0.038916f
C1 A Y 0.001808f
C2 B VPWR 0.040822f
C3 B Y 0.003341f
C4 B A 0.23582f
C5 VPB VGND 0.005678f
C6 VPWR VPB 0.071773f
C7 VPWR VGND 0.066517f
C8 VPB Y 0.008778f
C9 A VPB 0.082204f
C10 Y VGND 0.038107f
C11 VPWR Y 0.107281f
C12 A VGND 0.063473f
C13 A VPWR 0.034894f
C14 B VPB 0.064326f
C15 VGND VNB 0.399812f
C16 Y VNB 0.078329f
C17 VPWR VNB 0.351939f
C18 A VNB 0.216579f
C19 B VNB 0.212328f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__tapvpwrvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VPWR VGND
C0 VPWR VGND 0.358072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__tapvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvgnd_1 VPB VGND VPWR
C0 VPB VPWR 0.076141f
C1 VPWR VGND 0.094626f
C2 VPB VGND 0.270365f
.ends

* NGSPICE file created from sky130_fd_sc_hd__tapvgnd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvgnd2_1 VPB VGND VPWR
C0 VPB VPWR 0.067324f
C1 VPWR VGND 0.094626f
C2 VPB VGND 0.27175f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297.t1 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47.t1 A.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_470_297.t1 A.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t0 A.t3 a_470_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47.t5 B.t0 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_470_47.t3 B.t1 X.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X6 VGND.t3 A.t4 a_112_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_112_47.t0 A.t5 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X8 VGND.t4 B.t2 a_112_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t2 A.t6 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297.t2 B.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X11 X.t1 a_112_47.t6 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR.t5 B.t4 a_470_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND.t7 a_112_47.t7 X.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t0 A.t7 a_470_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297.t2 B.t5 a_112_47.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X.t3 a_112_47.t8 a_470_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297.t5 a_112_47.t9 X.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X.t4 B.t6 a_470_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_112_47.t2 B.t7 a_27_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n3 A.t0 212.081
R1 A.n4 A.t6 212.081
R2 A.n0 A.t2 212.081
R3 A.n1 A.t3 212.081
R4 A A.n2 197.637
R5 A A.n5 189.966
R6 A.n3 A.t4 139.78
R7 A.n4 A.t5 139.78
R8 A.n0 A.t1 139.78
R9 A.n1 A.t7 139.78
R10 A.n5 A.n4 32.8641
R11 A.n2 A.n0 28.8284
R12 A.n5 A.n3 28.4823
R13 A.n2 A.n1 25.95
R14 VPWR.n4 VPWR.n3 607.784
R15 VPWR.n13 VPWR.n1 606.505
R16 VPWR.n6 VPWR.n5 606.505
R17 VPWR.n3 VPWR.t5 37.4305
R18 VPWR.n7 VPWR.n2 34.6358
R19 VPWR.n11 VPWR.n2 34.6358
R20 VPWR.n12 VPWR.n11 34.6358
R21 VPWR.n1 VPWR.t3 26.5955
R22 VPWR.n1 VPWR.t2 26.5955
R23 VPWR.n5 VPWR.t1 26.5955
R24 VPWR.n5 VPWR.t0 26.5955
R25 VPWR.n3 VPWR.t4 26.5955
R26 VPWR.n13 VPWR.n12 24.8476
R27 VPWR.n7 VPWR.n6 18.0711
R28 VPWR.n8 VPWR.n7 9.3005
R29 VPWR.n9 VPWR.n2 9.3005
R30 VPWR.n11 VPWR.n10 9.3005
R31 VPWR.n12 VPWR.n0 9.3005
R32 VPWR.n14 VPWR.n13 7.32436
R33 VPWR.n6 VPWR.n4 7.00251
R34 VPWR.n8 VPWR.n4 0.622014
R35 VPWR.n14 VPWR.n0 0.145929
R36 VPWR.n9 VPWR.n8 0.120292
R37 VPWR.n10 VPWR.n9 0.120292
R38 VPWR.n10 VPWR.n0 0.120292
R39 VPWR VPWR.n14 0.117466
R40 a_27_297.n0 a_27_297.t2 877.042
R41 a_27_297.n0 a_27_297.t0 838.697
R42 a_27_297.n1 a_27_297.n0 585
R43 a_27_297.n1 a_27_297.t3 26.5955
R44 a_27_297.t1 a_27_297.n1 26.5955
R45 VPB.t4 VPB.t8 556.386
R46 VPB.t6 VPB.t1 556.386
R47 VPB.t5 VPB.t4 281.154
R48 VPB.t8 VPB.t9 248.599
R49 VPB.t2 VPB.t5 248.599
R50 VPB.t1 VPB.t2 248.599
R51 VPB.t7 VPB.t6 248.599
R52 VPB.t3 VPB.t7 248.599
R53 VPB.t0 VPB.t3 248.599
R54 VPB VPB.t0 201.246
R55 VGND.n7 VGND.t7 298.56
R56 VGND.n8 VGND.t6 286.426
R57 VGND.n17 VGND.t4 286.426
R58 VGND.n25 VGND.t2 282.147
R59 VGND.n15 VGND.n4 207.965
R60 VGND.n23 VGND.n1 207.965
R61 VGND.n10 VGND.n9 34.6358
R62 VGND.n10 VGND.n5 34.6358
R63 VGND.n14 VGND.n5 34.6358
R64 VGND.n18 VGND.n16 34.6358
R65 VGND.n22 VGND.n2 34.6358
R66 VGND.n24 VGND.n23 32.0005
R67 VGND.n25 VGND.n24 31.2476
R68 VGND.n16 VGND.n15 27.4829
R69 VGND.n9 VGND.n8 27.1064
R70 VGND.n17 VGND.n2 25.977
R71 VGND.n4 VGND.t1 24.9236
R72 VGND.n4 VGND.t0 24.9236
R73 VGND.n1 VGND.t5 24.9236
R74 VGND.n1 VGND.t3 24.9236
R75 VGND.n8 VGND.n7 14.4172
R76 VGND.n26 VGND.n25 12.6887
R77 VGND.n9 VGND.n6 9.3005
R78 VGND.n11 VGND.n10 9.3005
R79 VGND.n12 VGND.n5 9.3005
R80 VGND.n14 VGND.n13 9.3005
R81 VGND.n16 VGND.n3 9.3005
R82 VGND.n19 VGND.n18 9.3005
R83 VGND.n20 VGND.n2 9.3005
R84 VGND.n22 VGND.n21 9.3005
R85 VGND.n24 VGND.n0 9.3005
R86 VGND.n18 VGND.n17 8.65932
R87 VGND.n15 VGND.n14 7.15344
R88 VGND.n23 VGND.n22 2.63579
R89 VGND.n7 VGND.n6 0.862225
R90 VGND.n11 VGND.n6 0.120292
R91 VGND.n12 VGND.n11 0.120292
R92 VGND.n13 VGND.n12 0.120292
R93 VGND.n13 VGND.n3 0.120292
R94 VGND.n19 VGND.n3 0.120292
R95 VGND.n20 VGND.n19 0.120292
R96 VGND.n21 VGND.n20 0.120292
R97 VGND.n21 VGND.n0 0.120292
R98 VGND.n26 VGND.n0 0.120292
R99 VGND VGND.n26 0.0226354
R100 a_470_47.n0 a_470_47.t3 319.55
R101 a_470_47.n0 a_470_47.t0 188.593
R102 a_470_47.n1 a_470_47.n0 185
R103 a_470_47.n1 a_470_47.t2 24.9236
R104 a_470_47.t1 a_470_47.n1 24.9236
R105 VNB.t7 VNB.t8 2677.02
R106 VNB.t4 VNB.t0 2677.02
R107 VNB.t5 VNB.t7 1352.75
R108 VNB.t8 VNB.t9 1196.12
R109 VNB.t3 VNB.t5 1196.12
R110 VNB.t0 VNB.t3 1196.12
R111 VNB.t6 VNB.t4 1196.12
R112 VNB.t2 VNB.t6 1196.12
R113 VNB.t1 VNB.t2 1196.12
R114 VNB VNB.t1 968.285
R115 a_470_297.n0 a_470_297.t5 374.257
R116 a_470_297.n2 a_470_297.t0 373.235
R117 a_470_297.n1 a_470_297.t2 319.096
R118 a_470_297.n0 a_470_297.t4 319.096
R119 a_470_297.n3 a_470_297.n2 301.397
R120 a_470_297.n2 a_470_297.n1 50.9181
R121 a_470_297.n3 a_470_297.t3 26.5955
R122 a_470_297.t1 a_470_297.n3 26.5955
R123 a_470_297.n1 a_470_297.n0 9.78874
R124 B.n4 B.t3 212.081
R125 B.n6 B.t4 212.081
R126 B.n0 B.t5 212.081
R127 B.n1 B.t7 212.081
R128 B.n3 B.n2 187.363
R129 B B.n7 167.361
R130 B.n5 B.n3 152.96
R131 B.n4 B.t1 139.78
R132 B.n6 B.t6 139.78
R133 B.n0 B.t2 139.78
R134 B.n1 B.t0 139.78
R135 B.n2 B.n0 54.0429
R136 B.n7 B.n5 49.6611
R137 B.n5 B.n4 10.955
R138 B.n7 B.n6 8.76414
R139 B.n2 B.n1 7.30353
R140 B B.n3 5.4405
R141 a_112_47.n7 a_112_47.n6 585
R142 a_112_47.n6 a_112_47.n2 444.329
R143 a_112_47.n0 a_112_47.t9 212.081
R144 a_112_47.n1 a_112_47.t8 212.081
R145 a_112_47.n6 a_112_47.n5 184.805
R146 a_112_47.n0 a_112_47.t7 139.78
R147 a_112_47.n1 a_112_47.t6 139.78
R148 a_112_47.n5 a_112_47.n3 135.249
R149 a_112_47.n5 a_112_47.n4 98.982
R150 a_112_47.n2 a_112_47.n0 36.5157
R151 a_112_47.t3 a_112_47.n7 26.5955
R152 a_112_47.n7 a_112_47.t2 26.5955
R153 a_112_47.n3 a_112_47.t4 24.9236
R154 a_112_47.n3 a_112_47.t5 24.9236
R155 a_112_47.n4 a_112_47.t1 24.9236
R156 a_112_47.n4 a_112_47.t0 24.9236
R157 a_112_47.n2 a_112_47.n1 24.8308
R158 X X.n0 317.051
R159 X.n3 X.n1 274.491
R160 X.n3 X.n2 185
R161 X X.n3 39.8808
R162 X.n1 X.t4 35.0774
R163 X.n0 X.t2 26.5955
R164 X.n0 X.t3 26.5955
R165 X.n2 X.t0 24.9236
R166 X.n2 X.t1 24.9236
R167 X.n1 X.t5 24.9236
C0 VPB X 0.013903f
C1 A B 0.313872f
C2 B VGND 0.168441f
C3 VPWR X 0.018034f
C4 VPB VPWR 0.120361f
C5 B X 0.060375f
C6 A VGND 0.073414f
C7 VPB B 0.123555f
C8 B VPWR 0.130416f
C9 A X 4.38e-19
C10 VPB A 0.125644f
C11 X VGND 0.111128f
C12 VPB VGND 0.006848f
C13 A VPWR 0.062291f
C14 VPWR VGND 0.039949f
C15 VGND VNB 0.716454f
C16 X VNB 0.071264f
C17 VPWR VNB 0.552562f
C18 B VNB 0.385103f
C19 A VNB 0.391494f
C20 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_4 VNB VPB VGND VPWR B X A
X0 a_27_297.t3 A.t0 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_806_47.t7 B.t0 X.t3 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_806_47.t6 B.t1 X.t2 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_112_47.t3 A.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t6 B.t2 a_112_47.t7 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_806_297.t3 a_112_47.t12 X.t9 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t15 a_112_47.t13 X.t10 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X.t1 B.t3 a_806_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X.t11 a_112_47.t14 a_806_297.t2 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_112_47.t6 B.t4 a_27_297.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_806_297.t11 B.t5 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t3 A.t2 a_806_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t0 B.t6 a_806_47.t4 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND.t2 A.t3 a_806_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_806_297.t1 a_112_47.t15 X.t4 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27245 ps=2.56 w=1 l=0.15
X15 VGND.t6 A.t4 a_112_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_112_47.t1 A.t5 VGND.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X17 VGND.t4 A.t6 a_112_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t2 A.t7 a_27_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X19 a_806_297.t10 B.t7 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t11 B.t8 a_806_297.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND.t11 B.t9 a_112_47.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND.t10 B.t10 a_112_47.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VPWR.t8 B.t11 a_806_297.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_806_47.t1 A.t8 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_806_47.t0 A.t9 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_27_297.t5 B.t12 a_112_47.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_112_47.t9 B.t13 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VGND.t12 a_112_47.t16 X.t5 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_806_297.t7 A.t10 VPWR.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2568 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 a_112_47.t8 B.t14 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_112_47.t4 B.t15 a_27_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR.t6 A.t11 a_806_297.t6 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_27_297.t1 A.t12 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X.t6 a_112_47.t17 a_806_297.t0 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 VPWR.t0 A.t13 a_27_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_806_297.t5 A.t14 VPWR.t5 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X.t7 a_112_47.t18 VGND.t13 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 X.t8 a_112_47.t19 VGND.t14 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VPWR.t4 A.t15 a_806_297.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n15 A.n14 355.125
R1 A.n3 A.t12 212.081
R2 A.n17 A.t13 212.081
R3 A.n19 A.t0 212.081
R4 A.n1 A.t7 212.081
R5 A.n6 A.t10 212.081
R6 A.n5 A.t11 212.081
R7 A.n11 A.t14 212.081
R8 A.n12 A.t15 212.081
R9 A.n8 A.n7 173.761
R10 A.n21 A.n2 173.761
R11 A.n14 A.n13 152
R12 A.n10 A.n4 152
R13 A.n9 A.n8 152
R14 A.n16 A.n15 152
R15 A.n18 A.n0 152
R16 A.n21 A.n20 152
R17 A.n3 A.t6 139.78
R18 A.n17 A.t1 139.78
R19 A.n19 A.t4 139.78
R20 A.n1 A.t5 139.78
R21 A.n6 A.t9 139.78
R22 A.n5 A.t3 139.78
R23 A.n11 A.t8 139.78
R24 A.n12 A.t2 139.78
R25 A.n20 A.n18 49.6611
R26 A.n10 A.n9 49.6611
R27 A.n19 A.n2 45.2793
R28 A.n7 A.n5 44.549
R29 A.n13 A.n11 43.0884
R30 A.n17 A.n16 42.3581
R31 A.n8 A.n4 21.7605
R32 A.n14 A.n4 21.7605
R33 A.n15 A.n0 21.7605
R34 A.n16 A.n3 18.9884
R35 A.n13 A.n12 18.2581
R36 A.n7 A.n6 16.7975
R37 A.n2 A.n1 16.0672
R38 A A.n0 13.4405
R39 A A.n21 8.3205
R40 A.n18 A.n17 7.30353
R41 A.n11 A.n10 6.57323
R42 A.n9 A.n5 5.11262
R43 A.n20 A.n19 4.38232
R44 VPWR.n12 VPWR.n11 610.095
R45 VPWR.n31 VPWR.n1 604.457
R46 VPWR.n29 VPWR.n3 604.457
R47 VPWR.n17 VPWR.n16 604.457
R48 VPWR.n15 VPWR.n8 604.457
R49 VPWR.n10 VPWR.n9 604.457
R50 VPWR.n22 VPWR.n6 34.6358
R51 VPWR.n23 VPWR.n22 34.6358
R52 VPWR.n24 VPWR.n23 34.6358
R53 VPWR.n24 VPWR.n4 34.6358
R54 VPWR.n28 VPWR.n4 34.6358
R55 VPWR.n18 VPWR.n15 34.6358
R56 VPWR.n29 VPWR.n28 30.8711
R57 VPWR.n14 VPWR.n10 28.6123
R58 VPWR.n1 VPWR.t3 26.5955
R59 VPWR.n1 VPWR.t2 26.5955
R60 VPWR.n3 VPWR.t1 26.5955
R61 VPWR.n3 VPWR.t0 26.5955
R62 VPWR.n16 VPWR.t10 26.5955
R63 VPWR.n16 VPWR.t8 26.5955
R64 VPWR.n8 VPWR.t9 26.5955
R65 VPWR.n8 VPWR.t11 26.5955
R66 VPWR.n9 VPWR.t5 26.5955
R67 VPWR.n9 VPWR.t4 26.5955
R68 VPWR.n11 VPWR.t7 26.5955
R69 VPWR.n11 VPWR.t6 26.5955
R70 VPWR.n31 VPWR.n30 24.8476
R71 VPWR.n30 VPWR.n29 19.577
R72 VPWR.n15 VPWR.n14 15.8123
R73 VPWR.n18 VPWR.n17 9.78874
R74 VPWR.n14 VPWR.n13 9.3005
R75 VPWR.n15 VPWR.n7 9.3005
R76 VPWR.n19 VPWR.n18 9.3005
R77 VPWR.n20 VPWR.n6 9.3005
R78 VPWR.n22 VPWR.n21 9.3005
R79 VPWR.n23 VPWR.n5 9.3005
R80 VPWR.n25 VPWR.n24 9.3005
R81 VPWR.n26 VPWR.n4 9.3005
R82 VPWR.n28 VPWR.n27 9.3005
R83 VPWR.n29 VPWR.n2 9.3005
R84 VPWR.n30 VPWR.n0 9.3005
R85 VPWR.n32 VPWR.n31 7.32436
R86 VPWR.n12 VPWR.n10 6.58811
R87 VPWR.n17 VPWR.n6 6.02403
R88 VPWR.n13 VPWR.n12 0.578987
R89 VPWR.n32 VPWR.n0 0.145929
R90 VPWR.n13 VPWR.n7 0.120292
R91 VPWR.n19 VPWR.n7 0.120292
R92 VPWR.n20 VPWR.n19 0.120292
R93 VPWR.n21 VPWR.n20 0.120292
R94 VPWR.n21 VPWR.n5 0.120292
R95 VPWR.n25 VPWR.n5 0.120292
R96 VPWR.n26 VPWR.n25 0.120292
R97 VPWR.n27 VPWR.n26 0.120292
R98 VPWR.n27 VPWR.n2 0.120292
R99 VPWR.n2 VPWR.n0 0.120292
R100 VPWR VPWR.n32 0.117466
R101 a_27_297.n1 a_27_297.n0 585
R102 a_27_297.n1 a_27_297.t6 376.611
R103 a_27_297.n4 a_27_297.t2 359.478
R104 a_27_297.n5 a_27_297.n4 300.116
R105 a_27_297.n3 a_27_297.n2 288.212
R106 a_27_297.n3 a_27_297.n1 61.8028
R107 a_27_297.n4 a_27_297.n3 46.2327
R108 a_27_297.n2 a_27_297.t4 26.5955
R109 a_27_297.n2 a_27_297.t1 26.5955
R110 a_27_297.n0 a_27_297.t7 26.5955
R111 a_27_297.n0 a_27_297.t5 26.5955
R112 a_27_297.n5 a_27_297.t0 26.5955
R113 a_27_297.t3 a_27_297.n5 26.5955
R114 VPB.t5 VPB.t16 562.306
R115 VPB.t14 VPB.t9 556.386
R116 VPB.t18 VPB.t17 248.599
R117 VPB.t19 VPB.t18 248.599
R118 VPB.t16 VPB.t19 248.599
R119 VPB.t4 VPB.t5 248.599
R120 VPB.t1 VPB.t4 248.599
R121 VPB.t0 VPB.t1 248.599
R122 VPB.t11 VPB.t0 248.599
R123 VPB.t13 VPB.t11 248.599
R124 VPB.t12 VPB.t13 248.599
R125 VPB.t9 VPB.t12 248.599
R126 VPB.t15 VPB.t14 248.599
R127 VPB.t10 VPB.t15 248.599
R128 VPB.t8 VPB.t10 248.599
R129 VPB.t3 VPB.t8 248.599
R130 VPB.t2 VPB.t3 248.599
R131 VPB.t7 VPB.t2 248.599
R132 VPB.t6 VPB.t7 248.599
R133 VPB VPB.t6 201.246
R134 B.n3 B.t5 212.081
R135 B.n4 B.t8 212.081
R136 B.n2 B.t7 212.081
R137 B.n8 B.t11 212.081
R138 B.n14 B.t2 212.081
R139 B.n12 B.t4 212.081
R140 B.n11 B.t12 212.081
R141 B.n10 B.t15 212.081
R142 B.n6 B.n5 173.761
R143 B.n13 B.n1 173.761
R144 B.n7 B.n6 152
R145 B.n9 B.n0 152
R146 B.n17 B.n16 152
R147 B.n15 B.n1 152
R148 B.n3 B.t0 139.78
R149 B.n4 B.t3 139.78
R150 B.n2 B.t1 139.78
R151 B.n8 B.t6 139.78
R152 B.n14 B.t10 139.78
R153 B.n12 B.t14 139.78
R154 B.n11 B.t9 139.78
R155 B.n10 B.t13 139.78
R156 B.n4 B.n3 61.346
R157 B.n12 B.n11 61.346
R158 B.n11 B.n10 61.346
R159 B.n5 B.n4 54.0429
R160 B.n16 B.n9 49.6611
R161 B.n16 B.n15 49.6611
R162 B.n7 B.n2 42.3581
R163 B.n14 B.n13 42.3581
R164 B.n9 B.n8 30.6732
R165 B.n6 B.n0 21.7605
R166 B.n17 B.n1 21.7605
R167 B B.n0 21.1205
R168 B.n8 B.n7 18.9884
R169 B.n13 B.n12 18.9884
R170 B.n5 B.n2 7.30353
R171 B.n15 B.n14 7.30353
R172 B B.n17 0.6405
R173 X.n1 X.t4 359.663
R174 X.n1 X.n0 300.116
R175 X.n10 X.t6 223.875
R176 X.n5 X.n4 219.488
R177 X.n5 X.n3 190.518
R178 X.n8 X.n7 99.1759
R179 X.n6 X.n2 98.982
R180 X.n9 X.n8 49.2684
R181 X.n9 X.n1 42.9801
R182 X.n8 X.n6 38.5935
R183 X.n6 X.n5 36.2016
R184 X.n0 X.t9 26.5955
R185 X.n0 X.t11 26.5955
R186 X.n2 X.t5 24.9236
R187 X.n2 X.t7 24.9236
R188 X.n3 X.t3 24.9236
R189 X.n3 X.t1 24.9236
R190 X.n4 X.t2 24.9236
R191 X.n4 X.t0 24.9236
R192 X.n7 X.t10 24.9236
R193 X.n7 X.t8 24.9236
R194 X.n10 X.n9 5.69353
R195 X X.n10 1.63831
R196 a_806_47.n4 a_806_47.t4 312.334
R197 a_806_47.n5 a_806_47.n4 185
R198 a_806_47.n1 a_806_47.t0 174.512
R199 a_806_47.n1 a_806_47.n0 98.982
R200 a_806_47.n3 a_806_47.n2 88.3446
R201 a_806_47.n4 a_806_47.n3 53.5212
R202 a_806_47.n3 a_806_47.n1 48.9326
R203 a_806_47.n2 a_806_47.t3 24.9236
R204 a_806_47.n2 a_806_47.t7 24.9236
R205 a_806_47.n0 a_806_47.t2 24.9236
R206 a_806_47.n0 a_806_47.t1 24.9236
R207 a_806_47.n5 a_806_47.t5 24.9236
R208 a_806_47.t6 a_806_47.n5 24.9236
R209 VNB.t0 VNB.t17 2705.5
R210 VNB.t10 VNB.t12 2677.02
R211 VNB.t18 VNB.t19 1196.12
R212 VNB.t16 VNB.t18 1196.12
R213 VNB.t17 VNB.t16 1196.12
R214 VNB.t5 VNB.t0 1196.12
R215 VNB.t1 VNB.t5 1196.12
R216 VNB.t6 VNB.t1 1196.12
R217 VNB.t15 VNB.t6 1196.12
R218 VNB.t13 VNB.t15 1196.12
R219 VNB.t14 VNB.t13 1196.12
R220 VNB.t12 VNB.t14 1196.12
R221 VNB.t8 VNB.t10 1196.12
R222 VNB.t11 VNB.t8 1196.12
R223 VNB.t9 VNB.t11 1196.12
R224 VNB.t2 VNB.t9 1196.12
R225 VNB.t7 VNB.t2 1196.12
R226 VNB.t4 VNB.t7 1196.12
R227 VNB.t3 VNB.t4 1196.12
R228 VNB VNB.t3 968.285
R229 VGND.n16 VGND.t15 292.841
R230 VGND.n20 VGND.t13 286.426
R231 VGND.n51 VGND.t5 277.336
R232 VGND.n15 VGND.n14 207.965
R233 VGND.n11 VGND.n10 207.965
R234 VGND.n26 VGND.n9 207.965
R235 VGND.n40 VGND.n4 207.965
R236 VGND.n43 VGND.n42 207.965
R237 VGND.n49 VGND.n1 207.965
R238 VGND.n34 VGND.t10 154.131
R239 VGND.n19 VGND.n13 34.6358
R240 VGND.n22 VGND.n21 34.6358
R241 VGND.n28 VGND.n27 34.6358
R242 VGND.n28 VGND.n7 34.6358
R243 VGND.n32 VGND.n7 34.6358
R244 VGND.n33 VGND.n32 34.6358
R245 VGND.n35 VGND.n33 34.6358
R246 VGND.n39 VGND.n5 34.6358
R247 VGND.n44 VGND.n41 34.6358
R248 VGND.n48 VGND.n2 34.6358
R249 VGND.n21 VGND.n20 34.2593
R250 VGND.n25 VGND.n11 32.0005
R251 VGND.n50 VGND.n49 32.0005
R252 VGND.n26 VGND.n25 31.2476
R253 VGND.n15 VGND.n13 28.2358
R254 VGND.n43 VGND.n2 25.977
R255 VGND.n14 VGND.t14 24.9236
R256 VGND.n14 VGND.t12 24.9236
R257 VGND.n10 VGND.t0 24.9236
R258 VGND.n10 VGND.t2 24.9236
R259 VGND.n9 VGND.t1 24.9236
R260 VGND.n9 VGND.t3 24.9236
R261 VGND.n4 VGND.t8 24.9236
R262 VGND.n4 VGND.t11 24.9236
R263 VGND.n42 VGND.t9 24.9236
R264 VGND.n42 VGND.t4 24.9236
R265 VGND.n1 VGND.t7 24.9236
R266 VGND.n1 VGND.t6 24.9236
R267 VGND.n51 VGND.n50 24.8476
R268 VGND.n41 VGND.n40 19.9534
R269 VGND.n40 VGND.n39 14.6829
R270 VGND.n16 VGND.n15 13.3232
R271 VGND.n52 VGND.n51 9.3005
R272 VGND.n50 VGND.n0 9.3005
R273 VGND.n48 VGND.n47 9.3005
R274 VGND.n46 VGND.n2 9.3005
R275 VGND.n45 VGND.n44 9.3005
R276 VGND.n41 VGND.n3 9.3005
R277 VGND.n39 VGND.n38 9.3005
R278 VGND.n37 VGND.n5 9.3005
R279 VGND.n17 VGND.n13 9.3005
R280 VGND.n19 VGND.n18 9.3005
R281 VGND.n21 VGND.n12 9.3005
R282 VGND.n23 VGND.n22 9.3005
R283 VGND.n25 VGND.n24 9.3005
R284 VGND.n27 VGND.n8 9.3005
R285 VGND.n29 VGND.n28 9.3005
R286 VGND.n30 VGND.n7 9.3005
R287 VGND.n32 VGND.n31 9.3005
R288 VGND.n33 VGND.n6 9.3005
R289 VGND.n36 VGND.n35 9.3005
R290 VGND.n44 VGND.n43 8.65932
R291 VGND.n34 VGND.n5 7.52991
R292 VGND.n35 VGND.n34 6.77697
R293 VGND.n27 VGND.n26 3.38874
R294 VGND.n22 VGND.n11 2.63579
R295 VGND.n49 VGND.n48 2.63579
R296 VGND.n17 VGND.n16 0.826837
R297 VGND.n20 VGND.n19 0.376971
R298 VGND.n18 VGND.n17 0.120292
R299 VGND.n18 VGND.n12 0.120292
R300 VGND.n23 VGND.n12 0.120292
R301 VGND.n24 VGND.n23 0.120292
R302 VGND.n24 VGND.n8 0.120292
R303 VGND.n29 VGND.n8 0.120292
R304 VGND.n30 VGND.n29 0.120292
R305 VGND.n31 VGND.n30 0.120292
R306 VGND.n31 VGND.n6 0.120292
R307 VGND.n36 VGND.n6 0.120292
R308 VGND.n37 VGND.n36 0.120292
R309 VGND.n38 VGND.n37 0.120292
R310 VGND.n38 VGND.n3 0.120292
R311 VGND.n45 VGND.n3 0.120292
R312 VGND.n46 VGND.n45 0.120292
R313 VGND.n47 VGND.n46 0.120292
R314 VGND.n47 VGND.n0 0.120292
R315 VGND.n52 VGND.n0 0.120292
R316 VGND VGND.n52 0.0226354
R317 a_112_47.n19 a_112_47.n18 634.13
R318 a_112_47.n18 a_112_47.n0 589.609
R319 a_112_47.n9 a_112_47.t17 212.081
R320 a_112_47.n11 a_112_47.t12 212.081
R321 a_112_47.n14 a_112_47.t14 212.081
R322 a_112_47.n13 a_112_47.t15 212.081
R323 a_112_47.n17 a_112_47.n7 211.018
R324 a_112_47.n10 a_112_47.n8 173.761
R325 a_112_47.n16 a_112_47.n15 152
R326 a_112_47.n12 a_112_47.n8 152
R327 a_112_47.n9 a_112_47.t13 139.78
R328 a_112_47.n11 a_112_47.t19 139.78
R329 a_112_47.n14 a_112_47.t16 139.78
R330 a_112_47.n13 a_112_47.t18 139.78
R331 a_112_47.n3 a_112_47.n1 135.249
R332 a_112_47.n17 a_112_47.n16 118.1
R333 a_112_47.n3 a_112_47.n2 98.982
R334 a_112_47.n5 a_112_47.n4 98.982
R335 a_112_47.n7 a_112_47.n6 98.982
R336 a_112_47.n14 a_112_47.n13 61.346
R337 a_112_47.n15 a_112_47.n12 49.6611
R338 a_112_47.n11 a_112_47.n10 42.3581
R339 a_112_47.n18 a_112_47.n17 37.1054
R340 a_112_47.n5 a_112_47.n3 36.2672
R341 a_112_47.n7 a_112_47.n5 36.2672
R342 a_112_47.n0 a_112_47.t5 26.5955
R343 a_112_47.n0 a_112_47.t4 26.5955
R344 a_112_47.t7 a_112_47.n19 26.5955
R345 a_112_47.n19 a_112_47.t6 26.5955
R346 a_112_47.n6 a_112_47.t2 24.9236
R347 a_112_47.n6 a_112_47.t1 24.9236
R348 a_112_47.n1 a_112_47.t10 24.9236
R349 a_112_47.n1 a_112_47.t8 24.9236
R350 a_112_47.n2 a_112_47.t11 24.9236
R351 a_112_47.n2 a_112_47.t9 24.9236
R352 a_112_47.n4 a_112_47.t0 24.9236
R353 a_112_47.n4 a_112_47.t3 24.9236
R354 a_112_47.n16 a_112_47.n8 21.7605
R355 a_112_47.n10 a_112_47.n9 18.9884
R356 a_112_47.n12 a_112_47.n11 7.30353
R357 a_112_47.n15 a_112_47.n14 4.38232
R358 a_806_297.n1 a_806_297.t8 361.039
R359 a_806_297.n9 a_806_297.n8 345.31
R360 a_806_297.n6 a_806_297.t7 319.957
R361 a_806_297.n1 a_806_297.n0 300.116
R362 a_806_297.n3 a_806_297.n2 300.116
R363 a_806_297.n8 a_806_297.n7 298.837
R364 a_806_297.n5 a_806_297.n4 199.951
R365 a_806_297.n8 a_806_297.n6 65.3793
R366 a_806_297.n6 a_806_297.n5 46.2327
R367 a_806_297.n3 a_806_297.n1 34.3278
R368 a_806_297.n5 a_806_297.n3 34.3278
R369 a_806_297.n0 a_806_297.t9 26.5955
R370 a_806_297.n0 a_806_297.t10 26.5955
R371 a_806_297.n2 a_806_297.t4 26.5955
R372 a_806_297.n2 a_806_297.t11 26.5955
R373 a_806_297.n4 a_806_297.t6 26.5955
R374 a_806_297.n4 a_806_297.t5 26.5955
R375 a_806_297.n7 a_806_297.t2 26.5955
R376 a_806_297.n7 a_806_297.t1 26.5955
R377 a_806_297.n9 a_806_297.t0 26.5955
R378 a_806_297.t3 a_806_297.n9 26.5955
C0 X B 0.167049f
C1 VGND A 0.110666f
C2 VPB B 0.277445f
C3 B VPWR 0.073916f
C4 X A 0.03715f
C5 VPB A 0.266328f
C6 X VGND 0.508897f
C7 VPB VGND 0.008234f
C8 A VPWR 0.143854f
C9 VGND VPWR 0.075216f
C10 VPB X 0.031084f
C11 A B 0.458625f
C12 VGND B 0.113419f
C13 X VPWR 0.095212f
C14 VPB VPWR 0.18434f
C15 VGND VNB 1.12322f
C16 X VNB 0.113613f
C17 VPWR VNB 0.886255f
C18 B VNB 0.783492f
C19 A VNB 0.748649f
C20 VPB VNB 2.0223f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_1 VNB VPB VGND VPWR X C B A
X0 a_112_21.t0 C.t0 a_404_49.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.04 as=0.1728 ps=1.82 w=0.64 l=0.15
X1 a_1198_49.t5 a_931_365.t6 VGND.t4 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1824 pd=1.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_386_325.t0 B.t0 a_1198_49.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.140825 pd=1.1 as=0.19265 ps=1.285 w=0.64 l=0.15
X3 a_404_49.t5 a_266_93.t2 a_112_21.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.441 pd=2.73 as=0.1596 ps=1.22 w=0.84 l=0.15
X4 a_931_365.t2 a_827_297.t2 a_404_49.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1715 pd=1.355 as=0.1458 ps=1.205 w=0.84 l=0.15
X5 VPWR.t2 a_112_21.t4 X.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.2115 pd=1.45 as=0.28 ps=2.56 w=1 l=0.15
X6 a_827_297.t1 B.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1653 pd=1.82 as=0.195 ps=1.9 w=0.65 l=0.15
X7 a_1198_49.t2 a_827_297.t3 a_404_49.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.19265 pd=1.285 as=0.18365 ps=1.25 w=0.42 l=0.15
X8 VGND.t3 A.t0 a_931_365.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.11 ps=0.99 w=0.64 l=0.15
X9 a_112_21.t1 C.t1 a_386_325.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1596 pd=1.22 as=0.2688 ps=2.32 w=0.84 l=0.15
X10 a_1198_49.t1 a_827_297.t4 a_386_325.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.246 pd=1.525 as=0.2452 ps=1.45 w=0.64 l=0.15
X11 a_266_93.t0 C.t2 VPWR.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1792 pd=1.84 as=0.2115 ps=1.45 w=0.64 l=0.15
X12 a_1198_49.t4 a_931_365.t7 VPWR.t4 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X13 a_931_365.t4 a_827_297.t5 a_386_325.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.11 pd=0.99 as=0.140825 ps=1.1 w=0.6 l=0.15
X14 VPWR.t1 A.t1 a_931_365.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1715 ps=1.355 w=1 l=0.15
X15 a_827_297.t0 B.t2 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2526 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X16 VGND.t1 a_112_21.t5 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.144125 pd=1.12 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_386_325.t1 B.t3 a_931_365.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2452 pd=1.45 as=0.3536 ps=2.53 w=0.84 l=0.15
X18 a_266_93.t1 C.t3 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1764 pd=1.68 as=0.144125 ps=1.12 w=0.42 l=0.15
X19 a_404_49.t2 B.t4 a_931_365.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.18365 pd=1.25 as=0.1628 ps=1.8 w=0.64 l=0.15
X20 a_386_325.t5 a_266_93.t3 a_112_21.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.3168 pd=2.27 as=0.128 ps=1.04 w=0.64 l=0.15
X21 a_404_49.t3 B.t5 a_1198_49.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1458 pd=1.205 as=0.246 ps=1.525 w=0.64 l=0.15
R0 C.n0 C.t1 229.136
R1 C.n1 C.t2 154.24
R2 C.n0 C.t0 140.992
R3 C.n2 C.n1 125.09
R4 C.n1 C.t3 102.828
R5 C C.n2 68.4649
R6 C.n2 C.n0 27.396
R7 a_404_49.n3 a_404_49.n2 783.902
R8 a_404_49.n1 a_404_49.t5 723.856
R9 a_404_49.n1 a_404_49.t4 500.06
R10 a_404_49.n2 a_404_49.n0 310.861
R11 a_404_49.n2 a_404_49.n1 115.954
R12 a_404_49.n0 a_404_49.t0 99.3755
R13 a_404_49.n3 a_404_49.t3 67.7193
R14 a_404_49.t1 a_404_49.n3 34.3691
R15 a_404_49.n0 a_404_49.t2 25.313
R16 a_112_21.n3 a_112_21.n2 780.408
R17 a_112_21.n2 a_112_21.n0 352.341
R18 a_112_21.n1 a_112_21.t4 231.478
R19 a_112_21.n1 a_112_21.t5 159.179
R20 a_112_21.n2 a_112_21.n1 152
R21 a_112_21.n0 a_112_21.t3 49.688
R22 a_112_21.n3 a_112_21.t2 46.9053
R23 a_112_21.t1 a_112_21.n3 42.2148
R24 a_112_21.n0 a_112_21.t0 25.313
R25 VNB.t9 VNB.t2 3730.74
R26 VNB.t6 VNB.t7 3161.17
R27 VNB.t2 VNB.t5 2648.54
R28 VNB.t3 VNB.t1 2264.08
R29 VNB.t5 VNB.t3 2164.4
R30 VNB.t4 VNB.t6 1765.7
R31 VNB.t1 VNB.t8 1708.74
R32 VNB.t7 VNB.t9 1566.34
R33 VNB.t8 VNB.t10 1423.95
R34 VNB VNB.t4 1395.47
R35 VNB.t10 VNB.t0 1196.12
R36 a_931_365.n1 a_931_365.t1 775.927
R37 a_931_365.n6 a_931_365.n5 641.726
R38 a_931_365.n4 a_931_365.t7 241.536
R39 a_931_365.n1 a_931_365.t3 222.323
R40 a_931_365.n3 a_931_365.n2 185
R41 a_931_365.n4 a_931_365.t6 170.843
R42 a_931_365.n5 a_931_365.n4 152
R43 a_931_365.n5 a_931_365.n3 56.4377
R44 a_931_365.n0 a_931_365.t2 50.4231
R45 a_931_365.n2 a_931_365.t4 43.0005
R46 a_931_365.n7 a_931_365.n6 38.6969
R47 a_931_365.n0 a_931_365.t0 28.8712
R48 a_931_365.n3 a_931_365.n1 26.8515
R49 a_931_365.n2 a_931_365.t5 23.0795
R50 a_931_365.n6 a_931_365.n0 17.5898
R51 VGND.n7 VGND.n6 217.561
R52 VGND.n1 VGND.n0 213.868
R53 VGND.n5 VGND.t0 153.607
R54 VGND.n0 VGND.t2 78.5719
R55 VGND.n0 VGND.t1 36.0005
R56 VGND.n10 VGND.n9 34.6358
R57 VGND.n11 VGND.n10 34.6358
R58 VGND.n11 VGND.n3 34.6358
R59 VGND.n15 VGND.n3 34.6358
R60 VGND.n16 VGND.n15 34.6358
R61 VGND.n17 VGND.n16 34.6358
R62 VGND.n7 VGND.n5 34.3305
R63 VGND.n6 VGND.t4 25.313
R64 VGND.n6 VGND.t3 25.313
R65 VGND.n19 VGND.n1 12.9297
R66 VGND.n17 VGND.n1 10.5417
R67 VGND.n9 VGND.n8 9.3005
R68 VGND.n10 VGND.n4 9.3005
R69 VGND.n12 VGND.n11 9.3005
R70 VGND.n13 VGND.n3 9.3005
R71 VGND.n15 VGND.n14 9.3005
R72 VGND.n16 VGND.n2 9.3005
R73 VGND.n18 VGND.n17 9.3005
R74 VGND.n9 VGND.n5 7.90638
R75 VGND.n8 VGND.n7 0.147198
R76 VGND.n19 VGND.n18 0.141672
R77 VGND VGND.n19 0.121778
R78 VGND.n8 VGND.n4 0.120292
R79 VGND.n12 VGND.n4 0.120292
R80 VGND.n13 VGND.n12 0.120292
R81 VGND.n14 VGND.n13 0.120292
R82 VGND.n14 VGND.n2 0.120292
R83 VGND.n18 VGND.n2 0.120292
R84 a_1198_49.n2 a_1198_49.n1 590.155
R85 a_1198_49.t4 a_1198_49.n3 323.08
R86 a_1198_49.n3 a_1198_49.t5 318.813
R87 a_1198_49.n2 a_1198_49.n0 284.765
R88 a_1198_49.n1 a_1198_49.t1 209.827
R89 a_1198_49.n3 a_1198_49.n2 130.951
R90 a_1198_49.n0 a_1198_49.t2 94.7773
R91 a_1198_49.n1 a_1198_49.t3 41.5557
R92 a_1198_49.n0 a_1198_49.t0 38.438
R93 B.t5 B.t3 865.994
R94 B.n1 B.n0 298.841
R95 B.n0 B.t2 294.021
R96 B.n2 B.t5 235.109
R97 B.t3 B.n1 215.293
R98 B B.n2 194.166
R99 B.n0 B.t1 168.701
R100 B.n2 B.t0 167.63
R101 B.n1 B.t4 167.094
R102 a_386_325.n1 a_386_325.t3 720.771
R103 a_386_325.n2 a_386_325.n0 342.616
R104 a_386_325.n1 a_386_325.t5 302.955
R105 a_386_325.n3 a_386_325.n2 297.875
R106 a_386_325.n3 a_386_325.t2 83.1099
R107 a_386_325.n0 a_386_325.t4 51.3868
R108 a_386_325.n4 a_386_325.t1 40.7642
R109 a_386_325.n5 a_386_325.n4 39.4005
R110 a_386_325.n4 a_386_325.n3 27.7036
R111 a_386_325.n0 a_386_325.t0 25.3226
R112 a_386_325.n2 a_386_325.n1 20.5528
R113 a_266_93.t0 a_266_93.n1 725.702
R114 a_266_93.n1 a_266_93.t1 321.925
R115 a_266_93.n1 a_266_93.n0 261.704
R116 a_266_93.n0 a_266_93.t2 260.817
R117 a_266_93.n0 a_266_93.t3 167.63
R118 VPB.t0 VPB.t3 713.24
R119 VPB.t3 VPB.t2 648.131
R120 VPB.t8 VPB.t9 633.333
R121 VPB.t4 VPB.t1 517.913
R122 VPB.t2 VPB.t4 449.844
R123 VPB.t7 VPB.t8 355.14
R124 VPB.t9 VPB.t0 313.707
R125 VPB.t1 VPB.t6 304.829
R126 VPB VPB.t7 301.87
R127 VPB.t6 VPB.t5 298.911
R128 VPB.t5 VPB.t10 248.599
R129 a_827_297.t0 a_827_297.n3 802.28
R130 a_827_297.n0 a_827_297.t2 283.257
R131 a_827_297.n2 a_827_297.n1 224.564
R132 a_827_297.n3 a_827_297.t1 219.297
R133 a_827_297.n2 a_827_297.n0 175.175
R134 a_827_297.n1 a_827_297.t3 173.52
R135 a_827_297.n0 a_827_297.t5 161.202
R136 a_827_297.n1 a_827_297.t4 154.24
R137 a_827_297.n4 a_827_297.t0 102.441
R138 a_827_297.n3 a_827_297.n2 10.4313
R139 X.n1 X.n0 585
R140 X X.n0 298.827
R141 X.n1 X.t1 244.49
R142 X.n0 X.t0 26.5955
R143 X X.n1 4.02336
R144 VPWR.n4 VPWR.t0 854.342
R145 VPWR.n16 VPWR.n1 620.202
R146 VPWR.n6 VPWR.n5 605.511
R147 VPWR.n1 VPWR.t3 81.5708
R148 VPWR.n1 VPWR.t2 36.4455
R149 VPWR.n9 VPWR.n8 34.6358
R150 VPWR.n10 VPWR.n9 34.6358
R151 VPWR.n10 VPWR.n2 34.6358
R152 VPWR.n14 VPWR.n2 34.6358
R153 VPWR.n15 VPWR.n14 34.6358
R154 VPWR.n5 VPWR.t4 26.5955
R155 VPWR.n5 VPWR.t1 26.5955
R156 VPWR.n8 VPWR.n4 17.6946
R157 VPWR.n17 VPWR.n16 14.4356
R158 VPWR.n8 VPWR.n7 9.3005
R159 VPWR.n9 VPWR.n3 9.3005
R160 VPWR.n11 VPWR.n10 9.3005
R161 VPWR.n12 VPWR.n2 9.3005
R162 VPWR.n14 VPWR.n13 9.3005
R163 VPWR.n15 VPWR.n0 9.3005
R164 VPWR.n6 VPWR.n4 7.29413
R165 VPWR.n16 VPWR.n15 2.63579
R166 VPWR.n7 VPWR.n6 0.151957
R167 VPWR.n17 VPWR.n0 0.141672
R168 VPWR VPWR.n17 0.121778
R169 VPWR.n7 VPWR.n3 0.120292
R170 VPWR.n11 VPWR.n3 0.120292
R171 VPWR.n12 VPWR.n11 0.120292
R172 VPWR.n13 VPWR.n12 0.120292
R173 VPWR.n13 VPWR.n0 0.120292
R174 A.n0 A.t1 239.505
R175 A.n0 A.t0 168.811
R176 A A.n0 163.52
C0 VPWR B 0.058835f
C1 X C 0.002594f
C2 VGND VPB 0.011484f
C3 X B 1.21e-20
C4 X VPWR 0.096872f
C5 A VGND 0.01316f
C6 C VGND 0.01954f
C7 A VPB 0.028102f
C8 C VPB 0.137768f
C9 B VGND 0.034605f
C10 VPWR VGND 0.084689f
C11 B VPB 0.296884f
C12 VPWR VPB 0.17396f
C13 B A 0.002172f
C14 X VGND 0.075093f
C15 C B 5.03e-19
C16 VPWR A 0.014124f
C17 VPWR C 0.020771f
C18 X VPB 0.019314f
C19 VGND VNB 0.968822f
C20 A VNB 0.092322f
C21 B VNB 0.423782f
C22 C VNB 0.262015f
C23 VPWR VNB 0.788863f
C24 X VNB 0.094793f
C25 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_2 VNB VPB VGND VPWR X C B A
X0 a_120_21.t2 C.t0 a_496_49.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.04 as=0.1728 ps=1.82 w=0.64 l=0.15
X1 a_1023_365.t3 a_919_297.t2 a_478_325.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.11 pd=0.99 as=0.140825 ps=1.1 w=0.6 l=0.15
X2 VGND.t3 a_120_21.t4 X.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.144125 pd=1.12 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_358_93.t0 C.t1 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1764 pd=1.68 as=0.144125 ps=1.12 w=0.42 l=0.15
X4 a_496_49.t1 B.t0 a_1023_365.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.18365 pd=1.25 as=0.1628 ps=1.8 w=0.64 l=0.15
X5 a_496_49.t2 B.t1 a_1290_49.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1458 pd=1.205 as=0.246 ps=1.525 w=0.64 l=0.15
X6 a_1290_49.t2 a_919_297.t3 a_496_49.t4 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.19265 pd=1.285 as=0.18365 ps=1.25 w=0.42 l=0.15
X7 a_496_49.t0 a_358_93.t2 a_120_21.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.441 pd=2.73 as=0.1596 ps=1.22 w=0.84 l=0.15
X8 a_1023_365.t2 a_919_297.t4 a_496_49.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1715 pd=1.355 as=0.1458 ps=1.205 w=0.84 l=0.15
X9 a_1290_49.t4 a_1023_365.t6 VGND.t4 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 VPWR.t3 a_120_21.t5 X.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.2115 pd=1.45 as=0.135 ps=1.27 w=1 l=0.15
X11 a_478_325.t0 B.t2 a_1290_49.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.140825 pd=1.1 as=0.19265 ps=1.285 w=0.64 l=0.15
X12 X.t0 a_120_21.t6 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_1290_49.t3 a_919_297.t5 a_478_325.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.246 pd=1.525 as=0.2452 ps=1.45 w=0.64 l=0.15
X14 a_919_297.t0 B.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1653 pd=1.82 as=0.195 ps=1.9 w=0.65 l=0.15
X15 a_120_21.t3 C.t2 a_478_325.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1596 pd=1.22 as=0.2688 ps=2.32 w=0.84 l=0.15
X16 a_358_93.t1 C.t3 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1792 pd=1.84 as=0.2115 ps=1.45 w=0.64 l=0.15
X17 a_1290_49.t5 a_1023_365.t7 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND.t1 A.t0 a_1023_365.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.11 ps=0.99 w=0.64 l=0.15
X19 X.t1 a_120_21.t7 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 VPWR.t0 A.t1 a_1023_365.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1715 ps=1.355 w=1 l=0.15
X21 a_919_297.t1 B.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2526 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 a_478_325.t1 B.t5 a_1023_365.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2452 pd=1.45 as=0.3536 ps=2.53 w=0.84 l=0.15
X23 a_478_325.t4 a_358_93.t3 a_120_21.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.3168 pd=2.27 as=0.128 ps=1.04 w=0.64 l=0.15
R0 C.n0 C.t2 229.136
R1 C.n1 C.t3 154.24
R2 C.n0 C.t0 140.992
R3 C.n2 C.n1 125.09
R4 C.n1 C.t1 102.828
R5 C C.n2 68.4649
R6 C.n2 C.n0 27.396
R7 a_496_49.n2 a_496_49.n1 783.902
R8 a_496_49.t0 a_496_49.n3 723.856
R9 a_496_49.n3 a_496_49.t3 500.06
R10 a_496_49.n2 a_496_49.n0 310.861
R11 a_496_49.n3 a_496_49.n2 115.954
R12 a_496_49.n0 a_496_49.t4 99.3755
R13 a_496_49.n1 a_496_49.t2 67.7193
R14 a_496_49.n1 a_496_49.t5 34.3691
R15 a_496_49.n0 a_496_49.t1 25.313
R16 a_120_21.n5 a_120_21.n4 780.408
R17 a_120_21.n4 a_120_21.n0 352.341
R18 a_120_21.n3 a_120_21.t5 212.081
R19 a_120_21.n1 a_120_21.t6 212.081
R20 a_120_21.n4 a_120_21.n3 178.292
R21 a_120_21.n1 a_120_21.t7 142.702
R22 a_120_21.n2 a_120_21.t4 139.78
R23 a_120_21.n2 a_120_21.n1 58.4247
R24 a_120_21.n0 a_120_21.t1 49.688
R25 a_120_21.t0 a_120_21.n5 46.9053
R26 a_120_21.n5 a_120_21.t3 42.2148
R27 a_120_21.n0 a_120_21.t2 25.313
R28 a_120_21.n3 a_120_21.n2 2.92171
R29 VNB.t2 VNB.t1 3730.74
R30 VNB.t7 VNB.t8 3161.17
R31 VNB.t1 VNB.t3 2648.54
R32 VNB.t10 VNB.t0 2264.08
R33 VNB.t3 VNB.t10 2164.4
R34 VNB.t6 VNB.t7 1765.7
R35 VNB.t0 VNB.t9 1708.74
R36 VNB.t8 VNB.t2 1566.34
R37 VNB VNB.t5 1509.39
R38 VNB.t9 VNB.t4 1423.95
R39 VNB.t4 VNB.t11 1196.12
R40 VNB.t5 VNB.t6 1196.12
R41 a_919_297.t1 a_919_297.n3 802.28
R42 a_919_297.n0 a_919_297.t4 283.257
R43 a_919_297.n2 a_919_297.n1 224.564
R44 a_919_297.n3 a_919_297.t0 219.297
R45 a_919_297.n2 a_919_297.n0 175.175
R46 a_919_297.n1 a_919_297.t3 173.52
R47 a_919_297.n0 a_919_297.t2 161.202
R48 a_919_297.n1 a_919_297.t5 154.24
R49 a_919_297.n4 a_919_297.t1 102.441
R50 a_919_297.n3 a_919_297.n2 10.4313
R51 a_478_325.n1 a_478_325.t5 720.771
R52 a_478_325.n2 a_478_325.n0 342.616
R53 a_478_325.n1 a_478_325.t4 302.955
R54 a_478_325.n3 a_478_325.n2 297.875
R55 a_478_325.n3 a_478_325.t3 83.1099
R56 a_478_325.n0 a_478_325.t2 51.3868
R57 a_478_325.n4 a_478_325.t1 40.7642
R58 a_478_325.n5 a_478_325.n4 39.4005
R59 a_478_325.n4 a_478_325.n3 27.7036
R60 a_478_325.n0 a_478_325.t0 25.3226
R61 a_478_325.n2 a_478_325.n1 20.5528
R62 a_1023_365.n1 a_1023_365.t0 775.927
R63 a_1023_365.n6 a_1023_365.n5 641.726
R64 a_1023_365.n4 a_1023_365.t7 241.536
R65 a_1023_365.n1 a_1023_365.t4 222.323
R66 a_1023_365.n3 a_1023_365.n2 185
R67 a_1023_365.n4 a_1023_365.t6 170.843
R68 a_1023_365.n5 a_1023_365.n4 152
R69 a_1023_365.n5 a_1023_365.n3 56.4377
R70 a_1023_365.n0 a_1023_365.t2 50.4231
R71 a_1023_365.n2 a_1023_365.t3 43.0005
R72 a_1023_365.n7 a_1023_365.n6 38.6969
R73 a_1023_365.n0 a_1023_365.t1 28.8712
R74 a_1023_365.n3 a_1023_365.n1 26.8515
R75 a_1023_365.n2 a_1023_365.t5 23.0795
R76 a_1023_365.n6 a_1023_365.n0 17.5898
R77 X.n2 X.n0 224.799
R78 X.n2 X.n1 197.626
R79 X.n1 X.t3 26.5955
R80 X.n1 X.t0 26.5955
R81 X.n0 X.t2 24.9236
R82 X.n0 X.t1 24.9236
R83 X X.n2 1.36001
R84 VGND.n23 VGND.t2 282.817
R85 VGND.n8 VGND.n7 217.561
R86 VGND.n2 VGND.n1 213.868
R87 VGND.n6 VGND.t0 153.607
R88 VGND.n1 VGND.t5 78.5719
R89 VGND.n1 VGND.t3 36.0005
R90 VGND.n11 VGND.n10 34.6358
R91 VGND.n12 VGND.n11 34.6358
R92 VGND.n12 VGND.n4 34.6358
R93 VGND.n16 VGND.n4 34.6358
R94 VGND.n17 VGND.n16 34.6358
R95 VGND.n18 VGND.n17 34.6358
R96 VGND.n22 VGND.n21 34.6358
R97 VGND.n8 VGND.n6 34.3305
R98 VGND.n7 VGND.t4 25.313
R99 VGND.n7 VGND.t1 25.313
R100 VGND.n24 VGND.n23 14.5711
R101 VGND.n18 VGND.n2 10.5417
R102 VGND.n10 VGND.n9 9.3005
R103 VGND.n11 VGND.n5 9.3005
R104 VGND.n13 VGND.n12 9.3005
R105 VGND.n14 VGND.n4 9.3005
R106 VGND.n16 VGND.n15 9.3005
R107 VGND.n17 VGND.n3 9.3005
R108 VGND.n19 VGND.n18 9.3005
R109 VGND.n21 VGND.n20 9.3005
R110 VGND.n22 VGND.n0 9.3005
R111 VGND.n10 VGND.n6 7.90638
R112 VGND.n21 VGND.n2 5.27109
R113 VGND.n23 VGND.n22 4.51815
R114 VGND.n9 VGND.n8 0.147198
R115 VGND.n9 VGND.n5 0.120292
R116 VGND.n13 VGND.n5 0.120292
R117 VGND.n14 VGND.n13 0.120292
R118 VGND.n15 VGND.n14 0.120292
R119 VGND.n15 VGND.n3 0.120292
R120 VGND.n19 VGND.n3 0.120292
R121 VGND.n20 VGND.n19 0.120292
R122 VGND.n20 VGND.n0 0.120292
R123 VGND.n24 VGND.n0 0.120292
R124 VGND VGND.n24 0.0226354
R125 a_358_93.t1 a_358_93.n1 725.702
R126 a_358_93.n1 a_358_93.t0 321.925
R127 a_358_93.n1 a_358_93.n0 261.704
R128 a_358_93.n0 a_358_93.t2 260.817
R129 a_358_93.n0 a_358_93.t3 167.63
R130 B.t1 B.t5 865.994
R131 B.n1 B.n0 298.841
R132 B.n0 B.t4 294.021
R133 B.n2 B.t1 235.109
R134 B.t5 B.n1 215.293
R135 B B.n2 194.166
R136 B.n0 B.t3 168.701
R137 B.n2 B.t2 167.63
R138 B.n1 B.t0 167.094
R139 a_1290_49.n2 a_1290_49.n1 590.155
R140 a_1290_49.t5 a_1290_49.n3 323.08
R141 a_1290_49.n3 a_1290_49.t4 318.813
R142 a_1290_49.n2 a_1290_49.n0 284.765
R143 a_1290_49.n1 a_1290_49.t3 209.827
R144 a_1290_49.n3 a_1290_49.n2 130.951
R145 a_1290_49.n0 a_1290_49.t2 94.7773
R146 a_1290_49.n1 a_1290_49.t0 41.5557
R147 a_1290_49.n0 a_1290_49.t1 38.438
R148 VPB.t11 VPB.t2 713.24
R149 VPB.t2 VPB.t1 648.131
R150 VPB.t9 VPB.t10 633.333
R151 VPB.t4 VPB.t3 517.913
R152 VPB.t1 VPB.t4 449.844
R153 VPB.t7 VPB.t9 355.14
R154 VPB VPB.t6 325.546
R155 VPB.t10 VPB.t11 313.707
R156 VPB.t3 VPB.t5 304.829
R157 VPB.t5 VPB.t0 298.911
R158 VPB.t0 VPB.t8 248.599
R159 VPB.t6 VPB.t7 248.599
R160 VPWR.n8 VPWR.t1 854.342
R161 VPWR.n21 VPWR.t2 839.034
R162 VPWR.n2 VPWR.n1 620.202
R163 VPWR.n7 VPWR.n6 605.511
R164 VPWR.n1 VPWR.t5 81.5708
R165 VPWR.n1 VPWR.t3 36.4455
R166 VPWR.n20 VPWR.n19 34.6358
R167 VPWR.n10 VPWR.n9 34.6358
R168 VPWR.n10 VPWR.n4 34.6358
R169 VPWR.n14 VPWR.n4 34.6358
R170 VPWR.n15 VPWR.n14 34.6358
R171 VPWR.n16 VPWR.n15 34.6358
R172 VPWR.n6 VPWR.t4 26.5955
R173 VPWR.n6 VPWR.t0 26.5955
R174 VPWR.n9 VPWR.n8 17.6946
R175 VPWR.n22 VPWR.n21 14.5711
R176 VPWR.n9 VPWR.n5 9.3005
R177 VPWR.n11 VPWR.n10 9.3005
R178 VPWR.n12 VPWR.n4 9.3005
R179 VPWR.n14 VPWR.n13 9.3005
R180 VPWR.n15 VPWR.n3 9.3005
R181 VPWR.n17 VPWR.n16 9.3005
R182 VPWR.n19 VPWR.n18 9.3005
R183 VPWR.n20 VPWR.n0 9.3005
R184 VPWR.n8 VPWR.n7 7.29413
R185 VPWR.n19 VPWR.n2 6.77697
R186 VPWR.n21 VPWR.n20 3.01226
R187 VPWR.n16 VPWR.n2 2.63579
R188 VPWR.n7 VPWR.n5 0.151957
R189 VPWR.n11 VPWR.n5 0.120292
R190 VPWR.n12 VPWR.n11 0.120292
R191 VPWR.n13 VPWR.n12 0.120292
R192 VPWR.n13 VPWR.n3 0.120292
R193 VPWR.n17 VPWR.n3 0.120292
R194 VPWR.n18 VPWR.n17 0.120292
R195 VPWR.n18 VPWR.n0 0.120292
R196 VPWR.n22 VPWR.n0 0.120292
R197 VPWR VPWR.n22 0.0226354
R198 A.n0 A.t1 239.505
R199 A.n0 A.t0 168.811
R200 A A.n0 163.52
C0 B VPWR 0.058841f
C1 VGND C 0.019768f
C2 VGND VPB 0.015331f
C3 C VPB 0.138744f
C4 A VGND 0.01316f
C5 VGND X 0.078805f
C6 A VPB 0.028102f
C7 X C 0.001816f
C8 X VPB 0.012482f
C9 B VGND 0.034605f
C10 VGND VPWR 0.101096f
C11 B C 5.03e-19
C12 B VPB 0.296899f
C13 VPWR C 0.021151f
C14 VPWR VPB 0.190599f
C15 B A 0.002172f
C16 A VPWR 0.014124f
C17 B X 7.16e-21
C18 VPWR X 0.108423f
C19 VGND VNB 1.0332f
C20 A VNB 0.092322f
C21 B VNB 0.423766f
C22 C VNB 0.261039f
C23 X VNB 0.06141f
C24 VPWR VNB 0.84504f
C25 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_4 VNB VPB X C B A
X0 a_602_325.t1 B.t0 a_1402_49.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.140825 pd=1.1 as=0.19265 ps=1.285 w=0.64 l=0.15
X1 a_1031_297.t0 B.t1 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.2526 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2 a_608_49.t2 B.t2 a_1402_49.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1458 pd=1.205 as=0.246 ps=1.525 w=0.64 l=0.15
X3 VGND.t7 A.t0 a_1135_365.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0992 pd=0.95 as=0.11 ps=0.99 w=0.64 l=0.15
X4 a_1402_49.t4 a_1031_297.t2 a_608_49.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.19265 pd=1.285 as=0.18365 ps=1.25 w=0.42 l=0.15
X5 a_480_297.t1 C.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2048 pd=1.92 as=0.1572 ps=1.345 w=0.64 l=0.15
X6 a_608_49.t0 a_480_297.t2 a_79_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.441 pd=2.73 as=0.1596 ps=1.22 w=0.84 l=0.15
X7 a_1135_365.t2 a_1031_297.t3 a_608_49.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1715 pd=1.355 as=0.1458 ps=1.205 w=0.84 l=0.15
X8 X.t7 a_79_21.t4 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_1135_365.t3 a_1031_297.t4 a_602_325.t4 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.11 pd=0.99 as=0.140825 ps=1.1 w=0.6 l=0.15
X10 VGND.t4 a_79_21.t5 X.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t5 a_79_21.t6 X.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.16525 pd=1.185 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_1031_297.t1 B.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1653 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_1402_49.t5 a_1031_297.t5 a_602_325.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.246 pd=1.525 as=0.2452 ps=1.45 w=0.64 l=0.15
X14 a_79_21.t3 C.t1 a_602_325.t2 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1596 pd=1.22 as=0.2184 ps=2.2 w=0.84 l=0.15
X15 a_480_297.t0 C.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.16525 ps=1.185 w=0.42 l=0.15
X16 a_608_49.t3 B.t4 a_1135_365.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.18365 pd=1.25 as=0.1628 ps=1.8 w=0.64 l=0.15
X17 VPWR.t4 A.t1 a_1135_365.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1715 ps=1.355 w=1 l=0.15
X18 a_1402_49.t3 a_1135_365.t6 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0992 ps=0.95 w=0.64 l=0.15
X19 X.t1 a_79_21.t7 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_602_325.t0 B.t5 a_1135_365.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2452 pd=1.45 as=0.3536 ps=2.53 w=0.84 l=0.15
X21 VPWR.t2 a_79_21.t8 X.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1572 pd=1.345 as=0.135 ps=1.27 w=1 l=0.15
X22 a_602_325.t3 a_480_297.t3 a_79_21.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.3168 pd=2.27 as=0.128 ps=1.04 w=0.64 l=0.15
X23 X.t5 a_79_21.t9 VPWR.t6 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_79_21.t2 C.t3 a_608_49.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.04 as=0.1728 ps=1.82 w=0.64 l=0.15
X25 VPWR.t7 a_79_21.t10 X.t4 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 X.t0 a_79_21.t11 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 a_1402_49.t2 a_1135_365.t7 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
R0 B.t2 B.t5 865.994
R1 B.n1 B.n0 298.841
R2 B.n0 B.t1 294.021
R3 B.n2 B.t2 235.109
R4 B.t5 B.n1 215.293
R5 B B.n2 194.166
R6 B.n0 B.t3 168.701
R7 B.n2 B.t0 167.63
R8 B.n1 B.t4 167.094
R9 a_1402_49.n2 a_1402_49.n1 590.155
R10 a_1402_49.t2 a_1402_49.n3 322.493
R11 a_1402_49.n3 a_1402_49.t3 320.478
R12 a_1402_49.n2 a_1402_49.n0 284.765
R13 a_1402_49.n1 a_1402_49.t5 209.827
R14 a_1402_49.n3 a_1402_49.n2 132.988
R15 a_1402_49.n0 a_1402_49.t4 94.7773
R16 a_1402_49.n1 a_1402_49.t1 41.5557
R17 a_1402_49.n0 a_1402_49.t0 38.438
R18 a_602_325.n1 a_602_325.t2 720.771
R19 a_602_325.n2 a_602_325.n0 342.616
R20 a_602_325.n1 a_602_325.t3 302.955
R21 a_602_325.n3 a_602_325.n2 297.875
R22 a_602_325.n3 a_602_325.t5 83.1099
R23 a_602_325.n0 a_602_325.t4 51.3868
R24 a_602_325.n4 a_602_325.t0 40.7642
R25 a_602_325.n5 a_602_325.n4 39.4005
R26 a_602_325.n4 a_602_325.n3 27.7036
R27 a_602_325.n0 a_602_325.t1 25.3226
R28 a_602_325.n2 a_602_325.n1 20.5528
R29 VNB.t9 VNB.t3 3730.74
R30 VNB.t0 VNB.t1 2762.46
R31 VNB.t3 VNB.t2 2648.54
R32 VNB.t12 VNB.t4 2264.08
R33 VNB.t2 VNB.t12 2164.4
R34 VNB.t11 VNB.t0 1950.81
R35 VNB.t4 VNB.t13 1708.74
R36 VNB.t1 VNB.t9 1566.34
R37 VNB.t13 VNB.t7 1423.95
R38 VNB.t7 VNB.t8 1310.03
R39 VNB.t5 VNB.t11 1196.12
R40 VNB.t10 VNB.t5 1196.12
R41 VNB.t6 VNB.t10 1196.12
R42 VNB VNB.t6 669.256
R43 VPWR.n7 VPWR.t0 848.898
R44 VPWR.n3 VPWR.n1 733.888
R45 VPWR VPWR.n2 605.532
R46 VPWR.n5 VPWR.n4 601.292
R47 VPWR.n1 VPWR.t3 66.1802
R48 VPWR VPWR.t1 859.981
R49 VPWR.n2 VPWR.t4 34.4755
R50 VPWR.n1 VPWR.t2 29.0556
R51 VPWR.n4 VPWR.t6 26.5955
R52 VPWR.n4 VPWR.t7 26.5955
R53 VPWR.n2 VPWR.t5 26.5955
R54 VPWR.n6 VPWR.n5 25.977
R55 VPWR.n7 VPWR.n6 24.8476
R56 VPWR.n3 VPWR 7.17429
R57 VPWR.n3 VPWR.n0 24.5847
R58 VPWR VPWR.n7 19.0887
R59 VPWR.n5 VPWR.n0 4.6318
R60 VPWR.n6 VPWR 9.3005
R61 VPWR.n0 VPWR 3.33203
R62 a_1031_297.t0 a_1031_297.n3 802.28
R63 a_1031_297.n0 a_1031_297.t3 283.257
R64 a_1031_297.n2 a_1031_297.n1 224.564
R65 a_1031_297.n3 a_1031_297.t1 219.297
R66 a_1031_297.n2 a_1031_297.n0 175.175
R67 a_1031_297.n1 a_1031_297.t2 173.52
R68 a_1031_297.n0 a_1031_297.t4 161.202
R69 a_1031_297.n1 a_1031_297.t5 154.24
R70 a_1031_297.n4 a_1031_297.t0 102.441
R71 a_1031_297.n3 a_1031_297.n2 10.4313
R72 VPB.t0 VPB.t4 713.24
R73 VPB.t4 VPB.t2 648.131
R74 VPB.t6 VPB.t11 603.739
R75 VPB.t7 VPB.t3 517.913
R76 VPB.t2 VPB.t7 449.844
R77 VPB.t11 VPB.t0 313.707
R78 VPB.t3 VPB.t8 304.829
R79 VPB.t8 VPB.t9 298.911
R80 VPB.t5 VPB.t6 292.991
R81 VPB.t9 VPB.t10 272.274
R82 VPB.t12 VPB.t5 248.599
R83 VPB.t13 VPB.t12 248.599
R84 VPB.t1 VPB.t13 248.599
R85 VPB VPB.t1 198.287
R86 a_608_49.n2 a_608_49.n1 782.395
R87 a_608_49.t0 a_608_49.n3 723.856
R88 a_608_49.n3 a_608_49.t1 640.187
R89 a_608_49.n2 a_608_49.n0 311.574
R90 a_608_49.n3 a_608_49.n2 117.46
R91 a_608_49.n0 a_608_49.t5 99.3755
R92 a_608_49.n1 a_608_49.t2 67.7193
R93 a_608_49.n1 a_608_49.t4 34.3691
R94 a_608_49.n0 a_608_49.t3 25.313
R95 A.n0 A.t1 239.505
R96 A.n0 A.t0 168.811
R97 A A.n0 163.52
R98 a_1135_365.n1 a_1135_365.t1 775.927
R99 a_1135_365.n6 a_1135_365.n5 641.726
R100 a_1135_365.n4 a_1135_365.t7 241.536
R101 a_1135_365.n1 a_1135_365.t0 222.323
R102 a_1135_365.n3 a_1135_365.n2 185
R103 a_1135_365.n4 a_1135_365.t6 170.843
R104 a_1135_365.n5 a_1135_365.n4 152
R105 a_1135_365.n5 a_1135_365.n3 56.4377
R106 a_1135_365.n0 a_1135_365.t2 50.4231
R107 a_1135_365.n2 a_1135_365.t3 43.0005
R108 a_1135_365.n7 a_1135_365.n6 38.6969
R109 a_1135_365.n0 a_1135_365.t4 28.8712
R110 a_1135_365.n3 a_1135_365.n1 26.8515
R111 a_1135_365.n2 a_1135_365.t5 23.0795
R112 a_1135_365.n6 a_1135_365.n0 17.5898
R113 VGND.n6 VGND.t3 290.289
R114 VGND.n2 VGND.t5 257.88
R115 VGND VGND.n3 220.472
R116 VGND.n4 VGND.n1 199.739
R117 VGND.t5 VGND.t0 51.4291
R118 VGND.n0 VGND 48.6521
R119 VGND.n2 VGND.n0 15.8399
R120 VGND.n3 VGND.t7 32.813
R121 VGND.n6 VGND.n5 32.377
R122 VGND.n4 VGND 5.42048
R123 VGND.n3 VGND.t6 25.313
R124 VGND.n1 VGND.t2 24.9236
R125 VGND.n1 VGND.t4 24.9236
R126 VGND VGND.n2 30.2675
R127 VGND.n5 VGND.n4 18.4476
R128 VGND VGND.t1 172.579
R129 VGND VGND.n6 11.5593
R130 VGND.n5 VGND 9.3005
R131 VGND VGND.n0 4.56757
R132 C.n0 C.t1 229.136
R133 C.n1 C.t0 167.386
R134 C.n0 C.t3 140.992
R135 C.n2 C.n1 104.641
R136 C.n1 C.t2 102.828
R137 C C.n2 68.4649
R138 C.n2 C.n0 27.396
R139 a_480_297.t1 a_480_297.n1 702.655
R140 a_480_297.n1 a_480_297.t0 281.925
R141 a_480_297.n0 a_480_297.t2 260.817
R142 a_480_297.n1 a_480_297.n0 259.733
R143 a_480_297.n0 a_480_297.t3 167.63
R144 a_79_21.n9 a_79_21.n8 773.587
R145 a_79_21.n8 a_79_21.n0 344.969
R146 a_79_21.n7 a_79_21.t8 212.081
R147 a_79_21.n5 a_79_21.t9 212.081
R148 a_79_21.n3 a_79_21.t10 212.081
R149 a_79_21.n1 a_79_21.t4 212.081
R150 a_79_21.n8 a_79_21.n7 162.956
R151 a_79_21.n1 a_79_21.t11 154.553
R152 a_79_21.n2 a_79_21.t5 139.78
R153 a_79_21.n4 a_79_21.t7 139.78
R154 a_79_21.n6 a_79_21.t6 139.78
R155 a_79_21.n0 a_79_21.t1 49.688
R156 a_79_21.t0 a_79_21.n9 46.9053
R157 a_79_21.n6 a_79_21.n5 46.7399
R158 a_79_21.n4 a_79_21.n3 46.7399
R159 a_79_21.n2 a_79_21.n1 46.7399
R160 a_79_21.n9 a_79_21.t3 42.2148
R161 a_79_21.n0 a_79_21.t2 25.313
R162 a_79_21.n7 a_79_21.n6 14.6066
R163 a_79_21.n5 a_79_21.n4 14.6066
R164 a_79_21.n3 a_79_21.n2 14.6066
R165 X.n2 X.n0 213.059
R166 X.n4 X.n3 205.662
R167 X.n2 X.n1 205.5
R168 X X.n5 205.233
R169 X.n5 X.t4 26.5955
R170 X.n5 X.t7 26.5955
R171 X.n3 X.t6 26.5955
R172 X.n3 X.t5 26.5955
R173 X.n4 X.n2 26.4132
R174 X.n1 X.t2 24.9236
R175 X.n1 X.t1 24.9236
R176 X.n0 X.t3 24.9236
R177 X.n0 X.t0 24.9236
R178 X X.n4 2.01042
C0 VPB VPWR 0.211838f
C1 C B 5.09e-19
C2 VGND A 0.012575f
C3 X B 1.01e-20
C4 VPB A 0.02873f
C5 VGND B 0.02969f
C6 X C 0.001873f
C7 VGND C 0.019689f
C8 VPWR A 0.014113f
C9 VPB B 0.297132f
C10 VPB C 0.136043f
C11 VGND X 0.147614f
C12 VPWR B 0.058394f
C13 C VPWR 0.022152f
C14 VPB X 0.010626f
C15 VGND VPB 0.019878f
C16 X VPWR 0.207144f
C17 VGND VPWR 0.124297f
C18 B A 0.002172f
C19 A VNB 0.092864f
C20 B VNB 0.423522f
C21 C VNB 0.255022f
C22 X VNB 0.064502f
C23 VPB VNB 2.0223f
C24 VGND VNB 1.1326f
C25 VPWR VNB 0.922638f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_4 VNB VPB VGND VPWR X B1 A4 A3 A2 A1
X0 a_467_47.t8 A4.t0 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_467_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t1 A1.t0 a_467_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.15275 ps=1.12 w=0.65 l=0.15
X3 a_467_47.t5 B1.t0 a_79_21.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_467_47.t3 A2.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.15275 pd=1.12 as=0.19825 ps=1.26 w=0.65 l=0.15
X5 a_79_21.t3 B1.t1 VPWR.t5 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t6 A1.t1 a_1083_297.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t0 a_79_21.t6 X.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1083_297.t1 A2.t1 a_889_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t8 A3.t1 a_467_47.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_79_21.t4 B1.t2 a_467_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 X.t6 a_79_21.t7 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_889_297.t2 A2.t2 a_1083_297.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X13 VPWR.t3 a_79_21.t8 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t4 a_79_21.t9 X.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t9 a_79_21.t10 X.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_639_297.t1 A3.t2 a_889_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t3 A2.t3 a_467_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.09425 ps=0.94 w=0.65 l=0.15
X18 a_889_297.t0 A3.t3 a_639_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X.t1 a_79_21.t11 VGND.t10 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_639_297.t3 A4.t1 a_79_21.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR.t4 B1.t3 a_79_21.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.145 ps=1.29 w=1 l=0.15
X22 VGND.t6 A4.t2 a_467_47.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X23 a_1083_297.t2 A1.t2 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.49 pd=2.98 as=0.135 ps=1.27 w=1 l=0.15
X24 a_79_21.t1 A4.t3 a_639_297.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 a_467_47.t6 A1.t3 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.3185 pd=2.28 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 X.t4 a_79_21.t12 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X.t0 a_79_21.t13 VGND.t11 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A4.n0 A4.t1 221.72
R1 A4.n1 A4.t3 221.72
R2 A4.n3 A4.n2 152
R3 A4.n0 A4.t0 149.421
R4 A4.n1 A4.t2 149.421
R5 A4.n2 A4.n0 37.4894
R6 A4.n2 A4.n1 37.4894
R7 A4 A4.n3 21.1205
R8 A4.n3 A4 8.3205
R9 VGND.n36 VGND.t11 286.786
R10 VGND.n8 VGND.n7 208.147
R11 VGND.n34 VGND.n1 207.213
R12 VGND.n22 VGND.n21 207.109
R13 VGND.n19 VGND.n18 203.016
R14 VGND.n12 VGND.n11 185
R15 VGND.n10 VGND.n9 185
R16 VGND.n29 VGND.t9 155.51
R17 VGND.n11 VGND.n10 62.7697
R18 VGND.n17 VGND.n6 34.6358
R19 VGND.n23 VGND.n20 34.6358
R20 VGND.n27 VGND.n4 34.6358
R21 VGND.n28 VGND.n27 34.6358
R22 VGND.n33 VGND.n2 34.6358
R23 VGND.n29 VGND.n28 32.0005
R24 VGND.n9 VGND.n8 31.3827
R25 VGND.n35 VGND.n34 30.8711
R26 VGND.n36 VGND.n35 25.977
R27 VGND.n10 VGND.t2 24.9236
R28 VGND.n11 VGND.t3 24.9236
R29 VGND.n7 VGND.t5 24.9236
R30 VGND.n7 VGND.t1 24.9236
R31 VGND.n18 VGND.t0 24.9236
R32 VGND.n18 VGND.t8 24.9236
R33 VGND.n21 VGND.t7 24.9236
R34 VGND.n21 VGND.t6 24.9236
R35 VGND.n1 VGND.t10 24.9236
R36 VGND.n1 VGND.t4 24.9236
R37 VGND.n29 VGND.n2 18.4476
R38 VGND.n22 VGND.n4 15.4358
R39 VGND.n37 VGND.n36 9.3005
R40 VGND.n35 VGND.n0 9.3005
R41 VGND.n33 VGND.n32 9.3005
R42 VGND.n31 VGND.n2 9.3005
R43 VGND.n14 VGND.n13 9.3005
R44 VGND.n15 VGND.n6 9.3005
R45 VGND.n17 VGND.n16 9.3005
R46 VGND.n20 VGND.n5 9.3005
R47 VGND.n24 VGND.n23 9.3005
R48 VGND.n25 VGND.n4 9.3005
R49 VGND.n27 VGND.n26 9.3005
R50 VGND.n28 VGND.n3 9.3005
R51 VGND.n30 VGND.n29 9.3005
R52 VGND.n19 VGND.n17 8.65932
R53 VGND.n13 VGND.n12 6.29891
R54 VGND.n20 VGND.n19 5.64756
R55 VGND.n12 VGND.n6 3.87277
R56 VGND.n34 VGND.n33 3.76521
R57 VGND.n23 VGND.n22 2.63579
R58 VGND.n14 VGND.n8 1.28449
R59 VGND.n13 VGND.n9 0.610024
R60 VGND.n15 VGND.n14 0.120292
R61 VGND.n16 VGND.n15 0.120292
R62 VGND.n16 VGND.n5 0.120292
R63 VGND.n24 VGND.n5 0.120292
R64 VGND.n25 VGND.n24 0.120292
R65 VGND.n26 VGND.n25 0.120292
R66 VGND.n26 VGND.n3 0.120292
R67 VGND.n30 VGND.n3 0.120292
R68 VGND.n31 VGND.n30 0.120292
R69 VGND.n32 VGND.n31 0.120292
R70 VGND.n32 VGND.n0 0.120292
R71 VGND.n37 VGND.n0 0.120292
R72 VGND VGND.n37 0.0213333
R73 a_467_47.n5 a_467_47.t1 324.652
R74 a_467_47.n2 a_467_47.t6 228.788
R75 a_467_47.n3 a_467_47.n2 99.7652
R76 a_467_47.n7 a_467_47.n6 98.0737
R77 a_467_47.n3 a_467_47.n0 98.0727
R78 a_467_47.n2 a_467_47.n1 98.0727
R79 a_467_47.n5 a_467_47.n4 88.3446
R80 a_467_47.n6 a_467_47.n5 64.2574
R81 a_467_47.n6 a_467_47.n3 63.2476
R82 a_467_47.n1 a_467_47.t3 48.0005
R83 a_467_47.n1 a_467_47.t2 38.7697
R84 a_467_47.n0 a_467_47.t4 28.6159
R85 a_467_47.n4 a_467_47.t5 28.6159
R86 a_467_47.n0 a_467_47.t0 24.9236
R87 a_467_47.n4 a_467_47.t7 24.9236
R88 a_467_47.n7 a_467_47.t9 24.9236
R89 a_467_47.t8 a_467_47.n7 24.9236
R90 VNB.t11 VNB.t1 2677.02
R91 VNB.t4 VNB.t3 2164.4
R92 VNB.t3 VNB.t2 1765.7
R93 VNB.t0 VNB.t4 1253.07
R94 VNB.t6 VNB.t8 1253.07
R95 VNB.t2 VNB.t7 1196.12
R96 VNB.t10 VNB.t0 1196.12
R97 VNB.t9 VNB.t10 1196.12
R98 VNB.t8 VNB.t9 1196.12
R99 VNB.t1 VNB.t6 1196.12
R100 VNB.t12 VNB.t11 1196.12
R101 VNB.t5 VNB.t12 1196.12
R102 VNB.t13 VNB.t5 1196.12
R103 VNB VNB.t13 911.327
R104 A3.n0 A3.t2 221.72
R105 A3.n1 A3.t3 221.72
R106 A3.n3 A3.n2 152
R107 A3.n0 A3.t0 149.421
R108 A3.n1 A3.t1 149.421
R109 A3.n2 A3.n0 37.4894
R110 A3.n2 A3.n1 37.4894
R111 A3 A3.n3 16.0005
R112 A3.n3 A3 13.4405
R113 A1.n1 A1.t2 221.72
R114 A1.n2 A1.t1 221.72
R115 A1.n1 A1.n0 202.879
R116 A1.n4 A1.n3 152
R117 A1.n1 A1.t3 149.421
R118 A1.n2 A1.t0 149.421
R119 A1.n3 A1.n2 40.1672
R120 A1.n3 A1.n1 34.8116
R121 A1.n4 A1 17.6005
R122 A1.n0 A1 15.0405
R123 A1.n0 A1 13.1205
R124 A1 A1.n4 11.8405
R125 B1.n0 B1.t1 300.269
R126 B1.n0 B1.t3 221.72
R127 B1.n2 B1.t0 165.488
R128 B1 B1.n2 156.481
R129 B1.n1 B1.t2 149.421
R130 B1.n2 B1.n1 58.9116
R131 B1.n1 B1.n0 14.282
R132 a_79_21.n11 a_79_21.n9 378.438
R133 a_79_21.n1 a_79_21.t6 221.72
R134 a_79_21.n6 a_79_21.t7 221.72
R135 a_79_21.n4 a_79_21.t8 221.72
R136 a_79_21.n2 a_79_21.t12 221.72
R137 a_79_21.n13 a_79_21.n12 215.143
R138 a_79_21.n11 a_79_21.n10 206.53
R139 a_79_21.n3 a_79_21.n0 176.436
R140 a_79_21.n5 a_79_21.n0 152
R141 a_79_21.n8 a_79_21.n7 152
R142 a_79_21.n1 a_79_21.t10 149.421
R143 a_79_21.n6 a_79_21.t11 149.421
R144 a_79_21.n4 a_79_21.t9 149.421
R145 a_79_21.n2 a_79_21.t13 149.421
R146 a_79_21.n12 a_79_21.n8 38.9823
R147 a_79_21.n7 a_79_21.n6 38.382
R148 a_79_21.n6 a_79_21.n5 37.4894
R149 a_79_21.n5 a_79_21.n4 37.4894
R150 a_79_21.n4 a_79_21.n3 37.4894
R151 a_79_21.n3 a_79_21.n2 37.4894
R152 a_79_21.n7 a_79_21.n1 36.5968
R153 a_79_21.n10 a_79_21.t3 30.5355
R154 a_79_21.n10 a_79_21.t2 26.5955
R155 a_79_21.n9 a_79_21.t0 26.5955
R156 a_79_21.n9 a_79_21.t1 26.5955
R157 a_79_21.t5 a_79_21.n13 24.9236
R158 a_79_21.n13 a_79_21.t4 24.9236
R159 a_79_21.n8 a_79_21.n0 24.7278
R160 a_79_21.n12 a_79_21.n11 12.6176
R161 A2.n2 A2.t1 229.754
R162 A2.n0 A2.t2 221.72
R163 A2.n6 A2.t3 164.595
R164 A2.n3 A2.n2 152
R165 A2.n5 A2.n4 152
R166 A2.n7 A2.n6 152
R167 A2.n1 A2.t0 149.421
R168 A2.n6 A2.n5 77.6561
R169 A2.n1 A2.n0 39.2746
R170 A2.n2 A2.n1 27.6709
R171 A2.n7 A2 26.5605
R172 A2.n4 A2.n3 25.2805
R173 A2.n5 A2.n0 3.57087
R174 A2.n3 A2 2.8805
R175 A2 A2.n7 2.8805
R176 A2.n4 A2 1.2805
R177 VPWR.n6 VPWR.t4 342.841
R178 VPWR.n17 VPWR.t1 341.928
R179 VPWR.n15 VPWR.n1 320.976
R180 VPWR.n5 VPWR.n4 318.738
R181 VPWR.n9 VPWR.n8 230.879
R182 VPWR.n10 VPWR.n7 34.6358
R183 VPWR.n14 VPWR.n2 34.6358
R184 VPWR.n16 VPWR.n15 30.8711
R185 VPWR.n1 VPWR.t2 26.5955
R186 VPWR.n1 VPWR.t3 26.5955
R187 VPWR.n8 VPWR.t5 26.5955
R188 VPWR.n8 VPWR.t0 26.5955
R189 VPWR.n4 VPWR.t7 26.5955
R190 VPWR.n4 VPWR.t6 26.5955
R191 VPWR.n17 VPWR.n16 25.977
R192 VPWR.n9 VPWR.n2 24.8476
R193 VPWR.n7 VPWR.n6 13.9299
R194 VPWR.n10 VPWR.n9 9.78874
R195 VPWR.n6 VPWR.n5 9.48347
R196 VPWR.n7 VPWR.n3 9.3005
R197 VPWR.n11 VPWR.n10 9.3005
R198 VPWR.n12 VPWR.n2 9.3005
R199 VPWR.n14 VPWR.n13 9.3005
R200 VPWR.n16 VPWR.n0 9.3005
R201 VPWR.n18 VPWR.n17 9.3005
R202 VPWR.n15 VPWR.n14 3.76521
R203 VPWR.n5 VPWR.n3 0.147194
R204 VPWR.n11 VPWR.n3 0.120292
R205 VPWR.n12 VPWR.n11 0.120292
R206 VPWR.n13 VPWR.n12 0.120292
R207 VPWR.n13 VPWR.n0 0.120292
R208 VPWR.n18 VPWR.n0 0.120292
R209 VPWR VPWR.n18 0.0213333
R210 VPB.t1 VPB.t6 580.062
R211 VPB.t10 VPB.t8 556.386
R212 VPB.t11 VPB.t10 260.437
R213 VPB.t13 VPB.t12 248.599
R214 VPB.t7 VPB.t13 248.599
R215 VPB.t6 VPB.t7 248.599
R216 VPB.t0 VPB.t1 248.599
R217 VPB.t9 VPB.t0 248.599
R218 VPB.t8 VPB.t9 248.599
R219 VPB.t5 VPB.t11 248.599
R220 VPB.t4 VPB.t5 248.599
R221 VPB.t3 VPB.t4 248.599
R222 VPB.t2 VPB.t3 248.599
R223 VPB VPB.t2 189.409
R224 a_1083_297.n1 a_1083_297.t0 384.327
R225 a_1083_297.t2 a_1083_297.n1 334.435
R226 a_1083_297.n1 a_1083_297.n0 208.511
R227 a_1083_297.n0 a_1083_297.t3 26.5955
R228 a_1083_297.n0 a_1083_297.t1 26.5955
R229 X.n5 X.n3 238.502
R230 X.n5 X.n4 205.863
R231 X.n2 X.n0 133.534
R232 X.n2 X.n1 99.1759
R233 X.n3 X.t7 26.5955
R234 X.n3 X.t6 26.5955
R235 X.n4 X.t5 26.5955
R236 X.n4 X.t4 26.5955
R237 X.n0 X.t2 24.9236
R238 X.n0 X.t1 24.9236
R239 X.n1 X.t3 24.9236
R240 X.n1 X.t0 24.9236
R241 X X.n5 16.7882
R242 X.n6 X 14.5236
R243 X.n6 X.n2 11.4531
R244 X X.n6 2.21588
R245 a_889_297.n1 a_889_297.n0 691.38
R246 a_889_297.n0 a_889_297.t1 26.5955
R247 a_889_297.n0 a_889_297.t0 26.5955
R248 a_889_297.n1 a_889_297.t3 26.5955
R249 a_889_297.t2 a_889_297.n1 26.5955
R250 a_639_297.n1 a_639_297.t2 385.779
R251 a_639_297.t1 a_639_297.n1 379.861
R252 a_639_297.n1 a_639_297.n0 189.28
R253 a_639_297.n0 a_639_297.t0 26.5955
R254 a_639_297.n0 a_639_297.t3 26.5955
C0 VPWR VPB 0.165561f
C1 VPB A3 0.057304f
C2 VPWR A3 0.014671f
C3 VGND A4 0.026584f
C4 VGND A1 0.037253f
C5 B1 A4 0.049737f
C6 VGND B1 0.020815f
C7 X VGND 0.28996f
C8 VGND A2 0.039639f
C9 A2 A1 0.060677f
C10 VPB A4 0.057014f
C11 VPWR A4 0.015655f
C12 VGND VPB 0.014305f
C13 X B1 1.55e-19
C14 VPWR VGND 0.15323f
C15 VPB A1 0.078233f
C16 A4 A3 0.06324f
C17 VPWR A1 0.042877f
C18 VGND A3 0.027804f
C19 VPB B1 0.080819f
C20 X VPB 0.012787f
C21 VPWR B1 0.030538f
C22 VPWR X 0.399995f
C23 VPB A2 0.088139f
C24 VPWR A2 0.017886f
C25 A3 A2 0.052155f
C26 VGND VNB 0.873567f
C27 X VNB 0.059924f
C28 VPWR VNB 0.742977f
C29 A1 VNB 0.245319f
C30 A2 VNB 0.237615f
C31 A3 VNB 0.171338f
C32 A4 VNB 0.171222f
C33 B1 VNB 0.223974f
C34 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_1 VNB VPB VGND VPWR A1 A2 A3 A4 Y B1
X0 a_348_297.t0 A3.t0 a_193_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3125 ps=1.625 w=1 l=0.15
X1 a_109_47.t2 A1.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.11375 ps=1 w=0.65 l=0.15
X2 a_193_297.t1 A4.t0 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t1 A1.t1 a_432_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.175 ps=1.35 w=1 l=0.15
X4 VGND.t3 A4.t1 a_109_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.203125 ps=1.275 w=0.65 l=0.15
X5 VGND.t0 A2.t0 a_109_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_47.t1 A3.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_432_297.t1 A2.t1 a_348_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47.t3 B1.t1 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A3.n0 A3.t0 241.536
R1 A3.n0 A3.t1 169.237
R2 A3.n1 A3.n0 152
R3 A3.n1 A3 11.4005
R4 A3 A3.n1 2.2005
R5 a_193_297.t0 a_193_297.t1 123.126
R6 a_348_297.t0 a_348_297.t1 53.1905
R7 VPB.t4 VPB.t1 458.724
R8 VPB.t3 VPB.t2 295.95
R9 VPB.t1 VPB.t3 248.599
R10 VPB.t0 VPB.t4 248.599
R11 VPB VPB.t0 189.409
R12 A1.n0 A1.t1 239.505
R13 A1.n0 A1.t0 167.204
R14 A1 A1.n0 164.544
R15 VGND.n2 VGND.n1 211.802
R16 VGND.n2 VGND.n0 211.542
R17 VGND.n1 VGND.t0 39.6928
R18 VGND.n1 VGND.t2 24.9236
R19 VGND.n0 VGND.t1 24.9236
R20 VGND.n0 VGND.t3 24.9236
R21 VGND VGND.n2 0.729154
R22 a_109_47.n1 a_109_47.t2 180.305
R23 a_109_47.n1 a_109_47.n0 145.388
R24 a_109_47.n2 a_109_47.n1 99.5638
R25 a_109_47.n0 a_109_47.t3 83.1525
R26 a_109_47.n0 a_109_47.t4 31.6937
R27 a_109_47.t0 a_109_47.n2 24.9236
R28 a_109_47.n2 a_109_47.t1 24.9236
R29 VNB.t3 VNB.t4 2207.12
R30 VNB.t0 VNB.t2 1423.95
R31 VNB.t1 VNB.t0 1196.12
R32 VNB.t4 VNB.t1 1196.12
R33 VNB VNB.t3 911.327
R34 A4.n0 A4.t0 269.027
R35 A4.n0 A4.t1 165.488
R36 A4.n1 A4.n0 152
R37 A4.n1 A4 11.9612
R38 A4 A4.n1 2.3087
R39 Y Y.n0 237.577
R40 Y.n1 Y.t1 129.381
R41 Y.n0 Y.t2 26.5955
R42 Y.n0 Y.t0 26.5955
R43 Y Y.n1 23.0214
R44 Y Y.n2 15.0593
R45 Y.n2 Y 10.5417
R46 Y.n2 Y 6.4005
R47 Y.n1 Y 5.55208
R48 a_432_297.t0 a_432_297.t1 68.9505
R49 VPWR.n0 VPWR.t0 256.62
R50 VPWR.n0 VPWR.t1 250.655
R51 VPWR VPWR.n0 0.0544237
R52 A2.n0 A2.t1 239.505
R53 A2.n0 A2.t0 167.204
R54 A2 A2.n0 163.02
R55 B1.n0 B1.t0 234.392
R56 B1.n0 B1.t1 162.091
R57 B1 B1.n0 160
C0 A4 VGND 0.018396f
C1 A3 Y 8.86e-19
C2 VPWR VGND 0.064559f
C3 A2 VPWR 0.090958f
C4 VPB A4 0.043344f
C5 VPWR VPB 0.089473f
C6 B1 VGND 0.013042f
C7 A4 Y 0.119702f
C8 VPWR Y 0.134142f
C9 A1 VGND 0.015418f
C10 A4 A3 0.148837f
C11 A2 A1 0.077463f
C12 VPWR A3 0.039458f
C13 VPB B1 0.037312f
C14 A1 VPB 0.036048f
C15 B1 Y 0.0837f
C16 A2 VGND 0.014196f
C17 A1 Y 2.46e-19
C18 VPWR A4 0.046241f
C19 VPB VGND 0.007325f
C20 A2 VPB 0.031734f
C21 Y VGND 0.060987f
C22 A2 Y 4.67e-19
C23 B1 A4 0.041875f
C24 A3 VGND 0.012777f
C25 A2 A3 0.162027f
C26 VPWR B1 0.045265f
C27 VPB Y 0.004443f
C28 A1 VPWR 0.054764f
C29 VPB A3 0.032059f
C30 VGND VNB 0.395518f
C31 Y VNB 0.050536f
C32 VPWR VNB 0.402763f
C33 A1 VNB 0.132284f
C34 A2 VNB 0.094882f
C35 A3 VNB 0.088406f
C36 A4 VNB 0.113993f
C37 B1 VNB 0.14431f
C38 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_2 VNB VPB VGND VPWR A1 A2 A3 A4 Y B1
X0 a_27_47.t5 A2.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t2 A4.t0 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t6 A3.t0 a_27_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t4 A2.t1 a_27_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4 VGND.t0 A1.t0 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47.t7 A3.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t3 B1.t0 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47.t8 B1.t1 Y.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_299_297.t1 A3.t2 a_549_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_549_297.t0 A3.t3 a_299_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_299_297.t3 A4.t1 Y.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y.t4 A4.t2 a_299_297.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_743_297.t3 A1.t1 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR.t1 A1.t2 a_743_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_743_297.t1 A2.t2 a_549_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47.t3 A4.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 Y.t2 B1.t2 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_27_47.t1 A1.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_549_297.t2 A2.t3 a_743_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 Y.t0 B1.t3 a_27_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n1 A2.t2 221.72
R1 A2.n3 A2.t3 221.72
R2 A2.n4 A2.n3 171.755
R3 A2.n2 A2.n0 152
R4 A2.n1 A2.t0 138.173
R5 A2.n3 A2.t1 138.173
R6 A2.n3 A2.n2 39.5087
R7 A2.n2 A2.n1 26.8661
R8 A2.n4 A2.n0 24.0005
R9 A2 A2.n4 4.8005
R10 A2.n0 A2 0.6405
R11 VGND.n16 VGND.t3 287.534
R12 VGND.n9 VGND.t6 282.841
R13 VGND.n6 VGND.n5 218.76
R14 VGND.n7 VGND.n4 207.213
R15 VGND.n14 VGND.n1 207.213
R16 VGND.n9 VGND.n8 34.6358
R17 VGND.n13 VGND.n2 34.6358
R18 VGND.n15 VGND.n14 29.3652
R19 VGND.n8 VGND.n7 27.8593
R20 VGND.n16 VGND.n15 27.4829
R21 VGND.n5 VGND.t1 24.9236
R22 VGND.n5 VGND.t0 24.9236
R23 VGND.n4 VGND.t5 24.9236
R24 VGND.n4 VGND.t4 24.9236
R25 VGND.n1 VGND.t7 24.9236
R26 VGND.n1 VGND.t2 24.9236
R27 VGND.n9 VGND.n2 16.9417
R28 VGND.n7 VGND.n6 13.7161
R29 VGND.n8 VGND.n3 9.3005
R30 VGND.n10 VGND.n9 9.3005
R31 VGND.n11 VGND.n2 9.3005
R32 VGND.n13 VGND.n12 9.3005
R33 VGND.n15 VGND.n0 9.3005
R34 VGND.n17 VGND.n16 7.10563
R35 VGND.n14 VGND.n13 5.27109
R36 VGND.n6 VGND.n3 0.80874
R37 VGND VGND.n17 0.348167
R38 VGND.n17 VGND.n0 0.154648
R39 VGND.n10 VGND.n3 0.120292
R40 VGND.n11 VGND.n10 0.120292
R41 VGND.n12 VGND.n11 0.120292
R42 VGND.n12 VGND.n0 0.120292
R43 a_27_47.n0 a_27_47.t9 187.311
R44 a_27_47.n6 a_27_47.t1 174.282
R45 a_27_47.n5 a_27_47.t4 135.882
R46 a_27_47.n0 a_27_47.t8 127.48
R47 a_27_47.n2 a_27_47.n1 99.5638
R48 a_27_47.n4 a_27_47.n3 99.5638
R49 a_27_47.n7 a_27_47.n6 99.5638
R50 a_27_47.n2 a_27_47.n0 59.3284
R51 a_27_47.n5 a_27_47.n4 48.9417
R52 a_27_47.n4 a_27_47.n2 38.4005
R53 a_27_47.n6 a_27_47.n5 38.4005
R54 a_27_47.n1 a_27_47.t2 24.9236
R55 a_27_47.n1 a_27_47.t3 24.9236
R56 a_27_47.n3 a_27_47.t6 24.9236
R57 a_27_47.n3 a_27_47.t7 24.9236
R58 a_27_47.n7 a_27_47.t0 24.9236
R59 a_27_47.t5 a_27_47.n7 24.9236
R60 VNB.t6 VNB.t4 2790.94
R61 VNB.t8 VNB.t3 2677.02
R62 VNB.t0 VNB.t1 1196.12
R63 VNB.t5 VNB.t0 1196.12
R64 VNB.t4 VNB.t5 1196.12
R65 VNB.t7 VNB.t6 1196.12
R66 VNB.t2 VNB.t7 1196.12
R67 VNB.t3 VNB.t2 1196.12
R68 VNB.t9 VNB.t8 1196.12
R69 VNB VNB.t9 911.327
R70 A4.n2 A4.t2 235.168
R71 A4.n0 A4.t1 218.507
R72 A4.n3 A4.t3 163.464
R73 A4 A4.n1 160.641
R74 A4.n4 A4.n3 152
R75 A4.n0 A4.t0 149.421
R76 A4.n2 A4.n1 41.3148
R77 A4 A4.n4 22.0805
R78 A4.n1 A4.n0 18.0755
R79 A4.n4 A4 7.3605
R80 A4.n3 A4.n2 0.595562
R81 A3.n2 A3.t2 216.9
R82 A3.n0 A3.t3 216.9
R83 A3.n3 A3.n2 166.46
R84 A3.n1 A3 162.881
R85 A3.n2 A3.t0 144.601
R86 A3.n0 A3.t1 144.601
R87 A3.n2 A3.n1 53.0205
R88 A3.n3 A3 16.0005
R89 A3.n1 A3.n0 14.4605
R90 A3 A3.n3 13.4405
R91 A1.n1 A1.t1 221.72
R92 A1.n2 A1.t2 221.72
R93 A1.n1 A1.n0 194.845
R94 A1.n4 A1.n3 152
R95 A1.n1 A1.t3 149.421
R96 A1.n2 A1.t0 149.421
R97 A1.n3 A1.n2 38.382
R98 A1.n3 A1.n1 36.5968
R99 A1 A1.n4 21.4405
R100 A1.n0 A1 20.4805
R101 A1.n0 A1 8.9605
R102 A1.n4 A1 8.0005
R103 B1.n0 B1.t0 216.9
R104 B1.n1 B1.t2 216.9
R105 B1 B1.n1 191.607
R106 B1.n0 B1.t1 141.387
R107 B1.n1 B1.t3 141.387
R108 B1.n1 B1.n0 65.3037
R109 Y.n2 Y.n0 359.76
R110 Y.n2 Y.n1 210.714
R111 Y Y.n3 186.745
R112 Y.n1 Y.t3 26.5955
R113 Y.n1 Y.t2 26.5955
R114 Y.n0 Y.t5 26.5955
R115 Y.n0 Y.t4 26.5955
R116 Y.n3 Y.t1 24.9236
R117 Y.n3 Y.t0 24.9236
R118 Y Y.n4 11.9835
R119 Y.n4 Y 6.53667
R120 Y Y.n2 5.99199
R121 Y.n4 Y 4.65505
R122 VPWR.n3 VPWR.t3 342.841
R123 VPWR.n2 VPWR.n1 316.94
R124 VPWR.n5 VPWR.t2 249.362
R125 VPWR.n1 VPWR.t0 26.5955
R126 VPWR.n1 VPWR.t1 26.5955
R127 VPWR.n5 VPWR.n4 25.977
R128 VPWR.n4 VPWR.n3 24.4711
R129 VPWR.n4 VPWR.n0 9.3005
R130 VPWR.n6 VPWR.n5 9.3005
R131 VPWR.n3 VPWR.n2 7.259
R132 VPWR.n2 VPWR.n0 0.152503
R133 VPWR.n6 VPWR.n0 0.120292
R134 VPWR VPWR.n6 0.0213333
R135 VPB.t1 VPB.t2 580.062
R136 VPB.t7 VPB.t8 556.386
R137 VPB.t4 VPB.t5 248.599
R138 VPB.t3 VPB.t4 248.599
R139 VPB.t2 VPB.t3 248.599
R140 VPB.t0 VPB.t1 248.599
R141 VPB.t9 VPB.t0 248.599
R142 VPB.t8 VPB.t9 248.599
R143 VPB.t6 VPB.t7 248.599
R144 VPB VPB.t6 189.409
R145 a_549_297.n1 a_549_297.n0 675.189
R146 a_549_297.n0 a_549_297.t3 26.5955
R147 a_549_297.n0 a_549_297.t2 26.5955
R148 a_549_297.n1 a_549_297.t1 26.5955
R149 a_549_297.t0 a_549_297.n1 26.5955
R150 a_299_297.t1 a_299_297.n1 409.63
R151 a_299_297.n1 a_299_297.t2 406.575
R152 a_299_297.n1 a_299_297.n0 184.215
R153 a_299_297.n0 a_299_297.t0 26.5955
R154 a_299_297.n0 a_299_297.t3 26.5955
R155 a_743_297.n0 a_743_297.t0 384.327
R156 a_743_297.n0 a_743_297.t3 291.95
R157 a_743_297.n1 a_743_297.n0 208.511
R158 a_743_297.n1 a_743_297.t2 26.5955
R159 a_743_297.t1 a_743_297.n1 26.5955
C0 Y VGND 0.01201f
C1 A3 Y 5.75e-19
C2 A2 VPWR 0.021194f
C3 A4 Y 0.093785f
C4 B1 VGND 0.019659f
C5 VPB A2 0.067179f
C6 B1 A4 0.02088f
C7 A2 A1 0.06778f
C8 VPWR VGND 0.115735f
C9 A3 VPWR 0.020037f
C10 B1 Y 0.085823f
C11 VPB VGND 0.013233f
C12 A4 VPWR 0.018469f
C13 VPB A3 0.068016f
C14 VPB A4 0.069214f
C15 A1 VGND 0.031061f
C16 VPWR Y 0.227127f
C17 VPB Y 0.019354f
C18 B1 VPWR 0.058575f
C19 VPB B1 0.074492f
C20 A1 Y 1.33e-19
C21 A2 VGND 0.030035f
C22 A3 A2 0.037826f
C23 VPB VPWR 0.13675f
C24 A2 Y 2.32e-19
C25 A1 VPWR 0.041847f
C26 A3 VGND 0.02972f
C27 A4 VGND 0.031374f
C28 VPB A1 0.076236f
C29 A4 A3 0.063402f
C30 VGND VNB 0.681581f
C31 Y VNB 0.025872f
C32 VPWR VNB 0.59717f
C33 A1 VNB 0.240755f
C34 A2 VNB 0.197857f
C35 A3 VNB 0.197189f
C36 A4 VNB 0.203934f
C37 B1 VNB 0.239292f
C38 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_4 VNB VPB VGND VPWR B1 Y A4 A1 A2 A3
X0 VGND.t11 A2.t0 a_27_47.t13 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_467_297.t7 A4.t0 Y.t10 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t10 A2.t1 a_27_47.t12 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t4 A1.t0 a_1243_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t7 A1.t1 a_27_47.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47.t3 A4.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t9 A4.t2 a_467_297.t6 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47.t0 A4.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t7 B1.t0 Y.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47.t11 A2.t2 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47.t14 A2.t3 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t1 A4.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_27_47.t7 A1.t2 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t12 A3.t0 a_27_47.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t0 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1243_297.t2 A1.t3 VPWR.t3 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47.t17 A1.t4 VGND.t13 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t2 A4.t5 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t15 A3.t1 a_27_47.t19 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR.t5 B1.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t2 A1.t5 a_1243_297.t1 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_27_47.t4 B1.t3 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_27_47.t5 B1.t4 Y.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_467_297.t5 A4.t6 Y.t8 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1243_297.t5 A2.t4 a_885_297.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t11 A4.t7 a_467_297.t4 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_27_47.t8 A3.t2 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VGND.t14 A1.t6 a_27_47.t18 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_885_297.t2 A2.t5 a_1243_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_27_47.t9 A3.t3 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 Y.t4 B1.t5 a_27_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_1243_297.t7 A2.t6 a_885_297.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_467_297.t0 A3.t4 a_885_297.t7 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 a_885_297.t0 A2.t7 a_1243_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_885_297.t6 A3.t5 a_467_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_467_297.t2 A3.t6 a_885_297.t5 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y.t5 B1.t6 VPWR.t6 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X37 a_1243_297.t0 A1.t7 VPWR.t1 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X38 a_885_297.t4 A3.t7 a_467_297.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 Y.t7 B1.t7 a_27_47.t16 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n6 A2.t6 221.72
R1 A2.n1 A2.t4 221.72
R2 A2.n2 A2.t5 221.72
R3 A2.n7 A2.t7 221.72
R4 A2 A2.n3 166.4
R5 A2.n8 A2.n7 155.571
R6 A2.n4 A2.n0 152
R7 A2.n6 A2.n5 152
R8 A2.n6 A2.t2 149.421
R9 A2.n1 A2.t3 149.421
R10 A2.n2 A2.t1 149.421
R11 A2.n7 A2.t0 149.421
R12 A2.n7 A2.n6 74.9783
R13 A2.n6 A2.n0 71.4079
R14 A2.n3 A2.n2 68.7301
R15 A2 A2.n8 23.0405
R16 A2.n5 A2 21.7605
R17 A2 A2.n4 17.9205
R18 A2.n4 A2 11.5205
R19 A2.n5 A2 7.6805
R20 A2.n8 A2 6.4005
R21 A2.n3 A2.n1 6.24865
R22 A2.n2 A2.n0 3.57087
R23 a_27_47.n2 a_27_47.t5 268.077
R24 a_27_47.n1 a_27_47.n0 185
R25 a_27_47.n1 a_27_47.t16 182.894
R26 a_27_47.n7 a_27_47.t17 174.282
R27 a_27_47.n12 a_27_47.t13 138.675
R28 a_27_47.n13 a_27_47.t8 138.675
R29 a_27_47.n3 a_27_47.t1 127.852
R30 a_27_47.n7 a_27_47.n6 99.5638
R31 a_27_47.n9 a_27_47.n8 99.5638
R32 a_27_47.n11 a_27_47.n10 99.5638
R33 a_27_47.n15 a_27_47.n14 99.5638
R34 a_27_47.n5 a_27_47.n4 99.5638
R35 a_27_47.n17 a_27_47.n16 99.5638
R36 a_27_47.n2 a_27_47.n1 51.2005
R37 a_27_47.n5 a_27_47.n3 50.603
R38 a_27_47.n9 a_27_47.n7 38.4005
R39 a_27_47.n11 a_27_47.n9 38.4005
R40 a_27_47.n12 a_27_47.n11 38.4005
R41 a_27_47.n15 a_27_47.n13 38.4005
R42 a_27_47.n16 a_27_47.n5 38.4005
R43 a_27_47.n16 a_27_47.n15 38.4005
R44 a_27_47.n3 a_27_47.n2 33.739
R45 a_27_47.n6 a_27_47.t18 24.9236
R46 a_27_47.n6 a_27_47.t7 24.9236
R47 a_27_47.n8 a_27_47.t10 24.9236
R48 a_27_47.n8 a_27_47.t14 24.9236
R49 a_27_47.n10 a_27_47.t12 24.9236
R50 a_27_47.n10 a_27_47.t11 24.9236
R51 a_27_47.n14 a_27_47.t15 24.9236
R52 a_27_47.n14 a_27_47.t9 24.9236
R53 a_27_47.n0 a_27_47.t6 24.9236
R54 a_27_47.n0 a_27_47.t4 24.9236
R55 a_27_47.n4 a_27_47.t2 24.9236
R56 a_27_47.n4 a_27_47.t3 24.9236
R57 a_27_47.n17 a_27_47.t19 24.9236
R58 a_27_47.t0 a_27_47.n17 24.9236
R59 a_27_47.n13 a_27_47.n12 14.3064
R60 VGND.n13 VGND.n12 218.496
R61 VGND.n15 VGND.n14 207.213
R62 VGND.n11 VGND.n10 207.213
R63 VGND.n21 VGND.n9 207.213
R64 VGND.n27 VGND.n6 207.213
R65 VGND.n30 VGND.n29 207.213
R66 VGND.n36 VGND.n3 207.213
R67 VGND.n1 VGND.n0 207.213
R68 VGND.n20 VGND.n19 34.6358
R69 VGND.n22 VGND.n7 34.6358
R70 VGND.n26 VGND.n7 34.6358
R71 VGND.n31 VGND.n28 34.6358
R72 VGND.n35 VGND.n4 34.6358
R73 VGND.n38 VGND.n37 34.6358
R74 VGND.n40 VGND.n1 33.9541
R75 VGND.n16 VGND.n11 33.8829
R76 VGND.n16 VGND.n15 29.3652
R77 VGND.n21 VGND.n20 27.8593
R78 VGND.n27 VGND.n26 26.3534
R79 VGND.n12 VGND.t13 24.9236
R80 VGND.n12 VGND.t14 24.9236
R81 VGND.n14 VGND.t4 24.9236
R82 VGND.n14 VGND.t7 24.9236
R83 VGND.n10 VGND.t8 24.9236
R84 VGND.n10 VGND.t10 24.9236
R85 VGND.n9 VGND.t9 24.9236
R86 VGND.n9 VGND.t11 24.9236
R87 VGND.n6 VGND.t5 24.9236
R88 VGND.n6 VGND.t12 24.9236
R89 VGND.n29 VGND.t6 24.9236
R90 VGND.n29 VGND.t15 24.9236
R91 VGND.n3 VGND.t0 24.9236
R92 VGND.n3 VGND.t2 24.9236
R93 VGND.n0 VGND.t3 24.9236
R94 VGND.n0 VGND.t1 24.9236
R95 VGND.n31 VGND.n30 20.3299
R96 VGND.n37 VGND.n36 20.3299
R97 VGND.n30 VGND.n4 14.3064
R98 VGND.n36 VGND.n35 14.3064
R99 VGND.n15 VGND.n13 12.2589
R100 VGND.n17 VGND.n16 9.3005
R101 VGND.n19 VGND.n18 9.3005
R102 VGND.n20 VGND.n8 9.3005
R103 VGND.n23 VGND.n22 9.3005
R104 VGND.n24 VGND.n7 9.3005
R105 VGND.n26 VGND.n25 9.3005
R106 VGND.n28 VGND.n5 9.3005
R107 VGND.n32 VGND.n31 9.3005
R108 VGND.n33 VGND.n4 9.3005
R109 VGND.n35 VGND.n34 9.3005
R110 VGND.n37 VGND.n2 9.3005
R111 VGND.n39 VGND.n38 9.3005
R112 VGND.n28 VGND.n27 8.28285
R113 VGND.n38 VGND.n1 8.28285
R114 VGND.n22 VGND.n21 6.77697
R115 VGND.n17 VGND.n13 0.76003
R116 VGND.n19 VGND.n11 0.753441
R117 VGND VGND.n40 0.596506
R118 VGND.n40 VGND.n39 0.147181
R119 VGND.n18 VGND.n17 0.120292
R120 VGND.n18 VGND.n8 0.120292
R121 VGND.n23 VGND.n8 0.120292
R122 VGND.n24 VGND.n23 0.120292
R123 VGND.n25 VGND.n24 0.120292
R124 VGND.n25 VGND.n5 0.120292
R125 VGND.n32 VGND.n5 0.120292
R126 VGND.n33 VGND.n32 0.120292
R127 VGND.n34 VGND.n33 0.120292
R128 VGND.n34 VGND.n2 0.120292
R129 VGND.n39 VGND.n2 0.120292
R130 VNB.t8 VNB.t14 2677.02
R131 VNB.t5 VNB.t1 2677.02
R132 VNB.t18 VNB.t17 1196.12
R133 VNB.t7 VNB.t18 1196.12
R134 VNB.t10 VNB.t7 1196.12
R135 VNB.t11 VNB.t10 1196.12
R136 VNB.t13 VNB.t11 1196.12
R137 VNB.t12 VNB.t13 1196.12
R138 VNB.t14 VNB.t12 1196.12
R139 VNB.t15 VNB.t8 1196.12
R140 VNB.t9 VNB.t15 1196.12
R141 VNB.t19 VNB.t9 1196.12
R142 VNB.t0 VNB.t19 1196.12
R143 VNB.t2 VNB.t0 1196.12
R144 VNB.t3 VNB.t2 1196.12
R145 VNB.t1 VNB.t3 1196.12
R146 VNB.t6 VNB.t5 1196.12
R147 VNB.t4 VNB.t6 1196.12
R148 VNB.t16 VNB.t4 1196.12
R149 VNB VNB.t16 911.327
R150 A4.n9 A4.t7 232.214
R151 A4.n2 A4.t0 221.72
R152 A4.n1 A4.t2 221.72
R153 A4.n7 A4.t6 221.72
R154 A4.n9 A4.t4 159.915
R155 A4.n4 A4.n3 152
R156 A4.n6 A4.n5 152
R157 A4.n8 A4.n0 152
R158 A4.n10 A4.n9 152
R159 A4.n2 A4.t3 149.421
R160 A4.n1 A4.t5 149.421
R161 A4.n7 A4.t1 149.421
R162 A4.n3 A4.n2 37.4894
R163 A4.n3 A4.n1 37.4894
R164 A4.n6 A4.n1 37.4894
R165 A4.n7 A4.n6 37.4894
R166 A4.n8 A4.n7 36.5968
R167 A4.n9 A4.n8 24.9931
R168 A4.n5 A4 23.6805
R169 A4.n10 A4.n0 23.6805
R170 A4 A4.n4 21.1205
R171 A4.n4 A4 8.3205
R172 A4.n5 A4 5.7605
R173 A4 A4.n0 2.8805
R174 A4 A4.n10 2.8805
R175 Y.n6 Y.n4 339.204
R176 Y.n6 Y.n5 300.803
R177 Y.n10 Y.n8 224.822
R178 Y.n1 Y.n0 207.22
R179 Y.n3 Y.n2 207.22
R180 Y.n10 Y.n9 185
R181 Y.n7 Y.n6 41.7887
R182 Y.n4 Y.t10 26.5955
R183 Y.n4 Y.t9 26.5955
R184 Y.n5 Y.t8 26.5955
R185 Y.n5 Y.t11 26.5955
R186 Y.n0 Y.t1 26.5955
R187 Y.n0 Y.t5 26.5955
R188 Y.n2 Y.t6 26.5955
R189 Y.n2 Y.t0 26.5955
R190 Y.n8 Y.t2 24.9236
R191 Y.n8 Y.t7 24.9236
R192 Y.n9 Y.t3 24.9236
R193 Y.n9 Y.t4 24.9236
R194 Y.n3 Y 21.4593
R195 Y Y.n1 16.9417
R196 Y.n11 Y.n10 16.5931
R197 Y Y.n11 14.7867
R198 Y.n7 Y.n3 13.9299
R199 Y.n3 Y 11.6711
R200 Y Y.n7 3.75222
R201 Y.n1 Y 3.29747
R202 Y.n3 Y 3.29747
R203 Y.n11 Y 0.22119
R204 a_467_297.n4 a_467_297.t4 384.839
R205 a_467_297.n1 a_467_297.t0 365.798
R206 a_467_297.n1 a_467_297.n0 300.803
R207 a_467_297.n5 a_467_297.n4 299.14
R208 a_467_297.n3 a_467_297.n2 184.215
R209 a_467_297.n4 a_467_297.n3 88.0383
R210 a_467_297.n3 a_467_297.n1 75.1194
R211 a_467_297.n2 a_467_297.t3 26.5955
R212 a_467_297.n2 a_467_297.t7 26.5955
R213 a_467_297.n0 a_467_297.t1 26.5955
R214 a_467_297.n0 a_467_297.t2 26.5955
R215 a_467_297.t6 a_467_297.n5 26.5955
R216 a_467_297.n5 a_467_297.t5 26.5955
R217 VPB.t3 VPB.t6 556.386
R218 VPB.t10 VPB.t13 556.386
R219 VPB.t5 VPB.t19 248.599
R220 VPB.t17 VPB.t5 248.599
R221 VPB.t18 VPB.t17 248.599
R222 VPB.t9 VPB.t18 248.599
R223 VPB.t8 VPB.t9 248.599
R224 VPB.t7 VPB.t8 248.599
R225 VPB.t6 VPB.t7 248.599
R226 VPB.t4 VPB.t3 248.599
R227 VPB.t11 VPB.t4 248.599
R228 VPB.t12 VPB.t11 248.599
R229 VPB.t16 VPB.t12 248.599
R230 VPB.t15 VPB.t16 248.599
R231 VPB.t14 VPB.t15 248.599
R232 VPB.t13 VPB.t14 248.599
R233 VPB.t0 VPB.t10 248.599
R234 VPB.t1 VPB.t0 248.599
R235 VPB.t2 VPB.t1 248.599
R236 VPB VPB.t2 189.409
R237 A1.n1 A1.t7 221.72
R238 A1.n5 A1.t0 221.72
R239 A1.n7 A1.t3 221.72
R240 A1.n8 A1.t5 221.72
R241 A1 A1.n9 161.601
R242 A1.n2 A1.n1 160.034
R243 A1.n4 A1.n3 152
R244 A1.n6 A1.n0 152
R245 A1.n1 A1.t4 149.421
R246 A1.n5 A1.t6 149.421
R247 A1.n7 A1.t2 149.421
R248 A1.n8 A1.t1 149.421
R249 A1.n4 A1.n1 70.5153
R250 A1.n6 A1.n5 63.3746
R251 A1.n9 A1.n7 58.9116
R252 A1.n2 A1 20.1605
R253 A1.n3 A1 18.8805
R254 A1.n9 A1.n8 16.0672
R255 A1 A1.n0 15.6805
R256 A1 A1.n0 13.7605
R257 A1.n7 A1.n6 11.6042
R258 A1.n3 A1 10.5605
R259 A1 A1.n2 9.2805
R260 A1.n5 A1.n4 4.46346
R261 a_1243_297.n1 a_1243_297.t6 365.8
R262 a_1243_297.n1 a_1243_297.n0 300.803
R263 a_1243_297.t0 a_1243_297.n5 272.214
R264 a_1243_297.n3 a_1243_297.n2 207.22
R265 a_1243_297.n5 a_1243_297.n4 207.22
R266 a_1243_297.n3 a_1243_297.n1 38.4005
R267 a_1243_297.n5 a_1243_297.n3 38.4005
R268 a_1243_297.n0 a_1243_297.t4 26.5955
R269 a_1243_297.n0 a_1243_297.t7 26.5955
R270 a_1243_297.n2 a_1243_297.t1 26.5955
R271 a_1243_297.n2 a_1243_297.t5 26.5955
R272 a_1243_297.n4 a_1243_297.t3 26.5955
R273 a_1243_297.n4 a_1243_297.t2 26.5955
R274 VPWR.n33 VPWR.t7 342.841
R275 VPWR.n12 VPWR.n11 332.26
R276 VPWR.n38 VPWR.n1 320.976
R277 VPWR.n13 VPWR.n10 320.976
R278 VPWR.n40 VPWR.t6 249.362
R279 VPWR.n37 VPWR.n2 34.6358
R280 VPWR.n15 VPWR.n14 34.6358
R281 VPWR.n15 VPWR.n8 34.6358
R282 VPWR.n19 VPWR.n8 34.6358
R283 VPWR.n20 VPWR.n19 34.6358
R284 VPWR.n21 VPWR.n20 34.6358
R285 VPWR.n21 VPWR.n6 34.6358
R286 VPWR.n25 VPWR.n6 34.6358
R287 VPWR.n26 VPWR.n25 34.6358
R288 VPWR.n27 VPWR.n26 34.6358
R289 VPWR.n27 VPWR.n4 34.6358
R290 VPWR.n31 VPWR.n4 34.6358
R291 VPWR.n32 VPWR.n31 34.6358
R292 VPWR.n33 VPWR.n32 32.0005
R293 VPWR.n39 VPWR.n38 30.8711
R294 VPWR.n14 VPWR.n13 29.3652
R295 VPWR.n1 VPWR.t0 26.5955
R296 VPWR.n1 VPWR.t5 26.5955
R297 VPWR.n10 VPWR.t3 26.5955
R298 VPWR.n10 VPWR.t2 26.5955
R299 VPWR.n11 VPWR.t1 26.5955
R300 VPWR.n11 VPWR.t4 26.5955
R301 VPWR.n40 VPWR.n39 25.977
R302 VPWR.n33 VPWR.n2 18.4476
R303 VPWR.n13 VPWR.n12 12.2589
R304 VPWR.n14 VPWR.n9 9.3005
R305 VPWR.n16 VPWR.n15 9.3005
R306 VPWR.n17 VPWR.n8 9.3005
R307 VPWR.n19 VPWR.n18 9.3005
R308 VPWR.n20 VPWR.n7 9.3005
R309 VPWR.n22 VPWR.n21 9.3005
R310 VPWR.n23 VPWR.n6 9.3005
R311 VPWR.n25 VPWR.n24 9.3005
R312 VPWR.n26 VPWR.n5 9.3005
R313 VPWR.n28 VPWR.n27 9.3005
R314 VPWR.n29 VPWR.n4 9.3005
R315 VPWR.n31 VPWR.n30 9.3005
R316 VPWR.n32 VPWR.n3 9.3005
R317 VPWR.n34 VPWR.n33 9.3005
R318 VPWR.n35 VPWR.n2 9.3005
R319 VPWR.n37 VPWR.n36 9.3005
R320 VPWR.n39 VPWR.n0 9.3005
R321 VPWR.n41 VPWR.n40 9.3005
R322 VPWR.n38 VPWR.n37 3.76521
R323 VPWR.n12 VPWR.n9 0.76003
R324 VPWR.n16 VPWR.n9 0.120292
R325 VPWR.n17 VPWR.n16 0.120292
R326 VPWR.n18 VPWR.n17 0.120292
R327 VPWR.n18 VPWR.n7 0.120292
R328 VPWR.n22 VPWR.n7 0.120292
R329 VPWR.n23 VPWR.n22 0.120292
R330 VPWR.n24 VPWR.n23 0.120292
R331 VPWR.n24 VPWR.n5 0.120292
R332 VPWR.n28 VPWR.n5 0.120292
R333 VPWR.n29 VPWR.n28 0.120292
R334 VPWR.n30 VPWR.n29 0.120292
R335 VPWR.n30 VPWR.n3 0.120292
R336 VPWR.n34 VPWR.n3 0.120292
R337 VPWR.n35 VPWR.n34 0.120292
R338 VPWR.n36 VPWR.n35 0.120292
R339 VPWR.n36 VPWR.n0 0.120292
R340 VPWR.n41 VPWR.n0 0.120292
R341 VPWR VPWR.n41 0.0213333
R342 B1.n9 B1.t6 234.392
R343 B1.n2 B1.t0 221.72
R344 B1.n4 B1.t1 221.72
R345 B1.n0 B1.t2 221.72
R346 B1.n9 B1.t7 162.091
R347 B1.n3 B1.n1 152
R348 B1.n6 B1.n5 152
R349 B1.n8 B1.n7 152
R350 B1.n10 B1.n9 152
R351 B1.n2 B1.t4 149.421
R352 B1.n4 B1.t5 149.421
R353 B1.n0 B1.t3 149.421
R354 B1.n3 B1.n2 37.4894
R355 B1.n4 B1.n3 37.4894
R356 B1.n5 B1.n4 37.4894
R357 B1.n5 B1.n0 37.4894
R358 B1.n8 B1.n0 37.4894
R359 B1.n6 B1.n1 26.8805
R360 B1.n7 B1 24.9605
R361 B1.n9 B1.n8 24.1005
R362 B1.n10 B1 21.4405
R363 B1 B1.n10 8.0005
R364 B1.n7 B1 4.4805
R365 B1 B1.n6 1.9205
R366 B1.n1 B1 0.6405
R367 A3.n1 A3.t4 221.72
R368 A3.n0 A3.t5 221.72
R369 A3.n6 A3.t6 221.72
R370 A3.n7 A3.t7 221.72
R371 A3.n1 A3 196.596
R372 A3.n3 A3.n2 152
R373 A3.n5 A3.n4 152
R374 A3.n9 A3.n8 152
R375 A3.n1 A3.t2 149.421
R376 A3.n0 A3.t0 149.421
R377 A3.n6 A3.t3 149.421
R378 A3.n7 A3.t1 149.421
R379 A3.n5 A3.n0 38.382
R380 A3.n2 A3.n1 37.4894
R381 A3.n2 A3.n0 37.4894
R382 A3.n8 A3.n6 37.4894
R383 A3.n8 A3.n7 37.4894
R384 A3.n6 A3.n5 36.5968
R385 A3.n3 A3 18.5605
R386 A3.n4 A3 16.3205
R387 A3 A3.n9 16.0005
R388 A3.n9 A3 13.4405
R389 A3.n4 A3 13.1205
R390 A3 A3.n3 10.8805
R391 a_885_297.n5 a_885_297.n4 362.389
R392 a_885_297.n3 a_885_297.n2 358.243
R393 a_885_297.n3 a_885_297.n1 299.14
R394 a_885_297.n4 a_885_297.n0 299.14
R395 a_885_297.n4 a_885_297.n3 102.4
R396 a_885_297.n2 a_885_297.t5 26.5955
R397 a_885_297.n2 a_885_297.t4 26.5955
R398 a_885_297.n1 a_885_297.t7 26.5955
R399 a_885_297.n1 a_885_297.t6 26.5955
R400 a_885_297.n0 a_885_297.t1 26.5955
R401 a_885_297.n0 a_885_297.t0 26.5955
R402 a_885_297.t3 a_885_297.n5 26.5955
R403 a_885_297.n5 a_885_297.t2 26.5955
C0 A3 VPB 0.136268f
C1 VPB A2 0.129161f
C2 A4 A3 0.06324f
C3 A1 VPWR 0.063311f
C4 VGND VPB 0.016353f
C5 A4 VGND 0.053242f
C6 A3 Y 6.25e-19
C7 Y A2 1.93e-19
C8 A4 VPB 0.132843f
C9 A3 VPWR 0.031933f
C10 A2 VPWR 0.037819f
C11 Y VGND 0.03121f
C12 Y VPB 0.025274f
C13 A4 Y 0.211015f
C14 B1 VGND 0.036195f
C15 VGND VPWR 0.194389f
C16 B1 VPB 0.138748f
C17 B1 A4 0.020422f
C18 VPB VPWR 0.203352f
C19 A4 VPWR 0.03246f
C20 A2 A1 0.069422f
C21 B1 Y 0.336515f
C22 VGND A1 0.060492f
C23 Y VPWR 0.418158f
C24 VPB A1 0.130687f
C25 B1 VPWR 0.096065f
C26 A3 A2 0.041097f
C27 A3 VGND 0.053712f
C28 Y A1 1.05e-19
C29 VGND A2 0.059778f
C30 VGND VNB 1.08979f
C31 Y VNB 0.027565f
C32 VPWR VNB 0.946477f
C33 A1 VNB 0.40703f
C34 A2 VNB 0.37861f
C35 A3 VNB 0.392114f
C36 A4 VNB 0.386906f
C37 B1 VNB 0.425176f
C38 VPB VNB 2.0223f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211a_1 VNB VPB VGND VPWR X A1 A2 B1 C1
X0 VGND.t1 A1.t0 a_215_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47.t1 B1.t0 a_215_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21.t1 C1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR.t2 B1.t1 a_79_21.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21.t3 A2.t0 a_297_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297.t1 A1.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21.t0 C1.t1 a_510_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR.t1 a_79_21.t4 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND.t0 a_79_21.t5 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47.t2 A2.t1 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
R0 A1.n0 A1.t1 241.536
R1 A1.n0 A1.t0 169.237
R2 A1 A1.n0 157.44
R3 a_215_47.t0 a_215_47.n0 280.779
R4 a_215_47.n0 a_215_47.t1 56.3082
R5 a_215_47.n0 a_215_47.t2 24.9236
R6 VGND.n1 VGND.n0 212.492
R7 VGND.n1 VGND.t0 161.15
R8 VGND.n0 VGND.t1 30.462
R9 VGND.n0 VGND.t2 29.539
R10 VGND VGND.n1 0.436086
R11 VNB.t0 VNB.t2 2677.02
R12 VNB.t4 VNB.t3 1680.26
R13 VNB.t3 VNB.t1 1423.95
R14 VNB.t2 VNB.t4 1352.75
R15 VNB VNB.t0 911.327
R16 B1.n0 B1.t1 239.505
R17 B1.n0 B1.t0 167.204
R18 B1 B1.n0 157.44
R19 a_510_47.t0 a_510_47.t1 64.6159
R20 C1 C1.n0 217.548
R21 C1.n0 C1.t0 212.081
R22 C1.n0 C1.t1 139.78
R23 VPWR.n3 VPWR.t3 342.841
R24 VPWR.n2 VPWR.n1 316.767
R25 VPWR.n5 VPWR.t1 257.474
R26 VPWR.n6 VPWR.n5 43.1829
R27 VPWR.n1 VPWR.t0 34.4755
R28 VPWR.n1 VPWR.t2 34.4755
R29 VPWR.n4 VPWR.n3 25.977
R30 VPWR.n4 VPWR.n0 9.3005
R31 VPWR.n3 VPWR.n2 7.14534
R32 VPWR.n5 VPWR.n4 0.753441
R33 VPWR.n2 VPWR.n0 0.193172
R34 VPWR.n6 VPWR.n0 0.120292
R35 VPWR VPWR.n6 0.0213333
R36 a_79_21.n2 a_79_21.n0 271.341
R37 a_79_21.t1 a_79_21.n3 246.155
R38 a_79_21.n0 a_79_21.t4 239.548
R39 a_79_21.n2 a_79_21.n1 205.28
R40 a_79_21.n3 a_79_21.t0 178.083
R41 a_79_21.n0 a_79_21.t5 167.248
R42 a_79_21.n1 a_79_21.t2 60.0855
R43 a_79_21.n3 a_79_21.n2 53.8358
R44 a_79_21.n1 a_79_21.t3 26.5955
R45 VPB.t1 VPB.t4 556.386
R46 VPB.t3 VPB.t2 349.221
R47 VPB.t2 VPB.t0 295.95
R48 VPB.t4 VPB.t3 281.154
R49 VPB VPB.t1 189.409
R50 A2.n0 A2.t0 233.01
R51 A2.n0 A2.t1 160.709
R52 A2 A2.n0 154.133
R53 a_297_297.t0 a_297_297.t1 64.0255
R54 X.n2 X 593.095
R55 X.n2 X.n0 585
R56 X.n3 X.n2 585
R57 X.n1 X.t0 129.381
R58 X.n3 X.n1 62.368
R59 X.n2 X.t1 26.5955
R60 X X.n0 8.09462
R61 X.n1 X 5.55208
R62 X X.n0 4.70638
R63 X X.n3 4.70638
C0 VPWR VGND 0.073222f
C1 X A2 2.44e-19
C2 VGND C1 0.013287f
C3 VPB VGND 0.010817f
C4 A1 VPWR 0.018399f
C5 A2 B1 0.061079f
C6 VPB A1 0.032154f
C7 X VGND 0.099278f
C8 VPWR C1 0.020287f
C9 VGND B1 0.018554f
C10 A1 X 3.68e-19
C11 VPB VPWR 0.094379f
C12 VPB C1 0.055253f
C13 X VPWR 0.128521f
C14 VGND A2 0.015871f
C15 VPWR B1 0.018452f
C16 VPB X 0.01253f
C17 B1 C1 0.049531f
C18 VPB B1 0.029836f
C19 A1 A2 0.069292f
C20 X B1 1.2e-19
C21 VPWR A2 0.014254f
C22 A1 VGND 0.017007f
C23 VPB A2 0.033967f
C24 VGND VNB 0.449857f
C25 VPWR VNB 0.376877f
C26 X VNB 0.095064f
C27 C1 VNB 0.167477f
C28 B1 VNB 0.095044f
C29 A2 VNB 0.100735f
C30 A1 VNB 0.098893f
C31 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211a_2 VNB VPB VPWR VGND A2 A1 X C1 B1
X0 a_27_47.t1 B1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND.t3 a_27_47.t4 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.23075 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR.t2 C1.t0 a_27_47.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR.t0 A1.t0 a_373_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47.t1 A2.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 X.t3 a_27_47.t5 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47.t2 B1.t1 a_110_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.16535 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 X.t0 a_27_47.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297.t1 A2.t1 a_27_47.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3675 ps=1.735 w=1 l=0.15
X9 a_110_47.t0 C1.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 VPWR.t4 a_27_47.t7 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND.t1 A1.t1 a_182_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
R0 B1.n0 B1.t0 235.471
R1 B1.n0 B1.t1 163.172
R2 B1 B1.n0 156.073
R3 VPWR.n5 VPWR.t4 869.639
R4 VPWR.n10 VPWR.n1 309.724
R5 VPWR.n4 VPWR.n3 305.726
R6 VPWR.n3 VPWR.t3 39.4005
R7 VPWR.n3 VPWR.t0 37.4305
R8 VPWR.n8 VPWR.n2 34.6358
R9 VPWR.n9 VPWR.n8 34.6358
R10 VPWR.n1 VPWR.t1 27.5805
R11 VPWR.n1 VPWR.t2 27.5805
R12 VPWR.n10 VPWR.n9 22.2123
R13 VPWR.n4 VPWR.n2 9.78874
R14 VPWR.n6 VPWR.n2 9.3005
R15 VPWR.n8 VPWR.n7 9.3005
R16 VPWR.n9 VPWR.n0 9.3005
R17 VPWR.n11 VPWR.n10 7.16074
R18 VPWR.n5 VPWR.n4 6.68542
R19 VPWR.n6 VPWR.n5 0.731811
R20 VPWR.n11 VPWR.n0 0.148009
R21 VPWR.n7 VPWR.n6 0.120292
R22 VPWR.n7 VPWR.n0 0.120292
R23 VPWR VPWR.n11 0.114057
R24 a_27_47.n5 a_27_47.t3 406.817
R25 a_27_47.n7 a_27_47.n6 292.5
R26 a_27_47.n4 a_27_47.n0 292.5
R27 a_27_47.n1 a_27_47.t7 216.654
R28 a_27_47.n2 a_27_47.t5 213.688
R29 a_27_47.n5 a_27_47.t0 183.719
R30 a_27_47.n2 a_27_47.t6 142.746
R31 a_27_47.n1 a_27_47.t4 139.78
R32 a_27_47.n4 a_27_47.n3 135.462
R33 a_27_47.n7 a_27_47.n0 66.9805
R34 a_27_47.t1 a_27_47.n7 41.3705
R35 a_27_47.n0 a_27_47.t2 36.4455
R36 a_27_47.n3 a_27_47.n2 29.749
R37 a_27_47.n3 a_27_47.n1 24.1425
R38 a_27_47.n6 a_27_47.n5 22.5414
R39 a_27_47.n6 a_27_47.n4 4.55757
R40 VPB.t1 VPB.t2 523.832
R41 VPB.t0 VPB.t5 319.627
R42 VPB.t5 VPB.t4 254.518
R43 VPB.t3 VPB.t1 254.518
R44 VPB.t2 VPB.t0 213.084
R45 VPB VPB.t3 192.369
R46 X X.n0 712.271
R47 X X.n1 122.163
R48 X.n0 X.t2 27.5805
R49 X.n0 X.t3 27.5805
R50 X.n1 X.t1 25.8467
R51 X.n1 X.t0 25.8467
R52 VGND.n1 VGND.t3 244.201
R53 VGND.n5 VGND.t0 226.808
R54 VGND.n3 VGND.n2 204.609
R55 VGND.n2 VGND.t2 29.539
R56 VGND.n2 VGND.t1 29.539
R57 VGND.n5 VGND.n4 25.977
R58 VGND.n4 VGND.n3 18.4476
R59 VGND.n4 VGND.n0 9.3005
R60 VGND.n3 VGND.n1 7.07217
R61 VGND.n6 VGND.n5 6.7997
R62 VGND.n1 VGND.n0 0.600593
R63 VGND VGND.n6 0.343375
R64 VGND.n6 VGND.n0 0.159366
R65 VNB.t2 VNB.t1 2662.78
R66 VNB.t3 VNB.t4 1338.51
R67 VNB.t4 VNB.t5 1224.6
R68 VNB.t1 VNB.t3 1224.6
R69 VNB.t0 VNB.t2 1025.24
R70 VNB VNB.t0 925.567
R71 C1.n0 C1.t0 220.367
R72 C1.n0 C1.t1 157.653
R73 C1 C1.n0 156.849
R74 A1.n0 A1.t0 237.736
R75 A1.n0 A1.t1 165.435
R76 A1 A1.n0 161.697
R77 a_373_297.t0 a_373_297.t1 41.3705
R78 A2.n0 A2.t1 220.608
R79 A2.n0 A2.t0 160.173
R80 A2 A2.n0 158.012
R81 a_182_47.n0 a_182_47.t2 460.615
R82 a_182_47.t0 a_182_47.n0 25.8467
R83 a_182_47.n0 a_182_47.t1 25.8467
R84 a_110_47.t0 a_110_47.t1 38.7697
C0 A1 VPWR 0.01765f
C1 VGND VPWR 0.074137f
C2 C1 VPWR 0.019442f
C3 B1 VGND 0.016263f
C4 C1 B1 0.06f
C5 A2 VPWR 0.017479f
C6 VGND A1 0.025124f
C7 X VPWR 0.144258f
C8 B1 A2 0.047441f
C9 VPB VPWR 0.079237f
C10 C1 VGND 0.011308f
C11 B1 X 1.43e-19
C12 VPB B1 0.033915f
C13 X A1 0.001799f
C14 A2 A1 0.089722f
C15 VGND A2 0.019127f
C16 X VGND 0.13482f
C17 VPB A1 0.028091f
C18 VPB VGND 0.007904f
C19 VPB C1 0.038768f
C20 X A2 6.03e-19
C21 VPB X 0.012847f
C22 VPB A2 0.036003f
C23 B1 VPWR 0.020338f
C24 VGND VNB 0.45041f
C25 X VNB 0.071998f
C26 VPWR VNB 0.371183f
C27 A1 VNB 0.093059f
C28 A2 VNB 0.106828f
C29 B1 VNB 0.102823f
C30 C1 VNB 0.146137f
C31 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211a_4 VNB VPB VGND VPWR X C1 B1 A2 A1
X0 VGND.t1 A1.t0 a_474_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.104 ps=0.97 w=0.65 l=0.15
X1 VPWR.t6 a_79_21.t8 X.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR.t2 A1.t1 a_1122_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X.t0 a_79_21.t9 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 a_79_21.t6 B1.t0 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.2525 pd=1.505 as=0.14 ps=1.28 w=1 l=0.15
X5 VGND.t3 a_79_21.t10 X.t7 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND.t4 a_79_21.t11 X.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t7 C1.t0 a_79_21.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2525 ps=1.505 w=1 l=0.15
X8 a_950_297.t0 A1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X9 a_557_47.t0 B1.t1 a_474_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 a_474_47.t4 B1.t2 a_748_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND.t7 A2.t0 a_474_47.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 VPWR.t4 a_79_21.t12 X.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 X.t5 a_79_21.t13 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_79_21.t3 C1.t1 a_557_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.144625 pd=1.095 as=0.06825 ps=0.86 w=0.65 l=0.15
X15 a_474_47.t0 A1.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_79_21.t4 C1.t2 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X17 a_748_47.t1 C1.t3 a_79_21.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.144625 ps=1.095 w=0.65 l=0.15
X18 a_474_47.t2 A2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X19 VPWR.t0 B1.t3 a_79_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.195 ps=1.39 w=1 l=0.15
X20 a_79_21.t5 A2.t2 a_950_297.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 a_1122_297.t1 A2.t3 a_79_21.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 X.t2 a_79_21.t14 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 X.t4 a_79_21.t15 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1 A1.n0 242.544
R1 A1.n0 A1.t2 236.18
R2 A1.n1 A1.t1 231.963
R3 A1.n0 A1.t0 163.881
R4 A1 A1.n1 161.12
R5 A1.n1 A1.t3 159.663
R6 a_474_47.n1 a_474_47.t3 377.3
R7 a_474_47.t0 a_474_47.n3 176.292
R8 a_474_47.n3 a_474_47.n2 98.788
R9 a_474_47.n1 a_474_47.n0 89.3175
R10 a_474_47.n3 a_474_47.n1 56.4614
R11 a_474_47.n0 a_474_47.t4 30.462
R12 a_474_47.n0 a_474_47.t1 28.6159
R13 a_474_47.n2 a_474_47.t5 25.8467
R14 a_474_47.n2 a_474_47.t2 25.8467
R15 VGND.n23 VGND.t6 282.817
R16 VGND.n17 VGND.t4 271.546
R17 VGND.n7 VGND.n6 215.166
R18 VGND.n9 VGND.n8 199.63
R19 VGND.n21 VGND.n2 198.964
R20 VGND.n8 VGND.t2 38.7697
R21 VGND.n11 VGND.n10 34.6358
R22 VGND.n11 VGND.n4 34.6358
R23 VGND.n15 VGND.n4 34.6358
R24 VGND.n16 VGND.n15 34.6358
R25 VGND.n8 VGND.t1 33.2313
R26 VGND.n17 VGND.n16 29.3652
R27 VGND.n21 VGND.n1 25.977
R28 VGND.n6 VGND.t0 25.8467
R29 VGND.n6 VGND.t7 25.8467
R30 VGND.n2 VGND.t5 24.9236
R31 VGND.n2 VGND.t3 24.9236
R32 VGND.n10 VGND.n9 22.5887
R33 VGND.n23 VGND.n22 19.9534
R34 VGND.n22 VGND.n21 18.4476
R35 VGND.n17 VGND.n1 12.424
R36 VGND.n24 VGND.n23 9.3005
R37 VGND.n10 VGND.n5 9.3005
R38 VGND.n12 VGND.n11 9.3005
R39 VGND.n13 VGND.n4 9.3005
R40 VGND.n15 VGND.n14 9.3005
R41 VGND.n16 VGND.n3 9.3005
R42 VGND.n18 VGND.n17 9.3005
R43 VGND.n19 VGND.n1 9.3005
R44 VGND.n21 VGND.n20 9.3005
R45 VGND.n22 VGND.n0 9.3005
R46 VGND.n9 VGND.n7 6.72553
R47 VGND.n7 VGND.n5 0.519559
R48 VGND.n12 VGND.n5 0.120292
R49 VGND.n13 VGND.n12 0.120292
R50 VGND.n14 VGND.n13 0.120292
R51 VGND.n14 VGND.n3 0.120292
R52 VGND.n18 VGND.n3 0.120292
R53 VGND.n19 VGND.n18 0.120292
R54 VGND.n20 VGND.n19 0.120292
R55 VGND.n20 VGND.n0 0.120292
R56 VGND.n24 VGND.n0 0.120292
R57 VGND VGND.n24 0.0226354
R58 VNB.t7 VNB.t3 2790.94
R59 VNB.t5 VNB.t11 1694.5
R60 VNB.t1 VNB.t2 1537.86
R61 VNB.t4 VNB.t1 1338.51
R62 VNB.t10 VNB.t0 1224.6
R63 VNB.t2 VNB.t10 1224.6
R64 VNB.t11 VNB.t4 1224.6
R65 VNB.t8 VNB.t7 1196.12
R66 VNB.t6 VNB.t8 1196.12
R67 VNB.t9 VNB.t6 1196.12
R68 VNB.t3 VNB.t5 1025.24
R69 VNB VNB.t9 925.567
R70 a_79_21.n20 a_79_21.n19 598.755
R71 a_79_21.n17 a_79_21.n16 585
R72 a_79_21.n19 a_79_21.n18 376.793
R73 a_79_21.n15 a_79_21.n0 279.913
R74 a_79_21.n13 a_79_21.t8 225.226
R75 a_79_21.n11 a_79_21.t14 212.081
R76 a_79_21.n4 a_79_21.t12 212.081
R77 a_79_21.n5 a_79_21.t9 212.081
R78 a_79_21.n8 a_79_21.n3 173.761
R79 a_79_21.n3 a_79_21.t15 173.375
R80 a_79_21.n8 a_79_21.n7 152
R81 a_79_21.n10 a_79_21.n9 152
R82 a_79_21.n11 a_79_21.n1 152
R83 a_79_21.n14 a_79_21.n13 152
R84 a_79_21.n6 a_79_21.t10 139.78
R85 a_79_21.n2 a_79_21.t13 139.78
R86 a_79_21.n12 a_79_21.t11 139.78
R87 a_79_21.n17 a_79_21.n15 79.7629
R88 a_79_21.n19 a_79_21.n17 58.051
R89 a_79_21.n16 a_79_21.t2 52.2055
R90 a_79_21.n11 a_79_21.n10 49.6611
R91 a_79_21.n13 a_79_21.n12 48.2005
R92 a_79_21.n16 a_79_21.t6 47.2805
R93 a_79_21.n0 a_79_21.t7 43.3851
R94 a_79_21.n20 a_79_21.t4 41.3705
R95 a_79_21.n0 a_79_21.t3 38.7697
R96 a_79_21.n7 a_79_21.n4 36.5157
R97 a_79_21.t0 a_79_21.n20 35.4605
R98 a_79_21.n18 a_79_21.t1 27.5805
R99 a_79_21.n18 a_79_21.t5 27.5805
R100 a_79_21.n5 a_79_21.n3 23.3702
R101 a_79_21.n7 a_79_21.n6 21.9096
R102 a_79_21.n14 a_79_21.n1 21.7605
R103 a_79_21.n9 a_79_21.n1 21.7605
R104 a_79_21.n9 a_79_21.n8 21.7605
R105 a_79_21.n15 a_79_21.n14 14.4005
R106 a_79_21.n10 a_79_21.n2 10.2247
R107 a_79_21.n6 a_79_21.n5 4.38232
R108 a_79_21.n4 a_79_21.n2 2.92171
R109 a_79_21.n12 a_79_21.n11 1.46111
R110 X.n2 X.n1 351.517
R111 X.n2 X.n0 310.683
R112 X.n5 X.n4 256.272
R113 X.n5 X.n3 199.683
R114 X X.n2 70.6248
R115 X.n1 X.t1 27.5805
R116 X.n1 X.t2 27.5805
R117 X.n0 X.t3 27.5805
R118 X.n0 X.t0 27.5805
R119 X X.n5 25.1016
R120 X.n3 X.t7 24.9236
R121 X.n3 X.t4 24.9236
R122 X.n4 X.t6 24.9236
R123 X.n4 X.t5 24.9236
R124 VPWR.n8 VPWR.n7 602.389
R125 VPWR.n4 VPWR.n3 600.515
R126 VPWR.n12 VPWR.n6 598.965
R127 VPWR.n9 VPWR.t2 345.397
R128 VPWR.n20 VPWR.t5 338.507
R129 VPWR.n18 VPWR.n2 310.928
R130 VPWR.n7 VPWR.t1 35.4605
R131 VPWR.n13 VPWR.n4 34.6358
R132 VPWR.n18 VPWR.n17 30.1181
R133 VPWR.n11 VPWR.n8 28.6123
R134 VPWR.n2 VPWR.t3 27.5805
R135 VPWR.n2 VPWR.t4 27.5805
R136 VPWR.n3 VPWR.t9 27.5805
R137 VPWR.n3 VPWR.t6 27.5805
R138 VPWR.n6 VPWR.t8 27.5805
R139 VPWR.n6 VPWR.t7 27.5805
R140 VPWR.n7 VPWR.t0 27.5805
R141 VPWR.n20 VPWR.n19 25.6005
R142 VPWR.n13 VPWR.n12 22.2123
R143 VPWR.n12 VPWR.n11 22.2123
R144 VPWR.n19 VPWR.n18 14.3064
R145 VPWR.n17 VPWR.n4 9.78874
R146 VPWR.n11 VPWR.n10 9.3005
R147 VPWR.n12 VPWR.n5 9.3005
R148 VPWR.n14 VPWR.n13 9.3005
R149 VPWR.n15 VPWR.n4 9.3005
R150 VPWR.n17 VPWR.n16 9.3005
R151 VPWR.n18 VPWR.n1 9.3005
R152 VPWR.n19 VPWR.n0 9.3005
R153 VPWR.n21 VPWR.n20 6.96759
R154 VPWR.n9 VPWR.n8 6.95582
R155 VPWR.n10 VPWR.n9 0.175003
R156 VPWR.n21 VPWR.n0 0.150466
R157 VPWR.n10 VPWR.n5 0.120292
R158 VPWR.n14 VPWR.n5 0.120292
R159 VPWR.n15 VPWR.n14 0.120292
R160 VPWR.n16 VPWR.n15 0.120292
R161 VPWR.n16 VPWR.n1 0.120292
R162 VPWR.n1 VPWR.n0 0.120292
R163 VPWR VPWR.n21 0.112871
R164 VPB VPB.t6 423.209
R165 VPB.t11 VPB.t8 387.695
R166 VPB.t9 VPB.t0 319.627
R167 VPB.t0 VPB.t1 278.193
R168 VPB.t3 VPB.t2 254.518
R169 VPB.t10 VPB.t3 254.518
R170 VPB.t1 VPB.t10 254.518
R171 VPB.t8 VPB.t9 254.518
R172 VPB.t7 VPB.t11 254.518
R173 VPB.t4 VPB.t7 254.518
R174 VPB.t5 VPB.t4 254.518
R175 VPB.t6 VPB.t5 254.518
R176 a_1122_297.t0 a_1122_297.t1 55.1605
R177 B1.n0 B1.t0 239.04
R178 B1.n1 B1.t3 236.18
R179 B1 B1.n0 222.677
R180 B1.n0 B1.t1 166.739
R181 B1.n1 B1.t2 163.881
R182 B1 B1.n1 163.055
R183 C1.n1 C1.t0 212.081
R184 C1.n0 C1.t2 212.081
R185 C1.n1 C1.t1 163.881
R186 C1.n0 C1.t3 139.78
R187 C1 C1.n2 69.762
R188 C1.n2 C1.n0 34.9807
R189 C1.n2 C1.n1 21.1941
R190 a_950_297.t0 a_950_297.t1 55.1605
R191 a_557_47.t0 a_557_47.t1 38.7697
R192 a_748_47.t0 a_748_47.t1 51.6928
R193 A2.n0 A2.t3 212.081
R194 A2.n1 A2.t2 212.081
R195 A2.n0 A2.t0 139.78
R196 A2.n1 A2.t1 139.78
R197 A2 A2.n2 68.8661
R198 A2.n2 A2.n1 33.651
R199 A2.n2 A2.n0 22.4676
C0 X VGND 0.223508f
C1 B1 VGND 0.023384f
C2 VPB VGND 0.010036f
C3 A1 A2 0.228421f
C4 C1 VPWR 0.032396f
C5 B1 X 0.001071f
C6 VPB X 0.023952f
C7 B1 VPB 0.06927f
C8 VPWR VGND 0.127718f
C9 VPWR X 0.326777f
C10 B1 VPWR 0.043555f
C11 VPB VPWR 0.142104f
C12 A2 VGND 0.031935f
C13 B1 A2 6.95e-20
C14 VPB A2 0.056085f
C15 A1 VGND 0.036559f
C16 B1 A1 0.099515f
C17 A1 VPB 0.076448f
C18 A2 VPWR 0.027478f
C19 C1 VGND 0.018299f
C20 C1 X 2.17e-19
C21 A1 VPWR 0.083379f
C22 B1 C1 0.221164f
C23 C1 VPB 0.064626f
C24 VGND VNB 0.723618f
C25 X VNB 0.068448f
C26 VPWR VNB 0.629562f
C27 A2 VNB 0.177039f
C28 A1 VNB 0.251402f
C29 C1 VNB 0.187493f
C30 B1 VNB 0.193148f
C31 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_1 VPB VNB VGND VPWR A1 Y C1 B1 A2
X0 a_110_297.t1 A1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND.t0 A1.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X2 Y.t1 A2.t0 a_110_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR.t2 B1.t0 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47.t2 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_326_47.t0 B1.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 Y.t0 C1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y.t3 C1.t1 a_326_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
R0 A1.n0 A1.t0 233.288
R1 A1.n0 A1.t1 160.988
R2 A1 A1.n0 158.4
R3 VPWR.n1 VPWR.n0 604.893
R4 VPWR.n1 VPWR.t1 251.344
R5 VPWR.n0 VPWR.t0 45.3105
R6 VPWR.n0 VPWR.t2 31.5205
R7 VPWR VPWR.n1 0.138192
R8 a_110_297.t0 a_110_297.t1 41.3705
R9 VPB.t3 VPB.t0 319.627
R10 VPB.t1 VPB.t3 319.627
R11 VPB.t2 VPB.t1 213.084
R12 VPB VPB.t2 195.327
R13 a_27_47.n0 a_27_47.t1 272.409
R14 a_27_47.n0 a_27_47.t2 36.9236
R15 a_27_47.t0 a_27_47.n0 35.0774
R16 VGND VGND.n0 204.78
R17 VGND.n0 VGND.t0 38.7697
R18 VGND.n0 VGND.t1 33.2313
R19 VNB.t2 VNB.t0 1537.86
R20 VNB.t1 VNB.t2 1537.86
R21 VNB.t0 VNB.t3 1025.24
R22 VNB VNB.t1 939.807
R23 A2.n0 A2.t0 236.18
R24 A2 A2.n0 168.988
R25 A2.n0 A2.t1 163.881
R26 Y.n1 Y.n0 244.631
R27 Y.n1 Y.t0 209.291
R28 Y.n2 Y.t3 103.481
R29 Y.n2 Y.n1 71.0047
R30 Y.n0 Y.t1 39.4005
R31 Y.n0 Y.t2 37.4305
R32 Y Y.n2 2.25402
R33 B1.n0 B1.t0 230.923
R34 B1.n0 B1.t1 163.881
R35 B1 B1.n0 153.423
R36 a_326_47.t0 a_326_47.t1 38.7697
R37 C1.n0 C1.t0 230.576
R38 C1 C1.n0 163.055
R39 C1.n0 C1.t1 158.275
C0 VGND Y 0.100793f
C1 C1 Y 0.132967f
C2 VGND B1 0.021486f
C3 C1 B1 0.108739f
C4 Y A1 9.85e-19
C5 VPWR A2 0.087669f
C6 VGND VPWR 0.05511f
C7 C1 VPWR 0.017106f
C8 VGND A2 0.018293f
C9 VPWR A1 0.04837f
C10 A1 A2 0.09342f
C11 VPB Y 0.014362f
C12 VPB B1 0.034654f
C13 VGND C1 0.016045f
C14 VGND A1 0.01599f
C15 Y B1 0.058586f
C16 VPB VPWR 0.065014f
C17 VPB A2 0.033538f
C18 VPWR Y 0.235943f
C19 Y A2 0.068242f
C20 VGND VPB 0.004938f
C21 VPWR B1 0.022673f
C22 VPB C1 0.042819f
C23 A2 B1 0.077303f
C24 VPB A1 0.034077f
C25 VGND VNB 0.342128f
C26 Y VNB 0.103729f
C27 VPWR VNB 0.319183f
C28 C1 VNB 0.128953f
C29 B1 VNB 0.096625f
C30 A2 VNB 0.105185f
C31 A1 VNB 0.142014f
C32 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_2 VNB VPB VGND VPWR Y B1 A2 A1 C1
X0 a_286_47.t5 A1.t0 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR.t3 B1.t0 Y.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47.t2 A2.t0 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y.t3 A2.t1 a_487_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND.t2 A1.t1 a_286_47.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y.t4 C1.t0 a_27_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND.t1 A2.t2 a_286_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297.t0 A2.t3 Y.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47.t1 B1.t1 a_286_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR.t0 C1.t1 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR.t5 A1.t2 a_487_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47.t2 C1.t2 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y.t2 C1.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297.t2 A1.t3 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47.t1 B1.t2 a_27_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y.t6 B1.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A1.n1 A1.t3 212.081
R1 A1.n0 A1.t2 212.081
R2 A1.n1 A1.t1 139.78
R3 A1.n0 A1.t0 139.78
R4 A1 A1.n2 91.8412
R5 A1.n2 A1.n1 28.2474
R6 A1.n2 A1.n0 27.9568
R7 VGND.n1 VGND.t2 289.327
R8 VGND.n5 VGND.t0 283.175
R9 VGND.n3 VGND.n2 198.964
R10 VGND.n2 VGND.t3 25.8467
R11 VGND.n2 VGND.t1 25.8467
R12 VGND.n4 VGND.n3 19.9534
R13 VGND.n5 VGND.n4 19.9534
R14 VGND.n4 VGND.n0 9.3005
R15 VGND.n6 VGND.n5 7.18495
R16 VGND.n3 VGND.n1 6.55962
R17 VGND.n1 VGND.n0 0.734976
R18 VGND VGND.n6 0.591245
R19 VGND.n6 VGND.n0 0.153642
R20 a_286_47.n2 a_286_47.n0 271.553
R21 a_286_47.n3 a_286_47.n2 237.419
R22 a_286_47.n2 a_286_47.n1 185
R23 a_286_47.n0 a_286_47.t0 25.8467
R24 a_286_47.n0 a_286_47.t1 25.8467
R25 a_286_47.n1 a_286_47.t3 25.8467
R26 a_286_47.n1 a_286_47.t2 25.8467
R27 a_286_47.t4 a_286_47.n3 25.8467
R28 a_286_47.n3 a_286_47.t5 25.8467
R29 VNB.t1 VNB.t3 2819.42
R30 VNB.t7 VNB.t6 1224.6
R31 VNB.t5 VNB.t7 1224.6
R32 VNB.t3 VNB.t5 1224.6
R33 VNB.t2 VNB.t1 1224.6
R34 VNB.t0 VNB.t2 1224.6
R35 VNB.t4 VNB.t0 1224.6
R36 VNB VNB.t4 996.764
R37 B1.n0 B1.t0 212.081
R38 B1.n1 B1.t3 212.081
R39 B1.n0 B1.t1 139.78
R40 B1.n1 B1.t2 139.78
R41 B1 B1.n2 69.6396
R42 B1.n2 B1.n0 35.403
R43 B1.n2 B1.n1 21.1033
R44 Y.n2 Y.n0 386.01
R45 Y.n2 Y.n1 314.789
R46 Y.n4 Y.n3 307.005
R47 Y Y.n5 185.195
R48 Y.n4 Y.n2 45.177
R49 Y Y.n4 33.3581
R50 Y.n0 Y.t5 27.5805
R51 Y.n0 Y.t3 27.5805
R52 Y.n1 Y.t7 27.5805
R53 Y.n1 Y.t6 27.5805
R54 Y.n3 Y.t0 27.5805
R55 Y.n3 Y.t2 27.5805
R56 Y.n5 Y.t1 25.8467
R57 Y.n5 Y.t4 25.8467
R58 VPWR.n10 VPWR.t1 867.614
R59 VPWR.n3 VPWR.t3 338.082
R60 VPWR.n5 VPWR.n4 317.075
R61 VPWR.n8 VPWR.n2 310.502
R62 VPWR.n2 VPWR.t2 27.5805
R63 VPWR.n2 VPWR.t0 27.5805
R64 VPWR.n4 VPWR.t4 27.5805
R65 VPWR.n4 VPWR.t5 27.5805
R66 VPWR.n10 VPWR.n9 23.7181
R67 VPWR.n8 VPWR.n7 22.9652
R68 VPWR.n9 VPWR.n8 21.4593
R69 VPWR.n7 VPWR.n3 16.9417
R70 VPWR.n7 VPWR.n6 9.3005
R71 VPWR.n8 VPWR.n1 9.3005
R72 VPWR.n9 VPWR.n0 9.3005
R73 VPWR.n11 VPWR.n10 9.3005
R74 VPWR.n5 VPWR.n3 7.31426
R75 VPWR.n6 VPWR.n5 0.165196
R76 VPWR.n6 VPWR.n1 0.120292
R77 VPWR.n1 VPWR.n0 0.120292
R78 VPWR.n11 VPWR.n0 0.120292
R79 VPWR VPWR.n11 0.0226354
R80 VPB.t5 VPB.t2 585.981
R81 VPB.t7 VPB.t6 254.518
R82 VPB.t3 VPB.t7 254.518
R83 VPB.t2 VPB.t3 254.518
R84 VPB.t4 VPB.t5 254.518
R85 VPB.t0 VPB.t4 254.518
R86 VPB.t1 VPB.t0 254.518
R87 VPB VPB.t1 207.166
R88 A2.n1 A2.t3 212.081
R89 A2.n0 A2.t1 212.081
R90 A2.n1 A2.t2 139.78
R91 A2.n0 A2.t0 139.78
R92 A2 A2.n2 86.5779
R93 A2.n2 A2.n0 28.4795
R94 A2.n2 A2.n1 27.6489
R95 a_487_297.t1 a_487_297.n1 893.913
R96 a_487_297.n1 a_487_297.t2 421.942
R97 a_487_297.n1 a_487_297.n0 284.714
R98 a_487_297.n0 a_487_297.t3 27.5805
R99 a_487_297.n0 a_487_297.t0 27.5805
R100 C1.n0 C1.t1 212.081
R101 C1.n1 C1.t3 212.081
R102 C1 C1.n1 201.826
R103 C1.n0 C1.t2 139.78
R104 C1.n1 C1.t0 139.78
R105 C1.n1 C1.n0 62.8066
R106 a_27_47.n1 a_27_47.t3 326.538
R107 a_27_47.t1 a_27_47.n1 321.63
R108 a_27_47.n1 a_27_47.n0 96.3734
R109 a_27_47.n0 a_27_47.t0 25.8467
R110 a_27_47.n0 a_27_47.t2 25.8467
C0 VPWR VPB 0.105496f
C1 B1 VPB 0.063555f
C2 VPWR Y 0.333303f
C3 B1 Y 0.130573f
C4 A2 VPWR 0.020626f
C5 B1 A2 0.02957f
C6 B1 VPWR 0.041766f
C7 VGND C1 0.020559f
C8 A1 C1 3.91e-20
C9 A1 VGND 0.06615f
C10 VPB C1 0.07739f
C11 VGND VPB 0.009876f
C12 Y C1 0.147072f
C13 A1 VPB 0.059742f
C14 Y VGND 0.014562f
C15 A2 VGND 0.035398f
C16 A1 Y 0.001638f
C17 A2 A1 0.07322f
C18 Y VPB 0.02119f
C19 VPWR C1 0.07083f
C20 A2 VPB 0.06259f
C21 B1 C1 0.05901f
C22 VPWR VGND 0.091116f
C23 A1 VPWR 0.043112f
C24 A2 Y 0.084235f
C25 B1 VGND 0.019943f
C26 B1 A1 2.66e-19
C27 VGND VNB 0.537836f
C28 Y VNB 0.027292f
C29 VPWR VNB 0.448395f
C30 A1 VNB 0.231963f
C31 A2 VNB 0.190869f
C32 B1 VNB 0.191845f
C33 C1 VNB 0.263095f
C34 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_4 VNB VPB VGND VPWR C1 A2 A1 Y B1
X0 VPWR.t7 A1.t0 a_110_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y.t7 A2.t0 a_110_297.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_806_47.t3 B1.t0 a_27_47.t8 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_110_297.t0 A2.t1 Y.t6 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_297.t3 A1.t1 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND.t7 A1.t2 a_27_47.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VPWR.t0 B1.t1 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_110_297.t2 A1.t3 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47.t3 A2.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR.t4 A1.t4 a_110_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR.t10 C1.t0 Y.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47.t11 B1.t2 a_1314_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=2.09 as=0.104 ps=0.97 w=0.65 l=0.15
X12 Y.t8 C1.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47.t6 A1.t5 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 VPWR.t9 C1.t2 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y.t15 B1.t3 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND.t5 A1.t6 a_27_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X17 Y.t5 A2.t3 a_110_297.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_27_47.t4 A1.t7 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.09425 ps=0.94 w=0.65 l=0.15
X19 Y.t12 C1.t3 a_978_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y.t14 C1.t4 a_806_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_27_47.t2 A2.t4 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_27_47.t9 B1.t4 a_806_47.t2 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_110_297.t7 A2.t5 Y.t4 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 a_806_47.t0 C1.t5 Y.t13 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VPWR.t1 B1.t5 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.675 pd=3.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND.t1 A2.t6 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.091 ps=0.93 w=0.65 l=0.15
X27 a_978_47.t1 B1.t6 a_27_47.t10 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_1314_47.t0 C1.t6 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t9 C1.t7 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y.t3 B1.t7 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X31 VGND.t0 A2.t7 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 A1.n1 A1.n0 321.647
R1 A1.n0 A1.t4 236.18
R2 A1.n5 A1.t0 212.081
R3 A1.n3 A1.t3 212.081
R4 A1.n2 A1.t1 212.081
R5 A1.n0 A1.t7 163.881
R6 A1.n4 A1.n1 152
R7 A1.n5 A1.t5 139.78
R8 A1.n3 A1.t2 139.78
R9 A1.n2 A1.t6 139.78
R10 A1 A1.n6 74.5342
R11 A1.n5 A1.n4 49.6611
R12 A1.n6 A1.n2 35.7937
R13 A1.n6 A1.n5 20.3621
R14 A1.n4 A1.n3 13.146
R15 A1 A1.n1 3.67263
R16 a_110_297.n2 a_110_297.n0 649.453
R17 a_110_297.n5 a_110_297.n4 642.938
R18 a_110_297.n2 a_110_297.n1 585
R19 a_110_297.n4 a_110_297.n3 585
R20 a_110_297.n4 a_110_297.n2 66.452
R21 a_110_297.n3 a_110_297.t5 27.5805
R22 a_110_297.n3 a_110_297.t7 27.5805
R23 a_110_297.n1 a_110_297.t6 27.5805
R24 a_110_297.n1 a_110_297.t2 27.5805
R25 a_110_297.n0 a_110_297.t4 27.5805
R26 a_110_297.n0 a_110_297.t3 27.5805
R27 a_110_297.n5 a_110_297.t1 27.5805
R28 a_110_297.t0 a_110_297.n5 27.5805
R29 VPWR.n11 VPWR.t1 710.241
R30 VPWR.n6 VPWR.n5 602.067
R31 VPWR.n31 VPWR.n2 598.965
R32 VPWR.n19 VPWR.n8 598.965
R33 VPWR.n10 VPWR.n9 598.965
R34 VPWR.n13 VPWR.n12 598.755
R35 VPWR.n33 VPWR.t6 406.757
R36 VPWR.n25 VPWR.n24 34.6358
R37 VPWR.n26 VPWR.n25 34.6358
R38 VPWR.n26 VPWR.n3 34.6358
R39 VPWR.n30 VPWR.n3 34.6358
R40 VPWR.n21 VPWR.n20 34.6358
R41 VPWR.n18 VPWR.n10 33.8829
R42 VPWR.n5 VPWR.t2 31.5205
R43 VPWR.n5 VPWR.t4 31.5205
R44 VPWR.n14 VPWR.n13 27.8593
R45 VPWR.n2 VPWR.t5 27.5805
R46 VPWR.n2 VPWR.t7 27.5805
R47 VPWR.n8 VPWR.t11 27.5805
R48 VPWR.n8 VPWR.t0 27.5805
R49 VPWR.n9 VPWR.t3 26.5955
R50 VPWR.n9 VPWR.t9 26.5955
R51 VPWR.n12 VPWR.t8 26.5955
R52 VPWR.n12 VPWR.t10 26.5955
R53 VPWR.n31 VPWR.n30 24.4711
R54 VPWR.n33 VPWR.n32 22.9652
R55 VPWR.n32 VPWR.n31 19.9534
R56 VPWR.n24 VPWR.n6 12.424
R57 VPWR.n14 VPWR.n10 10.5417
R58 VPWR.n15 VPWR.n14 9.3005
R59 VPWR.n16 VPWR.n10 9.3005
R60 VPWR.n18 VPWR.n17 9.3005
R61 VPWR.n20 VPWR.n7 9.3005
R62 VPWR.n22 VPWR.n21 9.3005
R63 VPWR.n24 VPWR.n23 9.3005
R64 VPWR.n25 VPWR.n4 9.3005
R65 VPWR.n27 VPWR.n26 9.3005
R66 VPWR.n28 VPWR.n3 9.3005
R67 VPWR.n30 VPWR.n29 9.3005
R68 VPWR.n31 VPWR.n1 9.3005
R69 VPWR.n32 VPWR.n0 9.3005
R70 VPWR.n34 VPWR.n33 9.3005
R71 VPWR.n13 VPWR.n11 6.53128
R72 VPWR.n20 VPWR.n19 4.89462
R73 VPWR.n19 VPWR.n18 4.89462
R74 VPWR.n21 VPWR.n6 1.88285
R75 VPWR.n15 VPWR.n11 0.286241
R76 VPWR.n16 VPWR.n15 0.120292
R77 VPWR.n17 VPWR.n16 0.120292
R78 VPWR.n17 VPWR.n7 0.120292
R79 VPWR.n22 VPWR.n7 0.120292
R80 VPWR.n23 VPWR.n22 0.120292
R81 VPWR.n23 VPWR.n4 0.120292
R82 VPWR.n27 VPWR.n4 0.120292
R83 VPWR.n28 VPWR.n27 0.120292
R84 VPWR.n29 VPWR.n28 0.120292
R85 VPWR.n29 VPWR.n1 0.120292
R86 VPWR.n1 VPWR.n0 0.120292
R87 VPWR.n34 VPWR.n0 0.120292
R88 VPWR VPWR.n34 0.0213333
R89 VPB.t5 VPB.t2 278.193
R90 VPB.t0 VPB.t15 254.518
R91 VPB.t2 VPB.t0 254.518
R92 VPB.t3 VPB.t5 254.518
R93 VPB.t12 VPB.t3 254.518
R94 VPB.t14 VPB.t12 254.518
R95 VPB.t13 VPB.t14 254.518
R96 VPB.t6 VPB.t13 254.518
R97 VPB.t8 VPB.t6 254.518
R98 VPB.t7 VPB.t8 254.518
R99 VPB.t9 VPB.t1 248.599
R100 VPB.t11 VPB.t9 248.599
R101 VPB.t4 VPB.t11 248.599
R102 VPB.t10 VPB.t4 248.599
R103 VPB.t15 VPB.t10 248.599
R104 VPB VPB.t7 192.369
R105 A2.n2 A2.t1 196.013
R106 A2.n1 A2.t0 196.013
R107 A2.n7 A2.t5 196.013
R108 A2.n8 A2.t3 196.013
R109 A2.n4 A2.n3 168.119
R110 A2 A2.n9 157.69
R111 A2.n5 A2.n4 152
R112 A2.n6 A2.n0 152
R113 A2.n2 A2.t6 139.78
R114 A2.n1 A2.t4 139.78
R115 A2.n7 A2.t7 139.78
R116 A2.n8 A2.t2 139.78
R117 A2.n6 A2.n5 43.1268
R118 A2.n9 A2.n7 41.2242
R119 A2.n3 A2.n1 33.6137
R120 A2.n3 A2.n2 20.9294
R121 A2.n4 A2.n0 16.119
R122 A2.n9 A2.n8 13.3189
R123 A2 A2.n0 10.4301
R124 A2.n5 A2.n1 9.51366
R125 A2.n7 A2.n6 1.90313
R126 Y.n2 Y.n0 629.033
R127 Y.n2 Y.n1 585
R128 Y.n10 Y.n9 585
R129 Y.n8 Y.n7 585
R130 Y.n6 Y.n5 585
R131 Y.n4 Y.n3 585
R132 Y.n13 Y.n11 244.733
R133 Y.n13 Y.n12 185
R134 Y Y.n13 134.38
R135 Y.n4 Y.n2 81.9506
R136 Y.n6 Y.n4 43.7765
R137 Y.n10 Y.n8 43.0085
R138 Y.n8 Y.n6 43.0085
R139 Y Y.n10 28.7026
R140 Y.n3 Y.t0 27.5805
R141 Y.n3 Y.t3 27.5805
R142 Y.n0 Y.t4 27.5805
R143 Y.n0 Y.t5 27.5805
R144 Y.n1 Y.t6 27.5805
R145 Y.n1 Y.t7 27.5805
R146 Y.n5 Y.t10 26.5955
R147 Y.n5 Y.t15 26.5955
R148 Y.n7 Y.t11 26.5955
R149 Y.n7 Y.t8 26.5955
R150 Y.n9 Y.t2 26.5955
R151 Y.n9 Y.t9 26.5955
R152 Y.n11 Y.t13 24.9236
R153 Y.n11 Y.t12 24.9236
R154 Y.n12 Y.t1 24.9236
R155 Y.n12 Y.t14 24.9236
R156 B1 B1.n0 328.974
R157 B1.n0 B1.t5 241.536
R158 B1.n4 B1.t1 212.081
R159 B1.n3 B1.t3 212.081
R160 B1.n1 B1.t7 212.081
R161 B1.n0 B1.t2 169.237
R162 B1.n6 B1.n5 152
R163 B1.n4 B1.t4 139.78
R164 B1.n3 B1.t6 139.78
R165 B1.n1 B1.t0 139.78
R166 B1.n6 B1.n2 73.7757
R167 B1.n5 B1.n4 49.6611
R168 B1.n2 B1.n1 35.189
R169 B1.n4 B1.n2 20.8178
R170 B1.n5 B1.n3 13.146
R171 B1 B1.n6 0.464268
R172 a_27_47.n0 a_27_47.t11 299.728
R173 a_27_47.n0 a_27_47.t5 250.161
R174 a_27_47.n3 a_27_47.n1 241.751
R175 a_27_47.n0 a_27_47.n6 185
R176 a_27_47.n3 a_27_47.n2 185
R177 a_27_47.n5 a_27_47.n4 185
R178 a_27_47.n8 a_27_47.n7 185
R179 a_27_47.n7 a_27_47.n0 83.1624
R180 a_27_47.n5 a_27_47.n3 63.1971
R181 a_27_47.n7 a_27_47.n5 45.8672
R182 a_27_47.n2 a_27_47.t8 29.539
R183 a_27_47.n2 a_27_47.t4 27.6928
R184 a_27_47.n4 a_27_47.t1 25.8467
R185 a_27_47.n4 a_27_47.t2 25.8467
R186 a_27_47.n6 a_27_47.t7 25.8467
R187 a_27_47.n6 a_27_47.t6 25.8467
R188 a_27_47.n1 a_27_47.t10 25.8467
R189 a_27_47.n1 a_27_47.t9 25.8467
R190 a_27_47.t0 a_27_47.n8 25.8467
R191 a_27_47.n8 a_27_47.t3 25.8467
R192 a_806_47.n1 a_806_47.n0 490.534
R193 a_806_47.t2 a_806_47.n1 25.8467
R194 a_806_47.n1 a_806_47.t3 25.8467
R195 a_806_47.n0 a_806_47.t1 24.9236
R196 a_806_47.n0 a_806_47.t0 24.9236
R197 VNB.t0 VNB.t14 1338.51
R198 VNB.t5 VNB.t15 1310.03
R199 VNB.t2 VNB.t5 1253.07
R200 VNB.t13 VNB.t12 1224.6
R201 VNB.t15 VNB.t13 1224.6
R202 VNB.t3 VNB.t2 1224.6
R203 VNB.t1 VNB.t3 1224.6
R204 VNB.t4 VNB.t1 1224.6
R205 VNB.t8 VNB.t4 1224.6
R206 VNB.t7 VNB.t8 1224.6
R207 VNB.t6 VNB.t7 1224.6
R208 VNB.t11 VNB.t0 1196.12
R209 VNB.t10 VNB.t11 1196.12
R210 VNB.t9 VNB.t10 1196.12
R211 VNB.t12 VNB.t9 1196.12
R212 VNB VNB.t6 925.567
R213 VGND.n10 VGND.n1 205.707
R214 VGND.n6 VGND.n5 204.171
R215 VGND.n4 VGND.n3 198.964
R216 VGND.n13 VGND.n12 198.964
R217 VGND.n9 VGND.n2 34.6358
R218 VGND.n11 VGND.n10 30.1181
R219 VGND.n5 VGND.t4 27.6928
R220 VGND.n5 VGND.t1 25.8467
R221 VGND.n3 VGND.t2 25.8467
R222 VGND.n3 VGND.t0 25.8467
R223 VGND.n1 VGND.t3 25.8467
R224 VGND.n1 VGND.t7 25.8467
R225 VGND.n12 VGND.t6 25.8467
R226 VGND.n12 VGND.t5 25.8467
R227 VGND.n13 VGND.n11 22.2123
R228 VGND.n4 VGND.n2 13.177
R229 VGND.n7 VGND.n2 9.3005
R230 VGND.n9 VGND.n8 9.3005
R231 VGND.n11 VGND.n0 9.3005
R232 VGND.n14 VGND.n13 7.16074
R233 VGND.n6 VGND.n4 6.81482
R234 VGND.n10 VGND.n9 4.51815
R235 VGND.n7 VGND.n6 0.75671
R236 VGND.n14 VGND.n0 0.148009
R237 VGND.n8 VGND.n7 0.120292
R238 VGND.n8 VGND.n0 0.120292
R239 VGND VGND.n14 0.114057
R240 C1.n0 C1.t7 212.081
R241 C1.n4 C1.t0 212.081
R242 C1.n5 C1.t1 212.081
R243 C1.n2 C1.t2 212.081
R244 C1.n7 C1.n3 168.119
R245 C1 C1.n1 158.875
R246 C1.n7 C1.n6 152
R247 C1.n0 C1.t6 139.78
R248 C1.n4 C1.t4 139.78
R249 C1.n5 C1.t5 139.78
R250 C1.n2 C1.t3 139.78
R251 C1.n3 C1.n2 52.5823
R252 C1.n6 C1.n5 40.8975
R253 C1.n1 C1.n0 32.1338
R254 C1.n4 C1.n1 29.2126
R255 C1.n6 C1.n4 20.449
R256 C1 C1.n7 9.24494
R257 C1.n5 C1.n3 8.76414
R258 a_1314_47.t0 a_1314_47.t1 59.0774
R259 a_978_47.t0 a_978_47.t1 49.8467
C0 VPWR VPB 0.155187f
C1 VPWR VGND 0.025729f
C2 A1 VPB 0.131463f
C3 VGND A1 0.05327f
C4 Y A2 0.026527f
C5 VPWR B1 0.080681f
C6 A1 B1 0.099043f
C7 VPWR Y 0.401975f
C8 C1 VPB 0.115837f
C9 VPWR A2 0.0322f
C10 Y A1 0.170649f
C11 VGND C1 0.018441f
C12 A1 A2 0.301027f
C13 B1 C1 0.265455f
C14 VGND VPB 0.004845f
C15 B1 VPB 0.1299f
C16 VPWR A1 0.089511f
C17 Y C1 0.079193f
C18 VGND B1 0.01819f
C19 Y VPB 0.016005f
C20 Y VGND 0.155128f
C21 A2 VPB 0.116508f
C22 Y B1 0.403708f
C23 VPWR C1 0.058222f
C24 VGND A2 0.046492f
C25 VGND VNB 0.846099f
C26 Y VNB 0.08135f
C27 VPWR VNB 0.743981f
C28 C1 VNB 0.353893f
C29 B1 VNB 0.382855f
C30 A2 VNB 0.357989f
C31 A1 VNB 0.407226f
C32 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221a_1 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 a_240_47.t0 A2.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X.t1 a_51_297.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t2 A1.t0 a_240_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297.t1 B2.t0 a_245_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47.t0 C1.t0 a_51_297.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47.t2 B1.t0 a_149_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X6 VPWR.t3 A1.t1 a_512_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X.t0 a_51_297.t5 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47.t2 B2.t1 a_240_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297.t0 B1.t1 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR.t0 C1.t1 a_51_297.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297.t0 A2.t1 a_51_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
R0 A2.n0 A2.t1 233.576
R1 A2.n0 A2.t0 161.275
R2 A2 A2.n0 158.502
R3 VGND.n1 VGND.t1 298.283
R4 VGND.n1 VGND.n0 132.353
R5 VGND.n0 VGND.t0 24.9236
R6 VGND.n0 VGND.t2 24.9236
R7 VGND VGND.n1 1.04774
R8 a_240_47.n1 a_240_47.n0 368.68
R9 a_240_47.n0 a_240_47.t1 24.9236
R10 a_240_47.n0 a_240_47.t2 24.9236
R11 a_240_47.n1 a_240_47.t3 24.9236
R12 a_240_47.t0 a_240_47.n1 24.9236
R13 VNB.t2 VNB.t1 2677.02
R14 VNB VNB.t3 1495.15
R15 VNB.t3 VNB.t4 1295.79
R16 VNB.t5 VNB.t0 1196.12
R17 VNB.t1 VNB.t5 1196.12
R18 VNB.t4 VNB.t2 1196.12
R19 a_51_297.n3 a_51_297.n0 292.5
R20 a_51_297.n5 a_51_297.n4 292.5
R21 a_51_297.n4 a_51_297.n1 266.349
R22 a_51_297.n2 a_51_297.t3 243.661
R23 a_51_297.n1 a_51_297.t5 234.483
R24 a_51_297.n2 a_51_297.t2 184.224
R25 a_51_297.n1 a_51_297.t4 162.184
R26 a_51_297.n5 a_51_297.n0 109.335
R27 a_51_297.n3 a_51_297.n2 90.111
R28 a_51_297.t0 a_51_297.n5 26.5955
R29 a_51_297.n0 a_51_297.t1 26.5955
R30 a_51_297.n4 a_51_297.n3 12.0412
R31 X.n0 X.t0 326.3
R32 X X.t1 178.826
R33 X.n0 X 4.6085
R34 X X.n0 1.73283
R35 A1.n0 A1.t1 241.536
R36 A1.n0 A1.t0 169.237
R37 A1 A1.n0 153.565
R38 B2.n0 B2.t0 234.804
R39 B2.n0 B2.t1 162.504
R40 B2.n1 B2.n0 152
R41 B2 B2.n1 11.4005
R42 B2.n1 B2 2.2005
R43 a_245_297.t0 a_245_297.t1 41.3705
R44 VPB.t3 VPB.t1 577.104
R45 VPB VPB.t2 310.748
R46 VPB.t5 VPB.t4 284.113
R47 VPB.t2 VPB.t0 284.113
R48 VPB.t1 VPB.t5 213.084
R49 VPB.t0 VPB.t3 213.084
R50 C1 C1.n0 217.981
R51 C1.n0 C1.t1 212.081
R52 C1.n0 C1.t0 139.78
R53 a_149_47.n0 a_149_47.t2 512.086
R54 a_149_47.t0 a_149_47.n0 30.462
R55 a_149_47.n0 a_149_47.t1 25.8467
R56 B1.n0 B1.t1 241.536
R57 B1.n0 B1.t0 169.237
R58 B1 B1.n0 154.133
R59 a_512_297.t0 a_512_297.t1 41.3705
R60 VPWR.n2 VPWR.n0 325.372
R61 VPWR.n2 VPWR.n1 318.245
R62 VPWR.n1 VPWR.t2 38.4155
R63 VPWR.n0 VPWR.t1 34.4755
R64 VPWR.n0 VPWR.t0 30.5355
R65 VPWR.n1 VPWR.t3 26.5955
R66 VPWR VPWR.n2 0.184733
C0 B2 B1 0.079688f
C1 A1 VPB 0.02547f
C2 VPB C1 0.05148f
C3 B2 X 1.41e-19
C4 A2 VPWR 0.015093f
C5 VPWR VPB 0.087901f
C6 A2 VPB 0.038559f
C7 VGND B1 0.007938f
C8 B2 VPWR 0.013541f
C9 X VGND 0.143614f
C10 B2 A2 0.074588f
C11 A1 VGND 0.027709f
C12 B2 VPB 0.036569f
C13 X B1 8.13e-20
C14 VGND C1 0.014106f
C15 C1 B1 0.051961f
C16 VPWR VGND 0.079939f
C17 A2 VGND 0.015861f
C18 A1 X 9.4e-19
C19 VGND VPB 0.00816f
C20 VPWR B1 0.011497f
C21 VPB B1 0.025127f
C22 VPWR X 0.143364f
C23 A2 X 3.43e-19
C24 A1 VPWR 0.021536f
C25 B2 VGND 0.010662f
C26 VPWR C1 0.020061f
C27 X VPB 0.026158f
C28 A2 A1 0.080079f
C29 VGND VNB 0.493685f
C30 X VNB 0.106807f
C31 VPWR VNB 0.408842f
C32 A1 VNB 0.090821f
C33 A2 VNB 0.106876f
C34 B2 VNB 0.103396f
C35 B1 VNB 0.089709f
C36 C1 VNB 0.163785f
C37 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221a_2 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 VPWR.t3 a_38_47.t4 X.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t0 A1.t0 a_497_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X.t1 a_38_47.t5 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47.t2 B2.t0 a_225_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_497_297.t0 A2.t0 a_38_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3875 ps=1.775 w=1 l=0.15
X5 VGND.t3 A1.t1 a_225_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t1 C1.t0 a_38_47.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297.t0 B1.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47.t2 B2.t1 a_237_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3875 pd=1.775 as=0.1125 ps=1.225 w=1 l=0.15
X9 a_225_47.t1 A2.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X.t0 a_38_47.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_141_47.t1 C1.t1 a_38_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23725 ps=2.03 w=0.65 l=0.15
X12 VGND.t1 a_38_47.t7 X.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_225_47.t0 B1.t1 a_141_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_38_47.n5 a_38_47.n0 292.5
R1 a_38_47.n7 a_38_47.n6 292.5
R2 a_38_47.n4 a_38_47.t1 273.132
R3 a_38_47.n6 a_38_47.n3 267.926
R4 a_38_47.n4 a_38_47.t3 266.959
R5 a_38_47.n1 a_38_47.t4 212.081
R6 a_38_47.n2 a_38_47.t5 212.081
R7 a_38_47.n1 a_38_47.t7 139.78
R8 a_38_47.n2 a_38_47.t6 139.78
R9 a_38_47.n7 a_38_47.n0 99.4855
R10 a_38_47.n5 a_38_47.n4 64.2205
R11 a_38_47.n3 a_38_47.n1 37.9763
R12 a_38_47.t0 a_38_47.n7 26.5955
R13 a_38_47.n0 a_38_47.t2 26.5955
R14 a_38_47.n3 a_38_47.n2 23.3702
R15 a_38_47.n6 a_38_47.n5 10.9564
R16 X X.n0 319.075
R17 X X.n1 148.056
R18 X.n0 X.t2 26.5955
R19 X.n0 X.t1 26.5955
R20 X.n1 X.t3 24.9236
R21 X.n1 X.t0 24.9236
R22 VPWR.n3 VPWR.t3 846.052
R23 VPWR.n12 VPWR.n1 316.432
R24 VPWR.n5 VPWR.n4 312.053
R25 VPWR.n4 VPWR.t2 38.4155
R26 VPWR.n6 VPWR.n2 34.6358
R27 VPWR.n10 VPWR.n2 34.6358
R28 VPWR.n11 VPWR.n10 34.6358
R29 VPWR.n1 VPWR.t1 33.4905
R30 VPWR.n1 VPWR.t4 31.5205
R31 VPWR.n4 VPWR.t0 26.5955
R32 VPWR.n6 VPWR.n5 19.9534
R33 VPWR.n13 VPWR.n12 12.1767
R34 VPWR.n12 VPWR.n11 12.0476
R35 VPWR.n7 VPWR.n6 9.3005
R36 VPWR.n8 VPWR.n2 9.3005
R37 VPWR.n10 VPWR.n9 9.3005
R38 VPWR.n11 VPWR.n0 9.3005
R39 VPWR.n5 VPWR.n3 6.64746
R40 VPWR.n7 VPWR.n3 0.662502
R41 VPWR.n13 VPWR.n0 0.141672
R42 VPWR VPWR.n13 0.12308
R43 VPWR.n8 VPWR.n7 0.120292
R44 VPWR.n9 VPWR.n8 0.120292
R45 VPWR.n9 VPWR.n0 0.120292
R46 VPB.t2 VPB.t0 547.509
R47 VPB VPB.t3 290.031
R48 VPB.t1 VPB.t4 284.113
R49 VPB.t3 VPB.t6 284.113
R50 VPB.t4 VPB.t5 248.599
R51 VPB.t6 VPB.t2 221.964
R52 VPB.t0 VPB.t1 213.084
R53 A1.n0 A1.t0 241.536
R54 A1.n0 A1.t1 169.237
R55 A1 A1.n0 156.268
R56 a_497_297.t0 a_497_297.t1 41.3705
R57 B2.n0 B2.t1 233.869
R58 B2.n0 B2.t0 161.57
R59 B2.n1 B2.n0 152
R60 B2.n1 B2 12.5798
R61 B2 B2.n1 2.42809
R62 a_225_47.n1 a_225_47.n0 368.68
R63 a_225_47.n0 a_225_47.t2 24.9236
R64 a_225_47.n0 a_225_47.t1 24.9236
R65 a_225_47.n1 a_225_47.t3 24.9236
R66 a_225_47.t0 a_225_47.n1 24.9236
R67 a_141_47.n0 a_141_47.t2 516.324
R68 a_141_47.t0 a_141_47.n0 24.9236
R69 a_141_47.n0 a_141_47.t1 24.9236
R70 VNB.t6 VNB.t1 2677.02
R71 VNB VNB.t2 1452.43
R72 VNB.t4 VNB.t3 1196.12
R73 VNB.t5 VNB.t4 1196.12
R74 VNB.t1 VNB.t5 1196.12
R75 VNB.t0 VNB.t6 1196.12
R76 VNB.t2 VNB.t0 1196.12
R77 A2.n0 A2.t0 233.576
R78 A2.n0 A2.t1 161.275
R79 A2.n1 A2.n0 152
R80 A2.n1 A2 11.9612
R81 A2 A2.n1 2.3087
R82 VGND.n3 VGND.t1 293.514
R83 VGND.n0 VGND.t0 286.426
R84 VGND.n4 VGND.n2 121.451
R85 VGND.n4 VGND.n3 36.5149
R86 VGND.n6 VGND.n5 34.6358
R87 VGND.n2 VGND.t2 24.9236
R88 VGND.n2 VGND.t3 24.9236
R89 VGND.n6 VGND.n0 24.8476
R90 VGND.n8 VGND.n0 17.3894
R91 VGND.n5 VGND.n1 9.3005
R92 VGND.n7 VGND.n6 9.3005
R93 VGND.n5 VGND.n4 3.76521
R94 VGND.n3 VGND.n1 2.15642
R95 VGND VGND.n8 0.48397
R96 VGND.n8 VGND.n7 0.147154
R97 VGND.n7 VGND.n1 0.120292
R98 C1.n0 C1.t0 212.081
R99 C1 C1.n0 208.075
R100 C1.n0 C1.t1 133.353
R101 B1.n0 B1.t0 241.536
R102 B1.n0 B1.t1 169.237
R103 B1 B1.n0 154.042
R104 a_237_297.t0 a_237_297.t1 44.3255
C0 VPWR X 0.162381f
C1 B2 X 1.47e-19
C2 A2 VPWR 0.016485f
C3 VPWR C1 0.018502f
C4 X VPB 0.009512f
C5 B2 A2 0.076479f
C6 A2 VPB 0.037893f
C7 VPB C1 0.048821f
C8 B2 VPWR 0.015192f
C9 VPWR VPB 0.087549f
C10 B2 VPB 0.037167f
C11 A1 VGND 0.031803f
C12 VGND B1 0.008841f
C13 X VGND 0.156731f
C14 A2 VGND 0.017441f
C15 A1 X 9.18e-19
C16 X B1 8.17e-20
C17 VGND C1 0.012628f
C18 A2 A1 0.080308f
C19 C1 B1 0.053585f
C20 VPWR VGND 0.081242f
C21 A2 X 3.36e-19
C22 A1 VPWR 0.021111f
C23 B2 VGND 0.011586f
C24 VPWR B1 0.015821f
C25 VGND VPB 0.007384f
C26 A1 VPB 0.025441f
C27 B2 B1 0.077957f
C28 VPB B1 0.0254f
C29 VGND VNB 0.503191f
C30 X VNB 0.07188f
C31 VPWR VNB 0.413944f
C32 A1 VNB 0.090746f
C33 A2 VNB 0.105707f
C34 B2 VNB 0.104083f
C35 B1 VNB 0.089083f
C36 C1 VNB 0.161446f
C37 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221a_4 VNB VPB VGND VPWR B1 B2 A2 A1 X C1
X0 a_27_47.t3 B1.t0 a_277_47.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_109_47.t6 A2.t0 a_717_297.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_717_297.t1 A1.t0 VPWR.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3 VGND.t7 A2.t1 a_277_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_277_297.t3 B2.t0 a_109_47.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_47.t0 B2.t1 a_277_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t6 a_109_47.t8 X.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t7 a_109_47.t9 VGND.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_277_297.t1 B1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t2 a_109_47.t10 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_277_47.t5 A1.t1 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_277_47.t7 A2.t2 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t6 a_109_47.t11 VGND.t2 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR.t9 C1.t0 a_109_47.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_47.t1 C1.t1 a_109_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_27_47.t4 B2.t2 a_277_47.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t5 a_109_47.t12 X.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t0 A1.t2 a_277_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t4 a_109_47.t13 X.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_277_47.t3 B1.t2 a_27_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_277_47.t0 B2.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR.t8 a_109_47.t14 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t3 B1.t3 a_277_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X23 X.t0 a_109_47.t15 VPWR.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t0 A1.t3 a_717_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_109_47.t2 C1.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_717_297.t2 A2.t3 a_109_47.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_109_47.t7 C1.t3 a_27_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n1 B1.t1 241.536
R1 B1.n0 B1.t3 241.536
R2 B1.n2 B1.n0 238.719
R3 B1.n1 B1.t2 169.237
R4 B1.n0 B1.t0 169.237
R5 B1.n2 B1.n1 152
R6 B1 B1.n2 5.68939
R7 a_277_47.n4 a_277_47.n3 226.355
R8 a_277_47.n5 a_277_47.n4 185
R9 a_277_47.n2 a_277_47.n0 135.442
R10 a_277_47.n2 a_277_47.n1 97.6244
R11 a_277_47.n4 a_277_47.n2 77.3317
R12 a_277_47.n3 a_277_47.t6 24.9236
R13 a_277_47.n3 a_277_47.t3 24.9236
R14 a_277_47.n1 a_277_47.t1 24.9236
R15 a_277_47.n1 a_277_47.t5 24.9236
R16 a_277_47.n0 a_277_47.t2 24.9236
R17 a_277_47.n0 a_277_47.t7 24.9236
R18 a_277_47.n5 a_277_47.t4 24.9236
R19 a_277_47.t0 a_277_47.n5 24.9236
R20 a_27_47.t3 a_27_47.n3 316.95
R21 a_27_47.n3 a_27_47.n2 185
R22 a_27_47.n1 a_27_47.t5 180.946
R23 a_27_47.n1 a_27_47.n0 97.0637
R24 a_27_47.n3 a_27_47.n1 48.8732
R25 a_27_47.n0 a_27_47.t2 24.9236
R26 a_27_47.n0 a_27_47.t1 24.9236
R27 a_27_47.n2 a_27_47.t0 24.9236
R28 a_27_47.n2 a_27_47.t4 24.9236
R29 VNB.t5 VNB.t6 2677.02
R30 VNB.t12 VNB.t8 1196.12
R31 VNB.t7 VNB.t12 1196.12
R32 VNB.t11 VNB.t7 1196.12
R33 VNB.t2 VNB.t11 1196.12
R34 VNB.t10 VNB.t2 1196.12
R35 VNB.t1 VNB.t10 1196.12
R36 VNB.t6 VNB.t1 1196.12
R37 VNB.t0 VNB.t5 1196.12
R38 VNB.t9 VNB.t0 1196.12
R39 VNB.t4 VNB.t9 1196.12
R40 VNB.t3 VNB.t4 1196.12
R41 VNB.t13 VNB.t3 1196.12
R42 VNB VNB.t13 911.327
R43 A2.n0 A2.t3 212.081
R44 A2.n1 A2.t0 212.081
R45 A2 A2.n2 171.201
R46 A2.n0 A2.t2 139.78
R47 A2.n1 A2.t1 139.78
R48 A2.n2 A2.n0 30.6732
R49 A2.n2 A2.n1 30.6732
R50 a_717_297.n1 a_717_297.n0 1223.84
R51 a_717_297.n0 a_717_297.t3 26.5955
R52 a_717_297.n0 a_717_297.t1 26.5955
R53 a_717_297.t0 a_717_297.n1 26.5955
R54 a_717_297.n1 a_717_297.t2 26.5955
R55 a_109_47.n13 a_109_47.n12 585
R56 a_109_47.n15 a_109_47.n14 585
R57 a_109_47.n11 a_109_47.n10 239.397
R58 a_109_47.n1 a_109_47.t8 212.081
R59 a_109_47.n3 a_109_47.t10 212.081
R60 a_109_47.n5 a_109_47.t14 212.081
R61 a_109_47.n6 a_109_47.t15 212.081
R62 a_109_47.n11 a_109_47.n9 196.181
R63 a_109_47.n2 a_109_47.n0 180.8
R64 a_109_47.n14 a_109_47.n13 155.859
R65 a_109_47.n8 a_109_47.n7 152
R66 a_109_47.n4 a_109_47.n0 152
R67 a_109_47.n1 a_109_47.t13 139.78
R68 a_109_47.n3 a_109_47.t11 139.78
R69 a_109_47.n5 a_109_47.t12 139.78
R70 a_109_47.n6 a_109_47.t9 139.78
R71 a_109_47.n14 a_109_47.n8 114.522
R72 a_109_47.n13 a_109_47.n11 81.9512
R73 a_109_47.n4 a_109_47.n3 35.055
R74 a_109_47.n2 a_109_47.n1 30.6732
R75 a_109_47.n3 a_109_47.n2 30.6732
R76 a_109_47.n7 a_109_47.n5 30.6732
R77 a_109_47.n7 a_109_47.n6 30.6732
R78 a_109_47.n12 a_109_47.t4 26.5955
R79 a_109_47.n12 a_109_47.t0 26.5955
R80 a_109_47.n9 a_109_47.t3 26.5955
R81 a_109_47.n9 a_109_47.t2 26.5955
R82 a_109_47.n15 a_109_47.t5 26.5955
R83 a_109_47.t6 a_109_47.n15 26.5955
R84 a_109_47.n5 a_109_47.n4 26.2914
R85 a_109_47.n8 a_109_47.n0 24.9605
R86 a_109_47.n10 a_109_47.t1 24.9236
R87 a_109_47.n10 a_109_47.t7 24.9236
R88 VPB.t2 VPB.t9 556.386
R89 VPB.t7 VPB.t8 248.599
R90 VPB.t6 VPB.t7 248.599
R91 VPB.t5 VPB.t6 248.599
R92 VPB.t1 VPB.t5 248.599
R93 VPB.t12 VPB.t1 248.599
R94 VPB.t13 VPB.t12 248.599
R95 VPB.t9 VPB.t13 248.599
R96 VPB.t11 VPB.t2 248.599
R97 VPB.t0 VPB.t11 248.599
R98 VPB.t3 VPB.t0 248.599
R99 VPB.t10 VPB.t3 248.599
R100 VPB.t4 VPB.t10 248.599
R101 VPB VPB.t4 189.409
R102 A1.n3 A1.n0 247.34
R103 A1.n1 A1.t3 241.536
R104 A1.n0 A1.t0 240.484
R105 A1.n1 A1.t2 169.237
R106 A1.n0 A1.t1 168.185
R107 A1.n2 A1.n1 152
R108 A1 A1.n3 3.44665
R109 A1.n2 A1 2.8165
R110 A1.n3 A1.n2 0.7685
R111 VPWR.n30 VPWR.n2 606.505
R112 VPWR.n14 VPWR.n8 606.505
R113 VPWR.n10 VPWR.n9 606.505
R114 VPWR.n24 VPWR.n23 585
R115 VPWR.n22 VPWR.n21 585
R116 VPWR.n11 VPWR.t6 350.587
R117 VPWR.n32 VPWR.t4 250.975
R118 VPWR.n23 VPWR.n22 100.471
R119 VPWR.n25 VPWR.n3 34.6358
R120 VPWR.n29 VPWR.n3 34.6358
R121 VPWR.n16 VPWR.n15 34.6358
R122 VPWR.n16 VPWR.n6 34.6358
R123 VPWR.n20 VPWR.n6 34.6358
R124 VPWR.n13 VPWR.n10 30.4946
R125 VPWR.n23 VPWR.t3 28.5655
R126 VPWR.n30 VPWR.n29 28.2358
R127 VPWR.n22 VPWR.t1 26.5955
R128 VPWR.n2 VPWR.t2 26.5955
R129 VPWR.n2 VPWR.t9 26.5955
R130 VPWR.n8 VPWR.t7 26.5955
R131 VPWR.n8 VPWR.t0 26.5955
R132 VPWR.n9 VPWR.t5 26.5955
R133 VPWR.n9 VPWR.t8 26.5955
R134 VPWR.n31 VPWR.n30 22.2123
R135 VPWR.n32 VPWR.n31 22.2123
R136 VPWR.n14 VPWR.n13 13.9299
R137 VPWR.n25 VPWR.n24 12.5181
R138 VPWR.n13 VPWR.n12 9.3005
R139 VPWR.n15 VPWR.n7 9.3005
R140 VPWR.n17 VPWR.n16 9.3005
R141 VPWR.n18 VPWR.n6 9.3005
R142 VPWR.n20 VPWR.n19 9.3005
R143 VPWR.n5 VPWR.n4 9.3005
R144 VPWR.n26 VPWR.n25 9.3005
R145 VPWR.n27 VPWR.n3 9.3005
R146 VPWR.n29 VPWR.n28 9.3005
R147 VPWR.n30 VPWR.n1 9.3005
R148 VPWR.n31 VPWR.n0 9.3005
R149 VPWR.n33 VPWR.n32 9.3005
R150 VPWR.n11 VPWR.n10 6.47684
R151 VPWR.n21 VPWR.n5 5.83579
R152 VPWR.n21 VPWR.n20 4.23579
R153 VPWR.n24 VPWR.n5 3.76521
R154 VPWR.n15 VPWR.n14 1.88285
R155 VPWR.n12 VPWR.n11 0.58037
R156 VPWR.n12 VPWR.n7 0.120292
R157 VPWR.n17 VPWR.n7 0.120292
R158 VPWR.n18 VPWR.n17 0.120292
R159 VPWR.n19 VPWR.n18 0.120292
R160 VPWR.n19 VPWR.n4 0.120292
R161 VPWR.n26 VPWR.n4 0.120292
R162 VPWR.n27 VPWR.n26 0.120292
R163 VPWR.n28 VPWR.n27 0.120292
R164 VPWR.n28 VPWR.n1 0.120292
R165 VPWR.n1 VPWR.n0 0.120292
R166 VPWR.n33 VPWR.n0 0.120292
R167 VPWR VPWR.n33 0.0213333
R168 VGND.n0 VGND.t1 288.344
R169 VGND.n6 VGND.t4 287.603
R170 VGND.n7 VGND.n5 207.965
R171 VGND.n16 VGND.n2 207.965
R172 VGND.n10 VGND.n9 121.451
R173 VGND.n7 VGND.n6 35.1602
R174 VGND.n11 VGND.n8 34.6358
R175 VGND.n15 VGND.n3 34.6358
R176 VGND.n18 VGND.n17 34.6358
R177 VGND.n5 VGND.t2 24.9236
R178 VGND.n5 VGND.t5 24.9236
R179 VGND.n9 VGND.t3 24.9236
R180 VGND.n9 VGND.t0 24.9236
R181 VGND.n2 VGND.t6 24.9236
R182 VGND.n2 VGND.t7 24.9236
R183 VGND.n11 VGND.n10 23.3417
R184 VGND.n20 VGND.n0 19.2717
R185 VGND.n16 VGND.n15 17.3181
R186 VGND.n17 VGND.n16 17.3181
R187 VGND.n10 VGND.n3 11.2946
R188 VGND.n8 VGND.n4 9.3005
R189 VGND.n12 VGND.n11 9.3005
R190 VGND.n13 VGND.n3 9.3005
R191 VGND.n15 VGND.n14 9.3005
R192 VGND.n17 VGND.n1 9.3005
R193 VGND.n19 VGND.n18 9.3005
R194 VGND.n8 VGND.n7 5.27109
R195 VGND.n18 VGND.n0 4.89462
R196 VGND.n6 VGND.n4 1.66544
R197 VGND VGND.n20 0.716876
R198 VGND.n20 VGND.n19 0.147186
R199 VGND.n12 VGND.n4 0.120292
R200 VGND.n13 VGND.n12 0.120292
R201 VGND.n14 VGND.n13 0.120292
R202 VGND.n14 VGND.n1 0.120292
R203 VGND.n19 VGND.n1 0.120292
R204 B2.n0 B2.t0 212.081
R205 B2.n1 B2.t1 212.081
R206 B2 B2.n2 153.268
R207 B2.n0 B2.t3 139.78
R208 B2.n1 B2.t2 139.78
R209 B2.n2 B2.n0 30.6732
R210 B2.n2 B2.n1 30.6732
R211 a_277_297.n1 a_277_297.n0 1223.84
R212 a_277_297.n0 a_277_297.t0 26.5955
R213 a_277_297.n0 a_277_297.t3 26.5955
R214 a_277_297.n1 a_277_297.t2 26.5955
R215 a_277_297.t1 a_277_297.n1 26.5955
R216 X.n2 X.n0 360.301
R217 X.n2 X.n1 209.019
R218 X.n5 X.n3 135.249
R219 X.n5 X.n4 98.982
R220 X X.n5 36.1828
R221 X.n0 X.t1 26.5955
R222 X.n0 X.t0 26.5955
R223 X.n1 X.t3 26.5955
R224 X.n1 X.t2 26.5955
R225 X.n4 X.t4 24.9236
R226 X.n4 X.t6 24.9236
R227 X.n3 X.t5 24.9236
R228 X.n3 X.t7 24.9236
R229 X X.n2 18.9659
R230 C1.n0 C1.t0 212.081
R231 C1.n1 C1.t2 212.081
R232 C1 C1.n1 188.482
R233 C1.n0 C1.t1 139.78
R234 C1.n1 C1.t3 139.78
R235 C1.n1 C1.n0 61.346
C0 X VGND 0.297471f
C1 A2 VGND 0.022269f
C2 VPWR X 0.282599f
C3 A2 VPWR 0.014879f
C4 B2 VPB 0.051039f
C5 X B1 5.98e-20
C6 VGND C1 0.018754f
C7 VPWR C1 0.070491f
C8 C1 B1 0.062343f
C9 A2 X 3.82e-19
C10 A1 VGND 0.047133f
C11 A1 VPWR 0.043297f
C12 VGND VPB 0.013412f
C13 X C1 1.1e-20
C14 VPWR VPB 0.166158f
C15 A1 B1 0.056711f
C16 VPB B1 0.064515f
C17 B2 VGND 0.014797f
C18 A1 X 6.02e-19
C19 B2 VPWR 0.015813f
C20 A1 A2 0.210871f
C21 X VPB 0.016561f
C22 B2 B1 0.211961f
C23 A2 VPB 0.051257f
C24 VPB C1 0.069275f
C25 B2 X 5.87e-20
C26 VPWR VGND 0.148875f
C27 A1 VPB 0.067079f
C28 VGND B1 0.021015f
C29 VPWR B1 0.041286f
C30 VGND VNB 0.833326f
C31 X VNB 0.05941f
C32 VPWR VNB 0.719616f
C33 A2 VNB 0.168119f
C34 A1 VNB 0.196777f
C35 B2 VNB 0.166669f
C36 B1 VNB 0.191173f
C37 C1 VNB 0.230737f
C38 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221ai_1 VPB VNB VGND VPWR A1 A2 Y B2 C1 B1
X0 a_109_47.t2 B1.t0 a_213_123.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1652 ps=1.82 w=0.65 l=0.15
X1 Y.t3 B2.t0 a_295_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR.t1 A1.t0 a_493_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123.t0 B2.t1 a_109_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_295_297.t1 B1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297.t1 A2.t0 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR.t0 C1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND.t1 A2.t1 a_213_123.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123.t3 A1.t1 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_47.t0 C1.t1 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n0 B1.t1 235.471
R1 B1.n0 B1.t0 163.172
R2 B1 B1.n0 159.952
R3 a_213_123.n0 a_213_123.t1 272.211
R4 a_213_123.n0 a_213_123.t3 214.433
R5 a_213_123.n1 a_213_123.n0 185
R6 a_213_123.n1 a_213_123.t2 41.539
R7 a_213_123.t0 a_213_123.n1 24.9236
R8 a_109_47.t0 a_109_47.n0 456.844
R9 a_109_47.n1 a_109_47.t0 69.6005
R10 a_109_47.n0 a_109_47.t1 24.9236
R11 a_109_47.n0 a_109_47.t2 24.9236
R12 VNB.t0 VNB.t2 2648.54
R13 VNB.t1 VNB.t3 1452.43
R14 VNB.t3 VNB.t4 1196.12
R15 VNB.t2 VNB.t1 1196.12
R16 VNB VNB.t0 925.567
R17 B2.n0 B2.t0 241.536
R18 B2.n0 B2.t1 169.237
R19 B2 B2.n0 157.625
R20 a_295_297.t0 a_295_297.t1 47.2805
R21 Y.n0 Y 590.396
R22 Y.n1 Y.n0 291.928
R23 Y.n2 Y.t1 284.892
R24 Y.n2 Y.t0 253.489
R25 Y Y.n2 69.5598
R26 Y.n0 Y.t2 62.0555
R27 Y.n0 Y.t3 26.5955
R28 Y.n1 Y 5.81687
R29 Y Y.n1 2.69376
R30 VPB.t0 VPB.t3 538.63
R31 VPB.t2 VPB.t1 355.14
R32 VPB.t3 VPB.t2 230.841
R33 VPB.t1 VPB.t4 213.084
R34 VPB VPB.t0 204.207
R35 A1.n0 A1.t0 230.793
R36 A1.n0 A1.t1 158.494
R37 A1 A1.n0 153.53
R38 a_493_297.t0 a_493_297.t1 41.3705
R39 VPWR.n6 VPWR.n5 292.5
R40 VPWR.n4 VPWR.n3 292.5
R41 VPWR.n2 VPWR.t1 256.861
R42 VPWR.n5 VPWR.n4 90.6205
R43 VPWR.n3 VPWR.n2 30.1383
R44 VPWR.n4 VPWR.t2 29.5505
R45 VPWR.n5 VPWR.t0 29.5505
R46 VPWR.n1 VPWR.n0 9.3005
R47 VPWR.n7 VPWR.n6 7.68705
R48 VPWR.n6 VPWR.n1 5.9876
R49 VPWR.n3 VPWR.n1 0.344586
R50 VPWR.n2 VPWR.n0 0.210154
R51 VPWR.n7 VPWR.n0 0.145692
R52 VPWR VPWR.n7 0.117706
R53 A2.n0 A2.t0 241.536
R54 A2 A2.n0 192.534
R55 A2.n0 A2.t1 169.237
R56 C1.n0 C1.t0 236.934
R57 C1.n0 C1.t1 205.732
R58 C1 C1.n0 161.115
R59 VGND VGND.n0 213.309
R60 VGND.n0 VGND.t0 24.9236
R61 VGND.n0 VGND.t1 24.9236
C0 Y VPWR 0.292519f
C1 VPWR B2 0.008984f
C2 Y A2 0.080476f
C3 VPWR VPB 0.074602f
C4 Y C1 0.126655f
C5 B2 A2 0.066576f
C6 A2 VPB 0.032767f
C7 VPB C1 0.037968f
C8 Y B2 0.056881f
C9 Y VPB 0.020462f
C10 B2 VPB 0.027955f
C11 VGND A1 0.015109f
C12 VGND B1 0.010639f
C13 VPWR VGND 0.064475f
C14 VPWR A1 0.050257f
C15 VGND A2 0.016249f
C16 VGND C1 0.012757f
C17 VPWR B1 0.022234f
C18 A2 A1 0.089072f
C19 A2 B1 4.14e-19
C20 C1 B1 0.020871f
C21 Y VGND 0.045954f
C22 Y A1 3.82e-19
C23 VGND B2 0.011888f
C24 VPWR A2 0.115352f
C25 VGND VPB 0.006297f
C26 VPWR C1 0.021252f
C27 Y B1 0.076802f
C28 B2 A1 5.58e-19
C29 A1 VPB 0.03588f
C30 B2 B1 0.086799f
C31 VPB B1 0.034122f
C32 VGND VNB 0.390249f
C33 VPWR VNB 0.36154f
C34 Y VNB 0.085827f
C35 A1 VNB 0.139681f
C36 A2 VNB 0.096712f
C37 B2 VNB 0.093331f
C38 B1 VNB 0.105928f
C39 C1 VNB 0.144797f
C40 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221ai_2 VNB VPB VGND VPWR Y B1 B2 A2 A1 C1
X0 Y.t5 A2.t0 a_734_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_300_47.t1 B2.t0 a_28_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t3 C1.t0 VPWR.t5 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_300_47.t3 B1.t0 a_28_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_300_47.t6 A2.t1 VGND.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_300_47.t4 A1.t0 VGND.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_734_297.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7 a_28_47.t0 C1.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t1 C1.t2 a_28_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR.t4 C1.t3 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t2 B1.t1 a_382_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X11 a_382_297.t1 B2.t1 Y.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_28_47.t4 B1.t2 a_300_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_28_47.t2 B2.t2 a_300_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t3 A1.t2 a_300_47.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15 Y.t7 B2.t3 a_382_297.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR.t3 A1.t3 a_734_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t1 A2.t2 a_300_47.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_382_297.t2 B1.t3 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X19 a_734_297.t1 A2.t3 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A2.n0 A2.t3 212.081
R1 A2.n1 A2.t0 212.081
R2 A2 A2.n2 157.12
R3 A2.n0 A2.t2 139.78
R4 A2.n1 A2.t1 139.78
R5 A2.n2 A2.n0 30.6732
R6 A2.n2 A2.n1 30.6732
R7 a_734_297.n1 a_734_297.n0 935.015
R8 a_734_297.n0 a_734_297.t3 26.5955
R9 a_734_297.n0 a_734_297.t1 26.5955
R10 a_734_297.n1 a_734_297.t2 26.5955
R11 a_734_297.t0 a_734_297.n1 26.5955
R12 Y.n2 Y.n0 708.106
R13 Y.n2 Y.n1 585
R14 Y.n5 Y.n4 237.278
R15 Y.n5 Y.n3 196.209
R16 Y Y.n2 64.5652
R17 Y Y.n5 56.0314
R18 Y.n3 Y.t2 26.5955
R19 Y.n3 Y.t3 26.5955
R20 Y.n1 Y.t6 26.5955
R21 Y.n1 Y.t7 26.5955
R22 Y.n0 Y.t4 26.5955
R23 Y.n0 Y.t5 26.5955
R24 Y.n4 Y.t0 24.9236
R25 Y.n4 Y.t1 24.9236
R26 VPB.t1 VPB.t3 556.386
R27 VPB.t4 VPB.t0 295.95
R28 VPB.t5 VPB.t7 248.599
R29 VPB.t6 VPB.t5 248.599
R30 VPB.t0 VPB.t6 248.599
R31 VPB.t8 VPB.t4 248.599
R32 VPB.t9 VPB.t8 248.599
R33 VPB.t3 VPB.t9 248.599
R34 VPB.t2 VPB.t1 248.599
R35 VPB VPB.t2 195.327
R36 B2.n0 B2.t1 212.081
R37 B2.n1 B2.t3 212.081
R38 B2 B2.n2 153.268
R39 B2.n0 B2.t2 139.78
R40 B2.n1 B2.t0 139.78
R41 B2.n2 B2.n0 30.6732
R42 B2.n2 B2.n1 30.6732
R43 a_28_47.t0 a_28_47.n3 265.432
R44 a_28_47.t0 a_28_47.n4 263.462
R45 a_28_47.n2 a_28_47.n0 226.355
R46 a_28_47.n2 a_28_47.n1 185
R47 a_28_47.n4 a_28_47.t1 177.487
R48 a_28_47.n3 a_28_47.n2 44.3082
R49 a_28_47.n1 a_28_47.t3 24.9236
R50 a_28_47.n1 a_28_47.t4 24.9236
R51 a_28_47.n0 a_28_47.t5 24.9236
R52 a_28_47.n0 a_28_47.t2 24.9236
R53 a_28_47.n4 a_28_47.n3 13.0565
R54 a_300_47.n4 a_300_47.t2 312.334
R55 a_300_47.n5 a_300_47.n4 185
R56 a_300_47.n1 a_300_47.t4 174.512
R57 a_300_47.n1 a_300_47.n0 98.982
R58 a_300_47.n3 a_300_47.n2 89.3175
R59 a_300_47.n4 a_300_47.n3 51.265
R60 a_300_47.n3 a_300_47.n1 48.4528
R61 a_300_47.n2 a_300_47.t3 33.2313
R62 a_300_47.n2 a_300_47.t7 31.3851
R63 a_300_47.n0 a_300_47.t5 24.9236
R64 a_300_47.n0 a_300_47.t6 24.9236
R65 a_300_47.n5 a_300_47.t0 24.9236
R66 a_300_47.t1 a_300_47.n5 24.9236
R67 VNB.t0 VNB.t4 2677.02
R68 VNB.t5 VNB.t9 1423.95
R69 VNB.t7 VNB.t6 1196.12
R70 VNB.t8 VNB.t7 1196.12
R71 VNB.t9 VNB.t8 1196.12
R72 VNB.t2 VNB.t5 1196.12
R73 VNB.t3 VNB.t2 1196.12
R74 VNB.t4 VNB.t3 1196.12
R75 VNB.t1 VNB.t0 1196.12
R76 VNB VNB.t1 939.807
R77 C1.n0 C1.t3 212.081
R78 C1.n1 C1.t0 212.081
R79 C1 C1.n1 189.942
R80 C1.n0 C1.t1 139.78
R81 C1.n1 C1.t2 139.78
R82 C1.n1 C1.n0 61.346
R83 VPWR.n6 VPWR.n5 601.292
R84 VPWR.n17 VPWR.n16 585
R85 VPWR.n15 VPWR.n14 585
R86 VPWR.n4 VPWR.t3 269.519
R87 VPWR.n19 VPWR.t5 250.975
R88 VPWR.n16 VPWR.n15 102.441
R89 VPWR.n5 VPWR.t0 42.3555
R90 VPWR.n8 VPWR.n7 34.6358
R91 VPWR.n8 VPWR.n2 34.6358
R92 VPWR.n15 VPWR.t1 26.5955
R93 VPWR.n16 VPWR.t4 26.5955
R94 VPWR.n5 VPWR.t2 26.5955
R95 VPWR.n14 VPWR.n2 26.4476
R96 VPWR.n18 VPWR.n17 24.1887
R97 VPWR.n19 VPWR.n18 22.5887
R98 VPWR.n7 VPWR.n6 14.3064
R99 VPWR.n7 VPWR.n3 9.3005
R100 VPWR.n9 VPWR.n8 9.3005
R101 VPWR.n10 VPWR.n2 9.3005
R102 VPWR.n13 VPWR.n12 9.3005
R103 VPWR.n11 VPWR.n1 9.3005
R104 VPWR.n18 VPWR.n0 9.3005
R105 VPWR.n20 VPWR.n19 9.3005
R106 VPWR.n13 VPWR.n1 8.65932
R107 VPWR.n6 VPWR.n4 7.41157
R108 VPWR.n17 VPWR.n1 0.847559
R109 VPWR.n14 VPWR.n13 0.282853
R110 VPWR.n4 VPWR.n3 0.176425
R111 VPWR.n9 VPWR.n3 0.120292
R112 VPWR.n10 VPWR.n9 0.120292
R113 VPWR.n12 VPWR.n10 0.120292
R114 VPWR.n12 VPWR.n11 0.120292
R115 VPWR.n11 VPWR.n0 0.120292
R116 VPWR.n20 VPWR.n0 0.120292
R117 VPWR VPWR.n20 0.0226354
R118 B1.n1 B1.t3 241.536
R119 B1.n0 B1.t1 241.536
R120 B1.n2 B1.n0 238.481
R121 B1.n1 B1.t2 169.237
R122 B1.n0 B1.t0 169.237
R123 B1.n2 B1.n1 152
R124 B1 B1.n2 18.2524
R125 VGND.n2 VGND.n1 219.91
R126 VGND.n2 VGND.n0 218.131
R127 VGND.n1 VGND.t0 24.9236
R128 VGND.n1 VGND.t1 24.9236
R129 VGND.n0 VGND.t2 24.9236
R130 VGND.n0 VGND.t3 24.9236
R131 VGND VGND.n2 1.43742
R132 A1.n2 A1.n0 260.188
R133 A1.n1 A1.t3 241.536
R134 A1.n0 A1.t1 241.536
R135 A1.n1 A1.t0 169.237
R136 A1.n0 A1.t2 169.237
R137 A1.n2 A1.n1 152
R138 A1 A1.n2 23.6805
R139 a_382_297.n1 a_382_297.n0 1223.84
R140 a_382_297.n0 a_382_297.t0 26.5955
R141 a_382_297.n0 a_382_297.t2 26.5955
R142 a_382_297.n1 a_382_297.t3 26.5955
R143 a_382_297.t1 a_382_297.n1 26.5955
C0 Y A2 0.012855f
C1 VGND A1 0.033269f
C2 C1 B1 0.027476f
C3 VPB A1 0.071126f
C4 A1 A2 0.209888f
C5 VPWR VGND 0.109184f
C6 VPB VPWR 0.127604f
C7 B1 VGND 0.024364f
C8 VPWR A2 0.016891f
C9 VGND B2 0.01545f
C10 Y A1 0.089204f
C11 VPB B1 0.068932f
C12 VPB B2 0.050999f
C13 VPWR Y 0.323987f
C14 C1 VGND 0.019628f
C15 B1 Y 0.252756f
C16 VPWR A1 0.077937f
C17 Y B2 0.018876f
C18 VPB C1 0.075615f
C19 B1 A1 0.092645f
C20 VPB VGND 0.008367f
C21 B1 VPWR 0.052761f
C22 C1 Y 0.083591f
C23 VPWR B2 0.016799f
C24 VGND A2 0.02453f
C25 VPB A2 0.050973f
C26 B1 B2 0.212706f
C27 Y VGND 0.01334f
C28 C1 VPWR 0.07159f
C29 VPB Y 0.005053f
C30 VGND VNB 0.621597f
C31 Y VNB 0.019474f
C32 VPWR VNB 0.584493f
C33 A2 VNB 0.166288f
C34 A1 VNB 0.227657f
C35 B2 VNB 0.166404f
C36 B1 VNB 0.199244f
C37 C1 VNB 0.242462f
C38 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221ai_4 VNB VPB VGND VPWR B2 Y A2 A1 B1 C1
X0 a_471_47.t6 A2.t0 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_471_47.t7 B2.t0 a_27_47.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_471_47.t5 A2.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t11 C1.t0 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t0 A1.t0 a_1241_297.t7 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47.t15 B2.t1 a_27_47.t5 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_471_47.t1 A1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t7 C1.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t6 C1.t2 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1241_297.t6 A1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X10 a_27_47.t4 B2.t2 a_471_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t11 B1.t0 a_553_297.t7 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t3 A2.t2 a_471_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_553_297.t6 B1.t1 VPWR.t9 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X14 a_27_47.t3 B2.t3 a_471_47.t14 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t2 A2.t3 a_471_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47.t11 C1.t3 Y.t6 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t1 A1.t3 a_471_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t5 C1.t4 a_27_47.t7 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 a_27_47.t8 C1.t5 Y.t4 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_1241_297.t5 A1.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR.t8 B1.t2 a_553_297.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t3 A1.t5 a_1241_297.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y.t12 B2.t4 a_553_297.t3 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1241_297.t3 A2.t4 Y.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t9 C1.t6 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X26 a_553_297.t2 B2.t5 Y.t13 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_47.t8 A1.t6 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y.t2 A2.t5 a_1241_297.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_553_297.t1 B2.t6 Y.t15 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_47.t1 B1.t3 a_471_47.t10 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND.t7 A1.t7 a_471_47.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X32 Y.t14 B2.t7 a_553_297.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1241_297.t1 A2.t6 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_27_47.t2 B1.t4 a_471_47.t11 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_553_297.t4 B1.t5 VPWR.t10 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y.t0 A2.t7 a_1241_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR.t4 C1.t7 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_47.t12 B1.t6 a_27_47.t9 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_471_47.t13 B1.t7 a_27_47.t10 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A2.n3 A2.t4 212.081
R1 A2.n5 A2.t5 212.081
R2 A2.n7 A2.t6 212.081
R3 A2.n1 A2.t7 212.081
R4 A2.n4 A2.n0 173.761
R5 A2.n9 A2.n2 173.761
R6 A2.n6 A2.n0 152
R7 A2.n9 A2.n8 152
R8 A2.n3 A2.t3 139.78
R9 A2.n5 A2.t1 139.78
R10 A2.n7 A2.t2 139.78
R11 A2.n1 A2.t0 139.78
R12 A2.n8 A2.n6 49.6611
R13 A2.n7 A2.n2 48.2005
R14 A2.n5 A2.n4 39.4369
R15 A2.n4 A2.n3 21.9096
R16 A2 A2.n0 16.0005
R17 A2.n2 A2.n1 13.146
R18 A2.n6 A2.n5 10.2247
R19 A2 A2.n9 5.7605
R20 A2.n8 A2.n7 1.46111
R21 VGND.n7 VGND.n6 218.452
R22 VGND.n5 VGND.n4 207.965
R23 VGND.n10 VGND.n3 207.965
R24 VGND.n1 VGND.n0 207.965
R25 VGND.n12 VGND.n11 34.6358
R26 VGND.n9 VGND.n5 32.377
R27 VGND.n10 VGND.n9 30.8711
R28 VGND.n6 VGND.t6 24.9236
R29 VGND.n6 VGND.t1 24.9236
R30 VGND.n4 VGND.t0 24.9236
R31 VGND.n4 VGND.t2 24.9236
R32 VGND.n3 VGND.t4 24.9236
R33 VGND.n3 VGND.t3 24.9236
R34 VGND.n0 VGND.t5 24.9236
R35 VGND.n0 VGND.t7 24.9236
R36 VGND.n12 VGND.n1 24.8476
R37 VGND.n14 VGND.n1 17.3894
R38 VGND.n7 VGND.n5 9.34458
R39 VGND.n9 VGND.n8 9.3005
R40 VGND.n11 VGND.n2 9.3005
R41 VGND.n13 VGND.n12 9.3005
R42 VGND.n11 VGND.n10 3.76521
R43 VGND VGND.n14 1.5595
R44 VGND.n8 VGND.n7 0.662609
R45 VGND.n14 VGND.n13 0.147187
R46 VGND.n8 VGND.n2 0.120292
R47 VGND.n13 VGND.n2 0.120292
R48 a_471_47.n5 a_471_47.t10 324.902
R49 a_471_47.n9 a_471_47.n8 185
R50 a_471_47.n7 a_471_47.n6 185
R51 a_471_47.n5 a_471_47.n4 185
R52 a_471_47.n1 a_471_47.t8 174.512
R53 a_471_47.n1 a_471_47.n0 98.982
R54 a_471_47.n3 a_471_47.n2 98.982
R55 a_471_47.n13 a_471_47.n12 98.982
R56 a_471_47.n11 a_471_47.n10 97.4305
R57 a_471_47.n9 a_471_47.n7 61.4405
R58 a_471_47.n7 a_471_47.n5 61.4405
R59 a_471_47.n11 a_471_47.n9 48.2889
R60 a_471_47.n12 a_471_47.n11 40.3399
R61 a_471_47.n10 a_471_47.t13 39.6928
R62 a_471_47.n3 a_471_47.n1 38.7884
R63 a_471_47.n12 a_471_47.n3 36.2672
R64 a_471_47.n10 a_471_47.t9 24.9236
R65 a_471_47.n4 a_471_47.t11 24.9236
R66 a_471_47.n4 a_471_47.t12 24.9236
R67 a_471_47.n6 a_471_47.t14 24.9236
R68 a_471_47.n6 a_471_47.t7 24.9236
R69 a_471_47.n8 a_471_47.t0 24.9236
R70 a_471_47.n8 a_471_47.t15 24.9236
R71 a_471_47.n2 a_471_47.t3 24.9236
R72 a_471_47.n2 a_471_47.t5 24.9236
R73 a_471_47.n0 a_471_47.t2 24.9236
R74 a_471_47.n0 a_471_47.t1 24.9236
R75 a_471_47.n13 a_471_47.t4 24.9236
R76 a_471_47.t6 a_471_47.n13 24.9236
R77 VNB.t14 VNB.t11 2677.02
R78 VNB.t16 VNB.t10 1423.95
R79 VNB.t2 VNB.t9 1196.12
R80 VNB.t1 VNB.t2 1196.12
R81 VNB.t3 VNB.t1 1196.12
R82 VNB.t5 VNB.t3 1196.12
R83 VNB.t4 VNB.t5 1196.12
R84 VNB.t6 VNB.t4 1196.12
R85 VNB.t10 VNB.t6 1196.12
R86 VNB.t0 VNB.t16 1196.12
R87 VNB.t18 VNB.t0 1196.12
R88 VNB.t17 VNB.t18 1196.12
R89 VNB.t8 VNB.t17 1196.12
R90 VNB.t12 VNB.t8 1196.12
R91 VNB.t15 VNB.t12 1196.12
R92 VNB.t11 VNB.t15 1196.12
R93 VNB.t7 VNB.t14 1196.12
R94 VNB.t19 VNB.t7 1196.12
R95 VNB.t13 VNB.t19 1196.12
R96 VNB VNB.t13 968.285
R97 B2.n3 B2.t5 212.081
R98 B2.n2 B2.t4 212.081
R99 B2.n1 B2.t6 212.081
R100 B2.n0 B2.t7 212.081
R101 B2.n3 B2.t2 139.78
R102 B2.n2 B2.t1 139.78
R103 B2.n1 B2.t3 139.78
R104 B2.n0 B2.t0 139.78
R105 B2 B2.n4 69.9965
R106 B2.n2 B2.n1 61.346
R107 B2.n1 B2.n0 61.346
R108 B2.n4 B2.n3 31.1263
R109 B2.n4 B2.n2 23.4986
R110 a_27_47.n5 a_27_47.t8 263.462
R111 a_27_47.n2 a_27_47.n0 233.874
R112 a_27_47.n2 a_27_47.n1 185
R113 a_27_47.n7 a_27_47.n6 185
R114 a_27_47.n4 a_27_47.n3 185
R115 a_27_47.n9 a_27_47.n8 185
R116 a_27_47.n4 a_27_47.t7 178.347
R117 a_27_47.n7 a_27_47.n5 54.6914
R118 a_27_47.n8 a_27_47.n2 48.8732
R119 a_27_47.n8 a_27_47.n7 48.8732
R120 a_27_47.n5 a_27_47.n4 48.8732
R121 a_27_47.n3 a_27_47.t0 24.9236
R122 a_27_47.n3 a_27_47.t11 24.9236
R123 a_27_47.n6 a_27_47.t9 24.9236
R124 a_27_47.n6 a_27_47.t1 24.9236
R125 a_27_47.n1 a_27_47.t5 24.9236
R126 a_27_47.n1 a_27_47.t3 24.9236
R127 a_27_47.n0 a_27_47.t10 24.9236
R128 a_27_47.n0 a_27_47.t4 24.9236
R129 a_27_47.t6 a_27_47.n9 24.9236
R130 a_27_47.n9 a_27_47.t2 24.9236
R131 C1.n1 C1.t6 212.081
R132 C1.n2 C1.t7 212.081
R133 C1.n4 C1.t0 212.081
R134 C1.n6 C1.t2 212.081
R135 C1.n3 C1.n0 173.761
R136 C1.n5 C1.n0 152
R137 C1.n1 C1.t4 139.78
R138 C1.n2 C1.t5 139.78
R139 C1.n4 C1.t1 139.78
R140 C1.n6 C1.t3 139.78
R141 C1 C1.n7 85.7128
R142 C1.n6 C1.n5 37.9763
R143 C1.n3 C1.n2 35.055
R144 C1.n7 C1.n6 31.7924
R145 C1.n4 C1.n3 26.2914
R146 C1.n5 C1.n4 23.3702
R147 C1.n7 C1.n1 22.986
R148 C1 C1.n0 6.4005
R149 VPWR.n6 VPWR.n5 606.505
R150 VPWR.n14 VPWR.n13 606.505
R151 VPWR.n24 VPWR.n10 603.944
R152 VPWR.n37 VPWR.n3 585
R153 VPWR.n39 VPWR.n38 585
R154 VPWR.n44 VPWR.n2 316.757
R155 VPWR.n15 VPWR.t0 259.39
R156 VPWR.n46 VPWR.t5 250.975
R157 VPWR.n38 VPWR.n37 102.441
R158 VPWR.n26 VPWR.n25 34.6358
R159 VPWR.n26 VPWR.n8 34.6358
R160 VPWR.n30 VPWR.n8 34.6358
R161 VPWR.n31 VPWR.n30 34.6358
R162 VPWR.n32 VPWR.n31 34.6358
R163 VPWR.n18 VPWR.n17 34.6358
R164 VPWR.n19 VPWR.n18 34.6358
R165 VPWR.n19 VPWR.n11 34.6358
R166 VPWR.n23 VPWR.n11 34.6358
R167 VPWR.n10 VPWR.t1 34.4755
R168 VPWR.n10 VPWR.t8 34.4755
R169 VPWR.n36 VPWR.n35 30.4005
R170 VPWR.n44 VPWR.n43 27.4829
R171 VPWR.n38 VPWR.t9 26.5955
R172 VPWR.n37 VPWR.t4 26.5955
R173 VPWR.n2 VPWR.t7 26.5955
R174 VPWR.n2 VPWR.t6 26.5955
R175 VPWR.n5 VPWR.t10 26.5955
R176 VPWR.n5 VPWR.t11 26.5955
R177 VPWR.n13 VPWR.t2 26.5955
R178 VPWR.n13 VPWR.t3 26.5955
R179 VPWR.n45 VPWR.n44 22.9652
R180 VPWR.n46 VPWR.n45 21.4593
R181 VPWR.n17 VPWR.n14 19.9534
R182 VPWR.n43 VPWR.n3 19.2946
R183 VPWR.n35 VPWR.n6 15.4358
R184 VPWR.n24 VPWR.n23 15.4358
R185 VPWR.n17 VPWR.n16 9.3005
R186 VPWR.n18 VPWR.n12 9.3005
R187 VPWR.n20 VPWR.n19 9.3005
R188 VPWR.n21 VPWR.n11 9.3005
R189 VPWR.n23 VPWR.n22 9.3005
R190 VPWR.n25 VPWR.n9 9.3005
R191 VPWR.n27 VPWR.n26 9.3005
R192 VPWR.n28 VPWR.n8 9.3005
R193 VPWR.n30 VPWR.n29 9.3005
R194 VPWR.n31 VPWR.n7 9.3005
R195 VPWR.n33 VPWR.n32 9.3005
R196 VPWR.n35 VPWR.n34 9.3005
R197 VPWR.n36 VPWR.n4 9.3005
R198 VPWR.n41 VPWR.n40 9.3005
R199 VPWR.n43 VPWR.n42 9.3005
R200 VPWR.n44 VPWR.n1 9.3005
R201 VPWR.n45 VPWR.n0 9.3005
R202 VPWR.n47 VPWR.n46 9.3005
R203 VPWR.n40 VPWR.n39 7.71815
R204 VPWR.n15 VPWR.n14 6.81939
R205 VPWR.n40 VPWR.n3 2.07109
R206 VPWR.n39 VPWR.n36 0.941676
R207 VPWR.n16 VPWR.n15 0.750778
R208 VPWR.n25 VPWR.n24 0.376971
R209 VPWR.n32 VPWR.n6 0.376971
R210 VPWR.n16 VPWR.n12 0.120292
R211 VPWR.n20 VPWR.n12 0.120292
R212 VPWR.n21 VPWR.n20 0.120292
R213 VPWR.n22 VPWR.n21 0.120292
R214 VPWR.n22 VPWR.n9 0.120292
R215 VPWR.n27 VPWR.n9 0.120292
R216 VPWR.n28 VPWR.n27 0.120292
R217 VPWR.n29 VPWR.n28 0.120292
R218 VPWR.n29 VPWR.n7 0.120292
R219 VPWR.n33 VPWR.n7 0.120292
R220 VPWR.n34 VPWR.n33 0.120292
R221 VPWR.n34 VPWR.n4 0.120292
R222 VPWR.n41 VPWR.n4 0.120292
R223 VPWR.n42 VPWR.n41 0.120292
R224 VPWR.n42 VPWR.n1 0.120292
R225 VPWR.n1 VPWR.n0 0.120292
R226 VPWR.n47 VPWR.n0 0.120292
R227 VPWR VPWR.n47 0.0213333
R228 Y.n2 Y.n0 641.403
R229 Y.n11 Y.n10 585
R230 Y.n13 Y.n12 585
R231 Y.n2 Y.n1 585
R232 Y.n8 Y.n7 256.58
R233 Y.n5 Y.n3 233.874
R234 Y.n8 Y.n6 197.011
R235 Y.n5 Y.n4 185
R236 Y.n11 Y.n9 169.931
R237 Y Y.n13 80.7747
R238 Y.n9 Y.n5 64.1424
R239 Y.n13 Y.n11 55.4585
R240 Y Y.n2 35.4914
R241 Y.n1 Y.t1 26.5955
R242 Y.n1 Y.t0 26.5955
R243 Y.n12 Y.t13 26.5955
R244 Y.n12 Y.t12 26.5955
R245 Y.n10 Y.t15 26.5955
R246 Y.n10 Y.t14 26.5955
R247 Y.n6 Y.t8 26.5955
R248 Y.n6 Y.t11 26.5955
R249 Y.n7 Y.t10 26.5955
R250 Y.n7 Y.t9 26.5955
R251 Y.n0 Y.t3 26.5955
R252 Y.n0 Y.t2 26.5955
R253 Y.n3 Y.t6 24.9236
R254 Y.n3 Y.t5 24.9236
R255 Y.n4 Y.t4 24.9236
R256 Y.n4 Y.t7 24.9236
R257 Y.n9 Y.n8 12.0476
R258 VPB.t8 VPB.t17 556.386
R259 VPB.t12 VPB.t1 295.95
R260 VPB.t2 VPB.t0 248.599
R261 VPB.t7 VPB.t2 248.599
R262 VPB.t6 VPB.t7 248.599
R263 VPB.t5 VPB.t6 248.599
R264 VPB.t4 VPB.t5 248.599
R265 VPB.t3 VPB.t4 248.599
R266 VPB.t1 VPB.t3 248.599
R267 VPB.t15 VPB.t12 248.599
R268 VPB.t16 VPB.t15 248.599
R269 VPB.t14 VPB.t16 248.599
R270 VPB.t13 VPB.t14 248.599
R271 VPB.t18 VPB.t13 248.599
R272 VPB.t19 VPB.t18 248.599
R273 VPB.t17 VPB.t19 248.599
R274 VPB.t11 VPB.t8 248.599
R275 VPB.t10 VPB.t11 248.599
R276 VPB.t9 VPB.t10 248.599
R277 VPB VPB.t9 201.246
R278 A1.n6 A1.n2 323.546
R279 A1.n2 A1.t2 241.536
R280 A1.n0 A1.t0 212.081
R281 A1.n3 A1.t4 212.081
R282 A1.n4 A1.t5 212.081
R283 A1.n2 A1.t7 169.237
R284 A1.n6 A1.n5 152.726
R285 A1.n0 A1.t6 139.78
R286 A1.n3 A1.t3 139.78
R287 A1.n4 A1.t1 139.78
R288 A1 A1.n1 83.7928
R289 A1.n5 A1.n3 48.2005
R290 A1.n1 A1.n0 33.2102
R291 A1.n3 A1.n1 21.5682
R292 A1.n5 A1.n4 13.146
R293 A1 A1.n6 1.9205
R294 a_1241_297.n3 a_1241_297.n1 638.4
R295 a_1241_297.n3 a_1241_297.n2 585
R296 a_1241_297.n5 a_1241_297.n4 288.212
R297 a_1241_297.n4 a_1241_297.n0 257.983
R298 a_1241_297.n4 a_1241_297.n3 61.8028
R299 a_1241_297.n2 a_1241_297.t2 26.5955
R300 a_1241_297.n2 a_1241_297.t1 26.5955
R301 a_1241_297.n1 a_1241_297.t0 26.5955
R302 a_1241_297.n1 a_1241_297.t6 26.5955
R303 a_1241_297.n0 a_1241_297.t7 26.5955
R304 a_1241_297.n0 a_1241_297.t5 26.5955
R305 a_1241_297.n5 a_1241_297.t4 26.5955
R306 a_1241_297.t3 a_1241_297.n5 26.5955
R307 B1.n3 B1.n2 327.858
R308 B1.n2 B1.t2 241.536
R309 B1.n1 B1.t5 212.081
R310 B1.n5 B1.t0 212.081
R311 B1.n7 B1.t1 212.081
R312 B1.n2 B1.t7 169.237
R313 B1 B1.n8 164.481
R314 B1.n4 B1.n3 152
R315 B1.n6 B1.n0 152
R316 B1.n1 B1.t4 139.78
R317 B1.n5 B1.t6 139.78
R318 B1.n7 B1.t3 139.78
R319 B1.n8 B1.n6 49.6611
R320 B1.n5 B1.n4 44.549
R321 B1.n3 B1.n0 21.7605
R322 B1.n4 B1.n1 16.7975
R323 B1 B1.n0 9.2805
R324 B1.n8 B1.n7 6.57323
R325 B1.n6 B1.n5 5.11262
R326 a_553_297.n4 a_553_297.n0 639.212
R327 a_553_297.n5 a_553_297.n4 585
R328 a_553_297.n3 a_553_297.n1 361.488
R329 a_553_297.n3 a_553_297.n2 287.411
R330 a_553_297.n4 a_553_297.n3 68.0113
R331 a_553_297.n2 a_553_297.t0 26.5955
R332 a_553_297.n2 a_553_297.t4 26.5955
R333 a_553_297.n1 a_553_297.t7 26.5955
R334 a_553_297.n1 a_553_297.t6 26.5955
R335 a_553_297.n0 a_553_297.t5 26.5955
R336 a_553_297.n0 a_553_297.t2 26.5955
R337 a_553_297.t3 a_553_297.n5 26.5955
R338 a_553_297.n5 a_553_297.t1 26.5955
C0 Y A1 0.160979f
C1 VGND B2 0.027766f
C2 C1 B1 0.018341f
C3 A1 VPWR 0.111422f
C4 VPB Y 0.018946f
C5 B1 A1 0.093016f
C6 VPB VPWR 0.195845f
C7 Y VGND 0.033912f
C8 Y B2 0.046582f
C9 VPB B1 0.128911f
C10 VGND VPWR 0.188013f
C11 A1 A2 0.291492f
C12 B2 VPWR 0.028127f
C13 B1 VGND 0.041438f
C14 VPB A2 0.114794f
C15 B1 B2 0.254097f
C16 VPB C1 0.130786f
C17 VGND A2 0.058403f
C18 Y VPWR 0.498232f
C19 B2 A2 5.76e-19
C20 B1 Y 0.360375f
C21 C1 VGND 0.037341f
C22 VPB A1 0.133283f
C23 B1 VPWR 0.073133f
C24 Y A2 0.032103f
C25 VGND A1 0.062783f
C26 B2 A1 5.11e-19
C27 A2 VPWR 0.034066f
C28 VPB VGND 0.01241f
C29 C1 Y 0.323787f
C30 VPB B2 0.113959f
C31 B1 A2 3.11e-19
C32 C1 VPWR 0.112123f
C33 VGND VNB 1.02648f
C34 Y VNB 0.029153f
C35 VPWR VNB 0.916885f
C36 A2 VNB 0.351925f
C37 A1 VNB 0.402829f
C38 B2 VNB 0.350721f
C39 B1 VNB 0.373349f
C40 C1 VNB 0.410473f
C41 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_4 VNB VPB VPWR VGND D1 B1 C1 A2 A1 X
X0 VGND.t3 A1.t0 a_361_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X1 X.t7 a_27_297.t10 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297.t9 A2.t0 a_852_297.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1775 ps=1.355 w=1 l=0.15
X3 VPWR.t2 a_27_297.t11 X.t6 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t0 a_27_297.t12 X.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.115375 ps=1.005 w=0.65 l=0.15
X5 VPWR.t6 B1.t0 a_27_297.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_852_297.t0 A1.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7 a_27_297.t2 B1.t1 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_361_47.t0 A1.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t10 C1.t0 a_27_297.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t7 A2.t1 a_361_47.t4 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.144625 pd=1.095 as=0.12025 ps=1.02 w=0.65 l=0.15
X11 a_27_297.t4 D1.t0 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X.t2 a_27_297.t13 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.144625 ps=1.095 w=0.65 l=0.15
X13 X.t5 a_27_297.t14 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 a_27_47.t3 D1.t1 a_27_297.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_361_47.t3 B1.t2 a_277_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_361_47.t2 A2.t2 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_277_47.t1 C1.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_445_47.t0 B1.t3 a_361_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X.t1 a_27_297.t15 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.092625 ps=0.935 w=0.65 l=0.15
X20 a_27_297.t7 C1.t2 VPWR.t11 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X21 a_681_297.t1 A2.t3 a_27_297.t6 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.305 ps=1.61 w=1 l=0.15
X22 a_27_47.t1 C1.t3 a_445_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X23 VGND.t5 a_27_297.t16 X.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.095875 ps=0.945 w=0.65 l=0.15
X24 VPWR.t7 D1.t2 a_27_297.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 VPWR.t0 a_27_297.t17 X.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR.t4 A1.t3 a_681_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X27 a_27_297.t8 D1.t3 a_27_47.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t3 218.079
R1 A1.n0 A1.t1 194.782
R2 A1.n1 A1.t2 171.913
R3 A1 A1.n2 165.745
R4 A1.n1 A1.t0 145.957
R5 A1.n2 A1.n0 21.2836
R6 A1.n2 A1.n1 12.52
R7 a_361_47.n2 a_361_47.n0 284.502
R8 a_361_47.n3 a_361_47.n2 141.91
R9 a_361_47.n2 a_361_47.n1 95.5251
R10 a_361_47.n3 a_361_47.t4 34.1543
R11 a_361_47.t0 a_361_47.n3 34.1543
R12 a_361_47.n1 a_361_47.t2 33.2313
R13 a_361_47.n0 a_361_47.t5 24.9236
R14 a_361_47.n0 a_361_47.t3 24.9236
R15 a_361_47.n1 a_361_47.t1 24.9236
R16 VGND.n0 VGND.t6 282.817
R17 VGND.n4 VGND.t5 282.053
R18 VGND.n9 VGND.n8 203.356
R19 VGND.n6 VGND.n5 200.361
R20 VGND.n15 VGND.n14 198.147
R21 VGND.n8 VGND.t1 48.0005
R22 VGND.n13 VGND.n2 34.6358
R23 VGND.n17 VGND.n16 34.6358
R24 VGND.n8 VGND.t7 34.1543
R25 VGND.n9 VGND.n7 33.8829
R26 VGND.n5 VGND.t0 26.7697
R27 VGND.n5 VGND.t4 25.8467
R28 VGND.n14 VGND.t2 24.9236
R29 VGND.n14 VGND.t3 24.9236
R30 VGND.n7 VGND.n6 24.4711
R31 VGND.n19 VGND.n0 16.6364
R32 VGND.n9 VGND.n2 15.4358
R33 VGND.n7 VGND.n3 9.3005
R34 VGND.n10 VGND.n9 9.3005
R35 VGND.n11 VGND.n2 9.3005
R36 VGND.n13 VGND.n12 9.3005
R37 VGND.n16 VGND.n1 9.3005
R38 VGND.n18 VGND.n17 9.3005
R39 VGND.n6 VGND.n4 6.46386
R40 VGND.n16 VGND.n15 6.4005
R41 VGND.n17 VGND.n0 0.753441
R42 VGND VGND.n19 0.718178
R43 VGND.n4 VGND.n3 0.717579
R44 VGND.n15 VGND.n13 0.376971
R45 VGND.n19 VGND.n18 0.147186
R46 VGND.n10 VGND.n3 0.120292
R47 VGND.n11 VGND.n10 0.120292
R48 VGND.n12 VGND.n11 0.120292
R49 VGND.n12 VGND.n1 0.120292
R50 VGND.n18 VGND.n1 0.120292
R51 VNB.t9 VNB.t8 2776.7
R52 VNB.t12 VNB.t1 1694.5
R53 VNB.t2 VNB.t12 1480.91
R54 VNB.t1 VNB.t0 1438.19
R55 VNB.t8 VNB.t3 1324.27
R56 VNB.t6 VNB.t7 1267.31
R57 VNB.t0 VNB.t6 1238.83
R58 VNB.t3 VNB.t2 1196.12
R59 VNB.t11 VNB.t13 1196.12
R60 VNB.t4 VNB.t11 1196.12
R61 VNB.t5 VNB.t4 1196.12
R62 VNB.t10 VNB.t5 1196.12
R63 VNB.t13 VNB.t9 1025.24
R64 VNB VNB.t10 925.567
R65 a_27_297.n23 a_27_297.n22 606.427
R66 a_27_297.n21 a_27_297.n20 585
R67 a_27_297.n1 a_27_297.t1 338.296
R68 a_27_297.n17 a_27_297.t9 324.786
R69 a_27_297.n3 a_27_297.n2 300.154
R70 a_27_297.n19 a_27_297.n18 292.5
R71 a_27_297.n1 a_27_297.n0 227.852
R72 a_27_297.n6 a_27_297.t17 225.291
R73 a_27_297.n7 a_27_297.t10 221.72
R74 a_27_297.n11 a_27_297.t11 221.72
R75 a_27_297.n14 a_27_297.t14 221.72
R76 a_27_297.n9 a_27_297.n8 169.763
R77 a_27_297.n15 a_27_297.t13 165.488
R78 a_27_297.n16 a_27_297.n15 152
R79 a_27_297.n13 a_27_297.n4 152
R80 a_27_297.n10 a_27_297.n9 152
R81 a_27_297.n12 a_27_297.t12 149.421
R82 a_27_297.n5 a_27_297.t15 149.421
R83 a_27_297.n6 a_27_297.t16 149.421
R84 a_27_297.n18 a_27_297.n17 112.309
R85 a_27_297.n17 a_27_297.n16 74.2651
R86 a_27_297.n20 a_27_297.n19 66.9805
R87 a_27_297.n14 a_27_297.n13 50.8783
R88 a_27_297.n22 a_27_297.n21 50.7196
R89 a_27_297.n8 a_27_297.n6 49.0931
R90 a_27_297.n22 a_27_297.n3 41.3262
R91 a_27_297.n11 a_27_297.n10 36.5968
R92 a_27_297.n10 a_27_297.n5 30.3486
R93 a_27_297.n19 a_27_297.t6 26.5955
R94 a_27_297.n20 a_27_297.t7 26.5955
R95 a_27_297.n2 a_27_297.t5 26.5955
R96 a_27_297.n2 a_27_297.t4 26.5955
R97 a_27_297.t0 a_27_297.n23 26.5955
R98 a_27_297.n23 a_27_297.t2 26.5955
R99 a_27_297.n0 a_27_297.t3 24.9236
R100 a_27_297.n0 a_27_297.t8 24.9236
R101 a_27_297.n8 a_27_297.n7 22.3153
R102 a_27_297.n9 a_27_297.n4 17.7638
R103 a_27_297.n16 a_27_297.n4 17.7638
R104 a_27_297.n13 a_27_297.n12 13.3894
R105 a_27_297.n3 a_27_297.n1 11.3376
R106 a_27_297.n12 a_27_297.n11 10.7116
R107 a_27_297.n15 a_27_297.n14 9.81902
R108 a_27_297.n7 a_27_297.n5 8.03383
R109 a_27_297.n21 a_27_297.n18 6.85404
R110 VPWR.n16 VPWR.t1 868.288
R111 VPWR.n28 VPWR.n3 605.481
R112 VPWR.n30 VPWR.n1 599.74
R113 VPWR.n5 VPWR.n4 598.965
R114 VPWR.n8 VPWR.n7 598.965
R115 VPWR.n13 VPWR.t0 343.899
R116 VPWR.n12 VPWR.n11 311.062
R117 VPWR.n23 VPWR.n22 34.6358
R118 VPWR.n24 VPWR.n23 34.6358
R119 VPWR.n18 VPWR.n17 34.6358
R120 VPWR.n28 VPWR.n27 33.5064
R121 VPWR.n17 VPWR.n16 31.2476
R122 VPWR.n7 VPWR.t5 27.5805
R123 VPWR.n7 VPWR.t4 27.5805
R124 VPWR.n22 VPWR.n8 26.7299
R125 VPWR.n1 VPWR.t9 26.5955
R126 VPWR.n1 VPWR.t7 26.5955
R127 VPWR.n3 VPWR.t8 26.5955
R128 VPWR.n3 VPWR.t10 26.5955
R129 VPWR.n4 VPWR.t11 26.5955
R130 VPWR.n4 VPWR.t6 26.5955
R131 VPWR.n11 VPWR.t3 26.5955
R132 VPWR.n11 VPWR.t2 26.5955
R133 VPWR.n15 VPWR.n12 25.977
R134 VPWR.n30 VPWR.n29 22.9652
R135 VPWR.n29 VPWR.n28 18.824
R136 VPWR.n18 VPWR.n8 17.6946
R137 VPWR.n16 VPWR.n15 12.424
R138 VPWR.n27 VPWR.n5 9.41227
R139 VPWR.n15 VPWR.n14 9.3005
R140 VPWR.n16 VPWR.n10 9.3005
R141 VPWR.n17 VPWR.n9 9.3005
R142 VPWR.n19 VPWR.n18 9.3005
R143 VPWR.n20 VPWR.n8 9.3005
R144 VPWR.n22 VPWR.n21 9.3005
R145 VPWR.n23 VPWR.n6 9.3005
R146 VPWR.n25 VPWR.n24 9.3005
R147 VPWR.n27 VPWR.n26 9.3005
R148 VPWR.n28 VPWR.n2 9.3005
R149 VPWR.n29 VPWR.n0 9.3005
R150 VPWR.n31 VPWR.n30 7.12063
R151 VPWR.n13 VPWR.n12 6.27043
R152 VPWR.n14 VPWR.n13 0.730508
R153 VPWR.n24 VPWR.n5 0.376971
R154 VPWR.n31 VPWR.n0 0.148519
R155 VPWR.n14 VPWR.n10 0.120292
R156 VPWR.n10 VPWR.n9 0.120292
R157 VPWR.n19 VPWR.n9 0.120292
R158 VPWR.n20 VPWR.n19 0.120292
R159 VPWR.n21 VPWR.n20 0.120292
R160 VPWR.n21 VPWR.n6 0.120292
R161 VPWR.n25 VPWR.n6 0.120292
R162 VPWR.n26 VPWR.n25 0.120292
R163 VPWR.n26 VPWR.n2 0.120292
R164 VPWR.n2 VPWR.n0 0.120292
R165 VPWR VPWR.n31 0.114842
R166 X.n5 X.n3 377.07
R167 X.n5 X.n4 323.716
R168 X.n2 X.n0 255.928
R169 X.n2 X.n1 208.041
R170 X.n0 X.t2 40.6159
R171 X.n1 X.t0 28.6159
R172 X.n3 X.t6 26.5955
R173 X.n3 X.t5 26.5955
R174 X.n4 X.t4 26.5955
R175 X.n4 X.t7 26.5955
R176 X.n1 X.t1 25.8467
R177 X.n0 X.t3 24.9236
R178 X X.n5 23.7181
R179 X.n6 X.n2 19.577
R180 X.n6 X 15.4079
R181 X X.n6 0.711611
R182 VPB.t13 VPB.t1 556.386
R183 VPB.t12 VPB.t11 449.844
R184 VPB.t5 VPB.t13 298.911
R185 VPB.t4 VPB.t5 254.518
R186 VPB.t11 VPB.t4 251.559
R187 VPB.t3 VPB.t0 248.599
R188 VPB.t2 VPB.t3 248.599
R189 VPB.t1 VPB.t2 248.599
R190 VPB.t6 VPB.t12 248.599
R191 VPB.t8 VPB.t6 248.599
R192 VPB.t10 VPB.t8 248.599
R193 VPB.t9 VPB.t10 248.599
R194 VPB.t7 VPB.t9 248.599
R195 VPB VPB.t7 192.369
R196 A2.n2 A2.n1 273.329
R197 A2.n0 A2.t3 242.054
R198 A2.n1 A2.t0 234.012
R199 A2.n1 A2.t1 169.138
R200 A2.n0 A2.t2 160.357
R201 A2.n2 A2.n0 152.262
R202 A2 A2.n2 3.90558
R203 a_852_297.t0 a_852_297.t1 69.9355
R204 B1.n0 B1.t0 221.72
R205 B1.n1 B1.t1 221.72
R206 B1 B1.n2 153.601
R207 B1.n0 B1.t3 149.421
R208 B1.n1 B1.t2 149.421
R209 B1.n2 B1.n0 37.4894
R210 B1.n2 B1.n1 37.4894
R211 C1.n1 C1.t2 645.109
R212 C1.n2 C1.n0 273.384
R213 C1.n0 C1.t0 241.536
R214 C1.n0 C1.t1 169.237
R215 C1.n1 C1.t3 164.361
R216 C1.n2 C1.n1 152
R217 C1 C1.n2 1.87783
R218 D1.n1 D1.t2 230.793
R219 D1.n0 D1.t0 221.72
R220 D1.n1 D1.t3 158.494
R221 D1 D1.n1 154.133
R222 D1.n0 D1.t1 149.421
R223 D1.n1 D1.n0 61.5894
R224 a_27_47.n1 a_27_47.t1 358.233
R225 a_27_47.t2 a_27_47.n1 293.543
R226 a_27_47.n1 a_27_47.n0 185
R227 a_27_47.n0 a_27_47.t0 24.9236
R228 a_27_47.n0 a_27_47.t3 24.9236
R229 a_277_47.t0 a_277_47.t1 49.8467
R230 a_445_47.t0 a_445_47.t1 38.7697
R231 a_681_297.t0 a_681_297.t1 54.1755
C0 X D1 5.41e-21
C1 VPWR C1 0.042531f
C2 A1 X 1.72e-19
C3 VPB A1 0.059199f
C4 VPB D1 0.070924f
C5 VGND A2 0.038965f
C6 A1 VPWR 0.032428f
C7 A1 C1 1.02e-19
C8 D1 C1 0.060728f
C9 VPWR D1 0.03313f
C10 X VGND 0.247343f
C11 VGND B1 0.014917f
C12 X A2 0.001206f
C13 VPB A2 0.082943f
C14 VPB VGND 0.012728f
C15 VPWR VGND 0.144116f
C16 VPWR A2 0.03629f
C17 X B1 4.79e-20
C18 VGND C1 0.019416f
C19 C1 A2 0.053702f
C20 VPB B1 0.051554f
C21 VPB X 0.011896f
C22 A1 A2 0.18946f
C23 VPWR B1 0.027832f
C24 VGND D1 0.017912f
C25 VPWR X 0.322571f
C26 X C1 4.03e-19
C27 A1 VGND 0.027022f
C28 C1 B1 0.202654f
C29 VPB VPWR 0.149929f
C30 VPB C1 0.069585f
C31 VGND VNB 0.816291f
C32 X VNB 0.06354f
C33 VPWR VNB 0.686543f
C34 A1 VNB 0.187864f
C35 A2 VNB 0.2243f
C36 B1 VNB 0.166822f
C37 C1 VNB 0.197445f
C38 D1 VNB 0.246793f
C39 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_2 VPB VNB VGND VPWR X D1 C1 B1 A2 A1
X0 VPWR.t3 a_80_21.t5 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.14 ps=1.28 w=1 l=0.15
X1 X.t0 a_80_21.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 a_80_21.t2 D1.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.365 ps=1.73 w=1 l=0.15
X3 VGND.t2 a_80_21.t7 X.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR.t0 C1.t0 a_80_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X5 X.t2 a_80_21.t8 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_80_21.t1 B1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7 a_674_297.t1 A2.t0 a_80_21.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X8 a_386_47.t0 D1.t1 a_80_21.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X9 VPWR.t4 A1.t0 a_674_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X10 a_566_47.t1 B1.t1 a_458_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 VGND.t0 A2.t1 a_566_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 a_566_47.t0 A1.t1 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X13 a_458_47.t1 C1.t1 a_386_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
R0 a_80_21.n4 a_80_21.n3 335.526
R1 a_80_21.n5 a_80_21.n4 297.183
R2 a_80_21.n1 a_80_21.t5 212.081
R3 a_80_21.n0 a_80_21.t6 212.081
R4 a_80_21.n2 a_80_21.n1 182.673
R5 a_80_21.n2 a_80_21.t3 166.165
R6 a_80_21.n1 a_80_21.t7 139.78
R7 a_80_21.n0 a_80_21.t8 139.78
R8 a_80_21.n4 a_80_21.n2 64.2769
R9 a_80_21.n1 a_80_21.n0 62.8066
R10 a_80_21.n3 a_80_21.t1 39.4005
R11 a_80_21.n3 a_80_21.t4 37.4305
R12 a_80_21.t0 a_80_21.n5 27.5805
R13 a_80_21.n5 a_80_21.t2 27.5805
R14 X.n0 X 593.095
R15 X.n1 X.n0 289.336
R16 X X.n3 185.189
R17 X.n3 X.n2 185
R18 X.n2 X.n1 40.2141
R19 X.n0 X.t1 27.5805
R20 X.n0 X.t0 27.5805
R21 X.n3 X.t3 25.8467
R22 X.n3 X.t2 25.8467
R23 X X.n2 12.6123
R24 X.n1 X 11.0376
R25 VPWR.n4 VPWR.n3 599.74
R26 VPWR.n13 VPWR.n12 585
R27 VPWR.n11 VPWR.n10 585
R28 VPWR.n5 VPWR.t4 257.017
R29 VPWR.n15 VPWR.t2 256.889
R30 VPWR.n12 VPWR.n11 88.6505
R31 VPWR.n3 VPWR.t0 39.4005
R32 VPWR.n3 VPWR.t1 37.4305
R33 VPWR.n9 VPWR.n2 32.1918
R34 VPWR.n14 VPWR.n13 27.7606
R35 VPWR.n11 VPWR.t5 27.5805
R36 VPWR.n12 VPWR.t3 27.5805
R37 VPWR.n15 VPWR.n14 25.977
R38 VPWR.n4 VPWR.n2 19.2005
R39 VPWR.n6 VPWR.n2 9.3005
R40 VPWR.n9 VPWR.n8 9.3005
R41 VPWR.n7 VPWR.n1 9.3005
R42 VPWR.n14 VPWR.n0 9.3005
R43 VPWR.n16 VPWR.n15 9.3005
R44 VPWR.n10 VPWR.n1 8.81362
R45 VPWR.n5 VPWR.n4 7.17077
R46 VPWR.n10 VPWR.n9 0.839844
R47 VPWR.n13 VPWR.n1 0.630008
R48 VPWR.n6 VPWR.n5 0.204792
R49 VPWR.n8 VPWR.n6 0.120292
R50 VPWR.n8 VPWR.n7 0.120292
R51 VPWR.n7 VPWR.n0 0.120292
R52 VPWR.n16 VPWR.n0 0.120292
R53 VPWR VPWR.n16 0.0213333
R54 VPB.t3 VPB.t5 520.872
R55 VPB.t6 VPB.t4 319.627
R56 VPB.t1 VPB.t6 319.627
R57 VPB.t0 VPB.t1 319.627
R58 VPB.t5 VPB.t0 254.518
R59 VPB.t2 VPB.t3 254.518
R60 VPB VPB.t2 192.369
R61 D1.n0 D1.t0 230.793
R62 D1.n0 D1.t1 158.494
R63 D1 D1.n0 154.845
R64 VGND.n3 VGND.t2 285.966
R65 VGND.n2 VGND.n1 205.471
R66 VGND.n5 VGND.t1 159.273
R67 VGND.n1 VGND.t3 38.7697
R68 VGND.n1 VGND.t0 33.2313
R69 VGND.n4 VGND.n3 25.977
R70 VGND.n5 VGND.n4 25.977
R71 VGND.n6 VGND.n5 9.3005
R72 VGND.n4 VGND.n0 9.3005
R73 VGND.n3 VGND.n2 7.18319
R74 VGND.n2 VGND.n0 0.155401
R75 VGND.n6 VGND.n0 0.120292
R76 VGND VGND.n6 0.0213333
R77 VNB.t3 VNB.t4 2705.5
R78 VNB.t0 VNB.t6 1537.86
R79 VNB.t5 VNB.t0 1537.86
R80 VNB.t1 VNB.t5 1537.86
R81 VNB.t2 VNB.t3 1224.6
R82 VNB.t4 VNB.t1 1025.24
R83 VNB VNB.t2 925.567
R84 C1.n0 C1.t0 241.439
R85 C1 C1.n0 176.436
R86 C1.n0 C1.t1 169.138
R87 B1.n0 B1.t0 241.439
R88 B1.n0 B1.t1 169.138
R89 B1 B1.n0 154.016
R90 A2.n0 A2.t0 241.439
R91 A2.n0 A2.t1 169.138
R92 A2.n1 A2.n0 152
R93 A2.n1 A2 41.1775
R94 A2 A2.n1 1.95606
R95 a_674_297.t0 a_674_297.t1 76.8305
R96 a_386_47.t0 a_386_47.t1 38.7697
R97 A1.n0 A1.t0 236.022
R98 A1.n0 A1.t1 163.721
R99 A1.n1 A1.n0 152
R100 A1 A1.n1 10.736
R101 A1.n1 A1 8.25856
R102 a_458_47.t0 a_458_47.t1 72.0005
R103 a_566_47.t0 a_566_47.n0 274.149
R104 a_566_47.n0 a_566_47.t1 36.9236
R105 a_566_47.n0 a_566_47.t2 35.0774
C0 VGND D1 0.016542f
C1 VPWR B1 0.018374f
C2 A1 A2 0.087542f
C3 VPB D1 0.039539f
C4 VPWR VGND 0.106139f
C5 VPWR VPB 0.107888f
C6 D1 C1 0.115599f
C7 X D1 3.91e-19
C8 VPWR C1 0.020249f
C9 B1 A2 0.088285f
C10 A1 VGND 0.025113f
C11 VPWR X 0.155541f
C12 VGND A2 0.019732f
C13 A1 VPB 0.062872f
C14 VPB A2 0.035689f
C15 VPWR D1 0.02075f
C16 A1 C1 1.89e-19
C17 C1 A2 0.002803f
C18 VGND B1 0.019995f
C19 VPB B1 0.034184f
C20 VGND VPB 0.009192f
C21 D1 A2 1.6e-19
C22 C1 B1 0.083881f
C23 A1 VPWR 0.14498f
C24 VPWR A2 0.110679f
C25 VGND C1 0.058866f
C26 VPB C1 0.032235f
C27 X VGND 0.126316f
C28 X VPB 0.004531f
C29 VGND VNB 0.571881f
C30 X VNB 0.02426f
C31 VPWR VNB 0.47858f
C32 A1 VNB 0.190086f
C33 A2 VNB 0.098744f
C34 B1 VNB 0.099056f
C35 C1 VNB 0.103335f
C36 D1 VNB 0.106929f
C37 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_1 VNB VPB VPWR VGND X D1 C1 B1 A2 A1
X0 a_676_297.t0 A2.t0 a_79_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X1 a_512_47.t2 B1.t0 a_409_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X2 a_306_47.t1 D1.t0 a_79_21.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VGND.t0 A2.t1 a_512_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X4 VPWR.t2 C1.t0 a_79_21.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X5 a_79_21.t3 B1.t1 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR.t1 A1.t0 a_676_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47.t1 A1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_409_47.t1 C1.t1 a_306_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X9 VPWR.t4 a_79_21.t5 X.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21.t4 D1.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X11 VGND.t2 a_79_21.t6 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t0 241.439
R1 A2.n0 A2.t1 169.138
R2 A2 A2.n0 159.68
R3 a_79_21.n4 a_79_21.n3 387.012
R4 a_79_21.n3 a_79_21.n2 310.502
R5 a_79_21.n0 a_79_21.t5 234.804
R6 a_79_21.n1 a_79_21.t2 164.025
R7 a_79_21.n0 a_79_21.t6 162.504
R8 a_79_21.n1 a_79_21.n0 152
R9 a_79_21.n3 a_79_21.n1 73.6005
R10 a_79_21.n4 a_79_21.t3 57.1305
R11 a_79_21.n2 a_79_21.t1 44.3255
R12 a_79_21.n2 a_79_21.t4 41.3705
R13 a_79_21.t0 a_79_21.n4 26.5955
R14 a_676_297.t0 a_676_297.t1 41.3705
R15 VPB.t5 VPB.t3 541.59
R16 VPB.t1 VPB.t2 449.844
R17 VPB.t3 VPB.t1 346.262
R18 VPB.t2 VPB.t0 340.344
R19 VPB.t0 VPB.t4 213.084
R20 VPB VPB.t5 192.369
R21 B1.n0 B1.t1 238.194
R22 B1.n0 B1.t0 165.893
R23 B1 B1.n0 158.788
R24 a_409_47.t0 a_409_47.t1 67.3851
R25 a_512_47.n0 a_512_47.t1 411.134
R26 a_512_47.n0 a_512_47.t2 87.6928
R27 a_512_47.t0 a_512_47.n0 24.9236
R28 VNB.t5 VNB.t1 2805.18
R29 VNB.t3 VNB.t0 2164.4
R30 VNB.t4 VNB.t3 1466.67
R31 VNB.t1 VNB.t4 1466.67
R32 VNB.t0 VNB.t2 1196.12
R33 VNB VNB.t5 925.567
R34 D1.n0 D1.t1 241.439
R35 D1.n0 D1.t0 169.138
R36 D1 D1.n0 156.864
R37 a_306_47.t0 a_306_47.t1 67.3851
R38 VGND.n1 VGND.t2 289.567
R39 VGND.n1 VGND.n0 207.894
R40 VGND.n0 VGND.t1 24.9236
R41 VGND.n0 VGND.t0 24.9236
R42 VGND VGND.n1 0.149674
R43 C1.n0 C1.t0 241.439
R44 C1.n0 C1.t1 169.138
R45 C1 C1.n0 154.607
R46 VPWR.n5 VPWR.t1 344.557
R47 VPWR.n12 VPWR.n11 292.5
R48 VPWR.n10 VPWR.n9 292.5
R49 VPWR.n4 VPWR.n3 146.25
R50 VPWR.n11 VPWR.n10 94.5605
R51 VPWR.n3 VPWR.t0 60.0855
R52 VPWR.n3 VPWR.t2 60.0855
R53 VPWR.n8 VPWR.n2 31.5309
R54 VPWR.n11 VPWR.t4 28.5655
R55 VPWR.n10 VPWR.t3 27.5805
R56 VPWR.n9 VPWR.n8 22.8837
R57 VPWR.n6 VPWR.n2 9.3005
R58 VPWR.n8 VPWR.n7 9.3005
R59 VPWR.n1 VPWR.n0 9.3005
R60 VPWR.n5 VPWR.n4 9.22783
R61 VPWR.n13 VPWR.n12 7.26884
R62 VPWR.n12 VPWR.n1 6.0706
R63 VPWR.n4 VPWR.n2 3.69535
R64 VPWR.n9 VPWR.n1 0.264418
R65 VPWR.n6 VPWR.n5 0.255643
R66 VPWR.n13 VPWR.n0 0.146635
R67 VPWR.n7 VPWR.n6 0.120292
R68 VPWR.n7 VPWR.n0 0.120292
R69 VPWR VPWR.n13 0.116751
R70 A1.n0 A1.t0 234.213
R71 A1.n0 A1.t1 161.912
R72 A1.n1 A1.n0 152
R73 A1.n1 A1 11.055
R74 A1 A1.n1 2.13383
R75 X.n0 X 593.615
R76 X.n1 X.n0 585
R77 X X.t1 249.863
R78 X.n0 X.t0 26.5955
R79 X X.n1 8.61589
R80 X.n1 X 8.12358
C0 C1 B1 0.103764f
C1 D1 A2 1.08e-19
C2 VPWR VPB 0.088082f
C3 B1 A1 6.19e-19
C4 D1 VPWR 0.02327f
C5 A2 VGND 0.019125f
C6 B1 VPB 0.037747f
C7 VPWR VGND 0.086487f
C8 X VPB 0.010766f
C9 D1 X 3.34e-19
C10 A2 VPWR 0.084842f
C11 B1 VGND 0.032502f
C12 C1 VPB 0.034717f
C13 X VGND 0.065417f
C14 A1 VPB 0.040014f
C15 D1 C1 0.118164f
C16 B1 A2 0.053374f
C17 B1 VPWR 0.021829f
C18 C1 VGND 0.034208f
C19 D1 VPB 0.036506f
C20 X VPWR 0.094894f
C21 A1 VGND 0.018355f
C22 C1 A2 2.05e-19
C23 VGND VPB 0.007973f
C24 D1 VGND 0.038682f
C25 A2 A1 0.121151f
C26 C1 VPWR 0.021694f
C27 A2 VPB 0.035254f
C28 A1 VPWR 0.054995f
C29 VGND VNB 0.490847f
C30 VPWR VNB 0.414323f
C31 X VNB 0.090669f
C32 A1 VNB 0.153752f
C33 A2 VNB 0.104137f
C34 B1 VNB 0.113872f
C35 C1 VNB 0.098766f
C36 D1 VNB 0.112426f
C37 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_4 VGND VPWR VPB VNB A1 A2 A3 B1 C1 Y
X0 a_39_297.t7 A1.t0 VPWR.t9 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t11 C1.t0 VPWR.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t8 A1.t1 a_39_297.t6 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t11 B1.t0 Y.t14 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X4 a_125_47.t5 A3.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X5 a_125_47.t9 A1.t2 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_125_47.t10 A2.t0 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_1163_47.t7 B1.t1 a_125_47.t14 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_39_297.t5 A1.t3 VPWR.t7 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1163_47.t6 B1.t2 a_125_47.t13 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t4 A3.t1 a_125_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t5 C1.t1 Y.t10 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t8 A1.t4 a_125_47.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t3 A3.t2 a_125_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_39_297.t3 A2.t1 a_461_297.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t7 A1.t5 a_125_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_125_47.t12 B1.t3 a_1163_47.t5 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X17 Y.t9 C1.t2 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_125_47.t6 A1.t6 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 VGND.t11 A2.t2 a_125_47.t11 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_125_47.t15 B1.t4 a_1163_47.t4 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t0 A2.t3 a_125_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t13 C1.t3 a_1163_47.t3 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y.t12 C1.t4 a_1163_47.t2 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_461_297.t6 A2.t4 a_39_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t5 A3.t3 a_461_297.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR.t10 C1.t5 Y.t8 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t0 A3.t4 a_461_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y.t2 B1.t5 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_125_47.t2 A3.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR.t6 A1.t7 a_39_297.t4 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X31 a_461_297.t1 A3.t6 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_461_297.t0 A3.t7 Y.t15 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 VPWR.t2 B1.t6 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_125_47.t1 A2.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_1163_47.t1 C1.t6 Y.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 a_1163_47.t0 C1.t7 Y.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 Y.t4 B1.t7 VPWR.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 a_39_297.t1 A2.t6 a_461_297.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 a_461_297.t4 A2.t7 a_39_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A1.n1 A1.t0 221.72
R1 A1.n3 A1.t1 221.72
R2 A1.n0 A1.t3 221.72
R3 A1.n8 A1.t7 221.72
R4 A1.n2 A1 156.431
R5 A1.n5 A1.n4 152
R6 A1.n7 A1.n6 152
R7 A1.n10 A1.n9 152
R8 A1.n1 A1.t5 149.421
R9 A1.n3 A1.t2 149.421
R10 A1.n0 A1.t4 149.421
R11 A1.n8 A1.t6 149.421
R12 A1.n9 A1.n7 60.6968
R13 A1.n4 A1.n0 50.8783
R14 A1.n2 A1.n1 38.382
R15 A1.n3 A1.n2 36.5968
R16 A1.n4 A1.n3 24.1005
R17 A1 A1.n10 22.1543
R18 A1.n6 A1 16.2467
R19 A1.n5 A1 12.3082
R20 A1 A1.n5 10.339
R21 A1.n7 A1.n0 9.81902
R22 A1.n6 A1 6.4005
R23 A1.n9 A1.n8 4.46346
R24 A1.n10 A1 0.492808
R25 VPWR.n15 VPWR.n14 314.904
R26 VPWR.n36 VPWR.n3 309.726
R27 VPWR.n9 VPWR.n8 309.726
R28 VPWR.n18 VPWR.n11 309.726
R29 VPWR.n13 VPWR.n12 309.726
R30 VPWR.n38 VPWR.n1 309.724
R31 VPWR.n24 VPWR.n23 34.6358
R32 VPWR.n25 VPWR.n24 34.6358
R33 VPWR.n25 VPWR.n6 34.6358
R34 VPWR.n29 VPWR.n6 34.6358
R35 VPWR.n30 VPWR.n29 34.6358
R36 VPWR.n31 VPWR.n30 34.6358
R37 VPWR.n31 VPWR.n4 34.6358
R38 VPWR.n35 VPWR.n4 34.6358
R39 VPWR.n23 VPWR.n9 32.0005
R40 VPWR.n1 VPWR.t7 26.5955
R41 VPWR.n1 VPWR.t6 26.5955
R42 VPWR.n3 VPWR.t9 26.5955
R43 VPWR.n3 VPWR.t8 26.5955
R44 VPWR.n8 VPWR.t3 26.5955
R45 VPWR.n8 VPWR.t11 26.5955
R46 VPWR.n11 VPWR.t1 26.5955
R47 VPWR.n11 VPWR.t2 26.5955
R48 VPWR.n12 VPWR.t0 26.5955
R49 VPWR.n12 VPWR.t10 26.5955
R50 VPWR.n14 VPWR.t4 26.5955
R51 VPWR.n14 VPWR.t5 26.5955
R52 VPWR.n19 VPWR.n18 25.977
R53 VPWR.n36 VPWR.n35 22.9652
R54 VPWR.n37 VPWR.n36 21.4593
R55 VPWR.n17 VPWR.n13 19.9534
R56 VPWR.n18 VPWR.n17 18.4476
R57 VPWR.n38 VPWR.n37 16.9417
R58 VPWR.n19 VPWR.n9 12.424
R59 VPWR.n17 VPWR.n16 9.3005
R60 VPWR.n18 VPWR.n10 9.3005
R61 VPWR.n20 VPWR.n19 9.3005
R62 VPWR.n21 VPWR.n9 9.3005
R63 VPWR.n23 VPWR.n22 9.3005
R64 VPWR.n24 VPWR.n7 9.3005
R65 VPWR.n26 VPWR.n25 9.3005
R66 VPWR.n27 VPWR.n6 9.3005
R67 VPWR.n29 VPWR.n28 9.3005
R68 VPWR.n30 VPWR.n5 9.3005
R69 VPWR.n32 VPWR.n31 9.3005
R70 VPWR.n33 VPWR.n4 9.3005
R71 VPWR.n35 VPWR.n34 9.3005
R72 VPWR.n36 VPWR.n2 9.3005
R73 VPWR.n37 VPWR.n0 9.3005
R74 VPWR.n39 VPWR.n38 7.4049
R75 VPWR.n15 VPWR.n13 6.60089
R76 VPWR.n16 VPWR.n15 0.679611
R77 VPWR.n39 VPWR.n0 0.144904
R78 VPWR VPWR.n39 0.123712
R79 VPWR.n16 VPWR.n10 0.120292
R80 VPWR.n20 VPWR.n10 0.120292
R81 VPWR.n21 VPWR.n20 0.120292
R82 VPWR.n22 VPWR.n21 0.120292
R83 VPWR.n22 VPWR.n7 0.120292
R84 VPWR.n26 VPWR.n7 0.120292
R85 VPWR.n27 VPWR.n26 0.120292
R86 VPWR.n28 VPWR.n27 0.120292
R87 VPWR.n28 VPWR.n5 0.120292
R88 VPWR.n32 VPWR.n5 0.120292
R89 VPWR.n33 VPWR.n32 0.120292
R90 VPWR.n34 VPWR.n33 0.120292
R91 VPWR.n34 VPWR.n2 0.120292
R92 VPWR.n2 VPWR.n0 0.120292
R93 a_39_297.n2 a_39_297.t3 764.827
R94 a_39_297.n2 a_39_297.n1 591.777
R95 a_39_297.n4 a_39_297.t4 405.406
R96 a_39_297.n3 a_39_297.n0 305.539
R97 a_39_297.n5 a_39_297.n4 305.539
R98 a_39_297.n3 a_39_297.n2 44.8005
R99 a_39_297.n4 a_39_297.n3 44.8005
R100 a_39_297.n1 a_39_297.t0 26.5955
R101 a_39_297.n1 a_39_297.t1 26.5955
R102 a_39_297.n0 a_39_297.t2 26.5955
R103 a_39_297.n0 a_39_297.t7 26.5955
R104 a_39_297.t6 a_39_297.n5 26.5955
R105 a_39_297.n5 a_39_297.t5 26.5955
R106 VPB.t9 VPB.t19 556.386
R107 VPB.t10 VPB.t18 260.437
R108 VPB VPB.t13 251.559
R109 VPB.t12 VPB.t11 248.599
R110 VPB.t5 VPB.t12 248.599
R111 VPB.t17 VPB.t5 248.599
R112 VPB.t6 VPB.t17 248.599
R113 VPB.t7 VPB.t6 248.599
R114 VPB.t8 VPB.t7 248.599
R115 VPB.t18 VPB.t8 248.599
R116 VPB.t1 VPB.t10 248.599
R117 VPB.t0 VPB.t1 248.599
R118 VPB.t19 VPB.t0 248.599
R119 VPB.t2 VPB.t9 248.599
R120 VPB.t3 VPB.t2 248.599
R121 VPB.t4 VPB.t3 248.599
R122 VPB.t16 VPB.t4 248.599
R123 VPB.t15 VPB.t16 248.599
R124 VPB.t14 VPB.t15 248.599
R125 VPB.t13 VPB.t14 248.599
R126 C1.n9 C1.t5 228.862
R127 C1.n1 C1.t0 221.72
R128 C1.n5 C1.t1 221.72
R129 C1.n8 C1.t2 221.72
R130 C1.n1 C1.t7 156.561
R131 C1.n3 C1.n2 152
R132 C1.n6 C1.n0 152
R133 C1.n11 C1.n10 152
R134 C1.n9 C1.t3 149.421
R135 C1.n7 C1.t6 149.421
R136 C1.n4 C1.t4 149.421
R137 C1.n3 C1.n1 64.2672
R138 C1.n6 C1.n5 49.9857
R139 C1.n10 C1.n8 35.7042
R140 C1.n10 C1.n9 32.1338
R141 C1.n7 C1.n6 17.8524
R142 C1.n11 C1.n0 16.739
R143 C1.n2 C1 13.0467
R144 C1.n2 C1 9.6005
R145 C1.n5 C1.n4 7.14124
R146 C1.n8 C1.n7 7.14124
R147 C1 C1.n0 3.69281
R148 C1.n4 C1.n3 3.57087
R149 C1 C1.n11 2.21588
R150 Y.n9 Y.t15 764.827
R151 Y.n9 Y.n8 591.777
R152 Y.n14 Y.t11 354.565
R153 Y.n13 Y.n4 305.539
R154 Y.n12 Y.n5 305.539
R155 Y.n11 Y.n6 305.539
R156 Y.n10 Y.n7 304.18
R157 Y.n2 Y.n0 231.749
R158 Y.n2 Y.n1 185
R159 Y.n11 Y.n10 45.3338
R160 Y.n10 Y.n9 45.3338
R161 Y.n13 Y.n12 44.8005
R162 Y.n12 Y.n11 44.8005
R163 Y.n15 Y.n13 40.2672
R164 Y.n7 Y.t14 30.5355
R165 Y.n4 Y.t10 26.5955
R166 Y.n4 Y.t9 26.5955
R167 Y.n5 Y.t8 26.5955
R168 Y.n5 Y.t2 26.5955
R169 Y.n6 Y.t3 26.5955
R170 Y.n6 Y.t4 26.5955
R171 Y.n7 Y.t5 26.5955
R172 Y.n8 Y.t1 26.5955
R173 Y.n8 Y.t0 26.5955
R174 Y.n0 Y.t7 24.9236
R175 Y.n0 Y.t13 24.9236
R176 Y.n1 Y.t6 24.9236
R177 Y.n1 Y.t12 24.9236
R178 Y.n3 Y.n2 20.0353
R179 Y Y.n3 13.6132
R180 Y Y.n14 6.19103
R181 Y.n15 Y 6.06366
R182 Y.n14 Y 5.18783
R183 Y.n16 Y.n15 4.04261
R184 Y.n16 Y 1.6259
R185 Y Y.n16 1.34787
R186 Y.n3 Y 0.203675
R187 B1.n11 B1.t0 228.862
R188 B1.n1 B1.t5 221.72
R189 B1.n2 B1.t6 221.72
R190 B1.n10 B1.t7 221.72
R191 B1.n1 B1.t2 156.561
R192 B1.n5 B1.n4 152
R193 B1.n6 B1.n0 152
R194 B1.n8 B1.n7 152
R195 B1.n13 B1.n12 152
R196 B1.n11 B1.t3 149.421
R197 B1.n9 B1.t1 149.421
R198 B1.n3 B1.t4 149.421
R199 B1.n8 B1.n0 60.6968
R200 B1.n4 B1.n3 50.8783
R201 B1.n12 B1.n10 49.0931
R202 B1.n12 B1.n11 18.7449
R203 B1.n4 B1.n1 16.9598
R204 B1.n7 B1.n6 16.739
R205 B1.n13 B1 16.2467
R206 B1.n5 B1 11.3236
R207 B1 B1.n5 11.3236
R208 B1.n3 B1.n2 7.14124
R209 B1.n10 B1.n9 7.14124
R210 B1 B1.n13 6.4005
R211 B1.n6 B1 5.41588
R212 B1.n9 B1.n8 4.46346
R213 B1.n2 B1.n0 2.67828
R214 B1.n7 B1 0.492808
R215 A3.n3 A3.t3 277.062
R216 A3.n2 A3.t6 221.72
R217 A3.n7 A3.t4 221.72
R218 A3.n0 A3.t7 221.72
R219 A3.n14 A3.t0 165.488
R220 A3.n4 A3.n3 152
R221 A3.n6 A3.n5 152
R222 A3.n10 A3.n9 152
R223 A3.n12 A3.n11 152
R224 A3.n15 A3.n14 152
R225 A3.n13 A3.t2 149.421
R226 A3.n8 A3.t5 149.421
R227 A3.n1 A3.t1 149.421
R228 A3.n14 A3.n13 58.9116
R229 A3.n9 A3.n0 48.2005
R230 A3.n7 A3.n6 33.919
R231 A3.n6 A3.n1 26.7783
R232 A3.n3 A3.n2 19.6375
R233 A3.n11 A3.n10 16.739
R234 A3.n5 A3 14.5236
R235 A3.n2 A3.n1 14.282
R236 A3.n8 A3.n7 14.282
R237 A3.n4 A3 14.0313
R238 A3.n15 A3 13.0467
R239 A3.n9 A3.n8 12.4968
R240 A3.n12 A3.n0 12.4968
R241 A3 A3.n15 9.6005
R242 A3 A3.n4 8.61589
R243 A3.n5 A3 8.12358
R244 A3.n11 A3 3.69281
R245 A3.n10 A3 2.21588
R246 A3.n13 A3.n12 1.78569
R247 VGND.n7 VGND.t4 288.154
R248 VGND.n9 VGND.n8 198.964
R249 VGND.n17 VGND.n5 198.964
R250 VGND.n20 VGND.n19 198.964
R251 VGND.n24 VGND.n2 198.964
R252 VGND.n12 VGND.n11 198.167
R253 VGND.n26 VGND.t6 142.38
R254 VGND.n13 VGND.n10 34.6358
R255 VGND.n17 VGND.n4 32.0005
R256 VGND.n11 VGND.t0 28.6159
R257 VGND.n20 VGND.n18 25.977
R258 VGND.n8 VGND.t2 24.9236
R259 VGND.n8 VGND.t3 24.9236
R260 VGND.n11 VGND.t5 24.9236
R261 VGND.n5 VGND.t1 24.9236
R262 VGND.n5 VGND.t11 24.9236
R263 VGND.n19 VGND.t10 24.9236
R264 VGND.n19 VGND.t7 24.9236
R265 VGND.n2 VGND.t9 24.9236
R266 VGND.n2 VGND.t8 24.9236
R267 VGND.n25 VGND.n24 24.4711
R268 VGND.n24 VGND.n1 19.9534
R269 VGND.n20 VGND.n1 18.4476
R270 VGND.n9 VGND.n7 14.0348
R271 VGND.n26 VGND.n25 13.9299
R272 VGND.n18 VGND.n17 12.424
R273 VGND.n27 VGND.n26 9.3005
R274 VGND.n10 VGND.n6 9.3005
R275 VGND.n14 VGND.n13 9.3005
R276 VGND.n15 VGND.n4 9.3005
R277 VGND.n17 VGND.n16 9.3005
R278 VGND.n18 VGND.n3 9.3005
R279 VGND.n21 VGND.n20 9.3005
R280 VGND.n22 VGND.n1 9.3005
R281 VGND.n24 VGND.n23 9.3005
R282 VGND.n25 VGND.n0 9.3005
R283 VGND.n12 VGND.n4 6.4005
R284 VGND.n10 VGND.n9 1.88285
R285 VGND.n13 VGND.n12 1.88285
R286 VGND.n7 VGND.n6 1.42397
R287 VGND.n14 VGND.n6 0.120292
R288 VGND.n15 VGND.n14 0.120292
R289 VGND.n16 VGND.n15 0.120292
R290 VGND.n16 VGND.n3 0.120292
R291 VGND.n21 VGND.n3 0.120292
R292 VGND.n22 VGND.n21 0.120292
R293 VGND.n23 VGND.n22 0.120292
R294 VGND.n23 VGND.n0 0.120292
R295 VGND.n27 VGND.n0 0.120292
R296 VGND VGND.n27 0.0278438
R297 a_125_47.n9 a_125_47.n8 238.901
R298 a_125_47.n3 a_125_47.n1 231.749
R299 a_125_47.n9 a_125_47.n7 192.154
R300 a_125_47.n10 a_125_47.n6 192.154
R301 a_125_47.n11 a_125_47.n5 192.154
R302 a_125_47.n4 a_125_47.n0 192.154
R303 a_125_47.n13 a_125_47.n12 192.154
R304 a_125_47.n3 a_125_47.n2 185
R305 a_125_47.n4 a_125_47.n3 77.9135
R306 a_125_47.n12 a_125_47.n11 47.8614
R307 a_125_47.n12 a_125_47.n4 46.7483
R308 a_125_47.n11 a_125_47.n10 46.7483
R309 a_125_47.n10 a_125_47.n9 46.7483
R310 a_125_47.n2 a_125_47.t14 24.9236
R311 a_125_47.n2 a_125_47.t12 24.9236
R312 a_125_47.n1 a_125_47.t13 24.9236
R313 a_125_47.n1 a_125_47.t15 24.9236
R314 a_125_47.n8 a_125_47.t8 24.9236
R315 a_125_47.n8 a_125_47.t6 24.9236
R316 a_125_47.n7 a_125_47.t7 24.9236
R317 a_125_47.n7 a_125_47.t9 24.9236
R318 a_125_47.n6 a_125_47.t11 24.9236
R319 a_125_47.n6 a_125_47.t10 24.9236
R320 a_125_47.n5 a_125_47.t0 24.9236
R321 a_125_47.n5 a_125_47.t1 24.9236
R322 a_125_47.n0 a_125_47.t4 24.9236
R323 a_125_47.n0 a_125_47.t2 24.9236
R324 a_125_47.n13 a_125_47.t3 24.9236
R325 a_125_47.t5 a_125_47.n13 24.9236
R326 VNB.t4 VNB.t17 2790.94
R327 VNB.t0 VNB.t5 1253.07
R328 VNB VNB.t6 1210.36
R329 VNB.t13 VNB.t11 1196.12
R330 VNB.t12 VNB.t13 1196.12
R331 VNB.t14 VNB.t12 1196.12
R332 VNB.t18 VNB.t14 1196.12
R333 VNB.t16 VNB.t18 1196.12
R334 VNB.t19 VNB.t16 1196.12
R335 VNB.t17 VNB.t19 1196.12
R336 VNB.t2 VNB.t4 1196.12
R337 VNB.t3 VNB.t2 1196.12
R338 VNB.t5 VNB.t3 1196.12
R339 VNB.t1 VNB.t0 1196.12
R340 VNB.t15 VNB.t1 1196.12
R341 VNB.t10 VNB.t15 1196.12
R342 VNB.t7 VNB.t10 1196.12
R343 VNB.t9 VNB.t7 1196.12
R344 VNB.t8 VNB.t9 1196.12
R345 VNB.t6 VNB.t8 1196.12
R346 A2.n1 A2.t1 221.72
R347 A2.n2 A2.t4 221.72
R348 A2.n8 A2.t6 221.72
R349 A2.n9 A2.t7 221.72
R350 A2.n4 A2.n3 152
R351 A2.n5 A2.n0 152
R352 A2.n7 A2.n6 152
R353 A2.n11 A2.n10 152
R354 A2.n1 A2.t3 149.421
R355 A2.n2 A2.t5 149.421
R356 A2.n8 A2.t2 149.421
R357 A2.n9 A2.t0 149.421
R358 A2.n7 A2.n0 60.6968
R359 A2.n10 A2.n8 58.9116
R360 A2.n3 A2.n2 48.2005
R361 A2.n3 A2.n1 26.7783
R362 A2 A2.n11 17.4774
R363 A2.n5 A2.n4 16.739
R364 A2.n10 A2.n9 16.0672
R365 A2.n2 A2.n0 12.4968
R366 A2.n6 A2 11.5697
R367 A2.n6 A2 11.0774
R368 A2 A2.n5 5.66204
R369 A2.n11 A2 5.16973
R370 A2.n8 A2.n7 1.78569
R371 A2.n4 A2 0.246654
R372 a_1163_47.n3 a_1163_47.t5 317.462
R373 a_1163_47.n1 a_1163_47.t0 317.462
R374 a_1163_47.n1 a_1163_47.n0 185
R375 a_1163_47.n3 a_1163_47.n2 185
R376 a_1163_47.n5 a_1163_47.n4 96.3779
R377 a_1163_47.n4 a_1163_47.n1 46.7483
R378 a_1163_47.n4 a_1163_47.n3 46.7483
R379 a_1163_47.n2 a_1163_47.t4 24.9236
R380 a_1163_47.n2 a_1163_47.t7 24.9236
R381 a_1163_47.n0 a_1163_47.t2 24.9236
R382 a_1163_47.n0 a_1163_47.t1 24.9236
R383 a_1163_47.t3 a_1163_47.n5 24.9236
R384 a_1163_47.n5 a_1163_47.t6 24.9236
R385 a_461_297.n5 a_461_297.n4 334.938
R386 a_461_297.n2 a_461_297.n0 334.937
R387 a_461_297.n2 a_461_297.n1 296.538
R388 a_461_297.n4 a_461_297.n3 296.538
R389 a_461_297.n4 a_461_297.n2 77.5534
R390 a_461_297.n0 a_461_297.t5 26.5955
R391 a_461_297.n0 a_461_297.t4 26.5955
R392 a_461_297.n1 a_461_297.t7 26.5955
R393 a_461_297.n1 a_461_297.t6 26.5955
R394 a_461_297.n3 a_461_297.t2 26.5955
R395 a_461_297.n3 a_461_297.t0 26.5955
R396 a_461_297.t3 a_461_297.n5 26.5955
R397 a_461_297.n5 a_461_297.t1 26.5955
C0 VPB A2 0.122537f
C1 A3 Y 0.201311f
C2 B1 VPWR 0.077928f
C3 A1 A2 0.075533f
C4 A3 VGND 0.061197f
C5 B1 Y 0.193705f
C6 C1 VPWR 0.079176f
C7 B1 VGND 0.03403f
C8 C1 Y 0.320879f
C9 VPB VPWR 0.178593f
C10 A3 B1 0.059934f
C11 C1 VGND 0.033685f
C12 VPB Y 0.037472f
C13 A1 VPWR 0.081559f
C14 A1 Y 3.33e-20
C15 VPB VGND 0.014789f
C16 A2 VPWR 0.035056f
C17 B1 C1 0.078554f
C18 VPB A3 0.14912f
C19 A1 VGND 0.111166f
C20 A2 Y 9.85e-20
C21 VPB B1 0.118953f
C22 A2 VGND 0.059853f
C23 VPB C1 0.122801f
C24 A2 A3 0.057131f
C25 VPWR Y 0.739576f
C26 VPWR VGND 0.184622f
C27 VPB A1 0.125059f
C28 A3 VPWR 0.032442f
C29 Y VGND 0.037989f
C30 VGND VNB 1.04753f
C31 Y VNB 0.110271f
C32 VPWR VNB 0.850012f
C33 C1 VNB 0.382686f
C34 B1 VNB 0.364259f
C35 A3 VNB 0.411068f
C36 A2 VNB 0.357438f
C37 A1 VNB 0.400628f
C38 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_2 VGND VPWR VPB VNB Y B1 C1 A1 A2 A3
X0 VPWR.t2 A1.t0 a_51_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_55_47.t2 A1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t7 C1.t0 a_729_47.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t4 C1.t1 Y.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.205 ps=1.41 w=1 l=0.15
X4 Y.t4 C1.t2 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_55_47.t6 A3.t0 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23075 ps=1.36 w=0.65 l=0.15
X6 VGND.t1 A1.t2 a_55_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_55_47.t5 B1.t0 a_729_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND.t3 A2.t0 a_55_47.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t2 B1.t1 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.305 ps=1.61 w=1 l=0.15
X10 VGND.t0 A3.t1 a_55_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.23075 pd=1.36 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_729_47.t1 C1.t3 Y.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 a_51_297.t3 A2.t1 a_301_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_729_47.t0 B1.t2 a_55_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_301_297.t2 A2.t2 a_51_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_55_47.t7 A2.t3 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t0 B1.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X17 a_51_297.t1 A1.t3 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t0 A3.t2 a_301_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_301_297.t0 A3.t3 Y.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R0 A1.n3 A1.t0 223.506
R1 A1.n0 A1.t3 221.72
R2 A1 A1.n1 168.493
R3 A1.n0 A1.t1 152.99
R4 A1.n4 A1.n3 152
R5 A1.n2 A1.t2 149.421
R6 A1.n2 A1.n1 58.9116
R7 A1.n4 A1 22.4005
R8 A1.n1 A1.n0 12.4968
R9 A1.n3 A1.n2 1.78569
R10 A1 A1.n4 0.246654
R11 a_51_297.n0 a_51_297.t3 764.827
R12 a_51_297.n0 a_51_297.t2 407.087
R13 a_51_297.n1 a_51_297.n0 305.539
R14 a_51_297.t0 a_51_297.n1 26.5955
R15 a_51_297.n1 a_51_297.t1 26.5955
R16 VPWR.n8 VPWR.n5 314.938
R17 VPWR.n19 VPWR.n1 309.724
R18 VPWR.n7 VPWR.n6 146.25
R19 VPWR.n6 VPWR.t3 60.0855
R20 VPWR.n6 VPWR.t0 60.0855
R21 VPWR.n12 VPWR.n11 34.6358
R22 VPWR.n13 VPWR.n12 34.6358
R23 VPWR.n13 VPWR.n2 34.6358
R24 VPWR.n17 VPWR.n2 34.6358
R25 VPWR.n18 VPWR.n17 34.6358
R26 VPWR.n1 VPWR.t1 26.5955
R27 VPWR.n1 VPWR.t2 26.5955
R28 VPWR.n5 VPWR.t5 26.5955
R29 VPWR.n5 VPWR.t4 26.5955
R30 VPWR.n11 VPWR.n4 20.2472
R31 VPWR.n19 VPWR.n18 13.9299
R32 VPWR.n8 VPWR.n7 13.7082
R33 VPWR.n9 VPWR.n4 9.3005
R34 VPWR.n11 VPWR.n10 9.3005
R35 VPWR.n12 VPWR.n3 9.3005
R36 VPWR.n14 VPWR.n13 9.3005
R37 VPWR.n15 VPWR.n2 9.3005
R38 VPWR.n17 VPWR.n16 9.3005
R39 VPWR.n18 VPWR.n0 9.3005
R40 VPWR.n20 VPWR.n19 7.52093
R41 VPWR.n7 VPWR.n4 1.40709
R42 VPWR.n9 VPWR.n8 0.592533
R43 VPWR.n20 VPWR.n0 0.143429
R44 VPWR.n10 VPWR.n9 0.120292
R45 VPWR.n10 VPWR.n3 0.120292
R46 VPWR.n14 VPWR.n3 0.120292
R47 VPWR.n15 VPWR.n14 0.120292
R48 VPWR.n16 VPWR.n15 0.120292
R49 VPWR.n16 VPWR.n0 0.120292
R50 VPWR VPWR.n20 0.119998
R51 VPB.t7 VPB.t6 556.386
R52 VPB.t1 VPB.t5 449.844
R53 VPB.t5 VPB.t8 331.464
R54 VPB VPB.t4 263.397
R55 VPB.t8 VPB.t9 248.599
R56 VPB.t0 VPB.t1 248.599
R57 VPB.t6 VPB.t0 248.599
R58 VPB.t2 VPB.t7 248.599
R59 VPB.t3 VPB.t2 248.599
R60 VPB.t4 VPB.t3 248.599
R61 VGND.n11 VGND.n2 198.964
R62 VGND.n14 VGND.n13 198.964
R63 VGND.n6 VGND.n5 185
R64 VGND.n4 VGND.n3 185
R65 VGND.n5 VGND.n4 62.7697
R66 VGND.n4 VGND.t4 34.1543
R67 VGND.n5 VGND.t0 34.1543
R68 VGND.n12 VGND.n11 25.977
R69 VGND.n2 VGND.t5 24.9236
R70 VGND.n2 VGND.t3 24.9236
R71 VGND.n13 VGND.t2 24.9236
R72 VGND.n13 VGND.t1 24.9236
R73 VGND.n7 VGND.n1 24.3324
R74 VGND.n11 VGND.n1 18.4476
R75 VGND.n14 VGND.n12 12.424
R76 VGND.n8 VGND.n3 9.76941
R77 VGND.n8 VGND.n7 9.3005
R78 VGND.n9 VGND.n1 9.3005
R79 VGND.n11 VGND.n10 9.3005
R80 VGND.n12 VGND.n0 9.3005
R81 VGND.n6 VGND.n3 7.63559
R82 VGND.n15 VGND.n14 7.57378
R83 VGND.n7 VGND.n6 0.449623
R84 VGND.n15 VGND.n0 0.142757
R85 VGND VGND.n15 0.120679
R86 VGND.n9 VGND.n8 0.120292
R87 VGND.n10 VGND.n9 0.120292
R88 VGND.n10 VGND.n0 0.120292
R89 a_55_47.n2 a_55_47.t5 317.462
R90 a_55_47.n4 a_55_47.t1 258.661
R91 a_55_47.n3 a_55_47.n0 192.154
R92 a_55_47.n2 a_55_47.n1 192.154
R93 a_55_47.n5 a_55_47.n4 192.154
R94 a_55_47.n3 a_55_47.n2 71.2353
R95 a_55_47.n4 a_55_47.n3 46.7483
R96 a_55_47.n0 a_55_47.t0 24.9236
R97 a_55_47.n0 a_55_47.t7 24.9236
R98 a_55_47.n1 a_55_47.t3 24.9236
R99 a_55_47.n1 a_55_47.t6 24.9236
R100 a_55_47.n5 a_55_47.t4 24.9236
R101 a_55_47.t2 a_55_47.n5 24.9236
R102 VNB.t6 VNB.t4 2790.94
R103 VNB.t0 VNB.t7 2449.19
R104 VNB VNB.t1 1324.27
R105 VNB.t4 VNB.t8 1196.12
R106 VNB.t3 VNB.t6 1196.12
R107 VNB.t7 VNB.t3 1196.12
R108 VNB.t9 VNB.t0 1196.12
R109 VNB.t5 VNB.t9 1196.12
R110 VNB.t2 VNB.t5 1196.12
R111 VNB.t1 VNB.t2 1196.12
R112 C1.n3 C1.t1 225.291
R113 C1.n2 C1.t2 221.72
R114 C1.n1 C1.n0 187.704
R115 C1.n5 C1.n4 152
R116 C1.n3 C1.t3 149.421
R117 C1.n1 C1.t0 149.421
R118 C1.n4 C1.n3 49.9857
R119 C1.n4 C1.n2 21.4227
R120 C1.n5 C1.n0 16.739
R121 C1.n0 C1 3.69281
R122 C1.n2 C1.n1 3.57087
R123 C1 C1.n5 2.21588
R124 a_729_47.n1 a_729_47.n0 447.913
R125 a_729_47.n0 a_729_47.t2 24.9236
R126 a_729_47.n0 a_729_47.t1 24.9236
R127 a_729_47.n1 a_729_47.t3 24.9236
R128 a_729_47.t0 a_729_47.n1 24.9236
R129 Y.n4 Y.t3 713.808
R130 Y.n1 Y.t4 354.682
R131 Y.n5 Y.n3 305.539
R132 Y.n6 Y.n2 299.685
R133 Y Y.t6 270.892
R134 Y.n0 Y.t7 209.923
R135 Y.n6 Y.n5 66.6672
R136 Y.n5 Y.n4 41.9672
R137 Y.n8 Y.n0 40.4655
R138 Y.n2 Y.t5 40.3855
R139 Y.n2 Y.t2 40.3855
R140 Y.n3 Y.t1 26.5955
R141 Y.n3 Y.t0 26.5955
R142 Y.n8 Y 11.9116
R143 Y Y.n1 5.88349
R144 Y.n1 Y 4.93011
R145 Y.n0 Y 4.54787
R146 Y.n7 Y.n6 3.46717
R147 Y.n4 Y 2.7005
R148 Y Y.n7 1.42272
R149 Y.n7 Y 0.533833
R150 Y Y.n8 0.178278
R151 A3.n1 A3.t2 232.431
R152 A3.n3 A3.t3 221.72
R153 A3.n4 A3.t1 185.125
R154 A3.n2 A3.n0 152
R155 A3.n5 A3.n4 152
R156 A3.n1 A3.t0 149.421
R157 A3.n2 A3.n1 57.1264
R158 A3.n4 A3.n3 53.5561
R159 A3.n5 A3.n0 16.739
R160 A3.n3 A3.n2 7.14124
R161 A3.n0 A3 3.69281
R162 A3 A3.n5 2.21588
R163 B1.n0 B1.t1 291.342
R164 B1.n2 B1.t3 221.72
R165 B1.n0 B1 160.615
R166 B1.n2 B1.t2 160.131
R167 B1.n4 B1.n3 152
R168 B1.n1 B1.t0 149.421
R169 B1.n3 B1.n1 58.9116
R170 B1 B1.n4 14.5236
R171 B1.n4 B1 8.12358
R172 B1.n3 B1.n2 5.35606
R173 B1.n1 B1.n0 1.78569
R174 A2.n3 A2.t2 225.291
R175 A2.n1 A2.t1 221.72
R176 A2 A2.n4 154.215
R177 A2.n1 A2.t3 152.99
R178 A2.n2 A2.n0 152
R179 A2.n3 A2.t0 149.421
R180 A2.n4 A2.n2 60.6968
R181 A2 A2.n0 14.5236
R182 A2.n0 A2 8.12358
R183 A2.n2 A2.n1 5.35606
R184 A2.n4 A2.n3 5.35606
R185 a_301_297.n1 a_301_297.n0 670.626
R186 a_301_297.n0 a_301_297.t3 26.5955
R187 a_301_297.n0 a_301_297.t2 26.5955
R188 a_301_297.t1 a_301_297.n1 26.5955
R189 a_301_297.n1 a_301_297.t0 26.5955
C0 A2 Y 2.31e-19
C1 A3 VPWR 0.022579f
C2 A2 VPB 0.062709f
C3 C1 VGND 0.0203f
C4 VGND A1 0.031165f
C5 A2 VPWR 0.021152f
C6 A2 A3 0.065512f
C7 Y VGND 0.080228f
C8 C1 Y 0.22907f
C9 B1 VGND 0.021441f
C10 Y A1 1.39e-19
C11 B1 C1 0.028229f
C12 VGND VPB 0.011153f
C13 C1 VPB 0.074064f
C14 VPB A1 0.062674f
C15 VPWR VGND 0.115102f
C16 A3 VGND 0.037894f
C17 C1 VPWR 0.038127f
C18 B1 Y 0.146626f
C19 VPWR A1 0.038671f
C20 Y VPB 0.035032f
C21 B1 VPB 0.081954f
C22 VPWR Y 0.459897f
C23 B1 VPWR 0.041039f
C24 A3 Y 0.085144f
C25 A2 VGND 0.033179f
C26 VPWR VPB 0.117985f
C27 A3 B1 0.074874f
C28 A2 A1 0.077228f
C29 A3 VPB 0.08176f
C30 VGND VNB 0.653511f
C31 Y VNB 0.10744f
C32 VPWR VNB 0.549491f
C33 C1 VNB 0.243876f
C34 B1 VNB 0.215495f
C35 A3 VNB 0.224596f
C36 A2 VNB 0.179967f
C37 A1 VNB 0.21914f
C38 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_1 Y C1 B1 A3 A2 A1 VPB VNB VGND VPWR
X0 VGND.t2 A2.t0 a_138_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_138_47.t0 A1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 Y.t1 C1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.185 ps=1.37 w=1 l=0.15
X3 a_138_47.t1 A3.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t3 A3.t1 a_222_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t2 C1.t1 a_458_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 a_222_297.t0 A2.t1 a_138_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t0 B1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X8 a_458_47.t1 B1.t1 a_138_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.19825 ps=1.26 w=0.65 l=0.15
X9 a_138_297.t1 A1.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
R0 A2.n0 A2.t1 241.536
R1 A2.n0 A2.t0 169.237
R2 A2 A2.n0 154.272
R3 a_138_47.n1 a_138_47.n0 449.812
R4 a_138_47.n0 a_138_47.t3 87.6928
R5 a_138_47.n0 a_138_47.t1 24.9236
R6 a_138_47.n1 a_138_47.t2 24.9236
R7 a_138_47.t0 a_138_47.n1 24.9236
R8 VGND.n1 VGND.n0 204.189
R9 VGND.n1 VGND.t0 145.957
R10 VGND.n0 VGND.t1 24.9236
R11 VGND.n0 VGND.t2 24.9236
R12 VGND VGND.n1 0.562176
R13 VNB.t1 VNB.t3 2164.4
R14 VNB VNB.t0 1338.51
R15 VNB.t2 VNB.t1 1196.12
R16 VNB.t0 VNB.t2 1196.12
R17 VNB.t3 VNB.t4 1025.24
R18 A1.n0 A1.t1 231.017
R19 A1.n0 A1.t0 158.716
R20 A1.n1 A1.n0 152
R21 A1.n1 A1 10.0853
R22 A1 A1.n1 7.75808
R23 C1.n0 C1.t0 212.081
R24 C1 C1.n0 203.97
R25 C1.n0 C1.t1 139.78
R26 VPWR.n1 VPWR.n0 318.671
R27 VPWR.n1 VPWR.t2 236.828
R28 VPWR.n0 VPWR.t1 36.4455
R29 VPWR.n0 VPWR.t0 36.4455
R30 VPWR VPWR.n1 0.122103
R31 Y.n5 Y 589.073
R32 Y.n5 Y.n4 585
R33 Y.n6 Y.n5 585
R34 Y.n3 Y.n2 585
R35 Y.n2 Y.n1 292.567
R36 Y.n0 Y.t2 127.621
R37 Y.n5 Y.t0 44.3255
R38 Y.n5 Y.t3 44.3255
R39 Y Y.n6 35.9432
R40 Y.n2 Y.t1 32.5055
R41 Y.n7 Y.n3 19.9534
R42 Y.n8 Y 16.6703
R43 Y.n3 Y 8.81457
R44 Y.n7 Y 7.90638
R45 Y.n1 Y 6.7803
R46 Y.n4 Y 4.07323
R47 Y.n4 Y 3.8405
R48 Y.n6 Y 3.8405
R49 Y Y.n0 3.60106
R50 Y Y.n8 3.57259
R51 Y Y.n7 2.97724
R52 Y.n0 Y 2.65834
R53 Y.n1 Y 2.17881
R54 Y.n8 Y 1.11354
R55 VPB.t2 VPB.t0 355.14
R56 VPB.t0 VPB.t1 307.788
R57 VPB VPB.t4 278.193
R58 VPB.t3 VPB.t2 248.599
R59 VPB.t4 VPB.t3 248.599
R60 A3.n0 A3.t1 241.536
R61 A3.n0 A3.t0 169.237
R62 A3 A3.n0 154.012
R63 a_222_297.t0 a_222_297.t1 53.1905
R64 a_458_47.t0 a_458_47.t1 38.7697
R65 a_138_297.t0 a_138_297.t1 53.1905
R66 B1.n0 B1.t0 237.736
R67 B1.n0 B1.t1 165.435
R68 B1 B1.n0 153.656
C0 VPWR Y 0.292562f
C1 A3 Y 0.044876f
C2 A2 VGND 0.01743f
C3 B1 VPWR 0.017491f
C4 A3 B1 0.059175f
C5 A2 VPB 0.031106f
C6 VGND A1 0.067811f
C7 A3 VPWR 0.010151f
C8 A2 Y 0.08317f
C9 A2 B1 8.69e-19
C10 C1 VGND 0.007959f
C11 VPB A1 0.039018f
C12 VGND VPB 0.007288f
C13 C1 VPB 0.045822f
C14 B1 A1 2.07e-19
C15 A2 VPWR 0.128592f
C16 A2 A3 0.090297f
C17 Y VGND 0.10274f
C18 C1 Y 0.131277f
C19 B1 VGND 0.03582f
C20 B1 C1 0.055969f
C21 Y VPB 0.023565f
C22 VPWR A1 0.084905f
C23 B1 VPB 0.03109f
C24 VPWR VGND 0.066258f
C25 C1 VPWR 0.016966f
C26 A3 VGND 0.016402f
C27 B1 Y 0.112113f
C28 VPWR VPB 0.081179f
C29 A3 VPB 0.028351f
C30 A2 A1 0.086638f
C31 VGND VNB 0.416741f
C32 Y VNB 0.081773f
C33 VPWR VNB 0.361245f
C34 C1 VNB 0.155431f
C35 B1 VNB 0.102431f
C36 A3 VNB 0.09482f
C37 A2 VNB 0.092066f
C38 A1 VNB 0.146547f
C39 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_0 C1 A1 A2 Y B1 A3 VPB VNB VGND VPWR
X0 VGND.t2 A2.t0 a_138_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_138_369.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1792 ps=1.84 w=0.64 l=0.15
X2 a_138_47.t1 A1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3 a_138_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1281 pd=1.03 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 Y.t2 C1.t0 a_458_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 Y.t3 C1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1984 pd=1.9 as=0.1184 ps=1.01 w=0.64 l=0.15
X6 Y.t1 A3.t1 a_222_369.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.144 pd=1.09 as=0.0864 ps=0.91 w=0.64 l=0.15
X7 a_222_369.t0 A2.t1 a_138_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0864 ps=0.91 w=0.64 l=0.15
X8 a_458_47.t0 B1.t0 a_138_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 VPWR.t1 B1.t1 Y.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1184 pd=1.01 as=0.144 ps=1.09 w=0.64 l=0.15
R0 A2.n0 A2.t1 299.377
R1 A2.n0 A2.t0 206.19
R2 A2.n1 A2.n0 152
R3 A2.n1 A2 11.7682
R4 A2 A2.n1 2.27147
R5 a_138_47.n1 a_138_47.n0 464.872
R6 a_138_47.n1 a_138_47.t3 135.714
R7 a_138_47.n0 a_138_47.t2 38.5719
R8 a_138_47.n0 a_138_47.t1 38.5719
R9 a_138_47.t0 a_138_47.n1 38.5719
R10 VGND.n1 VGND.t1 230.663
R11 VGND.n1 VGND.n0 204.16
R12 VGND.n0 VGND.t0 38.5719
R13 VGND.n0 VGND.t2 38.5719
R14 VGND VGND.n1 0.608248
R15 VNB.t0 VNB.t4 2164.4
R16 VNB VNB.t1 1338.51
R17 VNB.t2 VNB.t0 1196.12
R18 VNB.t1 VNB.t2 1196.12
R19 VNB.t4 VNB.t3 1025.24
R20 A1.n0 A1.t0 288.856
R21 A1.n0 A1.t1 195.669
R22 A1.n1 A1.n0 152
R23 A1.n2 A1 6.0706
R24 A1.n1 A1 4.06399
R25 A1 A1.n2 3.65764
R26 A1.n2 A1.n1 1.6259
R27 VPWR.n1 VPWR.t0 365.007
R28 VPWR.n1 VPWR.n0 317.312
R29 VPWR.n0 VPWR.t2 56.9458
R30 VPWR.n0 VPWR.t1 56.9458
R31 VPWR VPWR.n1 0.122103
R32 a_138_369.t0 a_138_369.t1 83.1099
R33 VPB.t4 VPB.t2 355.14
R34 VPB.t2 VPB.t3 307.788
R35 VPB VPB.t0 278.193
R36 VPB.t1 VPB.t4 248.599
R37 VPB.t0 VPB.t1 248.599
R38 A3.n0 A3.t1 299.377
R39 A3.n0 A3.t0 206.19
R40 A3 A3.n0 154.012
R41 C1.n0 C1.t1 269.921
R42 C1 C1.n0 203.97
R43 C1.n0 C1.t0 176.733
R44 a_458_47.t0 a_458_47.t1 60.0005
R45 Y.n1 Y 589.888
R46 Y.n2 Y.n1 585
R47 Y.n0 Y.t3 347.041
R48 Y.n4 Y.t2 223.571
R49 Y.n1 Y.t0 69.2583
R50 Y.n1 Y.t1 69.2583
R51 Y.n3 Y 28.7675
R52 Y Y.n5 10.1214
R53 Y.n5 Y.n4 8.84756
R54 Y.n3 Y 7.90638
R55 Y Y.n0 7.2477
R56 Y Y.n2 4.88777
R57 Y.n4 Y 4.51815
R58 Y.n5 Y 3.95344
R59 Y.n2 Y 3.02595
R60 Y Y.n3 2.97724
R61 Y.n0 Y 1.71906
R62 a_222_369.t0 a_222_369.t1 83.1099
R63 B1.n0 B1.t1 295.575
R64 B1.n0 B1.t0 202.388
R65 B1 B1.n0 153.562
C0 VGND B1 0.039138f
C1 Y C1 0.153495f
C2 VPB B1 0.054925f
C3 A1 A3 4.21e-19
C4 A2 VPWR 0.103923f
C5 Y VGND 0.098221f
C6 VPB Y 0.040399f
C7 A1 A2 0.147954f
C8 Y B1 0.121857f
C9 VGND A3 0.016402f
C10 VPB A3 0.050379f
C11 A1 VPWR 0.083187f
C12 A2 VGND 0.017156f
C13 A3 B1 0.078546f
C14 VPB A2 0.054321f
C15 C1 VPWR 0.017478f
C16 Y A3 0.048739f
C17 VGND VPWR 0.063224f
C18 A2 B1 8.69e-19
C19 VPB VPWR 0.083306f
C20 A1 VGND 0.069118f
C21 A2 Y 0.083062f
C22 VPB A1 0.072628f
C23 B1 VPWR 0.01758f
C24 Y VPWR 0.282811f
C25 VGND C1 0.009918f
C26 A1 B1 0.002957f
C27 VPB C1 0.072878f
C28 A2 A3 0.126689f
C29 VPB VGND 0.008772f
C30 B1 C1 0.089061f
C31 A3 VPWR 0.010151f
C32 VGND VNB 0.410842f
C33 Y VNB 0.075178f
C34 VPWR VNB 0.353852f
C35 C1 VNB 0.194928f
C36 B1 VNB 0.117374f
C37 A3 VNB 0.110462f
C38 A2 VNB 0.104333f
C39 A1 VNB 0.200981f
C40 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311a_4 VPWR VGND VPB VNB X C1 B1 A3 A2 A1
X0 a_79_21.t6 C1.t0 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X1 a_467_47.t3 C1.t1 a_79_21.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t9 A2.t0 a_717_47.t7 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_467_47.t0 B1.t0 a_717_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND.t1 A1.t0 a_717_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t4 a_79_21.t8 X.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X6 a_79_21.t4 C1.t2 a_467_47.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X.t2 a_79_21.t9 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_717_47.t3 B1.t1 a_467_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t2 a_79_21.t10 X.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t4 a_79_21.t11 X.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t3 a_79_21.t12 X.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t7 A3.t0 a_717_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_1147_297.t1 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t0 A1.t2 a_1147_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 X.t5 a_79_21.t13 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_1147_297.t2 A2.t1 a_875_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR.t6 B1.t2 a_79_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21.t0 A3.t1 a_875_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_875_297.t0 A3.t2 a_79_21.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_79_21.t2 B1.t3 VPWR.t7 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_875_297.t2 A2.t2 a_1147_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_717_47.t4 A3.t3 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2015 ps=1.27 w=0.65 l=0.15
X23 a_717_47.t6 A2.t3 VGND.t8 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_717_47.t1 A1.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 X.t0 a_79_21.t14 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 VPWR.t8 C1.t3 a_79_21.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 X.t4 a_79_21.t15 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C1.n1 C1.t0 247.619
R1 C1.n0 C1.t3 221.72
R2 C1.n0 C1.t1 173.065
R3 C1.n3 C1.n2 152
R4 C1.n1 C1.t2 128.534
R5 C1.n2 C1.n1 21.5826
R6 C1 C1.n3 18.2159
R7 C1.n2 C1.n0 12.9498
R8 C1.n3 C1 4.43127
R9 VPWR.n6 VPWR.t6 656.058
R10 VPWR.n8 VPWR.n7 316.269
R11 VPWR.n19 VPWR.n2 309.726
R12 VPWR.n11 VPWR.n5 309.726
R13 VPWR.n21 VPWR.t3 242.871
R14 VPWR.n13 VPWR.n12 146.25
R15 VPWR.n12 VPWR.t9 60.0855
R16 VPWR.n12 VPWR.t4 60.0855
R17 VPWR.n14 VPWR.n11 32.0005
R18 VPWR.n10 VPWR.n6 30.4946
R19 VPWR.n2 VPWR.t5 26.5955
R20 VPWR.n2 VPWR.t2 26.5955
R21 VPWR.n5 VPWR.t7 26.5955
R22 VPWR.n5 VPWR.t8 26.5955
R23 VPWR.n7 VPWR.t1 26.5955
R24 VPWR.n7 VPWR.t0 26.5955
R25 VPWR.n19 VPWR.n18 25.977
R26 VPWR.n21 VPWR.n20 19.9534
R27 VPWR.n20 VPWR.n19 18.4476
R28 VPWR.n18 VPWR.n3 16.5735
R29 VPWR.n11 VPWR.n10 12.424
R30 VPWR.n14 VPWR.n13 11.1126
R31 VPWR.n10 VPWR.n9 9.3005
R32 VPWR.n11 VPWR.n4 9.3005
R33 VPWR.n15 VPWR.n14 9.3005
R34 VPWR.n16 VPWR.n3 9.3005
R35 VPWR.n18 VPWR.n17 9.3005
R36 VPWR.n19 VPWR.n1 9.3005
R37 VPWR.n20 VPWR.n0 9.3005
R38 VPWR.n22 VPWR.n21 9.3005
R39 VPWR.n8 VPWR.n6 7.18487
R40 VPWR.n13 VPWR.n3 0.563137
R41 VPWR.n9 VPWR.n8 0.153725
R42 VPWR.n9 VPWR.n4 0.120292
R43 VPWR.n15 VPWR.n4 0.120292
R44 VPWR.n16 VPWR.n15 0.120292
R45 VPWR.n17 VPWR.n16 0.120292
R46 VPWR.n17 VPWR.n1 0.120292
R47 VPWR.n1 VPWR.n0 0.120292
R48 VPWR.n22 VPWR.n0 0.120292
R49 VPWR VPWR.n22 0.0213333
R50 a_79_21.n2 a_79_21.n1 665.378
R51 a_79_21.n14 a_79_21.n13 305.541
R52 a_79_21.n2 a_79_21.n0 305.539
R53 a_79_21.n12 a_79_21.n3 264.776
R54 a_79_21.n10 a_79_21.t8 212.081
R55 a_79_21.n8 a_79_21.t9 212.081
R56 a_79_21.n6 a_79_21.t10 212.081
R57 a_79_21.n5 a_79_21.t14 212.081
R58 a_79_21.n7 a_79_21.n4 168.738
R59 a_79_21.n11 a_79_21.n10 159.304
R60 a_79_21.n9 a_79_21.n4 152
R61 a_79_21.n10 a_79_21.t12 139.78
R62 a_79_21.n8 a_79_21.t13 139.78
R63 a_79_21.n6 a_79_21.t11 139.78
R64 a_79_21.n5 a_79_21.t15 139.78
R65 a_79_21.n6 a_79_21.n5 61.346
R66 a_79_21.n13 a_79_21.n12 57.6005
R67 a_79_21.n13 a_79_21.n2 44.8005
R68 a_79_21.n10 a_79_21.n9 42.3581
R69 a_79_21.n8 a_79_21.n7 30.6732
R70 a_79_21.n7 a_79_21.n6 30.6732
R71 a_79_21.n1 a_79_21.t3 26.5955
R72 a_79_21.n1 a_79_21.t0 26.5955
R73 a_79_21.n0 a_79_21.t1 26.5955
R74 a_79_21.n0 a_79_21.t2 26.5955
R75 a_79_21.n14 a_79_21.t5 26.5955
R76 a_79_21.t6 a_79_21.n14 26.5955
R77 a_79_21.n3 a_79_21.t7 24.9236
R78 a_79_21.n3 a_79_21.t4 24.9236
R79 a_79_21.n9 a_79_21.n8 18.9884
R80 a_79_21.n11 a_79_21.n4 16.739
R81 a_79_21.n12 a_79_21.n11 3.93896
R82 VPB.t5 VPB.t2 568.225
R83 VPB.t11 VPB.t4 556.386
R84 VPB.t10 VPB.t13 449.844
R85 VPB.t0 VPB.t1 248.599
R86 VPB.t3 VPB.t0 248.599
R87 VPB.t4 VPB.t3 248.599
R88 VPB.t2 VPB.t11 248.599
R89 VPB.t6 VPB.t5 248.599
R90 VPB.t12 VPB.t6 248.599
R91 VPB.t13 VPB.t12 248.599
R92 VPB.t9 VPB.t10 248.599
R93 VPB.t8 VPB.t9 248.599
R94 VPB.t7 VPB.t8 248.599
R95 VPB VPB.t7 189.409
R96 a_467_47.n1 a_467_47.t0 311.086
R97 a_467_47.t2 a_467_47.n1 311.086
R98 a_467_47.n1 a_467_47.n0 96.031
R99 a_467_47.n0 a_467_47.t1 24.9236
R100 a_467_47.n0 a_467_47.t3 24.9236
R101 VNB.t0 VNB.t13 2705.5
R102 VNB.t8 VNB.t11 2677.02
R103 VNB.t13 VNB.t10 2192.88
R104 VNB.t2 VNB.t1 1196.12
R105 VNB.t4 VNB.t2 1196.12
R106 VNB.t3 VNB.t4 1196.12
R107 VNB.t10 VNB.t3 1196.12
R108 VNB.t5 VNB.t0 1196.12
R109 VNB.t12 VNB.t5 1196.12
R110 VNB.t11 VNB.t12 1196.12
R111 VNB.t7 VNB.t8 1196.12
R112 VNB.t9 VNB.t7 1196.12
R113 VNB.t6 VNB.t9 1196.12
R114 VNB VNB.t6 911.327
R115 A2.n0 A2.t1 221.72
R116 A2.n1 A2.t2 221.72
R117 A2.n3 A2.n2 152
R118 A2.n0 A2.t3 149.421
R119 A2.n1 A2.t0 149.421
R120 A2.n2 A2.n0 51.7709
R121 A2.n2 A2.n1 23.2079
R122 A2.n3 A2 19.2005
R123 A2 A2.n3 3.44665
R124 a_717_47.n1 a_717_47.t1 306.592
R125 a_717_47.n4 a_717_47.t5 258.846
R126 a_717_47.n5 a_717_47.n4 235.387
R127 a_717_47.n1 a_717_47.n0 185
R128 a_717_47.n3 a_717_47.n2 185
R129 a_717_47.n4 a_717_47.n3 69.0799
R130 a_717_47.n3 a_717_47.n1 51.2005
R131 a_717_47.n2 a_717_47.t7 24.9236
R132 a_717_47.n2 a_717_47.t4 24.9236
R133 a_717_47.n0 a_717_47.t2 24.9236
R134 a_717_47.n0 a_717_47.t6 24.9236
R135 a_717_47.t0 a_717_47.n5 24.9236
R136 a_717_47.n5 a_717_47.t3 24.9236
R137 VGND.n27 VGND.t3 287.534
R138 VGND.n9 VGND.n8 204.373
R139 VGND.n11 VGND.n10 198.964
R140 VGND.n32 VGND.n2 198.964
R141 VGND.n13 VGND.n6 185
R142 VGND.n15 VGND.n14 185
R143 VGND.n34 VGND.t5 149.232
R144 VGND.n14 VGND.n13 62.7697
R145 VGND.n20 VGND.n19 34.6358
R146 VGND.n21 VGND.n20 34.6358
R147 VGND.n21 VGND.n4 34.6358
R148 VGND.n25 VGND.n4 34.6358
R149 VGND.n26 VGND.n25 34.6358
R150 VGND.n28 VGND.n26 34.6358
R151 VGND.n12 VGND.n11 27.4829
R152 VGND.n32 VGND.n1 25.977
R153 VGND.n14 VGND.t6 25.8467
R154 VGND.n13 VGND.t7 25.8467
R155 VGND.n8 VGND.t0 24.9236
R156 VGND.n8 VGND.t1 24.9236
R157 VGND.n10 VGND.t8 24.9236
R158 VGND.n10 VGND.t9 24.9236
R159 VGND.n2 VGND.t2 24.9236
R160 VGND.n2 VGND.t4 24.9236
R161 VGND.n34 VGND.n33 19.9534
R162 VGND.n33 VGND.n32 18.4476
R163 VGND.n15 VGND.n12 14.6063
R164 VGND.n27 VGND.n1 12.424
R165 VGND.n19 VGND.n6 10.8416
R166 VGND.n35 VGND.n34 9.3005
R167 VGND.n12 VGND.n7 9.3005
R168 VGND.n17 VGND.n16 9.3005
R169 VGND.n19 VGND.n18 9.3005
R170 VGND.n20 VGND.n5 9.3005
R171 VGND.n22 VGND.n21 9.3005
R172 VGND.n23 VGND.n4 9.3005
R173 VGND.n25 VGND.n24 9.3005
R174 VGND.n26 VGND.n3 9.3005
R175 VGND.n29 VGND.n28 9.3005
R176 VGND.n30 VGND.n1 9.3005
R177 VGND.n32 VGND.n31 9.3005
R178 VGND.n33 VGND.n0 9.3005
R179 VGND.n11 VGND.n9 6.17809
R180 VGND.n16 VGND.n6 4.23101
R181 VGND.n28 VGND.n27 3.38874
R182 VGND.n16 VGND.n15 3.14626
R183 VGND.n9 VGND.n7 0.653571
R184 VGND.n17 VGND.n7 0.120292
R185 VGND.n18 VGND.n17 0.120292
R186 VGND.n18 VGND.n5 0.120292
R187 VGND.n22 VGND.n5 0.120292
R188 VGND.n23 VGND.n22 0.120292
R189 VGND.n24 VGND.n23 0.120292
R190 VGND.n24 VGND.n3 0.120292
R191 VGND.n29 VGND.n3 0.120292
R192 VGND.n30 VGND.n29 0.120292
R193 VGND.n31 VGND.n30 0.120292
R194 VGND.n31 VGND.n0 0.120292
R195 VGND.n35 VGND.n0 0.120292
R196 VGND VGND.n35 0.0213333
R197 B1.n1 B1.t3 229.907
R198 B1.n0 B1.t2 184.768
R199 B1.n0 B1.t0 180.661
R200 B1.n3 B1.n2 152
R201 B1.n1 B1.t1 139.78
R202 B1.n2 B1.n1 22.068
R203 B1 B1.n3 16.2467
R204 B1.n3 B1 6.4005
R205 B1.n2 B1.n0 5.80773
R206 A1.n1 A1.t1 237.655
R207 A1.n2 A1.t2 221.72
R208 A1.n1 A1.t3 165.356
R209 A1.n1 A1.n0 152
R210 A1.n4 A1.n3 152
R211 A1.n2 A1.t0 149.421
R212 A1.n3 A1.n2 36.5968
R213 A1.n3 A1.n1 24.9931
R214 A1.n4 A1.n0 16.739
R215 A1 A1.n4 3.2005
R216 A1.n0 A1 2.70819
R217 X.n2 X.n1 350.339
R218 X.n2 X.n0 305.541
R219 X.n5 X.n3 248.248
R220 X.n5 X.n4 185
R221 X.n0 X.t1 26.5955
R222 X.n0 X.t0 26.5955
R223 X.n1 X.t3 26.5955
R224 X.n1 X.t2 26.5955
R225 X X.n6 26.0928
R226 X.n4 X.t7 24.9236
R227 X.n4 X.t4 24.9236
R228 X.n3 X.t6 24.9236
R229 X.n3 X.t5 24.9236
R230 X.n6 X.n2 12.8005
R231 X.n6 X.n5 12.8005
R232 A3.n6 A3.t1 241.357
R233 A3.n4 A3.t2 221.72
R234 A3.n2 A3.t3 176.198
R235 A3.n2 A3.n1 152
R236 A3.n3 A3.n0 152
R237 A3.n7 A3.n6 152
R238 A3.n5 A3.t0 149.421
R239 A3.n3 A3.n2 60.6968
R240 A3.n5 A3.n4 44.6301
R241 A3.n7 A3.n0 16.739
R242 A3.n1 A3 14.2774
R243 A3.n6 A3.n5 10.7116
R244 A3.n1 A3 8.36973
R245 A3.n4 A3.n3 5.35606
R246 A3 A3.n7 3.44665
R247 A3 A3.n0 2.46204
R248 a_1147_297.n1 a_1147_297.t3 764.827
R249 a_1147_297.n1 a_1147_297.n0 591.777
R250 a_1147_297.t1 a_1147_297.n1 410.615
R251 a_1147_297.n0 a_1147_297.t0 26.5955
R252 a_1147_297.n0 a_1147_297.t2 26.5955
R253 a_875_297.n1 a_875_297.t0 748.644
R254 a_875_297.t1 a_875_297.n1 668.432
R255 a_875_297.n1 a_875_297.n0 340.962
R256 a_875_297.n0 a_875_297.t3 26.5955
R257 a_875_297.n0 a_875_297.t2 26.5955
C0 B1 VGND 0.018678f
C1 A1 VGND 0.034035f
C2 C1 VPWR 0.036732f
C3 VPB X 0.008844f
C4 A3 A2 0.06125f
C5 A2 VPWR 0.022022f
C6 C1 VGND 0.020341f
C7 A2 VGND 0.033167f
C8 VPB A3 0.090357f
C9 C1 B1 0.070079f
C10 VPB VPWR 0.164493f
C11 A2 A1 0.074892f
C12 VPWR X 0.356224f
C13 VPB VGND 0.014033f
C14 X VGND 0.262512f
C15 VPB B1 0.066826f
C16 VPB A1 0.066699f
C17 A3 VPWR 0.020228f
C18 VPWR VGND 0.154126f
C19 A3 VGND 0.035285f
C20 VPB C1 0.067237f
C21 VPB A2 0.057852f
C22 B1 A3 0.042298f
C23 B1 VPWR 0.041368f
C24 C1 X 2.75e-19
C25 A1 VPWR 0.040311f
C26 VGND VNB 0.873594f
C27 X VNB 0.043855f
C28 VPWR VNB 0.733649f
C29 A1 VNB 0.228877f
C30 A2 VNB 0.171608f
C31 A3 VNB 0.238367f
C32 B1 VNB 0.199521f
C33 C1 VNB 0.205918f
C34 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311a_2 VPWR VGND VPB VNB X A1 A2 A3 B1 C1
X0 X.t3 a_91_21.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_91_21.t1 C1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2 a_360_47.t1 A3.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR.t3 B1.t0 a_91_21.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X4 a_360_297.t0 A1.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X5 VGND.t2 A2.t0 a_360_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X6 a_360_47.t3 A1.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X7 VPWR.t0 a_91_21.t5 X.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t1 a_91_21.t6 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X.t0 a_91_21.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X10 a_677_47.t0 B1.t1 a_360_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X11 a_460_297.t0 A2.t1 a_360_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X12 a_91_21.t0 C1.t1 a_677_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X13 a_91_21.t3 A3.t1 a_460_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
R0 a_91_21.n3 a_91_21.n1 395.877
R1 a_91_21.t1 a_91_21.n4 386.803
R2 a_91_21.n1 a_91_21.t5 212.081
R3 a_91_21.n0 a_91_21.t4 212.081
R4 a_91_21.n3 a_91_21.n2 189.28
R5 a_91_21.n4 a_91_21.t0 185.898
R6 a_91_21.n1 a_91_21.t6 139.78
R7 a_91_21.n0 a_91_21.t7 139.78
R8 a_91_21.n1 a_91_21.n0 61.346
R9 a_91_21.n4 a_91_21.n3 45.389
R10 a_91_21.n2 a_91_21.t3 27.5805
R11 a_91_21.n2 a_91_21.t2 26.5955
R12 VPWR.n2 VPWR.n1 324.288
R13 VPWR.n4 VPWR.n3 306.897
R14 VPWR.n6 VPWR.t1 257.911
R15 VPWR.n3 VPWR.t4 69.9355
R16 VPWR.n3 VPWR.t0 53.1905
R17 VPWR.n1 VPWR.t2 29.5505
R18 VPWR.n1 VPWR.t3 29.5505
R19 VPWR.n5 VPWR.n4 28.9887
R20 VPWR.n6 VPWR.n5 23.3417
R21 VPWR.n5 VPWR.n0 9.3005
R22 VPWR.n7 VPWR.n6 9.3005
R23 VPWR.n4 VPWR.n2 6.11355
R24 VPWR.n2 VPWR.n0 0.173233
R25 VPWR.n7 VPWR.n0 0.120292
R26 VPWR VPWR.n7 0.0213333
R27 X.n1 X 592.753
R28 X.n1 X.n0 585
R29 X.n2 X.n1 585
R30 X.n5 X.n4 185
R31 X.n1 X.t2 26.5955
R32 X.n1 X.t3 26.5955
R33 X.n4 X.t1 24.9236
R34 X.n4 X.t0 24.9236
R35 X.n3 X 19.6928
R36 X.n3 X 9.37515
R37 X X.n5 8.61141
R38 X.n0 X 7.75261
R39 X X.n2 7.75261
R40 X.n5 X 7.21505
R41 X.n0 X 4.50754
R42 X.n2 X 4.50754
R43 X X.n3 2.88501
R44 VPB.t0 VPB.t6 458.724
R45 VPB.t3 VPB.t5 337.384
R46 VPB.t6 VPB.t3 295.95
R47 VPB.t4 VPB.t2 266.356
R48 VPB.t5 VPB.t4 251.559
R49 VPB.t1 VPB.t0 248.599
R50 VPB VPB.t1 224.923
R51 C1.n0 C1.t0 230.155
R52 C1.n0 C1.t1 157.856
R53 C1 C1.n0 154.91
R54 A3.n0 A3.t1 234.173
R55 A3.n0 A3.t0 161.873
R56 A3.n1 A3.n0 152
R57 A3 A3.n1 13.8194
R58 A3.n1 A3 2.42809
R59 VGND.n4 VGND.n3 190.963
R60 VGND.n8 VGND.t0 148.536
R61 VGND.n1 VGND.t4 59.0774
R62 VGND.n1 VGND.t1 56.3082
R63 VGND.n2 VGND.n1 46.2505
R64 VGND.n3 VGND.t3 38.7697
R65 VGND.n3 VGND.t2 38.7697
R66 VGND.n7 VGND.n6 25.1454
R67 VGND.n8 VGND.n7 23.3417
R68 VGND.n4 VGND.n2 11.0414
R69 VGND.n9 VGND.n8 9.3005
R70 VGND.n6 VGND.n5 9.3005
R71 VGND.n7 VGND.n0 9.3005
R72 VGND.n6 VGND.n2 2.53237
R73 VGND.n5 VGND.n4 0.50882
R74 VGND.n5 VGND.n0 0.120292
R75 VGND.n9 VGND.n0 0.120292
R76 VGND VGND.n9 0.0213333
R77 a_360_47.n1 a_360_47.n0 346.745
R78 a_360_47.n0 a_360_47.t1 34.1543
R79 a_360_47.n0 a_360_47.t2 33.2313
R80 a_360_47.t0 a_360_47.n1 33.2313
R81 a_360_47.n1 a_360_47.t3 31.3851
R82 VNB.t1 VNB.t5 2207.12
R83 VNB.t2 VNB.t3 1623.3
R84 VNB.t3 VNB.t4 1466.67
R85 VNB.t5 VNB.t2 1423.95
R86 VNB.t0 VNB.t1 1196.12
R87 VNB VNB.t0 1082.2
R88 VNB.t4 VNB.t6 1025.24
R89 B1.n0 B1.t0 238.155
R90 B1.n0 B1.t1 165.856
R91 B1 B1.n0 164.219
R92 A1.n0 A1.t0 241.536
R93 A1.n0 A1.t1 169.237
R94 A1 A1.n0 157.237
R95 a_360_297.t0 a_360_297.t1 68.9505
R96 A2.n0 A2.t1 241.536
R97 A2.n0 A2.t0 169.237
R98 A2.n1 A2.n0 152
R99 A2 A2.n1 12.0894
R100 A2.n1 A2 2.13383
R101 a_677_47.t0 a_677_47.t1 38.7697
R102 a_460_297.t0 a_460_297.t1 82.7405
C0 B1 VGND 0.016752f
C1 B1 VPB 0.027915f
C2 VGND A1 0.045341f
C3 C1 VPWR 0.02058f
C4 B1 X 6.93e-20
C5 VPB A1 0.031051f
C6 X A1 4.11e-19
C7 VPWR A2 0.013102f
C8 A2 A3 0.132989f
C9 VGND VPB 0.007138f
C10 B1 VPWR 0.016256f
C11 X VGND 0.177078f
C12 VPWR A1 0.008419f
C13 B1 A3 0.084907f
C14 X VPB 0.005974f
C15 B1 C1 0.058895f
C16 VPWR VGND 0.08862f
C17 VPWR VPB 0.090724f
C18 VGND A3 0.01939f
C19 VPWR X 0.218869f
C20 VPB A3 0.03464f
C21 A1 A2 0.078211f
C22 X A3 1.07e-19
C23 C1 VGND 0.008826f
C24 C1 VPB 0.038043f
C25 VGND A2 0.01833f
C26 VPB A2 0.031534f
C27 X A2 2e-19
C28 VPWR A3 0.013837f
C29 VGND VNB 0.502231f
C30 X VNB 0.031233f
C31 VPWR VNB 0.433132f
C32 C1 VNB 0.144887f
C33 B1 VNB 0.092815f
C34 A3 VNB 0.09991f
C35 A2 VNB 0.091862f
C36 A1 VNB 0.09397f
C37 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311a_1 X A1 A2 A3 B1 C1 VPB VNB VGND VPWR
X0 a_585_47.t0 B1.t0 a_266_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 VGND.t2 A2.t0 a_266_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR.t3 a_81_21.t4 X.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21.t2 C1.t0 a_585_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 VGND.t1 a_81_21.t5 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297.t1 A1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X6 a_368_297.t1 A2.t1 a_266_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47.t2 A3.t0 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X8 a_266_47.t3 A1.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X9 a_81_21.t0 A3.t1 a_368_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21.t3 C1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR.t0 B1.t1 a_81_21.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
R0 B1.n0 B1.t1 238.155
R1 B1.n0 B1.t0 165.856
R2 B1 B1.n0 164.219
R3 a_266_47.n1 a_266_47.n0 346.471
R4 a_266_47.n1 a_266_47.t2 34.1543
R5 a_266_47.n0 a_266_47.t1 33.2313
R6 a_266_47.n0 a_266_47.t3 33.2313
R7 a_266_47.t0 a_266_47.n1 33.2313
R8 a_585_47.t0 a_585_47.t1 38.7697
R9 VNB.t3 VNB.t5 2207.12
R10 VNB.t1 VNB.t2 1623.3
R11 VNB.t2 VNB.t0 1466.67
R12 VNB.t5 VNB.t1 1452.43
R13 VNB.t0 VNB.t4 1025.24
R14 VNB VNB.t3 968.285
R15 A2.n0 A2.t1 241.536
R16 A2.n0 A2.t0 169.237
R17 A2.n1 A2.n0 152
R18 A2 A2.n1 11.9012
R19 A2.n1 A2 2.07109
R20 VGND.n2 VGND.n1 191.246
R21 VGND.n0 VGND.t3 59.0774
R22 VGND.n0 VGND.t1 56.3082
R23 VGND.n2 VGND.n0 51.313
R24 VGND.n1 VGND.t0 38.7697
R25 VGND.n1 VGND.t2 38.7697
R26 VGND VGND.n2 0.357829
R27 a_81_21.n0 a_81_21.t3 386.803
R28 a_81_21.n2 a_81_21.n1 365.957
R29 a_81_21.n1 a_81_21.t4 231.017
R30 a_81_21.n3 a_81_21.n2 189.28
R31 a_81_21.n0 a_81_21.t2 185.898
R32 a_81_21.n1 a_81_21.t5 158.716
R33 a_81_21.n2 a_81_21.n0 45.389
R34 a_81_21.t0 a_81_21.n3 27.5805
R35 a_81_21.n3 a_81_21.t1 26.5955
R36 X.n1 X 592.864
R37 X.n1 X.n0 585
R38 X.n2 X.n1 585
R39 X.n3 X.t1 209.923
R40 X.n1 X.t0 26.5955
R41 X X.n3 8.77087
R42 X.n0 X 7.86336
R43 X X.n2 7.86336
R44 X.n3 X 7.34865
R45 X.n0 X 4.57193
R46 X.n2 X 4.57193
R47 VPWR.n2 VPWR.n0 324.312
R48 VPWR.n2 VPWR.n1 311.776
R49 VPWR.n1 VPWR.t2 69.9355
R50 VPWR.n1 VPWR.t3 53.1905
R51 VPWR.n0 VPWR.t1 29.5505
R52 VPWR.n0 VPWR.t0 29.5505
R53 VPWR VPWR.n2 0.172393
R54 VPB.t5 VPB.t4 458.724
R55 VPB.t3 VPB.t0 337.384
R56 VPB.t4 VPB.t3 301.87
R57 VPB.t1 VPB.t2 266.356
R58 VPB.t0 VPB.t1 251.559
R59 VPB VPB.t5 201.246
R60 C1.n0 C1.t1 230.155
R61 C1.n0 C1.t0 157.856
R62 C1 C1.n0 154.91
R63 A1.n0 A1.t0 241.536
R64 A1.n0 A1.t1 169.237
R65 A1 A1.n0 157.237
R66 a_266_297.t0 a_266_297.t1 70.9205
R67 a_368_297.t0 a_368_297.t1 82.7405
R68 A3.n0 A3.t1 234.173
R69 A3.n0 A3.t0 161.873
R70 A3.n1 A3.n0 152
R71 A3 A3.n1 13.8194
R72 A3.n1 A3 2.42809
C0 VPWR VPB 0.074178f
C1 VPB B1 0.027915f
C2 A2 X 1.97e-19
C3 VPWR B1 0.016256f
C4 VGND A3 0.01939f
C5 A1 A2 0.076636f
C6 VPB A3 0.03464f
C7 VGND A2 0.018378f
C8 A1 X 4.11e-19
C9 VPWR A3 0.013837f
C10 A3 B1 0.084907f
C11 VGND X 0.091215f
C12 VPB A2 0.031747f
C13 VPWR A2 0.013141f
C14 VGND A1 0.045005f
C15 VPB X 0.011438f
C16 VPWR X 0.105139f
C17 VGND C1 0.008826f
C18 B1 X 6.87e-20
C19 VPB A1 0.031201f
C20 VGND VPB 0.006542f
C21 VPWR A1 0.008378f
C22 VPB C1 0.038043f
C23 A2 A3 0.132989f
C24 VPWR VGND 0.07715f
C25 VGND B1 0.016752f
C26 VPWR C1 0.02058f
C27 B1 C1 0.058895f
C28 A3 X 1.06e-19
C29 VGND VNB 0.429376f
C30 VPWR VNB 0.361844f
C31 X VNB 0.093921f
C32 C1 VNB 0.144887f
C33 B1 VNB 0.092815f
C34 A3 VNB 0.09991f
C35 A2 VNB 0.092297f
C36 A1 VNB 0.09427f
C37 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_1 VPB VNB VGND VPWR Y A1 A2 C1 D1 B1
X0 VPWR.t2 C1.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X1 a_235_47.t1 C1.t1 a_163_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 a_343_47.t2 B1.t0 a_235_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.131625 pd=1.055 as=0.12675 ps=1.04 w=0.65 l=0.15
X3 Y.t0 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2025 pd=1.405 as=0.195 ps=1.39 w=1 l=0.15
X4 a_454_297.t1 A2.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.2025 ps=1.405 w=1 l=0.15
X5 Y.t2 D1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 VPWR.t3 A1.t0 a_454_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X7 a_163_47.t1 D1.t1 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X8 VGND.t1 A2.t1 a_343_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.131625 ps=1.055 w=0.65 l=0.15
X9 a_343_47.t1 A1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
R0 C1.n0 C1.t0 241.439
R1 C1 C1.n0 180.51
R2 C1.n0 C1.t1 169.138
R3 Y.n2 Y.n0 342.279
R4 Y.n2 Y.n1 295.932
R5 Y.n3 Y.t4 129.445
R6 Y.n3 Y.n2 93.5596
R7 Y.n0 Y.t0 42.3555
R8 Y.n0 Y.t1 37.4305
R9 Y.n1 Y.t3 27.5805
R10 Y.n1 Y.t2 27.5805
R11 Y Y.n3 3.23792
R12 VPWR.n7 VPWR.t1 863.645
R13 VPWR.n2 VPWR.n1 599.74
R14 VPWR.n3 VPWR.t3 346.313
R15 VPWR.n1 VPWR.t2 39.4005
R16 VPWR.n1 VPWR.t0 37.4305
R17 VPWR.n6 VPWR.n5 34.6358
R18 VPWR.n8 VPWR.n7 13.8181
R19 VPWR.n3 VPWR.n2 12.7961
R20 VPWR.n5 VPWR.n4 9.3005
R21 VPWR.n6 VPWR.n0 9.3005
R22 VPWR.n7 VPWR.n6 5.27109
R23 VPWR.n5 VPWR.n2 4.51815
R24 VPWR.n4 VPWR.n3 0.222113
R25 VPWR.n4 VPWR.n0 0.120292
R26 VPWR.n8 VPWR.n0 0.120292
R27 VPWR VPWR.n8 0.0226354
R28 VPB.t0 VPB.t1 328.505
R29 VPB.t1 VPB.t4 319.627
R30 VPB.t3 VPB.t0 319.627
R31 VPB VPB.t2 310.748
R32 VPB.t2 VPB.t3 254.518
R33 a_163_47.t0 a_163_47.t1 38.7697
R34 a_235_47.t0 a_235_47.t1 72.0005
R35 VNB VNB.t4 1694.5
R36 VNB.t2 VNB.t0 1580.58
R37 VNB.t0 VNB.t1 1537.86
R38 VNB.t3 VNB.t2 1537.86
R39 VNB.t4 VNB.t3 1025.24
R40 B1.n0 B1.t1 241.439
R41 B1.n0 B1.t0 169.138
R42 B1 B1.n0 156.232
R43 a_343_47.n0 a_343_47.t1 274.014
R44 a_343_47.n0 a_343_47.t2 39.6928
R45 a_343_47.t0 a_343_47.n0 35.0774
R46 A2.n0 A2.t0 241.439
R47 A2.n0 A2.t1 169.138
R48 A2 A2.n0 153.118
R49 a_454_297.t0 a_454_297.t1 76.8305
R50 D1.n0 D1.t0 241.439
R51 D1.n0 D1.t1 169.138
R52 D1 D1.n0 154.133
R53 A1.n0 A1.t0 233.868
R54 A1.n0 A1.t1 161.567
R55 A1 A1.n0 154.133
R56 VGND VGND.n0 205.594
R57 VGND.n0 VGND.t0 38.7697
R58 VGND.n0 VGND.t1 33.2313
C0 VPB Y 0.019469f
C1 D1 C1 0.104675f
C2 A1 VPB 0.043335f
C3 A2 D1 1.58e-19
C4 B1 C1 0.102954f
C5 B1 A2 0.097537f
C6 Y VGND 0.090585f
C7 VPWR Y 0.257894f
C8 A1 VGND 0.01688f
C9 A1 VPWR 0.055699f
C10 VPB C1 0.031796f
C11 A2 VPB 0.037148f
C12 C1 VGND 0.049665f
C13 A2 VGND 0.020705f
C14 A1 Y 3.09e-19
C15 VPWR C1 0.017521f
C16 A2 VPWR 0.105795f
C17 VPB D1 0.035528f
C18 B1 VPB 0.03329f
C19 D1 VGND 0.013293f
C20 C1 Y 0.082501f
C21 A2 Y 0.070186f
C22 B1 VGND 0.016455f
C23 A1 C1 2.05e-19
C24 VPWR D1 0.016012f
C25 A2 A1 0.108638f
C26 B1 VPWR 0.014301f
C27 D1 Y 0.116743f
C28 VPB VGND 0.006238f
C29 B1 Y 0.04151f
C30 VPWR VPB 0.076627f
C31 A2 C1 7.26e-19
C32 VPWR VGND 0.064777f
C33 VGND VNB 0.390697f
C34 Y VNB 0.094123f
C35 VPWR VNB 0.362327f
C36 A1 VNB 0.157525f
C37 A2 VNB 0.105404f
C38 B1 VNB 0.097563f
C39 C1 VNB 0.101559f
C40 D1 VNB 0.120188f
C41 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_2 VNB VPB VPWR VGND D1 Y C1 B1 A1 A2
X0 Y.t3 C1.t0 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_298_47.t1 C1.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND.t3 A1.t0 a_497_47.t5 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_664_297.t3 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND.t1 A2.t0 a_497_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VPWR.t3 C1.t2 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_298_47.t2 B1.t0 a_497_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.1755 ps=1.84 w=0.65 l=0.15
X7 a_497_47.t0 A2.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 Y.t7 D1.t0 a_27_47.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.22425 ps=1.99 w=0.65 l=0.15
X9 a_497_47.t2 B1.t1 a_298_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y.t1 B1.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 Y.t4 A2.t2 a_664_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.295 ps=2.59 w=1 l=0.15
X12 a_27_47.t1 C1.t3 a_298_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.091 ps=0.93 w=0.65 l=0.15
X13 VPWR.t6 D1.t1 Y.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 VPWR.t5 B1.t3 Y.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 a_27_47.t3 D1.t2 Y.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_497_47.t4 A1.t2 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.091 ps=0.93 w=0.65 l=0.15
X17 Y.t9 D1.t3 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 VPWR.t2 A1.t3 a_664_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_664_297.t0 A2.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 C1.n0 C1.t2 221.72
R1 C1.n1 C1.t0 221.72
R2 C1 C1.n2 157.12
R3 C1.n0 C1.t3 149.421
R4 C1.n1 C1.t1 149.421
R5 C1.n2 C1.n0 39.2746
R6 C1.n2 C1.n1 37.4894
R7 VPWR.n15 VPWR.t7 347.295
R8 VPWR.n7 VPWR.t5 338.082
R9 VPWR.n6 VPWR.n5 320.688
R10 VPWR.n13 VPWR.n2 310.502
R11 VPWR.n4 VPWR.n3 310.502
R12 VPWR.n2 VPWR.t4 27.5805
R13 VPWR.n2 VPWR.t6 27.5805
R14 VPWR.n3 VPWR.t0 27.5805
R15 VPWR.n3 VPWR.t3 27.5805
R16 VPWR.n5 VPWR.t1 27.5805
R17 VPWR.n5 VPWR.t2 27.5805
R18 VPWR.n14 VPWR.n13 25.977
R19 VPWR.n8 VPWR.n4 22.9652
R20 VPWR.n12 VPWR.n4 21.4593
R21 VPWR.n15 VPWR.n14 19.9534
R22 VPWR.n13 VPWR.n12 18.4476
R23 VPWR.n8 VPWR.n7 16.9417
R24 VPWR.n9 VPWR.n8 9.3005
R25 VPWR.n10 VPWR.n4 9.3005
R26 VPWR.n12 VPWR.n11 9.3005
R27 VPWR.n13 VPWR.n1 9.3005
R28 VPWR.n14 VPWR.n0 9.3005
R29 VPWR.n16 VPWR.n15 9.3005
R30 VPWR.n7 VPWR.n6 7.31606
R31 VPWR.n9 VPWR.n6 0.163403
R32 VPWR.n10 VPWR.n9 0.120292
R33 VPWR.n11 VPWR.n10 0.120292
R34 VPWR.n11 VPWR.n1 0.120292
R35 VPWR.n1 VPWR.n0 0.120292
R36 VPWR.n16 VPWR.n0 0.120292
R37 VPWR VPWR.n16 0.0226354
R38 Y.n4 Y.n2 699.923
R39 Y.n0 Y 593.615
R40 Y.n1 Y.n0 585
R41 Y.n4 Y.n3 319.216
R42 Y.n6 Y.n5 317.82
R43 Y Y.n7 188.201
R44 Y.n6 Y.n4 50.4476
R45 Y.n8 Y.n6 50.4476
R46 Y.n0 Y.t6 27.5805
R47 Y.n0 Y.t9 27.5805
R48 Y.n2 Y.t0 27.5805
R49 Y.n2 Y.t4 27.5805
R50 Y.n3 Y.t5 27.5805
R51 Y.n3 Y.t1 27.5805
R52 Y.n5 Y.t2 27.5805
R53 Y.n5 Y.t3 27.5805
R54 Y.n7 Y.t8 25.8467
R55 Y.n7 Y.t7 25.8467
R56 Y.n1 Y 14.2774
R57 Y Y.n8 10.0928
R58 Y.n8 Y 6.64665
R59 Y Y.n1 2.46204
R60 VPB.t7 VPB.t6 583.023
R61 VPB.t3 VPB.t2 254.518
R62 VPB.t0 VPB.t3 254.518
R63 VPB.t6 VPB.t0 254.518
R64 VPB.t1 VPB.t7 254.518
R65 VPB.t4 VPB.t1 254.518
R66 VPB.t5 VPB.t4 254.518
R67 VPB.t8 VPB.t5 254.518
R68 VPB.t9 VPB.t8 254.518
R69 VPB VPB.t9 242.679
R70 a_27_47.n0 a_27_47.t1 284.692
R71 a_27_47.n0 a_27_47.t2 188.227
R72 a_27_47.n1 a_27_47.n0 185
R73 a_27_47.n1 a_27_47.t3 26.7697
R74 a_27_47.t0 a_27_47.n1 24.9236
R75 a_298_47.n1 a_298_47.n0 492.92
R76 a_298_47.t1 a_298_47.n1 26.7697
R77 a_298_47.n0 a_298_47.t3 25.8467
R78 a_298_47.n0 a_298_47.t2 25.8467
R79 a_298_47.n1 a_298_47.t0 24.9236
R80 VNB.t3 VNB.t5 2805.18
R81 VNB.t0 VNB.t1 1224.6
R82 VNB.t2 VNB.t0 1224.6
R83 VNB.t7 VNB.t2 1224.6
R84 VNB.t6 VNB.t7 1224.6
R85 VNB.t5 VNB.t6 1224.6
R86 VNB.t4 VNB.t3 1224.6
R87 VNB.t9 VNB.t4 1224.6
R88 VNB.t8 VNB.t9 1224.6
R89 VNB VNB.t8 1167.64
R90 A1.n0 A1.t1 221.72
R91 A1.n1 A1.t3 221.72
R92 A1.n3 A1.n2 152
R93 A1.n0 A1.t2 149.421
R94 A1.n1 A1.t0 149.421
R95 A1.n2 A1.n1 44.6301
R96 A1.n2 A1.n0 32.1338
R97 A1.n3 A1 20.7365
R98 A1 A1.n3 2.8165
R99 a_497_47.n1 a_497_47.t1 320.356
R100 a_497_47.n2 a_497_47.t4 279.764
R101 a_497_47.n3 a_497_47.n2 190.054
R102 a_497_47.n1 a_497_47.n0 185
R103 a_497_47.n2 a_497_47.n1 55.452
R104 a_497_47.n0 a_497_47.t3 26.7697
R105 a_497_47.n3 a_497_47.t5 25.8467
R106 a_497_47.t0 a_497_47.n3 25.8467
R107 a_497_47.n0 a_497_47.t2 24.9236
R108 VGND.n2 VGND.n0 205.404
R109 VGND.n2 VGND.n1 205.194
R110 VGND.n0 VGND.t2 25.8467
R111 VGND.n0 VGND.t3 25.8467
R112 VGND.n1 VGND.t0 25.8467
R113 VGND.n1 VGND.t1 25.8467
R114 VGND VGND.n2 1.37576
R115 a_664_297.n0 a_664_297.t3 444.772
R116 a_664_297.n0 a_664_297.t1 386.841
R117 a_664_297.n1 a_664_297.n0 187.786
R118 a_664_297.t2 a_664_297.n1 27.5805
R119 a_664_297.n1 a_664_297.t0 27.5805
R120 A2.n0 A2.t3 221.72
R121 A2.n1 A2.t2 221.72
R122 A2 A2.n2 156.608
R123 A2.n0 A2.t1 149.421
R124 A2.n1 A2.t0 149.421
R125 A2.n2 A2.n1 40.1672
R126 A2.n2 A2.n0 36.5968
R127 B1.n3 B1.t2 237.787
R128 B1.n2 B1.t3 221.72
R129 B1.n0 B1.t1 192.264
R130 B1 B1.n0 157.888
R131 B1 B1.n3 156.096
R132 B1.n1 B1.t0 149.421
R133 B1.n3 B1.n2 60.6968
R134 B1.n1 B1.n0 33.919
R135 B1.n2 B1.n1 22.3153
R136 D1.n0 D1.t1 212.081
R137 D1.n1 D1.t3 212.081
R138 D1 D1.n1 200.345
R139 D1.n0 D1.t2 139.78
R140 D1.n1 D1.t0 139.78
R141 D1.n1 D1.n0 62.8066
C0 A1 VPB 0.059588f
C1 A1 Y 2.66e-19
C2 VPB C1 0.053867f
C3 VPWR B1 0.045786f
C4 Y C1 0.119921f
C5 A1 VGND 0.033971f
C6 VGND C1 0.021281f
C7 A2 VPB 0.060398f
C8 A1 VPWR 0.041522f
C9 A2 Y 0.073368f
C10 VPB D1 0.075862f
C11 VPWR C1 0.041648f
C12 Y D1 0.091394f
C13 C1 B1 0.0519f
C14 A2 VGND 0.034637f
C15 VGND D1 0.021535f
C16 A2 VPWR 0.020172f
C17 Y VPB 0.023049f
C18 VPWR D1 0.067513f
C19 A2 B1 0.060621f
C20 VGND VPB 0.011201f
C21 Y VGND 0.017161f
C22 A2 A1 0.073225f
C23 VPWR VPB 0.129744f
C24 VPWR Y 0.570858f
C25 D1 C1 0.054719f
C26 VPB B1 0.084837f
C27 Y B1 0.117265f
C28 VPWR VGND 0.108077f
C29 VGND B1 0.025101f
C30 VGND VNB 0.615058f
C31 Y VNB 0.024315f
C32 VPWR VNB 0.541254f
C33 A1 VNB 0.211674f
C34 A2 VNB 0.17669f
C35 B1 VNB 0.23225f
C36 C1 VNB 0.179265f
C37 D1 VNB 0.243601f
C38 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_4 VNB VPB VGND VPWR Y D1 C1 B1 A2 A1
X0 a_27_47.t4 C1.t0 a_445_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_803_47.t5 A2.t0 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_47.t3 C1.t1 a_445_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t2 A2.t1 a_803_47.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t9 C1.t2 Y.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t1 A2.t2 a_803_47.t3 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.095875 ps=0.945 w=0.65 l=0.15
X7 Y.t11 D1.t0 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1475 ps=1.295 w=1 l=0.15
X10 a_445_47.t7 B1.t0 a_803_47.t7 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t11 D1.t1 Y.t12 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47.t6 B1.t1 a_803_47.t6 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 Y.t13 D1.t2 VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t12 A1.t0 a_1163_297# VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47.t7 D1.t3 Y.t14 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47.t5 D1.t4 Y.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t14 B1.t2 Y.t15 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t0 B1.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.135 ps=1.27 w=1 l=0.15
X19 a_1163_297# A1.t1 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_803_47.t0 B1.t4 a_445_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t1 B1.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 Y.t7 C1.t3 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2375 pd=1.475 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t5 A1.t2 a_1163_297# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_803_47.t1 B1.t6 a_445_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 Y.t10 D1.t5 a_27_47.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t2 B1.t7 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2375 ps=1.475 w=1 l=0.15
X27 a_445_47.t5 C1.t4 a_27_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VPWR.t7 C1.t5 Y.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_1163_297# A1.t3 VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X30 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25335 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X31 a_445_47.t4 C1.t6 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 Y.t5 C1.t7 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_803_47.t2 A2.t3 VGND.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 VPWR.t3 D1.t6 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 Y.t4 D1.t7 a_27_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C1.n1 C1.t3 221.72
R1 C1.n2 C1.t5 221.72
R2 C1.n8 C1.t7 221.72
R3 C1.n9 C1.t2 221.72
R4 C1.n4 C1.n3 152
R5 C1.n5 C1.n0 152
R6 C1.n7 C1.n6 152
R7 C1.n11 C1.n10 152
R8 C1.n1 C1.t1 149.421
R9 C1.n2 C1.t6 149.421
R10 C1.n8 C1.t0 149.421
R11 C1.n9 C1.t4 149.421
R12 C1.n7 C1.n0 60.6968
R13 C1.n10 C1.n8 58.9116
R14 C1.n3 C1.n2 48.2005
R15 C1.n3 C1.n1 26.7783
R16 C1.n5 C1.n4 16.119
R17 C1.n10 C1.n9 16.0672
R18 C1.n6 C1 15.6449
R19 C1.n2 C1.n0 12.4968
R20 C1 C1.n11 11.8524
R21 C1.n11 C1 9.95606
R22 C1.n6 C1 6.16346
R23 C1.n4 C1 5.21532
R24 C1.n8 C1.n7 1.78569
R25 C1 C1.n5 0.474574
R26 a_445_47.n5 a_445_47.n4 241.589
R27 a_445_47.n2 a_445_47.n0 241.589
R28 a_445_47.n4 a_445_47.n3 185
R29 a_445_47.n2 a_445_47.n1 185
R30 a_445_47.n4 a_445_47.n2 91.6216
R31 a_445_47.n0 a_445_47.t3 24.9236
R32 a_445_47.n0 a_445_47.t5 24.9236
R33 a_445_47.n1 a_445_47.t2 24.9236
R34 a_445_47.n1 a_445_47.t4 24.9236
R35 a_445_47.n3 a_445_47.t1 24.9236
R36 a_445_47.n3 a_445_47.t6 24.9236
R37 a_445_47.t0 a_445_47.n5 24.9236
R38 a_445_47.n5 a_445_47.t7 24.9236
R39 a_27_47.n1 a_27_47.t0 320.051
R40 a_27_47.n4 a_27_47.t3 300.815
R41 a_27_47.n1 a_27_47.n0 185
R42 a_27_47.n3 a_27_47.n2 185
R43 a_27_47.n5 a_27_47.n4 185
R44 a_27_47.n3 a_27_47.n1 62.99
R45 a_27_47.n4 a_27_47.n3 55.3417
R46 a_27_47.n2 a_27_47.t2 24.9236
R47 a_27_47.n2 a_27_47.t5 24.9236
R48 a_27_47.n0 a_27_47.t6 24.9236
R49 a_27_47.n0 a_27_47.t7 24.9236
R50 a_27_47.n5 a_27_47.t1 24.9236
R51 a_27_47.t4 a_27_47.n5 24.9236
R52 VNB.t5 VNB.t13 2677.02
R53 VNB.t0 VNB.t15 1267.31
R54 VNB.t7 VNB.t8 1253.07
R55 VNB.t8 VNB.t11 1196.12
R56 VNB.t15 VNB.t7 1196.12
R57 VNB.t14 VNB.t0 1196.12
R58 VNB.t1 VNB.t14 1196.12
R59 VNB.t13 VNB.t1 1196.12
R60 VNB.t3 VNB.t5 1196.12
R61 VNB.t6 VNB.t3 1196.12
R62 VNB.t4 VNB.t6 1196.12
R63 VNB.t9 VNB.t4 1196.12
R64 VNB.t10 VNB.t9 1196.12
R65 VNB.t12 VNB.t10 1196.12
R66 VNB.t2 VNB.t12 1196.12
R67 VNB VNB.t2 911.327
R68 A2.n12 A2.n10 278.007
R69 A2.n3 A2.n2 221.72
R70 A2.n8 A2.n0 221.72
R71 A2.n3 A2.t3 209.225
R72 A2.n12 A2.n11 198.944
R73 A2.n13 A2.t2 174.939
R74 A2.n5 A2.n4 152
R75 A2.n7 A2.n6 152
R76 A2.n15 A2.n14 152
R77 A2.n9 A2.t0 149.421
R78 A2.n1 A2.t1 149.421
R79 A2.n7 A2.n1 46.4153
R80 A2.n13 A2.n12 33.0789
R81 A2.n14 A2.n9 28.5635
R82 A2.n9 A2.n8 18.7449
R83 A2.n6 A2.n5 16.119
R84 A2.n4 A2.n1 14.282
R85 A2.n14 A2.n13 14.282
R86 A2.n8 A2.n7 13.3894
R87 A2.n15 A2 12.8005
R88 A2 A2.n15 9.00791
R89 A2.n6 A2 3.31902
R90 A2.n5 A2 2.37087
R91 A2.n4 A2.n3 0.893093
R92 VGND.n2 VGND.n1 204.965
R93 VGND.n2 VGND.n0 204.618
R94 VGND.n0 VGND.t0 24.9236
R95 VGND.n0 VGND.t2 24.9236
R96 VGND.n1 VGND.t3 24.9236
R97 VGND.n1 VGND.t1 24.9236
R98 VGND VGND.n2 1.97903
R99 a_803_47.n1 a_803_47.t6 311.086
R100 a_803_47.n4 a_803_47.t2 303.533
R101 a_803_47.n3 a_803_47.n2 185
R102 a_803_47.n1 a_803_47.n0 185
R103 a_803_47.n5 a_803_47.n4 185
R104 a_803_47.n3 a_803_47.n1 44.2885
R105 a_803_47.n4 a_803_47.n3 43.0085
R106 a_803_47.n2 a_803_47.t0 29.539
R107 a_803_47.n5 a_803_47.t4 28.6159
R108 a_803_47.n0 a_803_47.t7 24.9236
R109 a_803_47.n0 a_803_47.t1 24.9236
R110 a_803_47.n2 a_803_47.t3 24.9236
R111 a_803_47.t5 a_803_47.n5 24.9236
R112 Y Y.n0 593.145
R113 Y.n15 Y.n0 585
R114 Y.n2 Y.t0 397.906
R115 Y.n10 Y.n9 324.022
R116 Y.n2 Y.n1 322.37
R117 Y.n4 Y.n3 322.37
R118 Y.n6 Y.n5 322.37
R119 Y.n8 Y.n7 322.37
R120 Y.n13 Y.n11 248.248
R121 Y.n13 Y.n12 185
R122 Y.n3 Y.t2 66.9805
R123 Y.n4 Y.n2 64.377
R124 Y.n6 Y.n4 48.9417
R125 Y.n8 Y.n6 48.9417
R126 Y.n10 Y.n8 48.9417
R127 Y.n14 Y.n10 48.1887
R128 Y.n0 Y.t3 26.5955
R129 Y.n1 Y.t15 26.5955
R130 Y.n1 Y.t1 26.5955
R131 Y.n3 Y.t7 26.5955
R132 Y.n5 Y.t6 26.5955
R133 Y.n5 Y.t5 26.5955
R134 Y.n7 Y.t8 26.5955
R135 Y.n7 Y.t11 26.5955
R136 Y.n9 Y.t12 26.5955
R137 Y.n9 Y.t13 26.5955
R138 Y.n12 Y.t14 24.9236
R139 Y.n12 Y.t4 24.9236
R140 Y.n11 Y.t9 24.9236
R141 Y.n11 Y.t10 24.9236
R142 Y Y.n13 24.51
R143 Y Y.n14 8.40677
R144 Y.n15 Y 8.14595
R145 Y Y.n15 7.6805
R146 Y.n14 Y 6.84188
R147 VPB.t0 VPB.t15 1559.66
R148 VPB.t8 VPB.t2 369.938
R149 VPB.t4 VPB.t12 248.599
R150 VPB.t5 VPB.t4 248.599
R151 VPB.t15 VPB.t5 248.599
R152 VPB.t14 VPB.t0 248.599
R153 VPB.t1 VPB.t14 248.599
R154 VPB.t2 VPB.t1 248.599
R155 VPB.t7 VPB.t8 248.599
R156 VPB.t6 VPB.t7 248.599
R157 VPB.t9 VPB.t6 248.599
R158 VPB.t10 VPB.t9 248.599
R159 VPB.t11 VPB.t10 248.599
R160 VPB.t13 VPB.t11 248.599
R161 VPB.t3 VPB.t13 248.599
R162 VPB VPB.t3 189.409
R163 VPWR.n14 VPWR.t15 788.865
R164 VPWR.n15 VPWR.t12 344.89
R165 VPWR.n42 VPWR.n3 312.438
R166 VPWR.n29 VPWR.n11 312.096
R167 VPWR.n5 VPWR.n4 310.834
R168 VPWR.n36 VPWR.n7 310.834
R169 VPWR.n17 VPWR.n16 310.834
R170 VPWR.n44 VPWR.n1 310.543
R171 VPWR.n31 VPWR.n10 309.99
R172 VPWR.n38 VPWR.n37 34.6358
R173 VPWR.n35 VPWR.n8 34.6358
R174 VPWR.n23 VPWR.n22 34.6358
R175 VPWR.n24 VPWR.n23 34.6358
R176 VPWR.n24 VPWR.n12 34.6358
R177 VPWR.n28 VPWR.n12 34.6358
R178 VPWR.n31 VPWR.n30 32.377
R179 VPWR.n22 VPWR.n14 32.0005
R180 VPWR.n42 VPWR.n41 29.7417
R181 VPWR.n18 VPWR.n17 27.1064
R182 VPWR.n1 VPWR.t13 26.5955
R183 VPWR.n1 VPWR.t3 26.5955
R184 VPWR.n3 VPWR.t10 26.5955
R185 VPWR.n3 VPWR.t11 26.5955
R186 VPWR.n4 VPWR.t6 26.5955
R187 VPWR.n4 VPWR.t9 26.5955
R188 VPWR.n7 VPWR.t8 26.5955
R189 VPWR.n7 VPWR.t7 26.5955
R190 VPWR.n10 VPWR.t1 26.5955
R191 VPWR.n10 VPWR.t2 26.5955
R192 VPWR.n11 VPWR.t0 26.5955
R193 VPWR.n11 VPWR.t14 26.5955
R194 VPWR.n16 VPWR.t4 26.5955
R195 VPWR.n16 VPWR.t5 26.5955
R196 VPWR.n44 VPWR.n43 22.9652
R197 VPWR.n43 VPWR.n42 18.0711
R198 VPWR.n31 VPWR.n8 12.424
R199 VPWR.n18 VPWR.n14 12.424
R200 VPWR.n41 VPWR.n5 10.1652
R201 VPWR.n19 VPWR.n18 9.3005
R202 VPWR.n20 VPWR.n14 9.3005
R203 VPWR.n22 VPWR.n21 9.3005
R204 VPWR.n23 VPWR.n13 9.3005
R205 VPWR.n25 VPWR.n24 9.3005
R206 VPWR.n26 VPWR.n12 9.3005
R207 VPWR.n28 VPWR.n27 9.3005
R208 VPWR.n30 VPWR.n9 9.3005
R209 VPWR.n32 VPWR.n31 9.3005
R210 VPWR.n33 VPWR.n8 9.3005
R211 VPWR.n35 VPWR.n34 9.3005
R212 VPWR.n37 VPWR.n6 9.3005
R213 VPWR.n39 VPWR.n38 9.3005
R214 VPWR.n41 VPWR.n40 9.3005
R215 VPWR.n42 VPWR.n2 9.3005
R216 VPWR.n43 VPWR.n0 9.3005
R217 VPWR.n30 VPWR.n29 7.52991
R218 VPWR.n45 VPWR.n44 7.18025
R219 VPWR.n36 VPWR.n35 7.15344
R220 VPWR.n17 VPWR.n15 6.26659
R221 VPWR.n29 VPWR.n28 5.27109
R222 VPWR.n37 VPWR.n36 4.14168
R223 VPWR.n38 VPWR.n5 1.12991
R224 VPWR.n19 VPWR.n15 0.71414
R225 VPWR.n45 VPWR.n0 0.147761
R226 VPWR.n20 VPWR.n19 0.120292
R227 VPWR.n21 VPWR.n20 0.120292
R228 VPWR.n21 VPWR.n13 0.120292
R229 VPWR.n25 VPWR.n13 0.120292
R230 VPWR.n26 VPWR.n25 0.120292
R231 VPWR.n27 VPWR.n26 0.120292
R232 VPWR.n27 VPWR.n9 0.120292
R233 VPWR.n32 VPWR.n9 0.120292
R234 VPWR.n33 VPWR.n32 0.120292
R235 VPWR.n34 VPWR.n33 0.120292
R236 VPWR.n34 VPWR.n6 0.120292
R237 VPWR.n39 VPWR.n6 0.120292
R238 VPWR.n40 VPWR.n39 0.120292
R239 VPWR.n40 VPWR.n2 0.120292
R240 VPWR.n2 VPWR.n0 0.120292
R241 VPWR VPWR.n45 0.114308
R242 D1.n1 D1.t0 192.8
R243 D1.n0 D1.t1 192.8
R244 D1.n5 D1.t2 192.8
R245 D1.n6 D1.t6 192.8
R246 D1 D1.n2 153.66
R247 D1.n4 D1.n3 152
R248 D1.n8 D1.n7 152
R249 D1.n1 D1.t4 149.421
R250 D1.n0 D1.t5 149.421
R251 D1.n5 D1.t3 149.421
R252 D1.n6 D1.t7 149.421
R253 D1.n2 D1.n0 34.1422
R254 D1.n7 D1.n6 32.1338
R255 D1.n5 D1.n4 30.7949
R256 D1.n4 D1.n0 25.4394
R257 D1.n7 D1.n5 24.1005
R258 D1.n2 D1.n1 22.0922
R259 D1.n3 D1 19.4375
R260 D1.n8 D1 17.0672
R261 D1 D1.n8 4.74124
R262 D1.n3 D1 2.37087
R263 B1.n10 B1.t7 260.281
R264 B1.n1 B1.t4 233.84
R265 B1.n1 B1.t3 222.718
R266 B1.n3 B1.t2 221.72
R267 B1.n8 B1.t5 221.72
R268 B1.n2 B1.t0 168.701
R269 B1.n5 B1.n4 152
R270 B1.n7 B1.n6 152
R271 B1.n11 B1.n10 152
R272 B1.n9 B1.t1 147.814
R273 B1.n0 B1.t6 147.814
R274 B1.n4 B1.n2 53.4587
R275 B1.n7 B1.n0 30.6732
R276 B1.n8 B1.n7 24.5387
R277 B1 B1.n11 20.3857
R278 B1.n3 B1.n0 18.4041
R279 B1.n9 B1.n8 18.4041
R280 B1.n10 B1.n9 16.6514
R281 B1.n6 B1 14.6968
R282 B1.n5 B1 12.8005
R283 B1.n4 B1.n3 10.5169
R284 B1 B1.n5 9.00791
R285 B1.n2 B1.n1 7.91443
R286 B1.n6 B1 7.11161
R287 B1.n11 B1 1.42272
R288 A1.n5 A1.t0 248.499
R289 A1.n3 A1.t1 221.72
R290 A1.n11 A1.t2 221.72
R291 A1.n15 A1.t3 221.72
R292 A1.n15 A1.n14 176.198
R293 A1.n7 A1.n6 152
R294 A1.n9 A1.n8 152
R295 A1.n12 A1.n0 152
R296 A1.n17 A1.n16 152
R297 A1.n13 A1.n1 149.421
R298 A1.n10 A1.n2 149.421
R299 A1.n5 A1.n4 149.421
R300 A1.n11 A1.n10 48.2005
R301 A1.n6 A1.n3 42.8449
R302 A1.n16 A1.n13 37.4894
R303 A1.n13 A1.n12 23.2079
R304 A1.n9 A1.n3 17.8524
R305 A1.n17 A1.n0 16.4231
R306 A1.n7 A1 16.1816
R307 A1.n8 A1 11.8345
R308 A1.n16 A1.n15 10.7116
R309 A1.n8 A1 10.3854
R310 A1.n10 A1.n9 8.92643
R311 A1 A1.n7 6.03824
R312 A1.n6 A1.n5 5.35606
R313 A1 A1.n0 4.58918
R314 A1.n12 A1.n11 3.57087
R315 A1 A1.n17 1.20805
C0 VPWR VPB 0.191367f
C1 a_1163_297# A1 0.156245f
C2 D1 VPWR 0.085953f
C3 C1 Y 0.201167f
C4 C1 VPB 0.120467f
C5 A2 VGND 0.068863f
C6 A1 VPWR 0.11276f
C7 Y VPB 0.032529f
C8 D1 C1 0.073873f
C9 a_1163_297# A2 0.046385f
C10 B1 A2 0.053855f
C11 D1 Y 0.311952f
C12 a_1163_297# VGND 0.008306f
C13 D1 VPB 0.117001f
C14 A2 VPWR 0.034752f
C15 B1 VGND 0.039194f
C16 A1 Y 0.001164f
C17 A1 VPB 0.134855f
C18 VPWR VGND 0.187416f
C19 a_1163_297# VPWR 0.517099f
C20 C1 VGND 0.032642f
C21 A2 Y 0.156195f
C22 B1 VPWR 0.074395f
C23 A2 VPB 0.136936f
C24 Y VGND 0.040514f
C25 VGND VPB 0.013113f
C26 C1 B1 0.04507f
C27 a_1163_297# Y 0.236313f
C28 a_1163_297# VPB 0.018264f
C29 D1 VGND 0.036444f
C30 B1 Y 0.205311f
C31 C1 VPWR 0.071563f
C32 A2 A1 0.048312f
C33 B1 VPB 0.134119f
C34 A1 VGND 0.071693f
C35 Y VPWR 1.0833f
C36 VGND VNB 1.02946f
C37 VPWR VNB 0.888625f
C38 Y VNB 0.090132f
C39 A1 VNB 0.414111f
C40 A2 VNB 0.382906f
C41 B1 VNB 0.402563f
C42 C1 VNB 0.365244f
C43 D1 VNB 0.381078f
C44 VPB VNB 1.9337f
C45 a_1163_297# VNB 0.004479f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_0 VNB VPB VGND VPWR B A X
X0 VGND.t1 A.t0 a_68_355.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_150_355.t1 B.t0 a_68_355.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_68_355.t1 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X.t0 a_68_355.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4 VPWR.t1 A.t1 a_150_355.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.09895 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 X.t1 a_68_355.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2176 pd=1.96 as=0.09895 ps=0.975 w=0.64 l=0.15
R0 A.n0 A.t1 241.536
R1 A A.n0 154.167
R2 A.n0 A.t0 132.282
R3 a_68_355.n1 a_68_355.t2 662.71
R4 a_68_355.n0 a_68_355.t4 271.527
R5 a_68_355.n2 a_68_355.n1 264.825
R6 a_68_355.n1 a_68_355.n0 263.435
R7 a_68_355.n0 a_68_355.t3 126.927
R8 a_68_355.t0 a_68_355.n2 38.5719
R9 a_68_355.n2 a_68_355.t1 38.5719
R10 VGND.n1 VGND.t2 265.688
R11 VGND.n1 VGND.n0 231.069
R12 VGND.n0 VGND.t1 55.7148
R13 VGND.n0 VGND.t0 40.0005
R14 VGND VGND.n1 0.437652
R15 VNB.t1 VNB.t0 1381.23
R16 VNB VNB.t2 1338.51
R17 VNB.t2 VNB.t1 1196.12
R18 B.n0 B.t0 227.987
R19 B B.n0 157.575
R20 B.n0 B.t1 118.734
R21 a_150_355.t0 a_150_355.t1 98.5005
R22 VPB VPB.t2 313.707
R23 VPB.t1 VPB.t0 287.072
R24 VPB.t2 VPB.t1 213.084
R25 X X.t1 673.548
R26 X X.t0 274.437
R27 VPWR VPWR.n0 614.836
R28 VPWR.n0 VPWR.t1 96.1553
R29 VPWR.n0 VPWR.t0 40.0161
C0 VPWR X 0.100569f
C1 VPWR VPB 0.071185f
C2 VGND A 0.033958f
C3 B A 0.083556f
C4 VGND B 0.039782f
C5 X A 0.001592f
C6 VPB A 0.049089f
C7 X VGND 0.071192f
C8 VPWR A 0.01077f
C9 X B 1.65e-19
C10 VGND VPB 0.010804f
C11 VPB B 0.070456f
C12 VPWR VGND 0.046086f
C13 VPWR B 0.010854f
C14 X VPB 0.023702f
C15 VGND VNB 0.360064f
C16 X VNB 0.091765f
C17 VPWR VNB 0.263522f
C18 A VNB 0.089905f
C19 B VNB 0.166389f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND.t0 A.t0 a_68_297.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297.t1 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X.t1 a_68_297.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR.t0 A.t1 a_150_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X.t0 a_68_297.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297.t1 B.t1 a_68_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A.n0 A.t0 206.19
R1 A A.n0 154.657
R2 A.n0 A.t1 148.35
R3 a_68_297.n1 a_68_297.t2 662.71
R4 a_68_297.n2 a_68_297.n1 260.308
R5 a_68_297.n1 a_68_297.n0 241.601
R6 a_68_297.n0 a_68_297.t4 236.18
R7 a_68_297.n0 a_68_297.t3 163.881
R8 a_68_297.t0 a_68_297.n2 38.5719
R9 a_68_297.n2 a_68_297.t1 38.5719
R10 VGND.n1 VGND.t2 253.421
R11 VGND.n1 VGND.n0 217.375
R12 VGND.n0 VGND.t0 55.7148
R13 VGND.n0 VGND.t1 26.8576
R14 VGND VGND.n1 0.437652
R15 VNB.t0 VNB.t1 1381.23
R16 VNB VNB.t2 1338.51
R17 VNB.t2 VNB.t0 1196.12
R18 B.n0 B.t0 192.639
R19 B B.n0 158.172
R20 B.n0 B.t1 134.799
R21 X.n0 X.t0 340.584
R22 X X.t1 174.464
R23 X.n0 X 2.4386
R24 X X.n0 1.43601
R25 a_150_297.t0 a_150_297.t1 98.5005
R26 VPWR VPWR.n0 320.877
R27 VPWR.n0 VPWR.t0 96.1553
R28 VPWR.n0 VPWR.t1 25.6105
R29 VPB VPB.t2 313.707
R30 VPB.t0 VPB.t1 287.072
R31 VPB.t2 VPB.t0 213.084
C0 B X 1.65e-19
C1 A VPB 0.030968f
C2 VGND VPWR 0.046447f
C3 B A 0.07509f
C4 VPWR X 0.128567f
C5 B VPB 0.046202f
C6 VGND X 0.113947f
C7 VPWR A 0.008464f
C8 VPWR VPB 0.080528f
C9 VGND A 0.034653f
C10 VGND VPB 0.011204f
C11 VPWR B 0.008552f
C12 A X 0.013051f
C13 X VPB 0.020902f
C14 VGND B 0.043653f
C15 VGND VNB 0.320425f
C16 X VNB 0.100952f
C17 A VNB 0.110717f
C18 B VNB 0.182719f
C19 VPWR VNB 0.268565f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297.t0 B.t0 a_39_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X.t2 a_39_297.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR.t1 a_39_297.t4 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X.t0 a_39_297.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND.t2 a_39_297.t6 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t2 A.t0 a_121_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND.t3 A.t1 a_39_297.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297.t1 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 B.n0 B.t1 193.303
R1 B B.n0 154.514
R2 B.n0 B.t0 135.463
R3 a_39_297.t0 a_39_297.n4 655.557
R4 a_39_297.n4 a_39_297.n3 262.327
R5 a_39_297.n4 a_39_297.n2 240.095
R6 a_39_297.n0 a_39_297.t4 212.081
R7 a_39_297.n1 a_39_297.t5 212.081
R8 a_39_297.n0 a_39_297.t6 139.78
R9 a_39_297.n1 a_39_297.t3 139.78
R10 a_39_297.n2 a_39_297.n0 41.6278
R11 a_39_297.n3 a_39_297.t2 38.5719
R12 a_39_297.n3 a_39_297.t1 38.5719
R13 a_39_297.n2 a_39_297.n1 19.7187
R14 a_121_297.t0 a_121_297.t1 98.5005
R15 VPB.t3 VPB.t1 298.911
R16 VPB.t1 VPB.t2 248.599
R17 VPB VPB.t0 224.923
R18 VPB.t0 VPB.t3 213.084
R19 VGND.n1 VGND.t2 284.966
R20 VGND.n5 VGND.t0 246.506
R21 VGND.n3 VGND.n2 202.474
R22 VGND.n2 VGND.t3 61.4291
R23 VGND.n4 VGND.n3 25.977
R24 VGND.n5 VGND.n4 25.977
R25 VGND.n2 VGND.t1 25.8467
R26 VGND.n6 VGND.n5 9.3005
R27 VGND.n4 VGND.n0 9.3005
R28 VGND.n3 VGND.n1 6.26408
R29 VGND.n1 VGND.n0 0.754779
R30 VGND.n6 VGND.n0 0.120292
R31 VGND VGND.n6 0.0213333
R32 X X.n0 304.012
R33 X X.n1 236.436
R34 X.n0 X.t3 26.5955
R35 X.n0 X.t0 26.5955
R36 X.n1 X.t1 24.9236
R37 X.n1 X.t2 24.9236
R38 VNB.t3 VNB.t2 1438.19
R39 VNB.t2 VNB.t1 1196.12
R40 VNB.t0 VNB.t3 1196.12
R41 VNB VNB.t0 911.327
R42 VPWR.n1 VPWR.t1 885.475
R43 VPWR.n1 VPWR.n0 328.57
R44 VPWR.n0 VPWR.t2 101.832
R45 VPWR.n0 VPWR.t0 26.596
R46 VPWR VPWR.n1 0.723344
R47 A.n0 A.t1 206.19
R48 A A.n0 154.744
R49 A.n0 A.t0 148.35
C0 VGND VPB 0.009551f
C1 X VPWR 0.165357f
C2 A B 0.07509f
C3 X VGND 0.098122f
C4 A VPWR 0.007338f
C5 X VPB 0.010843f
C6 VPWR B 0.005935f
C7 A VGND 0.050944f
C8 A VPB 0.031784f
C9 VGND B 0.03618f
C10 VPB B 0.041587f
C11 A X 0.014013f
C12 X B 1.51e-19
C13 VGND VPWR 0.047529f
C14 VPB VPWR 0.071364f
C15 VGND VNB 0.32269f
C16 X VNB 0.072361f
C17 A VNB 0.112463f
C18 B VNB 0.177703f
C19 VPWR VNB 0.283697f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_4 VNB VPB VGND VPWR B A X
X0 a_121_297.t0 B.t0 a_35_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1 VPWR.t4 a_35_297.t3 X.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2 X.t6 a_35_297.t4 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X.t3 a_35_297.t5 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4 X.t2 a_35_297.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t2 a_35_297.t7 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X.t4 a_35_297.t8 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X7 VGND.t2 a_35_297.t9 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t0 A.t0 a_121_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X9 VGND.t1 a_35_297.t10 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t5 A.t1 a_35_297.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_35_297.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t0 228.649
R1 B.n0 B.t1 156.35
R2 B B.n0 154.514
R3 a_35_297.t1 a_35_297.n10 229.608
R4 a_35_297.n1 a_35_297.t3 212.081
R5 a_35_297.n3 a_35_297.t4 212.081
R6 a_35_297.n5 a_35_297.t7 212.081
R7 a_35_297.n6 a_35_297.t8 212.081
R8 a_35_297.n2 a_35_297.n0 177.601
R9 a_35_297.n10 a_35_297.n9 152.671
R10 a_35_297.n4 a_35_297.n0 152
R11 a_35_297.n8 a_35_297.n7 152
R12 a_35_297.n1 a_35_297.t10 139.78
R13 a_35_297.n3 a_35_297.t6 139.78
R14 a_35_297.n5 a_35_297.t9 139.78
R15 a_35_297.n6 a_35_297.t5 139.78
R16 a_35_297.n10 a_35_297.n8 80.0602
R17 a_35_297.n2 a_35_297.n1 58.4247
R18 a_35_297.n4 a_35_297.n3 46.7399
R19 a_35_297.n7 a_35_297.n5 35.055
R20 a_35_297.n7 a_35_297.n6 26.2914
R21 a_35_297.n9 a_35_297.t2 24.9236
R22 a_35_297.n9 a_35_297.t0 24.9236
R23 a_35_297.n8 a_35_297.n0 22.5887
R24 a_35_297.n5 a_35_297.n4 14.6066
R25 a_35_297.n3 a_35_297.n2 2.92171
R26 a_121_297.t0 a_121_297.t1 41.3705
R27 VPB.t1 VPB.t2 298.911
R28 VPB.t4 VPB.t5 248.599
R29 VPB.t3 VPB.t4 248.599
R30 VPB.t2 VPB.t3 248.599
R31 VPB VPB.t0 224.923
R32 VPB.t0 VPB.t1 213.084
R33 X.n2 X.n0 340.637
R34 X.n2 X.n1 195.577
R35 X.n5 X.n3 137.189
R36 X.n5 X.n4 98.788
R37 X X.n5 36.7418
R38 X X.n2 28.2652
R39 X.n1 X.t7 26.5955
R40 X.n1 X.t6 26.5955
R41 X.n0 X.t5 26.5955
R42 X.n0 X.t4 26.5955
R43 X.n3 X.t1 24.9236
R44 X.n3 X.t3 24.9236
R45 X.n4 X.t0 24.9236
R46 X.n4 X.t2 24.9236
R47 VPWR.n3 VPWR.n2 607.212
R48 VPWR.n4 VPWR.t4 359.043
R49 VPWR.n8 VPWR.n1 320.223
R50 VPWR.n9 VPWR.n8 41.9179
R51 VPWR.n1 VPWR.t0 35.4605
R52 VPWR.n7 VPWR.n6 34.6358
R53 VPWR.n1 VPWR.t1 34.4755
R54 VPWR.n6 VPWR.n3 31.2476
R55 VPWR.n2 VPWR.t3 26.5955
R56 VPWR.n2 VPWR.t2 26.5955
R57 VPWR.n4 VPWR.n3 10.4058
R58 VPWR.n6 VPWR.n5 9.3005
R59 VPWR.n7 VPWR.n0 9.3005
R60 VPWR.n5 VPWR.n4 0.732469
R61 VPWR.n8 VPWR.n7 0.376971
R62 VPWR.n9 VPWR.n0 0.141672
R63 VPWR VPWR.n9 0.120476
R64 VPWR.n5 VPWR.n0 0.120292
R65 VGND.n5 VGND.t1 294.036
R66 VGND.n11 VGND.t0 276.098
R67 VGND.n9 VGND.n1 221.894
R68 VGND.n4 VGND.n3 208.719
R69 VGND.n8 VGND.n2 34.6358
R70 VGND.n10 VGND.n9 34.2593
R71 VGND.n1 VGND.t5 33.2313
R72 VGND.n1 VGND.t4 32.3082
R73 VGND.n4 VGND.n2 31.2476
R74 VGND.n11 VGND.n10 25.977
R75 VGND.n3 VGND.t3 24.9236
R76 VGND.n3 VGND.t2 24.9236
R77 VGND.n5 VGND.n4 10.4058
R78 VGND.n12 VGND.n11 9.3005
R79 VGND.n6 VGND.n2 9.3005
R80 VGND.n8 VGND.n7 9.3005
R81 VGND.n10 VGND.n0 9.3005
R82 VGND.n6 VGND.n5 0.732469
R83 VGND.n9 VGND.n8 0.376971
R84 VGND.n7 VGND.n6 0.120292
R85 VGND.n7 VGND.n0 0.120292
R86 VGND.n12 VGND.n0 0.120292
R87 VGND VGND.n12 0.0213333
R88 VNB.t5 VNB.t4 1438.19
R89 VNB.t3 VNB.t1 1196.12
R90 VNB.t2 VNB.t3 1196.12
R91 VNB.t4 VNB.t2 1196.12
R92 VNB.t0 VNB.t5 1196.12
R93 VNB VNB.t0 911.327
R94 A.n0 A.t0 241.536
R95 A.n0 A.t1 169.237
R96 A A.n0 156.655
C0 VGND B 0.043469f
C1 X A 0.001831f
C2 VPB B 0.040063f
C3 VPWR A 0.017354f
C4 VGND VPB 0.007212f
C5 X B 8.28e-20
C6 X VGND 0.279114f
C7 X VPB 0.014415f
C8 VPWR B 0.013865f
C9 B A 0.06146f
C10 VPWR VGND 0.067209f
C11 VPWR VPB 0.072286f
C12 VGND A 0.040051f
C13 VPB A 0.026073f
C14 VPWR X 0.3151f
C15 VGND VNB 0.420729f
C16 X VNB 0.061219f
C17 VPWR VNB 0.355695f
C18 A VNB 0.090802f
C19 B VNB 0.159752f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR VNB VPB A X B_N
X0 a_219_297.t2 a_27_53.t2 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X1 VGND.t2 B_N.t0 a_27_53.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t0 A.t0 a_301_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X.t1 a_219_297.t3 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_301_297.t1 a_27_53.t3 a_219_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X.t0 a_219_297.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6 a_27_53.t1 B_N.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND.t1 A.t1 a_219_297.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 a_27_53.n1 a_27_53.t1 672.086
R1 a_27_53.t0 a_27_53.n1 261.192
R2 a_27_53.n0 a_27_53.t2 186.03
R3 a_27_53.n1 a_27_53.n0 171.394
R4 a_27_53.n0 a_27_53.t3 137.829
R5 VGND.n3 VGND.n2 202.195
R6 VGND.n7 VGND.n6 185
R7 VGND.n9 VGND.n8 185
R8 VGND.n8 VGND.n7 137.143
R9 VGND.n2 VGND.t1 52.8576
R10 VGND.n7 VGND.t3 38.5719
R11 VGND.n8 VGND.t2 38.5719
R12 VGND.n10 VGND.n9 38.1787
R13 VGND.n6 VGND.n3 29.3949
R14 VGND.n2 VGND.t0 27.5691
R15 VGND.n1 VGND.n0 9.3005
R16 VGND.n5 VGND.n4 9.3005
R17 VGND.n5 VGND.n1 9.05896
R18 VGND.n4 VGND.n3 2.16256
R19 VGND.n6 VGND.n5 0.197423
R20 VGND.n9 VGND.n1 0.197423
R21 VGND.n4 VGND.n0 0.120292
R22 VGND.n10 VGND.n0 0.120292
R23 VGND VGND.n10 0.0213333
R24 a_219_297.n1 a_219_297.t1 731.812
R25 a_219_297.n2 a_219_297.n1 263.83
R26 a_219_297.n0 a_219_297.t4 240.484
R27 a_219_297.n0 a_219_297.t3 168.185
R28 a_219_297.n1 a_219_297.n0 152
R29 a_219_297.t0 a_219_297.n2 38.5719
R30 a_219_297.n2 a_219_297.t2 38.5719
R31 VNB.t1 VNB.t2 2563.11
R32 VNB.t0 VNB.t3 1395.47
R33 VNB.t2 VNB.t0 1196.12
R34 VNB VNB.t1 911.327
R35 B_N.n0 B_N.t0 185.376
R36 B_N B_N.n0 157.632
R37 B_N.n0 B_N.t1 137.177
R38 A A.t0 563.896
R39 A.t0 A.t1 392.027
R40 a_301_297.t0 a_301_297.t1 98.5005
R41 VPWR.n1 VPWR.t2 708.777
R42 VPWR.n1 VPWR.n0 321.704
R43 VPWR.n0 VPWR.t0 96.1553
R44 VPWR.n0 VPWR.t1 26.5955
R45 VPWR VPWR.n1 0.065704
R46 VPB.t3 VPB.t1 568.225
R47 VPB.t0 VPB.t2 290.031
R48 VPB.t1 VPB.t0 213.084
R49 VPB VPB.t3 189.409
R50 X X.t0 360.769
R51 X X.t1 287.072
C0 VGND VPWR 0.057039f
C1 VPB B_N 0.046613f
C2 A B_N 2.16e-19
C3 VPWR X 0.087835f
C4 VPB A 0.160525f
C5 VGND X 0.035406f
C6 VPWR B_N 0.037442f
C7 VPB VPWR 0.097059f
C8 VGND B_N 0.0173f
C9 VPWR A 0.194142f
C10 VPB VGND 0.009103f
C11 VGND A 0.01651f
C12 VPB X 0.010908f
C13 A X 0.002526f
C14 VGND VNB 0.353111f
C15 X VNB 0.08883f
C16 B_N VNB 0.169579f
C17 A VNB 0.135517f
C18 VPWR VNB 0.324987f
C19 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_2 VPWR VGND VNB VPB A B_N X
X0 VPWR.t2 A.t0 a_300_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297.t0 a_27_53.t2 VGND.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.15645 ps=1.165 w=0.42 l=0.15
X2 VGND.t4 B_N.t0 a_27_53.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.15645 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_300_297.t0 a_27_53.t3 a_218_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X.t1 a_218_297.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VPWR.t0 a_218_297.t4 X.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X.t2 a_218_297.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND.t0 a_218_297.t6 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_53.t0 B_N.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND.t3 A.t1 a_218_297.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 A A.t0 563.904
R1 A.t0 A.t1 392.027
R2 a_300_297.t0 a_300_297.t1 98.5005
R3 VPWR.n9 VPWR.t3 700.506
R4 VPWR.n3 VPWR.n2 315.406
R5 VPWR.n4 VPWR.t0 257.017
R6 VPWR.n2 VPWR.t2 96.1553
R7 VPWR.n7 VPWR.n1 34.6358
R8 VPWR.n8 VPWR.n7 34.6358
R9 VPWR.n2 VPWR.t1 26.5955
R10 VPWR.n9 VPWR.n8 25.977
R11 VPWR.n3 VPWR.n1 22.5887
R12 VPWR.n5 VPWR.n1 9.3005
R13 VPWR.n7 VPWR.n6 9.3005
R14 VPWR.n8 VPWR.n0 9.3005
R15 VPWR.n10 VPWR.n9 9.3005
R16 VPWR.n4 VPWR.n3 6.72481
R17 VPWR.n5 VPWR.n4 0.64287
R18 VPWR.n6 VPWR.n5 0.120292
R19 VPWR.n6 VPWR.n0 0.120292
R20 VPWR.n10 VPWR.n0 0.120292
R21 VPWR VPWR.n10 0.0213333
R22 VPB.t4 VPB.t2 565.265
R23 VPB.t3 VPB.t1 290.031
R24 VPB.t1 VPB.t0 248.599
R25 VPB.t2 VPB.t3 213.084
R26 VPB VPB.t4 189.409
R27 a_27_53.t0 a_27_53.n1 672.644
R28 a_27_53.n1 a_27_53.t1 261.13
R29 a_27_53.n0 a_27_53.t2 186.03
R30 a_27_53.n1 a_27_53.n0 171.394
R31 a_27_53.n0 a_27_53.t3 137.829
R32 VGND.n4 VGND.n3 198.475
R33 VGND.n10 VGND.n9 185
R34 VGND.n12 VGND.n11 185
R35 VGND.n5 VGND.t0 155.502
R36 VGND.n11 VGND.n10 135.714
R37 VGND.n3 VGND.t3 52.8576
R38 VGND.n10 VGND.t2 38.5719
R39 VGND.n11 VGND.t4 38.5719
R40 VGND.n13 VGND.n12 38.1787
R41 VGND.n3 VGND.t1 27.5691
R42 VGND.n9 VGND.n2 25.085
R43 VGND.n4 VGND.n2 16.5652
R44 VGND.n1 VGND.n0 9.3005
R45 VGND.n8 VGND.n7 9.3005
R46 VGND.n6 VGND.n2 9.3005
R47 VGND.n8 VGND.n1 9.05896
R48 VGND.n5 VGND.n4 6.62926
R49 VGND.n6 VGND.n5 0.662235
R50 VGND.n12 VGND.n1 0.197423
R51 VGND.n7 VGND.n6 0.120292
R52 VGND.n7 VGND.n0 0.120292
R53 VGND.n13 VGND.n0 0.120292
R54 VGND.n9 VGND.n8 0.0989615
R55 VGND VGND.n13 0.0226354
R56 a_218_297.n2 a_218_297.t1 731.812
R57 a_218_297.n3 a_218_297.n2 263.83
R58 a_218_297.n0 a_218_297.t4 212.081
R59 a_218_297.n1 a_218_297.t5 212.081
R60 a_218_297.n2 a_218_297.n1 162.225
R61 a_218_297.n0 a_218_297.t6 139.78
R62 a_218_297.n1 a_218_297.t3 139.78
R63 a_218_297.n1 a_218_297.n0 61.346
R64 a_218_297.n3 a_218_297.t2 38.5719
R65 a_218_297.t0 a_218_297.n3 38.5719
R66 VNB.t4 VNB.t0 2548.87
R67 VNB.t1 VNB.t3 1395.47
R68 VNB.t3 VNB.t2 1196.12
R69 VNB.t0 VNB.t1 1196.12
R70 VNB VNB.t4 925.567
R71 B_N.n0 B_N.t0 185.168
R72 B_N B_N.n0 157.632
R73 B_N.n0 B_N.t1 136.969
R74 X X.n0 300.495
R75 X X.n1 265.942
R76 X.n0 X.t3 26.5955
R77 X.n0 X.t2 26.5955
R78 X.n1 X.t0 24.9236
R79 X.n1 X.t1 24.9236
C0 VPB VPWR 0.11428f
C1 VPB A 0.162561f
C2 VPWR VGND 0.080505f
C3 A VGND 0.016862f
C4 VPWR X 0.166155f
C5 VPB VGND 0.011216f
C6 A X 0.002323f
C7 VPWR B_N 0.03796f
C8 VPB X 0.003951f
C9 A B_N 2.16e-19
C10 X VGND 0.075684f
C11 VPB B_N 0.046828f
C12 VPWR A 0.194451f
C13 B_N VGND 0.017333f
C14 VGND VNB 0.423661f
C15 X VNB 0.024711f
C16 B_N VNB 0.169989f
C17 A VNB 0.133481f
C18 VPWR VNB 0.398291f
C19 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_4 VNB VPB VGND VPWR X A B_N
X0 VPWR.t5 a_219_297.t3 X.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t6 B_N.t0 a_27_53.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.201775 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t0 A.t0 a_301_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.105 ps=1.21 w=1 l=0.15
X3 a_27_53.t0 B_N.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X.t7 a_219_297.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1105 ps=0.99 w=0.65 l=0.15
X5 a_301_297.t0 a_27_53.t2 a_219_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6 X.t3 a_219_297.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t1 A.t1 a_219_297.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t3 a_219_297.t6 X.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t4 a_219_297.t7 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X.t1 a_219_297.t8 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17 ps=1.34 w=1 l=0.15
X11 VGND.t3 a_219_297.t9 X.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_219_297.t0 a_27_53.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.201775 ps=1.4 w=0.65 l=0.15
X13 X.t0 a_219_297.t10 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_219_297.t2 a_219_297.n10 258.82
R1 a_219_297.n1 a_219_297.t3 212.081
R2 a_219_297.n3 a_219_297.t5 212.081
R3 a_219_297.n5 a_219_297.t6 212.081
R4 a_219_297.n6 a_219_297.t8 212.081
R5 a_219_297.n2 a_219_297.n0 177.601
R6 a_219_297.n10 a_219_297.n9 152.359
R7 a_219_297.n8 a_219_297.n7 152
R8 a_219_297.n4 a_219_297.n0 152
R9 a_219_297.n1 a_219_297.t9 139.78
R10 a_219_297.n3 a_219_297.t10 139.78
R11 a_219_297.n5 a_219_297.t7 139.78
R12 a_219_297.n6 a_219_297.t4 139.78
R13 a_219_297.n10 a_219_297.n8 105.035
R14 a_219_297.n7 a_219_297.n6 54.7732
R15 a_219_297.n5 a_219_297.n4 43.0884
R16 a_219_297.n3 a_219_297.n2 31.4035
R17 a_219_297.n2 a_219_297.n1 29.9429
R18 a_219_297.n8 a_219_297.n0 25.6005
R19 a_219_297.n9 a_219_297.t1 24.9236
R20 a_219_297.n9 a_219_297.t0 24.9236
R21 a_219_297.n4 a_219_297.n3 18.2581
R22 a_219_297.n7 a_219_297.n5 6.57323
R23 X.n2 X.n1 330.135
R24 X.n2 X.n0 197.011
R25 X.n5 X.n3 137.189
R26 X.n5 X.n4 98.788
R27 X X.n5 33.9562
R28 X.n0 X.t4 26.5955
R29 X.n0 X.t3 26.5955
R30 X.n1 X.t2 26.5955
R31 X.n1 X.t1 26.5955
R32 X.n3 X.t6 24.9236
R33 X.n3 X.t7 24.9236
R34 X.n4 X.t5 24.9236
R35 X.n4 X.t0 24.9236
R36 X X.n2 22.152
R37 VPWR.n14 VPWR.t1 669.907
R38 VPWR.n6 VPWR.n5 606.505
R39 VPWR.n4 VPWR.t5 351.957
R40 VPWR.n8 VPWR.n3 313.707
R41 VPWR.n3 VPWR.t0 39.4005
R42 VPWR.n12 VPWR.n1 34.6358
R43 VPWR.n13 VPWR.n12 34.6358
R44 VPWR.n3 VPWR.t2 27.5805
R45 VPWR.n5 VPWR.t4 26.5955
R46 VPWR.n5 VPWR.t3 26.5955
R47 VPWR.n14 VPWR.n13 25.977
R48 VPWR.n8 VPWR.n7 25.224
R49 VPWR.n8 VPWR.n1 22.9652
R50 VPWR.n7 VPWR.n6 19.2005
R51 VPWR.n7 VPWR.n2 9.3005
R52 VPWR.n9 VPWR.n8 9.3005
R53 VPWR.n10 VPWR.n1 9.3005
R54 VPWR.n12 VPWR.n11 9.3005
R55 VPWR.n13 VPWR.n0 9.3005
R56 VPWR.n15 VPWR.n14 9.3005
R57 VPWR.n6 VPWR.n4 6.81902
R58 VPWR.n4 VPWR.n2 0.780517
R59 VPWR.n9 VPWR.n2 0.120292
R60 VPWR.n10 VPWR.n9 0.120292
R61 VPWR.n11 VPWR.n10 0.120292
R62 VPWR.n11 VPWR.n0 0.120292
R63 VPWR.n15 VPWR.n0 0.120292
R64 VPWR VPWR.n15 0.0226354
R65 VPB.t1 VPB.t6 568.225
R66 VPB.t0 VPB.t2 290.031
R67 VPB.t4 VPB.t5 248.599
R68 VPB.t3 VPB.t4 248.599
R69 VPB.t2 VPB.t3 248.599
R70 VPB.t6 VPB.t0 213.084
R71 VPB VPB.t1 192.369
R72 B_N.n0 B_N.t1 323.55
R73 B_N.n0 B_N.t0 185.376
R74 B_N B_N.n0 153.673
R75 a_27_53.t0 a_27_53.n1 718.227
R76 a_27_53.n1 a_27_53.t1 265.216
R77 a_27_53.n0 a_27_53.t2 220.845
R78 a_27_53.n1 a_27_53.n0 205.312
R79 a_27_53.n0 a_27_53.t3 139.78
R80 VGND.n5 VGND.t3 283.193
R81 VGND.n6 VGND.n4 207.589
R82 VGND.n15 VGND.n14 191.169
R83 VGND.n17 VGND.n16 185
R84 VGND.n16 VGND.n15 128.234
R85 VGND.n9 VGND.n8 127.584
R86 VGND.n16 VGND.t6 38.5719
R87 VGND.n18 VGND.n17 38.1787
R88 VGND.n8 VGND.t1 37.8467
R89 VGND.n14 VGND.n2 29.1567
R90 VGND.n7 VGND.n6 28.6123
R91 VGND.n9 VGND.n7 28.2358
R92 VGND.n9 VGND.n2 27.8593
R93 VGND.n4 VGND.t2 24.9236
R94 VGND.n4 VGND.t4 24.9236
R95 VGND.n8 VGND.t5 24.9236
R96 VGND.n15 VGND.t0 18.5261
R97 VGND.n6 VGND.n5 12.9585
R98 VGND.n1 VGND.n0 9.3005
R99 VGND.n13 VGND.n12 9.3005
R100 VGND.n11 VGND.n2 9.3005
R101 VGND.n7 VGND.n3 9.3005
R102 VGND.n10 VGND.n9 9.3005
R103 VGND.n13 VGND.n1 9.05896
R104 VGND.n5 VGND.n3 0.815041
R105 VGND.n14 VGND.n13 0.197423
R106 VGND.n17 VGND.n1 0.197423
R107 VGND.n10 VGND.n3 0.120292
R108 VGND.n11 VGND.n10 0.120292
R109 VGND.n12 VGND.n11 0.120292
R110 VGND.n12 VGND.n0 0.120292
R111 VGND.n18 VGND.n0 0.120292
R112 VGND VGND.n18 0.0226354
R113 VNB.t6 VNB.t0 2563.11
R114 VNB.t1 VNB.t5 1395.47
R115 VNB.t2 VNB.t3 1196.12
R116 VNB.t4 VNB.t2 1196.12
R117 VNB.t5 VNB.t4 1196.12
R118 VNB.t0 VNB.t1 1196.12
R119 VNB VNB.t6 925.567
R120 A.n0 A.t0 241.536
R121 A.n0 A.t1 169.237
R122 A A.n0 160.641
R123 a_301_297.t0 a_301_297.t1 41.3705
C0 X VPB 0.014093f
C1 VGND VPWR 0.084798f
C2 B_N VPWR 0.048023f
C3 X VPWR 0.320016f
C4 VGND A 0.046099f
C5 VPB VPWR 0.100774f
C6 X A 7.12e-19
C7 VGND B_N 0.019357f
C8 VPB A 0.025902f
C9 X VGND 0.27702f
C10 X B_N 0.001049f
C11 VGND VPB 0.009008f
C12 VPB B_N 0.110915f
C13 A VPWR 0.021522f
C14 VGND VNB 0.49717f
C15 X VNB 0.059982f
C16 VPWR VNB 0.436103f
C17 A VNB 0.093384f
C18 B_N VNB 0.212799f
C19 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X.t0 a_29_53.t4 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297.t1 C.t0 a_29_53.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X.t1 a_29_53.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297.t0 B.t0 a_111_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR.t1 A.t0 a_183_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53.t3 B.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND.t2 C.t1 a_29_53.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND.t1 A.t1 a_29_53.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 a_29_53.t0 a_29_53.n3 779.24
R1 a_29_53.n1 a_29_53.t2 293.971
R2 a_29_53.n2 a_29_53.t4 241.536
R3 a_29_53.n1 a_29_53.n0 198.929
R4 a_29_53.n2 a_29_53.t5 169.237
R5 a_29_53.n3 a_29_53.n2 152
R6 a_29_53.n3 a_29_53.n1 63.3981
R7 a_29_53.n0 a_29_53.t1 38.5719
R8 a_29_53.n0 a_29_53.t3 38.5719
R9 VPWR VPWR.n0 321.644
R10 VPWR.n0 VPWR.t1 96.1553
R11 VPWR.n0 VPWR.t0 26.5955
R12 X X.t0 358.464
R13 X X.t1 286.675
R14 VPB.t3 VPB.t1 290.031
R15 VPB.t0 VPB.t3 284.113
R16 VPB.t2 VPB.t0 213.084
R17 VPB VPB.t2 201.246
R18 C.n0 C.t1 185.376
R19 C C.n0 156.462
R20 C.n0 C.t0 137.177
R21 a_111_297.t0 a_111_297.t1 98.5005
R22 VGND.n2 VGND.n1 205.815
R23 VGND.n2 VGND.n0 203.786
R24 VGND.n0 VGND.t1 52.8576
R25 VGND.n1 VGND.t3 38.5719
R26 VGND.n1 VGND.t2 38.5719
R27 VGND.n0 VGND.t0 27.5691
R28 VGND VGND.n2 0.56118
R29 VNB.t1 VNB.t0 1395.47
R30 VNB.t3 VNB.t1 1196.12
R31 VNB.t2 VNB.t3 1196.12
R32 VNB VNB.t2 968.285
R33 B.t0 B.t1 378.255
R34 B B.t0 329.56
R35 a_183_297.t0 a_183_297.t1 154.786
R36 A.n0 A.t1 196.549
R37 A A.n0 161.504
R38 A.n0 A.t0 148.35
R39 A A.n1 14.1581
R40 A.n1 A 7.87742
R41 A.n1 A 3.68535
C0 C VGND 0.016088f
C1 A X 0.001269f
C2 VPWR A 0.009364f
C3 B C 0.080229f
C4 B VGND 0.0152f
C5 A VPB 0.037711f
C6 X VGND 0.035971f
C7 VPWR C 0.004565f
C8 B X 6.52e-19
C9 VPWR VGND 0.045852f
C10 C VPB 0.039602f
C11 VGND VPB 0.007241f
C12 VPWR B 0.147145f
C13 VPWR X 0.088535f
C14 C A 0.034282f
C15 B VPB 0.096179f
C16 A VGND 0.018737f
C17 X VPB 0.010881f
C18 B A 0.07874f
C19 VPWR VPB 0.064885f
C20 VGND VNB 0.306355f
C21 X VNB 0.088191f
C22 A VNB 0.117495f
C23 C VNB 0.160014f
C24 B VNB 0.116674f
C25 VPWR VNB 0.252671f
C26 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR.t2 a_30_53.t4 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t3 a_30_53.t5 X.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X.t0 a_30_53.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297.t0 C.t0 a_30_53.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X.t2 a_30_53.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VGND.t0 A.t0 a_30_53.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53.t2 B.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND.t1 C.t1 a_30_53.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297.t0 B.t1 a_112_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR.t0 A.t1 a_184_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
R0 a_30_53.n2 a_30_53.t3 779.13
R1 a_30_53.n3 a_30_53.t1 293.971
R2 a_30_53.n0 a_30_53.t4 212.081
R3 a_30_53.n1 a_30_53.t6 212.081
R4 a_30_53.n4 a_30_53.n3 198.929
R5 a_30_53.n2 a_30_53.n1 155.653
R6 a_30_53.n0 a_30_53.t5 139.78
R7 a_30_53.n1 a_30_53.t7 139.78
R8 a_30_53.n3 a_30_53.n2 63.3981
R9 a_30_53.n1 a_30_53.n0 61.346
R10 a_30_53.t0 a_30_53.n4 38.5719
R11 a_30_53.n4 a_30_53.t2 38.5719
R12 X X.n0 299.197
R13 X X.n1 261.752
R14 X.n0 X.t1 26.5955
R15 X.n0 X.t0 26.5955
R16 X.n1 X.t3 24.9236
R17 X.n1 X.t2 24.9236
R18 VPWR.n1 VPWR.n0 320.846
R19 VPWR.n1 VPWR.t2 260.173
R20 VPWR.n0 VPWR.t0 96.1553
R21 VPWR.n0 VPWR.t1 26.5955
R22 VPWR VPWR.n1 0.741478
R23 VPB.t0 VPB.t1 290.031
R24 VPB.t3 VPB.t0 284.113
R25 VPB.t1 VPB.t2 248.599
R26 VPB.t4 VPB.t3 213.084
R27 VPB VPB.t4 201.246
R28 VGND.n6 VGND.n5 200.516
R29 VGND.n3 VGND.n2 198.475
R30 VGND.n1 VGND.t3 150.135
R31 VGND.n2 VGND.t0 52.8576
R32 VGND.n5 VGND.t4 38.5719
R33 VGND.n5 VGND.t1 38.5719
R34 VGND.n2 VGND.t2 27.5691
R35 VGND.n6 VGND.n4 21.8358
R36 VGND.n4 VGND.n3 16.5652
R37 VGND.n4 VGND.n0 9.3005
R38 VGND.n7 VGND.n6 7.18025
R39 VGND.n3 VGND.n1 6.6817
R40 VGND.n1 VGND.n0 0.619035
R41 VGND.n7 VGND.n0 0.147761
R42 VGND VGND.n7 0.11561
R43 VNB.t0 VNB.t2 1395.47
R44 VNB.t2 VNB.t3 1196.12
R45 VNB.t4 VNB.t0 1196.12
R46 VNB.t1 VNB.t4 1196.12
R47 VNB VNB.t1 968.285
R48 C.n0 C.t1 185.168
R49 C C.n0 156.268
R50 C.n0 C.t0 136.969
R51 a_112_297.t0 a_112_297.t1 98.5005
R52 A.n0 A.t0 196.549
R53 A A.n0 161.504
R54 A.n0 A.t1 148.35
R55 A.n1 A 13.5763
R56 A.n1 A 6.82717
R57 A A.n1 4.26717
R58 B.t1 B.t0 378.255
R59 B B.t1 329.56
R60 a_184_297.t0 a_184_297.t1 154.786
C0 VPWR X 0.176032f
C1 B A 0.078772f
C2 VPB VGND 0.008444f
C3 A VGND 0.019219f
C4 VPB VPWR 0.081821f
C5 B C 0.08024f
C6 VPB X 0.00385f
C7 VPWR A 0.009818f
C8 C VGND 0.016263f
C9 A X 0.001292f
C10 VPWR C 0.004588f
C11 VPB A 0.038249f
C12 B VGND 0.0151f
C13 VPB C 0.039896f
C14 VPWR B 0.14788f
C15 B X 6.52e-19
C16 VPWR VGND 0.071169f
C17 C A 0.034282f
C18 X VGND 0.078621f
C19 VPB B 0.097241f
C20 VGND VNB 0.380303f
C21 X VNB 0.024476f
C22 A VNB 0.116974f
C23 C VNB 0.16054f
C24 B VNB 0.115702f
C25 VPWR VNB 0.330061f
C26 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3_4 VPB VNB VPWR VGND B C A X
X0 X.t7 a_27_47.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X.t3 a_27_47.t5 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X.t6 a_27_47.t6 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t3 a_27_47.t7 X.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t4 A.t0 a_193_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297.t1 B.t0 a_109_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t2 a_27_47.t8 X.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t2 a_27_47.t9 X.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X.t1 a_27_47.t10 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR.t0 a_27_47.t11 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297.t0 C.t0 a_27_47.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND.t6 C.t1 a_27_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t2 a_27_47.n13 381.998
R1 a_27_47.n4 a_27_47.t8 212.081
R2 a_27_47.n5 a_27_47.t10 212.081
R3 a_27_47.n10 a_27_47.t11 212.081
R4 a_27_47.n12 a_27_47.t5 212.081
R5 a_27_47.n13 a_27_47.n12 180.482
R6 a_27_47.n7 a_27_47.n6 177.601
R7 a_27_47.n2 a_27_47.t3 174.017
R8 a_27_47.n11 a_27_47.n0 152
R9 a_27_47.n9 a_27_47.n8 152
R10 a_27_47.n7 a_27_47.n3 152
R11 a_27_47.n4 a_27_47.t7 139.78
R12 a_27_47.n5 a_27_47.t6 139.78
R13 a_27_47.n10 a_27_47.t9 139.78
R14 a_27_47.n12 a_27_47.t4 139.78
R15 a_27_47.n2 a_27_47.n1 98.5941
R16 a_27_47.n13 a_27_47.n2 63.0954
R17 a_27_47.n9 a_27_47.n3 49.6611
R18 a_27_47.n6 a_27_47.n5 47.4702
R19 a_27_47.n11 a_27_47.n10 40.1672
R20 a_27_47.n8 a_27_47.n7 25.6005
R21 a_27_47.n8 a_27_47.n0 25.6005
R22 a_27_47.n1 a_27_47.t1 24.9236
R23 a_27_47.n1 a_27_47.t0 24.9236
R24 a_27_47.n13 a_27_47.n0 23.7181
R25 a_27_47.n12 a_27_47.n11 21.1793
R26 a_27_47.n6 a_27_47.n4 13.8763
R27 a_27_47.n10 a_27_47.n9 9.49444
R28 a_27_47.n5 a_27_47.n3 2.19141
R29 VGND.n6 VGND.t3 284.86
R30 VGND.n5 VGND.n4 207.965
R31 VGND.n18 VGND.n1 207.965
R32 VGND.n10 VGND.n2 185
R33 VGND.n12 VGND.n11 185
R34 VGND.n11 VGND.n10 97.8467
R35 VGND.n19 VGND.n18 43.1829
R36 VGND.n17 VGND.n16 34.6358
R37 VGND.n9 VGND.n8 31.0417
R38 VGND.n8 VGND.n5 27.1064
R39 VGND.n11 VGND.t5 24.9236
R40 VGND.n10 VGND.t1 24.9236
R41 VGND.n4 VGND.t4 24.9236
R42 VGND.n4 VGND.t2 24.9236
R43 VGND.n1 VGND.t0 24.9236
R44 VGND.n1 VGND.t6 24.9236
R45 VGND.n16 VGND.n2 23.1593
R46 VGND.n6 VGND.n5 14.4172
R47 VGND.n17 VGND.n0 9.3005
R48 VGND.n16 VGND.n15 9.3005
R49 VGND.n14 VGND.n13 9.3005
R50 VGND.n8 VGND.n7 9.3005
R51 VGND.n9 VGND.n3 9.3005
R52 VGND.n13 VGND.n12 8.8005
R53 VGND.n13 VGND.n2 1.8005
R54 VGND.n7 VGND.n6 0.862225
R55 VGND.n18 VGND.n17 0.753441
R56 VGND.n12 VGND.n9 0.4005
R57 VGND.n7 VGND.n3 0.120292
R58 VGND.n14 VGND.n3 0.120292
R59 VGND.n15 VGND.n14 0.120292
R60 VGND.n15 VGND.n0 0.120292
R61 VGND.n19 VGND.n0 0.120292
R62 VGND VGND.n19 0.0213333
R63 X.n5 X.n3 252.931
R64 X.n5 X.n4 208.507
R65 X.n2 X.n0 137.576
R66 X.n2 X.n1 99.1759
R67 X.n6 X.n5 56.6269
R68 X.n3 X.t0 26.5955
R69 X.n3 X.t3 26.5955
R70 X.n4 X.t2 26.5955
R71 X.n4 X.t1 26.5955
R72 X.n0 X.t4 24.9236
R73 X.n0 X.t7 24.9236
R74 X.n1 X.t5 24.9236
R75 X.n1 X.t6 24.9236
R76 X.n6 X.n2 21.8358
R77 X X.n6 2.42809
R78 VNB.t1 VNB.t5 2705.5
R79 VNB.t4 VNB.t3 1196.12
R80 VNB.t2 VNB.t4 1196.12
R81 VNB.t5 VNB.t2 1196.12
R82 VNB.t0 VNB.t1 1196.12
R83 VNB.t6 VNB.t0 1196.12
R84 VNB VNB.t6 911.327
R85 VPWR.n3 VPWR.n1 585
R86 VPWR.n2 VPWR.n1 585
R87 VPWR.n6 VPWR.t2 352.238
R88 VPWR.n8 VPWR.n7 318.293
R89 VPWR.n5 VPWR.n4 271.262
R90 VPWR.n4 VPWR.n3 42.4778
R91 VPWR.n4 VPWR.n2 42.4778
R92 VPWR.n3 VPWR.t4 39.4005
R93 VPWR.n10 VPWR.n9 29.7417
R94 VPWR.n2 VPWR.t3 26.5955
R95 VPWR.n7 VPWR.t1 26.5955
R96 VPWR.n7 VPWR.t0 26.5955
R97 VPWR.n9 VPWR.n8 17.6946
R98 VPWR.n9 VPWR.n0 9.3005
R99 VPWR.n10 VPWR.n5 6.94907
R100 VPWR.n8 VPWR.n6 6.81832
R101 VPWR.n5 VPWR.n1 6.21764
R102 VPWR.n11 VPWR.n10 3.96366
R103 VPWR.n6 VPWR.n0 0.837252
R104 VPWR VPWR.n11 0.413273
R105 VPWR.n11 VPWR.n0 0.208849
R106 VPB.t5 VPB.t4 562.306
R107 VPB.t2 VPB.t3 248.599
R108 VPB.t1 VPB.t2 248.599
R109 VPB.t4 VPB.t1 248.599
R110 VPB.t6 VPB.t5 248.599
R111 VPB.t0 VPB.t6 248.599
R112 VPB VPB.t0 189.409
R113 A.n0 A.t0 239.505
R114 A.n0 A.t1 167.204
R115 A A.n0 159.168
R116 a_193_297.t0 a_193_297.t1 53.1905
R117 B.n0 B.t0 241.536
R118 B.n0 B.t1 169.237
R119 B B.n0 167.752
R120 a_109_297.t0 a_109_297.t1 53.1905
R121 C.n0 C.t0 231.017
R122 C.n0 C.t1 158.716
R123 C C.n0 157.632
C0 X VPB 0.014642f
C1 VPWR C 0.009207f
C2 VGND A 0.016419f
C3 VPB C 0.036876f
C4 B A 0.078254f
C5 VPWR VPB 0.08674f
C6 VGND B 0.016256f
C7 X A 5.59e-19
C8 X VGND 0.264606f
C9 VPWR A 0.019597f
C10 VGND C 0.014913f
C11 VPB A 0.032433f
C12 C B 0.086443f
C13 VPWR VGND 0.086422f
C14 VPWR B 0.013194f
C15 VGND VPB 0.006984f
C16 VPB B 0.030241f
C17 VPWR X 0.365404f
C18 VGND VNB 0.493458f
C19 X VNB 0.061057f
C20 VPWR VNB 0.417624f
C21 A VNB 0.098686f
C22 B VNB 0.093805f
C23 C VNB 0.140554f
C24 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93.t0 C_N.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53.t0 B.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND.t3 a_109_93.t2 a_215_53.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND.t0 A.t0 a_215_53.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR.t2 A.t1 a_369_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297.t0 B.t1 a_297_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X.t0 a_215_53.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297.t1 a_109_93.t3 a_215_53.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93.t1 C_N.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X.t1 a_215_53.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
R0 C_N C_N.n0 157.632
R1 C_N.n0 C_N.t1 137.177
R2 C_N.n0 C_N.t0 121.109
R3 VGND.n8 VGND.t2 259.51
R4 VGND.n4 VGND.n3 203.887
R5 VGND.n2 VGND.n1 200.516
R6 VGND.n3 VGND.t0 51.4291
R7 VGND.n1 VGND.t4 38.5719
R8 VGND.n1 VGND.t3 38.5719
R9 VGND.n7 VGND.n6 34.6358
R10 VGND.n3 VGND.t1 28.3801
R11 VGND.n8 VGND.n7 25.977
R12 VGND.n6 VGND.n2 22.9652
R13 VGND.n9 VGND.n8 9.3005
R14 VGND.n6 VGND.n5 9.3005
R15 VGND.n7 VGND.n0 9.3005
R16 VGND.n4 VGND.n2 6.46566
R17 VGND.n5 VGND.n4 0.656389
R18 VGND.n5 VGND.n0 0.120292
R19 VGND.n9 VGND.n0 0.120292
R20 VGND VGND.n9 0.0226354
R21 a_109_93.n1 a_109_93.t1 672.838
R22 a_109_93.t0 a_109_93.n1 234.579
R23 a_109_93.n0 a_109_93.t2 183.492
R24 a_109_93.n1 a_109_93.n0 168.097
R25 a_109_93.n0 a_109_93.t3 135.292
R26 VNB.t2 VNB.t3 2677.02
R27 VNB.t0 VNB.t1 1381.23
R28 VNB.t4 VNB.t0 1196.12
R29 VNB.t3 VNB.t4 1196.12
R30 VNB VNB.t2 925.567
R31 B.t1 B.t0 378.255
R32 B B.t1 318.055
R33 a_215_53.n1 a_215_53.t3 779.13
R34 a_215_53.n2 a_215_53.t2 296.173
R35 a_215_53.n0 a_215_53.t4 241.536
R36 a_215_53.n3 a_215_53.n2 198.929
R37 a_215_53.n0 a_215_53.t5 169.237
R38 a_215_53.n1 a_215_53.n0 152
R39 a_215_53.n2 a_215_53.n1 63.0217
R40 a_215_53.n3 a_215_53.t1 38.5719
R41 a_215_53.t0 a_215_53.n3 38.5719
R42 A.n0 A.t0 267.065
R43 A A.n0 161.504
R44 A.n0 A.t1 148.35
R45 A A.n1 13.1884
R46 A.n1 A 5.29705
R47 A.n1 A 4.65505
R48 a_369_297.t0 a_369_297.t1 152.44
R49 VPWR.n1 VPWR.t0 707.763
R50 VPWR.n1 VPWR.n0 321.83
R51 VPWR.n0 VPWR.t2 96.1553
R52 VPWR.n0 VPWR.t1 26.5955
R53 VPWR VPWR.n1 0.0570582
R54 VPB.t1 VPB.t3 556.386
R55 VPB.t4 VPB.t2 290.031
R56 VPB.t0 VPB.t4 281.154
R57 VPB.t3 VPB.t0 213.084
R58 VPB VPB.t1 192.369
R59 a_297_297.t0 a_297_297.t1 98.5005
R60 X X.t0 359.536
R61 X X.t1 286.675
C0 VGND A 0.018847f
C1 C_N VPWR 0.037773f
C2 A VPB 0.03757f
C3 A X 0.001274f
C4 VGND C_N 0.042739f
C5 C_N VPB 0.046442f
C6 B VPWR 0.234984f
C7 C_N X 1.86e-20
C8 VGND VPWR 0.06567f
C9 VGND B 0.015735f
C10 VPB VPWR 0.109107f
C11 B VPB 0.110475f
C12 X VPWR 0.088522f
C13 B X 6.53e-19
C14 VGND VPB 0.010346f
C15 VGND X 0.035902f
C16 A VPWR 0.009622f
C17 X VPB 0.010957f
C18 B A 0.079275f
C19 VGND VNB 0.439259f
C20 X VNB 0.08839f
C21 A VNB 0.112741f
C22 C_N VNB 0.150085f
C23 B VNB 0.103426f
C24 VPWR VNB 0.362977f
C25 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR.t1 C_N.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND.t4 a_176_21.t4 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X.t2 a_176_21.t5 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR.t2 a_176_21.t6 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t1 B.t0 a_176_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X.t0 a_176_21.t7 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21.t2 a_27_47.t2 a_472_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297.t0 B.t1 a_388_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21.t1 A.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10 a_176_21.t3 a_27_47.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND.t0 C_N.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A.n0 A.t1 196.549
R1 A A.n0 154.964
R2 A.n0 A.t0 148.35
R3 VPWR.n2 VPWR.n1 662.133
R4 VPWR.n2 VPWR.n0 610.341
R5 VPWR.n0 VPWR.t0 98.5005
R6 VPWR.n1 VPWR.t1 96.1553
R7 VPWR.n1 VPWR.t3 34.3058
R8 VPWR.n0 VPWR.t2 25.6105
R9 VPWR VPWR.n2 0.555057
R10 a_388_297.t0 a_388_297.t1 126.644
R11 VPB.t3 VPB.t0 290.031
R12 VPB.t2 VPB.t4 287.072
R13 VPB.t5 VPB.t1 248.599
R14 VPB.t0 VPB.t5 248.599
R15 VPB.t4 VPB.t3 248.599
R16 VPB VPB.t2 189.409
R17 C_N.n0 C_N.t0 238.397
R18 C_N.n0 C_N.t1 195.017
R19 C_N C_N.n0 154.493
R20 a_27_47.t0 a_27_47.n1 669.62
R21 a_27_47.n1 a_27_47.t1 334.906
R22 a_27_47.n1 a_27_47.n0 330.421
R23 a_27_47.n0 a_27_47.t3 196.549
R24 a_27_47.n0 a_27_47.t2 148.35
R25 a_176_21.n1 a_176_21.t2 712.27
R26 a_176_21.n1 a_176_21.t3 230.349
R27 a_176_21.n3 a_176_21.n0 221.07
R28 a_176_21.n0 a_176_21.t6 212.081
R29 a_176_21.n2 a_176_21.t7 212.081
R30 a_176_21.n4 a_176_21.n3 205.329
R31 a_176_21.n0 a_176_21.t4 139.78
R32 a_176_21.n2 a_176_21.t5 139.78
R33 a_176_21.n0 a_176_21.n2 61.346
R34 a_176_21.n3 a_176_21.n1 57.7203
R35 a_176_21.t0 a_176_21.n4 38.5719
R36 a_176_21.n4 a_176_21.t1 38.5719
R37 X.n2 X.n0 667.854
R38 X.n2 X.n1 185
R39 X.n0 X.t1 26.5955
R40 X.n0 X.t0 26.5955
R41 X.n1 X.t3 24.9236
R42 X.n1 X.t2 24.9236
R43 X X.n2 0.183357
R44 VGND.n3 VGND.n2 208.719
R45 VGND.n9 VGND.n1 208.719
R46 VGND.n5 VGND.n4 206.101
R47 VGND.n2 VGND.t2 52.8576
R48 VGND.n1 VGND.t3 44.0005
R49 VGND.n10 VGND.n9 43.1829
R50 VGND.n4 VGND.t5 38.5719
R51 VGND.n4 VGND.t1 38.5719
R52 VGND.n1 VGND.t0 38.5719
R53 VGND.n8 VGND.n7 34.6358
R54 VGND.n7 VGND.n3 34.2593
R55 VGND.n2 VGND.t4 28.3166
R56 VGND.n8 VGND.n0 9.3005
R57 VGND.n7 VGND.n6 9.3005
R58 VGND.n5 VGND.n3 7.61135
R59 VGND.n9 VGND.n8 0.753441
R60 VGND.n6 VGND.n5 0.490177
R61 VGND.n6 VGND.n0 0.120292
R62 VGND.n10 VGND.n0 0.120292
R63 VGND VGND.n10 0.0226354
R64 VNB.t4 VNB.t2 1395.47
R65 VNB.t0 VNB.t3 1381.23
R66 VNB.t1 VNB.t5 1196.12
R67 VNB.t2 VNB.t1 1196.12
R68 VNB.t3 VNB.t4 1196.12
R69 VNB VNB.t0 925.567
R70 B.t1 B.t0 392.027
R71 B B.t1 325.118
R72 a_472_297.t0 a_472_297.t1 126.644
C0 X A 0.013329f
C1 C_N VGND 0.017227f
C2 VPWR X 0.014357f
C3 B VPB 0.095043f
C4 A VGND 0.016504f
C5 VPWR VGND 0.064268f
C6 C_N A 0.002835f
C7 VPWR C_N 0.01171f
C8 X B 6.04e-19
C9 X VPB 0.00308f
C10 VPWR A 0.008235f
C11 B VGND 0.015106f
C12 VPB VGND 0.008614f
C13 C_N B 0.001496f
C14 C_N VPB 0.079431f
C15 B A 0.077538f
C16 X VGND 0.096191f
C17 VPB A 0.035979f
C18 C_N X 0.002709f
C19 VPWR B 0.121785f
C20 VPWR VPB 0.085809f
C21 VGND VNB 0.398057f
C22 A VNB 0.106442f
C23 B VNB 0.107892f
C24 X VNB 0.003804f
C25 C_N VNB 0.190285f
C26 VPWR VNB 0.33505f
C27 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_4 VNB VPB VGND VPWR C_N X A B
X0 a_176_21.t3 a_27_47.t2 a_626_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1 a_626_297.t0 B.t0 a_542_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 C_N.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND.t7 a_176_21.t4 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_542_297.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t2 a_176_21.t5 X.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X.t2 a_176_21.t6 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t6 a_176_21.t7 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X8 X.t5 a_176_21.t8 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_176_21.t1 A.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR.t3 a_176_21.t9 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 X.t0 a_176_21.t10 VPWR.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X12 a_176_21.t2 a_27_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X13 VGND.t4 a_176_21.t11 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t2 B.t1 a_176_21.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t0 C_N.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t0 a_27_47.n1 669.62
R1 a_27_47.n1 a_27_47.n0 396.721
R2 a_27_47.n1 a_27_47.t1 334.906
R3 a_27_47.n0 a_27_47.t2 241.536
R4 a_27_47.n0 a_27_47.t3 169.237
R5 a_626_297.t0 a_626_297.t1 65.0105
R6 a_176_21.t3 a_176_21.n9 928.168
R7 a_176_21.n9 a_176_21.t2 216.701
R8 a_176_21.n4 a_176_21.t5 212.081
R9 a_176_21.n5 a_176_21.t6 212.081
R10 a_176_21.n2 a_176_21.t9 212.081
R11 a_176_21.n1 a_176_21.t10 212.081
R12 a_176_21.n8 a_176_21.n0 198.929
R13 a_176_21.n7 a_176_21.n6 152
R14 a_176_21.n4 a_176_21.t11 139.78
R15 a_176_21.n5 a_176_21.t8 139.78
R16 a_176_21.n2 a_176_21.t4 139.78
R17 a_176_21.n1 a_176_21.t7 139.78
R18 a_176_21.n7 a_176_21.n3 96.7795
R19 a_176_21.n9 a_176_21.n8 68.6379
R20 a_176_21.n8 a_176_21.n7 65.4619
R21 a_176_21.n2 a_176_21.n1 61.346
R22 a_176_21.n6 a_176_21.n5 47.4702
R23 a_176_21.n3 a_176_21.n2 32.75
R24 a_176_21.n0 a_176_21.t0 24.9236
R25 a_176_21.n0 a_176_21.t1 24.9236
R26 a_176_21.n5 a_176_21.n3 22.0949
R27 a_176_21.n6 a_176_21.n4 13.8763
R28 VPB.t1 VPB.t4 287.072
R29 VPB.t2 VPB.t3 284.113
R30 VPB.t0 VPB.t2 248.599
R31 VPB.t7 VPB.t0 248.599
R32 VPB.t6 VPB.t7 248.599
R33 VPB.t5 VPB.t6 248.599
R34 VPB.t4 VPB.t5 248.599
R35 VPB VPB.t1 189.409
R36 B.n0 B.t0 241.536
R37 B.n0 B.t1 169.237
R38 B B.n0 155.722
R39 a_542_297.t0 a_542_297.t1 53.1905
R40 C_N.n0 C_N.t0 238.397
R41 C_N.n0 C_N.t1 195.017
R42 C_N C_N.n0 154.493
R43 VPWR.n7 VPWR.n1 656.938
R44 VPWR.n3 VPWR.n2 606.128
R45 VPWR.n5 VPWR.n4 601.486
R46 VPWR.n1 VPWR.t1 96.1553
R47 VPWR.n1 VPWR.t5 34.3058
R48 VPWR.n4 VPWR.t4 26.5955
R49 VPWR.n4 VPWR.t3 26.5955
R50 VPWR.n2 VPWR.t0 26.5955
R51 VPWR.n2 VPWR.t2 26.5955
R52 VPWR.n6 VPWR.n5 20.3299
R53 VPWR.n7 VPWR.n6 18.0711
R54 VPWR.n6 VPWR.n0 9.3005
R55 VPWR.n8 VPWR.n7 7.25484
R56 VPWR.n5 VPWR.n3 6.57973
R57 VPWR.n3 VPWR.n0 0.680178
R58 VPWR.n8 VPWR.n0 0.146813
R59 VPWR VPWR.n8 0.115269
R60 X X.n0 585.674
R61 X.n5 X.n4 585
R62 X.n3 X.n2 263.635
R63 X.n3 X.n1 95.684
R64 X.n5 X.n3 55.8304
R65 X X.n5 37.0531
R66 X.n4 X.t1 26.5955
R67 X.n4 X.t0 26.5955
R68 X.n0 X.t3 26.5955
R69 X.n0 X.t2 26.5955
R70 X.n1 X.t7 24.9236
R71 X.n1 X.t6 24.9236
R72 X.n2 X.t4 24.9236
R73 X.n2 X.t5 24.9236
R74 VGND.n11 VGND.n3 208.719
R75 VGND.n1 VGND.n0 208.719
R76 VGND.n7 VGND.n6 202.81
R77 VGND.n5 VGND.n4 200.516
R78 VGND.n0 VGND.t0 45.7148
R79 VGND.n0 VGND.t6 36.8576
R80 VGND.n6 VGND.t3 36.0005
R81 VGND.n10 VGND.n9 34.6358
R82 VGND.n12 VGND.n1 33.5064
R83 VGND.n12 VGND.n11 32.7534
R84 VGND.n6 VGND.t2 24.9236
R85 VGND.n4 VGND.t1 24.9236
R86 VGND.n4 VGND.t4 24.9236
R87 VGND.n3 VGND.t5 24.9236
R88 VGND.n3 VGND.t7 24.9236
R89 VGND.n9 VGND.n5 14.3064
R90 VGND.n13 VGND.n12 9.3005
R91 VGND.n10 VGND.n2 9.3005
R92 VGND.n9 VGND.n8 9.3005
R93 VGND.n14 VGND.n1 8.78851
R94 VGND.n7 VGND.n5 6.79197
R95 VGND.n11 VGND.n10 1.88285
R96 VGND.n8 VGND.n7 0.725498
R97 VGND.n14 VGND.n13 0.141672
R98 VGND VGND.n14 0.120476
R99 VGND.n8 VGND.n2 0.120292
R100 VGND.n13 VGND.n2 0.120292
R101 VNB.t0 VNB.t6 1381.23
R102 VNB.t2 VNB.t3 1366.99
R103 VNB.t1 VNB.t2 1196.12
R104 VNB.t4 VNB.t1 1196.12
R105 VNB.t5 VNB.t4 1196.12
R106 VNB.t7 VNB.t5 1196.12
R107 VNB.t6 VNB.t7 1196.12
R108 VNB VNB.t0 911.327
R109 A.n0 A.t0 241.536
R110 A A.n0 177.504
R111 A.n0 A.t1 169.237
C0 B VGND 0.015316f
C1 B VPWR 0.012007f
C2 A VGND 0.016192f
C3 VPWR A 0.018856f
C4 C_N VPB 0.080628f
C5 C_N X 0.004783f
C6 VPB VGND 0.006839f
C7 X VGND 0.207334f
C8 VPWR VPB 0.087194f
C9 B A 0.116718f
C10 VPWR X 0.032126f
C11 C_N VGND 0.017158f
C12 B VPB 0.0279f
C13 VPWR C_N 0.011811f
C14 VPB A 0.027687f
C15 X A 0.02614f
C16 VPWR VGND 0.082157f
C17 B C_N 8.7e-20
C18 C_N A 1.35e-19
C19 X VPB 0.005746f
C20 VGND VNB 0.486196f
C21 X VNB 0.008146f
C22 C_N VNB 0.192964f
C23 VPWR VNB 0.410093f
C24 B VNB 0.089115f
C25 A VNB 0.087932f
C26 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297.t3 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297.t1 D.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297.t1 B.t1 a_205_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR.t1 A.t0 a_277_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X.t1 a_27_297.t5 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297.t1 C.t0 a_109_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X.t0 a_27_297.t6 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND.t0 C.t1 a_27_297.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297.t1 D.t1 a_27_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND.t4 A.t1 a_27_297.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 B.t1 B.t0 618.109
R1 B B.t1 329.56
R2 VGND.n6 VGND.t1 242.965
R3 VGND.n2 VGND.n1 203.697
R4 VGND.n4 VGND.n3 200.516
R5 VGND.n1 VGND.t4 52.8576
R6 VGND.n3 VGND.t2 38.5719
R7 VGND.n3 VGND.t0 38.5719
R8 VGND.n1 VGND.t3 27.5691
R9 VGND.n5 VGND.n4 22.9652
R10 VGND.n6 VGND.n5 19.9534
R11 VGND.n7 VGND.n6 9.3005
R12 VGND.n5 VGND.n0 9.3005
R13 VGND.n4 VGND.n2 6.46652
R14 VGND.n2 VGND.n0 0.655453
R15 VGND.n7 VGND.n0 0.120292
R16 VGND VGND.n7 0.0213333
R17 a_27_297.n2 a_27_297.t2 816.391
R18 a_27_297.n4 a_27_297.n3 264.435
R19 a_27_297.n1 a_27_297.t6 241
R20 a_27_297.n3 a_27_297.n0 198.929
R21 a_27_297.n1 a_27_297.t5 168.701
R22 a_27_297.n2 a_27_297.n1 152
R23 a_27_297.n3 a_27_297.n2 63.5404
R24 a_27_297.t0 a_27_297.n4 47.1434
R25 a_27_297.n4 a_27_297.t1 47.1434
R26 a_27_297.n0 a_27_297.t4 38.5719
R27 a_27_297.n0 a_27_297.t3 38.5719
R28 VNB.t4 VNB.t3 1395.47
R29 VNB.t1 VNB.t0 1366.99
R30 VNB.t2 VNB.t4 1196.12
R31 VNB.t0 VNB.t2 1196.12
R32 VNB VNB.t1 911.327
R33 D.n0 D.t0 186.03
R34 D D.n0 154.012
R35 D.n0 D.t1 137.829
R36 a_205_297.t0 a_205_297.t1 98.5005
R37 a_277_297.t0 a_277_297.t1 154.786
R38 VPB.t1 VPB.t3 290.031
R39 VPB.t2 VPB.t1 284.113
R40 VPB.t0 VPB.t4 284.113
R41 VPB.t4 VPB.t2 213.084
R42 VPB VPB.t0 189.409
R43 A.n0 A.t1 196.549
R44 A A.n0 161.31
R45 A.n0 A.t0 148.35
R46 VPWR VPWR.n0 321.769
R47 VPWR.n0 VPWR.t1 96.1553
R48 VPWR.n0 VPWR.t0 26.5955
R49 X X.t0 360.769
R50 X X.t1 287.072
R51 C.n0 C.t1 196.549
R52 C.n1 C.n0 152
R53 C.n0 C.t0 148.35
R54 C C.n1 5.78114
R55 C.n1 C 3.71663
R56 a_109_297.t0 a_109_297.t1 154.786
C0 VPB D 0.04052f
C1 A X 0.00133f
C2 VPB A 0.032976f
C3 B C 0.091653f
C4 D A 2.13e-19
C5 B X 6.42e-19
C6 VPWR VGND 0.054645f
C7 VPB B 0.106123f
C8 VPWR C 0.007234f
C9 B D 0.002868f
C10 B A 0.063905f
C11 VPWR X 0.087835f
C12 C VGND 0.0191f
C13 VPB VPWR 0.074974f
C14 X VGND 0.035406f
C15 VPB VGND 0.007962f
C16 VPWR D 0.005033f
C17 VPWR A 0.007689f
C18 D VGND 0.051725f
C19 VPB C 0.033818f
C20 A VGND 0.015956f
C21 VPB X 0.010895f
C22 VPWR B 0.19276f
C23 D C 0.095434f
C24 B VGND 0.015869f
C25 C A 0.028036f
C26 VGND VNB 0.366967f
C27 X VNB 0.088347f
C28 A VNB 0.109286f
C29 C VNB 0.104884f
C30 D VNB 0.175262f
C31 B VNB 0.114665f
C32 VPWR VNB 0.289978f
C33 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297.t1 B.t0 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297.t2 D.t0 VGND.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297.t0 B.t1 a_205_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR.t0 A.t0 a_277_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X.t3 a_27_297.t5 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297.t1 C.t0 a_109_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR.t2 a_27_297.t6 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t2 a_27_297.t7 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X.t0 a_27_297.t8 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND.t0 C.t1 a_27_297.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297.t1 D.t1 a_27_297.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND.t5 A.t1 a_27_297.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 B.t1 B.t0 378.255
R1 B B.t1 329.56
R2 VGND.n10 VGND.t4 242.677
R3 VGND.n8 VGND.n2 200.516
R4 VGND.n4 VGND.n3 198.475
R5 VGND.n5 VGND.t2 161.261
R6 VGND.n3 VGND.t5 52.8576
R7 VGND.n2 VGND.t3 38.5719
R8 VGND.n2 VGND.t0 38.5719
R9 VGND.n3 VGND.t1 27.5691
R10 VGND.n9 VGND.n8 22.9652
R11 VGND.n8 VGND.n1 21.4593
R12 VGND.n10 VGND.n9 19.9534
R13 VGND.n4 VGND.n1 16.9417
R14 VGND.n11 VGND.n10 9.3005
R15 VGND.n6 VGND.n1 9.3005
R16 VGND.n8 VGND.n7 9.3005
R17 VGND.n9 VGND.n0 9.3005
R18 VGND.n5 VGND.n4 6.61608
R19 VGND.n6 VGND.n5 0.686761
R20 VGND.n7 VGND.n6 0.120292
R21 VGND.n7 VGND.n0 0.120292
R22 VGND.n11 VGND.n0 0.120292
R23 VGND VGND.n11 0.0213333
R24 a_27_297.n3 a_27_297.t3 816.135
R25 a_27_297.n5 a_27_297.n4 264.435
R26 a_27_297.n1 a_27_297.t6 212.081
R27 a_27_297.n2 a_27_297.t8 212.081
R28 a_27_297.n4 a_27_297.n0 198.929
R29 a_27_297.n3 a_27_297.n2 155.653
R30 a_27_297.n1 a_27_297.t7 139.78
R31 a_27_297.n2 a_27_297.t5 139.78
R32 a_27_297.n4 a_27_297.n3 63.3981
R33 a_27_297.n2 a_27_297.n1 61.346
R34 a_27_297.t0 a_27_297.n5 47.1434
R35 a_27_297.n5 a_27_297.t2 47.1434
R36 a_27_297.n0 a_27_297.t4 38.5719
R37 a_27_297.n0 a_27_297.t1 38.5719
R38 VNB.t3 VNB.t5 1395.47
R39 VNB.t2 VNB.t0 1366.99
R40 VNB.t5 VNB.t4 1196.12
R41 VNB.t1 VNB.t3 1196.12
R42 VNB.t0 VNB.t1 1196.12
R43 VNB VNB.t2 911.327
R44 D.n0 D.t0 186.03
R45 D D.n0 153.983
R46 D.n0 D.t1 137.829
R47 a_205_297.t0 a_205_297.t1 98.5005
R48 a_277_297.t0 a_277_297.t1 154.786
R49 VPB.t5 VPB.t2 290.031
R50 VPB.t1 VPB.t5 284.113
R51 VPB.t0 VPB.t4 284.113
R52 VPB.t2 VPB.t3 248.599
R53 VPB.t4 VPB.t1 213.084
R54 VPB VPB.t0 189.409
R55 A.n0 A.t1 196.549
R56 A A.n0 161.504
R57 A.n0 A.t0 148.35
R58 VPWR.n1 VPWR.n0 320.808
R59 VPWR.n1 VPWR.t2 272.065
R60 VPWR.n0 VPWR.t0 96.1553
R61 VPWR.n0 VPWR.t1 26.5955
R62 VPWR VPWR.n1 0.914166
R63 X X.n0 299.197
R64 X X.n1 261.752
R65 X.n0 X.t1 26.5955
R66 X.n0 X.t0 26.5955
R67 X.n1 X.t2 24.9236
R68 X.n1 X.t3 24.9236
R69 C.n0 C.t1 196.549
R70 C.n1 C.n0 152
R71 C.n0 C.t0 148.35
R72 C C.n1 5.78114
R73 C.n1 C 3.71663
R74 a_109_297.t0 a_109_297.t1 154.786
C0 VPWR D 0.005055f
C1 D VPB 0.040538f
C2 A X 0.001337f
C3 X VPWR 0.173976f
C4 A B 0.063526f
C5 X VPB 0.00408f
C6 VGND C 0.0191f
C7 VPWR B 0.193485f
C8 B VPB 0.107155f
C9 D C 0.095434f
C10 A VPWR 0.00784f
C11 A VPB 0.033504f
C12 VGND D 0.052207f
C13 VPWR VPB 0.089203f
C14 B C 0.091653f
C15 X VGND 0.085613f
C16 VGND B 0.015875f
C17 A C 0.028036f
C18 B D 0.002868f
C19 VPWR C 0.007234f
C20 C VPB 0.033818f
C21 A VGND 0.01624f
C22 A D 2.13e-19
C23 X B 6.52e-19
C24 VGND VPWR 0.076788f
C25 VGND VPB 0.010012f
C26 VGND VNB 0.44429f
C27 X VNB 0.02206f
C28 A VNB 0.108882f
C29 C VNB 0.104884f
C30 D VNB 0.175382f
C31 B VNB 0.11382f
C32 VPWR VNB 0.369371f
C33 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4_4 VNB VPB VPWR VGND D C B A X
X0 VPWR.t4 A.t0 a_304_297.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297.t0 B.t0 a_220_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t6 C.t0 a_32_297.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3 a_220_297.t1 C.t1 a_114_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297.t1 D.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297.t2 B.t1 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 a_32_297.t5 X.t7 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t6 a_32_297.t6 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t7 A.t1 a_32_297.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t2 a_32_297.t7 X.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X.t3 a_32_297.t8 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X.t2 a_32_297.t9 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t4 a_32_297.t10 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297.t0 D.t1 a_32_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND.t2 a_32_297.t11 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t3 a_32_297.t12 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n0 A.t0 241.536
R1 A A.n0 177.601
R2 A.n0 A.t1 169.237
R3 a_304_297.t0 a_304_297.t1 53.1905
R4 VPWR.n2 VPWR.t0 351.567
R5 VPWR.n4 VPWR.n3 318.293
R6 VPWR.n1 VPWR.n0 318.293
R7 VPWR.n0 VPWR.t3 37.4305
R8 VPWR.n0 VPWR.t4 37.4305
R9 VPWR.n5 VPWR.n4 27.8593
R10 VPWR.n3 VPWR.t1 26.5955
R11 VPWR.n3 VPWR.t2 26.5955
R12 VPWR.n5 VPWR.n1 20.7064
R13 VPWR.n6 VPWR.n5 9.3005
R14 VPWR.n7 VPWR.n1 7.42335
R15 VPWR.n4 VPWR.n2 6.55195
R16 VPWR.n6 VPWR.n2 0.662135
R17 VPWR VPWR.n7 0.475961
R18 VPWR.n7 VPWR.n6 0.149912
R19 VPB.t7 VPB.t5 313.707
R20 VPB.t0 VPB.t6 313.707
R21 VPB.t3 VPB.t2 248.599
R22 VPB.t4 VPB.t3 248.599
R23 VPB.t5 VPB.t4 248.599
R24 VPB.t1 VPB.t7 248.599
R25 VPB.t6 VPB.t1 248.599
R26 VPB VPB.t0 210.125
R27 B.n0 B.t0 241.536
R28 B B.n0 183.668
R29 B.n0 B.t1 169.237
R30 a_220_297.t0 a_220_297.t1 53.1905
R31 C.n0 C.t1 241.536
R32 C C.n0 192.671
R33 C.n0 C.t0 169.237
R34 a_32_297.t0 a_32_297.n14 307.396
R35 a_32_297.n4 a_32_297.t5 212.081
R36 a_32_297.n3 a_32_297.t6 212.081
R37 a_32_297.n8 a_32_297.t7 212.081
R38 a_32_297.n10 a_32_297.t10 212.081
R39 a_32_297.n14 a_32_297.n0 197.424
R40 a_32_297.n13 a_32_297.n1 197.424
R41 a_32_297.n6 a_32_297.n5 177.601
R42 a_32_297.n12 a_32_297.n11 152
R43 a_32_297.n9 a_32_297.n2 152
R44 a_32_297.n7 a_32_297.n6 152
R45 a_32_297.n4 a_32_297.t12 139.78
R46 a_32_297.n3 a_32_297.t9 139.78
R47 a_32_297.n8 a_32_297.t11 139.78
R48 a_32_297.n10 a_32_297.t8 139.78
R49 a_32_297.n13 a_32_297.n12 79.0593
R50 a_32_297.n14 a_32_297.n13 65.5064
R51 a_32_297.n11 a_32_297.n9 49.6611
R52 a_32_297.n8 a_32_297.n7 46.7399
R53 a_32_297.n0 a_32_297.t1 39.6928
R54 a_32_297.n5 a_32_297.n3 35.055
R55 a_32_297.n0 a_32_297.t3 30.462
R56 a_32_297.n5 a_32_297.n4 26.2914
R57 a_32_297.n6 a_32_297.n2 25.6005
R58 a_32_297.n12 a_32_297.n2 25.6005
R59 a_32_297.n1 a_32_297.t4 24.9236
R60 a_32_297.n1 a_32_297.t2 24.9236
R61 a_32_297.n7 a_32_297.n3 14.6066
R62 a_32_297.n11 a_32_297.n10 8.76414
R63 a_32_297.n9 a_32_297.n8 2.92171
R64 VGND.n6 VGND.t3 289.649
R65 VGND.n17 VGND.t0 271.12
R66 VGND.n5 VGND.n4 207.965
R67 VGND.n15 VGND.n2 200.516
R68 VGND.n11 VGND.n10 198.475
R69 VGND.n10 VGND.t7 43.3851
R70 VGND.n6 VGND.n5 37.4475
R71 VGND.n9 VGND.n8 34.6358
R72 VGND.n16 VGND.n15 28.6123
R73 VGND.n10 VGND.t4 26.7697
R74 VGND.n11 VGND.n1 26.3534
R75 VGND.n4 VGND.t1 24.9236
R76 VGND.n4 VGND.t2 24.9236
R77 VGND.n2 VGND.t5 24.9236
R78 VGND.n2 VGND.t6 24.9236
R79 VGND.n17 VGND.n16 24.0946
R80 VGND.n15 VGND.n1 15.8123
R81 VGND.n11 VGND.n9 14.3064
R82 VGND.n18 VGND.n17 9.3005
R83 VGND.n8 VGND.n7 9.3005
R84 VGND.n9 VGND.n3 9.3005
R85 VGND.n12 VGND.n11 9.3005
R86 VGND.n13 VGND.n1 9.3005
R87 VGND.n15 VGND.n14 9.3005
R88 VGND.n16 VGND.n0 9.3005
R89 VGND.n8 VGND.n5 2.63579
R90 VGND.n7 VGND.n6 2.35328
R91 VGND.n7 VGND.n3 0.120292
R92 VGND.n12 VGND.n3 0.120292
R93 VGND.n13 VGND.n12 0.120292
R94 VGND.n14 VGND.n13 0.120292
R95 VGND.n14 VGND.n0 0.120292
R96 VGND.n18 VGND.n0 0.120292
R97 VGND VGND.n18 0.0239375
R98 VNB.t7 VNB.t4 1509.39
R99 VNB.t0 VNB.t6 1509.39
R100 VNB.t3 VNB.t1 1196.12
R101 VNB.t2 VNB.t3 1196.12
R102 VNB.t4 VNB.t2 1196.12
R103 VNB.t5 VNB.t7 1196.12
R104 VNB.t6 VNB.t5 1196.12
R105 VNB VNB.t0 1011
R106 a_114_297.t0 a_114_297.t1 74.8605
R107 D.n0 D.t1 231.017
R108 D.n0 D.t0 158.716
R109 D D.n0 155.256
R110 X.n5 X.n3 252.931
R111 X.n2 X.n0 238.163
R112 X.n5 X.n4 208.507
R113 X.n2 X.n1 98.982
R114 X.n6 X.n5 55.9486
R115 X.n3 X.t5 26.5955
R116 X.n3 X.t4 26.5955
R117 X.n4 X.t7 26.5955
R118 X.n4 X.t6 26.5955
R119 X.n0 X.t1 24.9236
R120 X.n0 X.t3 24.9236
R121 X.n1 X.t0 24.9236
R122 X.n1 X.t2 24.9236
R123 X.n6 X.n2 14.2227
R124 X X.n6 2.61274
C0 C VGND 0.016852f
C1 VPB B 0.028231f
C2 C VPWR 0.043951f
C3 VGND X 0.245268f
C4 B A 0.10797f
C5 VPWR X 0.358476f
C6 VPB C 0.029146f
C7 D VGND 0.046879f
C8 D VPWR 0.013631f
C9 VPB X 0.012566f
C10 VGND VPWR 0.083527f
C11 A X 0.015701f
C12 VPB D 0.039214f
C13 VPB VGND 0.006824f
C14 C B 0.162549f
C15 VPB VPWR 0.086383f
C16 VGND A 0.018403f
C17 A VPWR 0.052513f
C18 B X 0.004605f
C19 VPB A 0.030992f
C20 VGND B 0.017696f
C21 B VPWR 0.082692f
C22 D C 0.046429f
C23 VGND VNB 0.509096f
C24 X VNB 0.058359f
C25 VPWR VNB 0.422751f
C26 A VNB 0.091075f
C27 B VNB 0.089178f
C28 C VNB 0.090691f
C29 D VNB 0.157668f
C30 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X.t1 a_215_297.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53.t0 D_N.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297.t3 a_109_53.t2 VGND.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X.t0 a_215_297.t6 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297.t0 C.t0 a_297_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297.t0 B.t0 a_392_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297.t0 B.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR.t2 A.t0 a_465_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297.t1 a_109_53.t3 a_215_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53.t1 D_N.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND.t2 C.t1 a_215_297.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND.t4 A.t1 a_215_297.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 a_215_297.n1 a_215_297.t4 814.366
R1 a_215_297.n3 a_215_297.n2 262.553
R2 a_215_297.n0 a_215_297.t5 241.536
R3 a_215_297.n4 a_215_297.n3 198.929
R4 a_215_297.n0 a_215_297.t6 169.237
R5 a_215_297.n1 a_215_297.n0 152
R6 a_215_297.n3 a_215_297.n1 63.3981
R7 a_215_297.n2 a_215_297.t3 47.1434
R8 a_215_297.n2 a_215_297.t1 40.0005
R9 a_215_297.n4 a_215_297.t2 38.5719
R10 a_215_297.t0 a_215_297.n4 38.5719
R11 VPWR.n1 VPWR.t1 692.894
R12 VPWR.n1 VPWR.n0 321.947
R13 VPWR.n0 VPWR.t2 96.1553
R14 VPWR.n0 VPWR.t0 26.5955
R15 VPWR VPWR.n1 0.0591666
R16 X X.t1 359.536
R17 X X.t0 286.675
R18 VPB.t2 VPB.t5 556.386
R19 VPB.t4 VPB.t0 290.031
R20 VPB.t5 VPB.t3 281.154
R21 VPB.t1 VPB.t4 269.315
R22 VPB.t3 VPB.t1 216.044
R23 VPB VPB.t2 189.409
R24 D_N.n0 D_N.t0 185.168
R25 D_N D_N.n0 154.071
R26 D_N.n0 D_N.t1 136.969
R27 VGND.n8 VGND.t5 242.965
R28 VGND.n10 VGND.t3 242.395
R29 VGND.n5 VGND.n2 203.686
R30 VGND.n4 VGND.n3 200.516
R31 VGND.n2 VGND.t4 52.8576
R32 VGND.n3 VGND.t1 38.5719
R33 VGND.n3 VGND.t2 38.5719
R34 VGND.n2 VGND.t0 27.5691
R35 VGND.n9 VGND.n8 25.977
R36 VGND.n4 VGND.n1 22.5887
R37 VGND.n10 VGND.n9 19.9534
R38 VGND.n8 VGND.n1 18.4476
R39 VGND.n11 VGND.n10 9.3005
R40 VGND.n6 VGND.n1 9.3005
R41 VGND.n8 VGND.n7 9.3005
R42 VGND.n9 VGND.n0 9.3005
R43 VGND.n5 VGND.n4 6.48594
R44 VGND.n6 VGND.n5 0.65716
R45 VGND.n7 VGND.n6 0.120292
R46 VGND.n7 VGND.n0 0.120292
R47 VGND.n11 VGND.n0 0.120292
R48 VGND VGND.n11 0.0213333
R49 a_109_53.n1 a_109_53.t1 669.389
R50 a_109_53.t0 a_109_53.n1 249.434
R51 a_109_53.n0 a_109_53.t2 184.572
R52 a_109_53.n1 a_109_53.n0 169.456
R53 a_109_53.n0 a_109_53.t3 136.373
R54 VNB.t4 VNB.t1 2677.02
R55 VNB.t5 VNB.t0 1395.47
R56 VNB.t1 VNB.t3 1295.79
R57 VNB.t2 VNB.t5 1196.12
R58 VNB.t3 VNB.t2 1196.12
R59 VNB VNB.t4 911.327
R60 C.n0 C.t1 196.549
R61 C.n1 C.n0 152
R62 C.n0 C.t0 148.35
R63 C.n1 C 6.29727
R64 C C.n1 3.2005
R65 a_297_297.t0 a_297_297.t1 152.44
R66 a_392_297.t0 a_392_297.t1 100.846
R67 B.t0 B.t1 382.909
R68 B B.t0 318.317
R69 a_465_297.t0 a_465_297.t1 143.06
R70 A.n0 A.t1 196.549
R71 A A.n0 161.504
R72 A.n0 A.t0 148.35
C0 C VPB 0.033675f
C1 X VPB 0.010957f
C2 B C 0.089339f
C3 VPWR VGND 0.074967f
C4 B X 6.65e-19
C5 D_N VPB 0.046076f
C6 A VPB 0.032495f
C7 VPWR C 0.007534f
C8 VPWR X 0.088522f
C9 B A 0.066627f
C10 C VGND 0.020222f
C11 X VGND 0.035904f
C12 B VPB 0.115837f
C13 VPWR D_N 0.041199f
C14 VPWR A 0.007304f
C15 D_N VGND 0.053053f
C16 A VGND 0.015787f
C17 VPWR VPB 0.122221f
C18 VGND VPB 0.011459f
C19 VPWR B 0.254723f
C20 B VGND 0.016065f
C21 C A 0.028079f
C22 A X 0.001269f
C23 VGND VNB 0.469379f
C24 X VNB 0.088401f
C25 A VNB 0.10846f
C26 C VNB 0.10053f
C27 D_N VNB 0.185426f
C28 B VNB 0.100557f
C29 VPWR VNB 0.398869f
C30 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C D_N X A B
X0 a_176_21.t4 C.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND.t6 D_N.t0 a_27_53.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND.t2 a_176_21.t5 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X.t2 a_176_21.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR.t2 a_176_21.t7 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.16835 pd=1.495 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297.t1 C.t1 a_483_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21.t0 a_27_53.t2 a_555_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X.t0 a_176_21.t8 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1693 ps=1.5 w=1 l=0.15
X8 a_387_297.t1 A.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.16835 ps=1.495 w=0.42 l=0.15
X9 a_483_297.t0 B.t0 a_387_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND.t1 B.t1 a_176_21.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND.t0 a_27_53.t3 a_176_21.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR.t0 D_N.t1 a_27_53.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1693 pd=1.5 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_176_21.t3 A.t1 VGND.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.10025 ps=0.985 w=0.42 l=0.15
R0 C.n0 C.t0 196.549
R1 C C.n0 161.28
R2 C.n0 C.t1 148.35
R3 VGND.n5 VGND.t0 249.263
R4 VGND.n1 VGND.n0 208.719
R5 VGND.n4 VGND.n3 200.516
R6 VGND.n9 VGND.n8 198.475
R7 VGND.n8 VGND.t4 52.8576
R8 VGND.n0 VGND.t6 48.5719
R9 VGND.n3 VGND.t5 38.5719
R10 VGND.n3 VGND.t1 38.5719
R11 VGND.n10 VGND.n1 32.7534
R12 VGND.n0 VGND.t3 31.2372
R13 VGND.n8 VGND.t2 26.9515
R14 VGND.n7 VGND.n4 23.7181
R15 VGND.n10 VGND.n9 21.4593
R16 VGND.n9 VGND.n7 19.2005
R17 VGND.n12 VGND.n1 9.54145
R18 VGND.n11 VGND.n10 9.3005
R19 VGND.n9 VGND.n2 9.3005
R20 VGND.n7 VGND.n6 9.3005
R21 VGND.n5 VGND.n4 6.33263
R22 VGND.n6 VGND.n5 0.754842
R23 VGND.n12 VGND.n11 0.141672
R24 VGND VGND.n12 0.120476
R25 VGND.n6 VGND.n2 0.120292
R26 VGND.n11 VGND.n2 0.120292
R27 a_176_21.t0 a_176_21.n5 811.324
R28 a_176_21.n2 a_176_21.n1 272.719
R29 a_176_21.n4 a_176_21.t7 212.081
R30 a_176_21.n3 a_176_21.t8 212.081
R31 a_176_21.n2 a_176_21.n0 204.953
R32 a_176_21.n5 a_176_21.n4 152
R33 a_176_21.n4 a_176_21.t5 139.78
R34 a_176_21.n3 a_176_21.t6 139.78
R35 a_176_21.n4 a_176_21.n3 61.346
R36 a_176_21.n5 a_176_21.n2 60.868
R37 a_176_21.n0 a_176_21.t2 55.7148
R38 a_176_21.n0 a_176_21.t3 38.5719
R39 a_176_21.n1 a_176_21.t1 38.5719
R40 a_176_21.n1 a_176_21.t4 38.5719
R41 VNB.t4 VNB.t2 1381.23
R42 VNB.t6 VNB.t3 1381.23
R43 VNB.t2 VNB.t1 1366.99
R44 VNB.t5 VNB.t0 1196.12
R45 VNB.t1 VNB.t5 1196.12
R46 VNB.t3 VNB.t4 1196.12
R47 VNB VNB.t6 911.327
R48 D_N.n0 D_N.t0 186.03
R49 D_N D_N.n0 155.911
R50 D_N.n0 D_N.t1 137.829
R51 a_27_53.t0 a_27_53.n0 665.164
R52 a_27_53.n0 a_27_53.t2 516.605
R53 a_27_53.t2 a_27_53.t3 392.027
R54 a_27_53.n0 a_27_53.t1 318.603
R55 X.n2 X.n0 707.843
R56 X.n2 X.n1 185
R57 X.n0 X.t1 26.5955
R58 X.n0 X.t0 26.5955
R59 X.n1 X.t3 24.9236
R60 X.n1 X.t2 24.9236
R61 X X.n2 4.11479
R62 VPWR.n2 VPWR.n0 727.775
R63 VPWR.n2 VPWR.n1 725.153
R64 VPWR.n0 VPWR.t3 96.1553
R65 VPWR.n1 VPWR.t0 96.1553
R66 VPWR.n0 VPWR.t2 27.8072
R67 VPWR.n1 VPWR.t1 27.7095
R68 VPWR VPWR.n2 0.395964
R69 VPB.t4 VPB.t6 287.072
R70 VPB.t2 VPB.t3 287.072
R71 VPB.t5 VPB.t0 284.113
R72 VPB.t6 VPB.t1 284.113
R73 VPB.t3 VPB.t4 248.599
R74 VPB.t1 VPB.t5 213.084
R75 VPB VPB.t2 189.409
R76 a_483_297.t0 a_483_297.t1 98.5005
R77 a_555_297.t0 a_555_297.t1 154.786
R78 A.n0 A.t1 196.549
R79 A A.n0 156.161
R80 A.n0 A.t0 148.35
R81 a_387_297.t0 a_387_297.t1 154.786
R82 B.t0 B.t1 392.027
R83 B B.t0 326.015
C0 C VPWR 0.004715f
C1 A D_N 0.004645f
C2 A VPB 0.033105f
C3 VGND B 0.01488f
C4 VPB B 0.086777f
C5 A C 0.013784f
C6 A VPWR 0.00421f
C7 C B 0.075313f
C8 VGND X 0.088568f
C9 VPWR B 0.081771f
C10 D_N X 0.001639f
C11 VPB X 0.002241f
C12 C X 4.42e-20
C13 A B 0.065423f
C14 VGND D_N 0.015284f
C15 VGND VPB 0.0117f
C16 VPWR X 0.01138f
C17 VPB D_N 0.044834f
C18 C VGND 0.035352f
C19 A X 0.001247f
C20 VGND VPWR 0.073077f
C21 C VPB 0.02921f
C22 VPWR D_N 0.005061f
C23 VPB VPWR 0.096981f
C24 X B 8.59e-19
C25 A VGND 0.016117f
C26 VGND VNB 0.461543f
C27 C VNB 0.110591f
C28 A VNB 0.106422f
C29 B VNB 0.098191f
C30 X VNB 0.008139f
C31 D_N VNB 0.16808f
C32 VPWR VNB 0.370944f
C33 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4b_4 VNB VPB VGND VPWR X D_N C B A
X0 X.t3 a_215_297.t5 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t4 a_215_297.t6 X.t7 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t3 a_215_297.t7 X.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93.t1 D_N.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 a_215_297.t2 a_109_93.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 VGND.t0 C.t0 a_215_297.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6 VGND.t7 A.t0 a_215_297.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X.t1 a_215_297.t8 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297.t4 B.t0 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_93.t0 D_N.t1 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR.t0 A.t1 a_487_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t3 a_215_297.t9 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_487_297.t0 B.t1 a_403_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297.t1 C.t1 a_297_297.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR.t1 a_215_297.t10 X.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X.t5 a_215_297.t11 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X16 X.t4 a_215_297.t12 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_297_297.t1 a_109_93.t3 a_215_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
R0 a_215_297.t1 a_215_297.n14 310.466
R1 a_215_297.n4 a_215_297.t10 212.081
R2 a_215_297.n3 a_215_297.t5 212.081
R3 a_215_297.n8 a_215_297.t7 212.081
R4 a_215_297.n10 a_215_297.t8 212.081
R5 a_215_297.n14 a_215_297.n0 197.424
R6 a_215_297.n13 a_215_297.n1 197.424
R7 a_215_297.n6 a_215_297.n5 177.601
R8 a_215_297.n12 a_215_297.n11 152
R9 a_215_297.n9 a_215_297.n2 152
R10 a_215_297.n7 a_215_297.n6 152
R11 a_215_297.n4 a_215_297.t6 139.78
R12 a_215_297.n3 a_215_297.t12 139.78
R13 a_215_297.n8 a_215_297.t9 139.78
R14 a_215_297.n10 a_215_297.t11 139.78
R15 a_215_297.n13 a_215_297.n12 79.0593
R16 a_215_297.n14 a_215_297.n13 65.5064
R17 a_215_297.n11 a_215_297.n9 49.6611
R18 a_215_297.n8 a_215_297.n7 46.7399
R19 a_215_297.n0 a_215_297.t2 39.6928
R20 a_215_297.n5 a_215_297.n3 35.055
R21 a_215_297.n0 a_215_297.t0 30.462
R22 a_215_297.n5 a_215_297.n4 26.2914
R23 a_215_297.n6 a_215_297.n2 25.6005
R24 a_215_297.n12 a_215_297.n2 25.6005
R25 a_215_297.n1 a_215_297.t3 24.9236
R26 a_215_297.n1 a_215_297.t4 24.9236
R27 a_215_297.n7 a_215_297.n3 14.6066
R28 a_215_297.n11 a_215_297.n10 8.76414
R29 a_215_297.n9 a_215_297.n8 2.92171
R30 VPWR.n18 VPWR.t5 667.521
R31 VPWR.n7 VPWR.t1 351.546
R32 VPWR.n10 VPWR.n4 318.293
R33 VPWR.n6 VPWR.n5 318.293
R34 VPWR.n4 VPWR.t2 37.4305
R35 VPWR.n4 VPWR.t0 37.4305
R36 VPWR.n12 VPWR.n11 34.6358
R37 VPWR.n12 VPWR.n1 34.6358
R38 VPWR.n16 VPWR.n1 34.6358
R39 VPWR.n17 VPWR.n16 34.6358
R40 VPWR.n11 VPWR.n10 29.3652
R41 VPWR.n9 VPWR.n6 27.4829
R42 VPWR.n5 VPWR.t4 26.5955
R43 VPWR.n5 VPWR.t3 26.5955
R44 VPWR.n18 VPWR.n17 24.4711
R45 VPWR.n10 VPWR.n9 21.0829
R46 VPWR.n9 VPWR.n8 9.3005
R47 VPWR.n10 VPWR.n3 9.3005
R48 VPWR.n11 VPWR.n2 9.3005
R49 VPWR.n13 VPWR.n12 9.3005
R50 VPWR.n14 VPWR.n1 9.3005
R51 VPWR.n16 VPWR.n15 9.3005
R52 VPWR.n17 VPWR.n0 9.3005
R53 VPWR.n19 VPWR.n18 9.3005
R54 VPWR.n7 VPWR.n6 6.57198
R55 VPWR.n8 VPWR.n7 0.662015
R56 VPWR.n8 VPWR.n3 0.120292
R57 VPWR.n3 VPWR.n2 0.120292
R58 VPWR.n13 VPWR.n2 0.120292
R59 VPWR.n14 VPWR.n13 0.120292
R60 VPWR.n15 VPWR.n14 0.120292
R61 VPWR.n15 VPWR.n0 0.120292
R62 VPWR.n19 VPWR.n0 0.120292
R63 VPWR VPWR.n19 0.0226354
R64 X.n5 X.n3 252.931
R65 X.n2 X.n0 238.163
R66 X.n5 X.n4 208.507
R67 X.n2 X.n1 98.982
R68 X.n6 X.n5 56.7378
R69 X.n3 X.t2 26.5955
R70 X.n3 X.t1 26.5955
R71 X.n4 X.t0 26.5955
R72 X.n4 X.t3 26.5955
R73 X.n0 X.t6 24.9236
R74 X.n0 X.t5 24.9236
R75 X.n1 X.t7 24.9236
R76 X.n1 X.t4 24.9236
R77 X.n6 X.n2 14.2227
R78 X X.n6 2.66717
R79 VPB.t8 VPB.t1 556.386
R80 VPB.t2 VPB.t4 313.707
R81 VPB.t1 VPB.t7 313.707
R82 VPB.t6 VPB.t3 248.599
R83 VPB.t5 VPB.t6 248.599
R84 VPB.t4 VPB.t5 248.599
R85 VPB.t0 VPB.t2 248.599
R86 VPB.t7 VPB.t0 248.599
R87 VPB VPB.t8 192.369
R88 VGND.n5 VGND.t4 289.776
R89 VGND.n21 VGND.t6 256.065
R90 VGND.n19 VGND.t5 231.744
R91 VGND.n7 VGND.n6 207.965
R92 VGND.n15 VGND.n14 200.516
R93 VGND.n12 VGND.n4 198.475
R94 VGND.n4 VGND.t7 43.3851
R95 VGND.n7 VGND.n5 37.7583
R96 VGND.n8 VGND.n3 34.6358
R97 VGND.n15 VGND.n1 28.2358
R98 VGND.n4 VGND.t2 26.7697
R99 VGND.n13 VGND.n12 25.977
R100 VGND.n20 VGND.n19 25.977
R101 VGND.n21 VGND.n20 25.977
R102 VGND.n6 VGND.t1 24.9236
R103 VGND.n6 VGND.t3 24.9236
R104 VGND.n14 VGND.t8 24.9236
R105 VGND.n14 VGND.t0 24.9236
R106 VGND.n19 VGND.n1 24.4711
R107 VGND.n15 VGND.n13 16.1887
R108 VGND.n12 VGND.n3 14.6829
R109 VGND.n22 VGND.n21 9.3005
R110 VGND.n9 VGND.n8 9.3005
R111 VGND.n10 VGND.n3 9.3005
R112 VGND.n12 VGND.n11 9.3005
R113 VGND.n13 VGND.n2 9.3005
R114 VGND.n16 VGND.n15 9.3005
R115 VGND.n17 VGND.n1 9.3005
R116 VGND.n19 VGND.n18 9.3005
R117 VGND.n20 VGND.n0 9.3005
R118 VGND.n9 VGND.n5 2.4189
R119 VGND.n8 VGND.n7 2.25932
R120 VGND.n10 VGND.n9 0.120292
R121 VGND.n11 VGND.n10 0.120292
R122 VGND.n11 VGND.n2 0.120292
R123 VGND.n16 VGND.n2 0.120292
R124 VGND.n17 VGND.n16 0.120292
R125 VGND.n18 VGND.n17 0.120292
R126 VGND.n18 VGND.n0 0.120292
R127 VGND.n22 VGND.n0 0.120292
R128 VGND VGND.n22 0.0226354
R129 VNB.t6 VNB.t5 2677.02
R130 VNB.t7 VNB.t2 1509.39
R131 VNB.t5 VNB.t0 1509.39
R132 VNB.t1 VNB.t4 1196.12
R133 VNB.t3 VNB.t1 1196.12
R134 VNB.t2 VNB.t3 1196.12
R135 VNB.t8 VNB.t7 1196.12
R136 VNB.t0 VNB.t8 1196.12
R137 VNB VNB.t6 925.567
R138 D_N.n0 D_N.t1 328.659
R139 D_N D_N.n0 154.868
R140 D_N.n0 D_N.t0 126.219
R141 a_109_93.t0 a_109_93.n1 718.187
R142 a_109_93.n1 a_109_93.t1 242.817
R143 a_109_93.n0 a_109_93.t3 228.311
R144 a_109_93.n1 a_109_93.n0 168.679
R145 a_109_93.n0 a_109_93.t2 156.012
R146 C.n0 C.t1 241.536
R147 C C.n0 192.502
R148 C.n0 C.t0 169.237
R149 A.n0 A.t1 241.536
R150 A A.n0 178.353
R151 A.n0 A.t0 169.237
R152 B.n0 B.t1 241.536
R153 B B.n0 185.817
R154 B.n0 B.t0 169.237
R155 a_487_297.t0 a_487_297.t1 53.1905
R156 a_403_297.t0 a_403_297.t1 53.1905
R157 a_297_297.t0 a_297_297.t1 74.8605
C0 D_N A 7.84e-20
C1 C B 0.161257f
C2 B VPWR 0.081928f
C3 D_N VGND 0.042627f
C4 VPWR X 0.357977f
C5 VPB B 0.028227f
C6 VPB X 0.012723f
C7 D_N B 3.04e-19
C8 C VPWR 0.045204f
C9 D_N X 3.65e-19
C10 A VGND 0.018403f
C11 VPB C 0.029208f
C12 VPB VPWR 0.116786f
C13 D_N C 6.87e-19
C14 D_N VPWR 0.048585f
C15 B A 0.10797f
C16 B VGND 0.017742f
C17 A X 0.015701f
C18 X VGND 0.245005f
C19 VPB D_N 0.107071f
C20 A VPWR 0.052581f
C21 B X 0.004605f
C22 C VGND 0.017002f
C23 VPWR VGND 0.10333f
C24 VPB A 0.030992f
C25 VPB VGND 0.010541f
C26 VGND VNB 0.630714f
C27 X VNB 0.058124f
C28 VPWR VNB 0.514749f
C29 A VNB 0.091075f
C30 B VNB 0.089178f
C31 C VNB 0.09076f
C32 D_N VNB 0.185891f
C33 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4bb_1 VPWR VGND VPB VNB B A X D_N C_N
X0 VGND.t4 A.t0 a_311_413.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR.t3 A.t1 a_561_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
X2 a_393_413.t1 a_205_93.t2 a_311_413.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND.t2 C_N.t0 a_27_410.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR.t1 C_N.t1 a_27_410.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X.t0 a_311_413.t5 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X6 VGND.t0 a_27_410.t2 a_311_413.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05985 ps=0.705 w=0.42 l=0.15
X7 a_561_297.t0 B.t0 a_489_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93.t1 D_N.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X9 a_205_93.t0 D_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X10 a_489_297.t1 a_27_410.t3 a_393_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X11 a_311_413.t2 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413.t4 a_205_93.t3 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 X.t1 a_311_413.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
R0 A.n0 A.t0 206.19
R1 A A.n0 161.504
R2 A.n0 A.t1 148.35
R3 a_311_413.n2 a_311_413.t1 835.578
R4 a_311_413.n4 a_311_413.n3 263.307
R5 a_311_413.n1 a_311_413.t5 241.536
R6 a_311_413.n3 a_311_413.n0 198.929
R7 a_311_413.n1 a_311_413.t6 169.237
R8 a_311_413.n2 a_311_413.n1 152
R9 a_311_413.n3 a_311_413.n2 63.3981
R10 a_311_413.t0 a_311_413.n4 42.8576
R11 a_311_413.n0 a_311_413.t3 38.5719
R12 a_311_413.n0 a_311_413.t2 38.5719
R13 a_311_413.n4 a_311_413.t4 38.5719
R14 VGND.n9 VGND.t6 237.226
R15 VGND.n1 VGND.n0 228.294
R16 VGND.n6 VGND.n5 203.686
R17 VGND.n4 VGND.n3 200.516
R18 VGND.n5 VGND.t4 52.8576
R19 VGND.n0 VGND.t2 45.7148
R20 VGND.n3 VGND.t1 38.5719
R21 VGND.n3 VGND.t0 38.5719
R22 VGND.n0 VGND.t5 38.5719
R23 VGND.n10 VGND.n1 30.8711
R24 VGND.n5 VGND.t3 30.6379
R25 VGND.n10 VGND.n9 24.0946
R26 VGND.n8 VGND.n4 22.5887
R27 VGND.n9 VGND.n8 16.9417
R28 VGND.n12 VGND.n1 11.4238
R29 VGND.n8 VGND.n7 9.3005
R30 VGND.n9 VGND.n2 9.3005
R31 VGND.n11 VGND.n10 9.3005
R32 VGND.n6 VGND.n4 6.48594
R33 VGND.n7 VGND.n6 0.65716
R34 VGND.n12 VGND.n11 0.141672
R35 VGND VGND.n12 0.121778
R36 VGND.n7 VGND.n2 0.120292
R37 VGND.n11 VGND.n2 0.120292
R38 VNB.t5 VNB.t6 2677.02
R39 VNB.t4 VNB.t3 1395.47
R40 VNB.t2 VNB.t5 1267.31
R41 VNB.t6 VNB.t0 1238.83
R42 VNB.t1 VNB.t4 1196.12
R43 VNB.t0 VNB.t1 1196.12
R44 VNB VNB.t2 1025.24
R45 a_561_297.t0 a_561_297.t1 133.679
R46 VPWR.n2 VPWR.n1 607.428
R47 VPWR.n1 VPWR.t0 327.592
R48 VPWR.n2 VPWR.n0 321.981
R49 VPWR.n0 VPWR.t3 96.1553
R50 VPWR.n1 VPWR.t1 63.3219
R51 VPWR.n0 VPWR.t2 26.5955
R52 VPWR VPWR.n2 0.14839
R53 VPB.t0 VPB.t2 553.428
R54 VPB.t6 VPB.t5 290.031
R55 VPB.t3 VPB.t0 287.072
R56 VPB.t2 VPB.t1 284.113
R57 VPB.t4 VPB.t6 257.478
R58 VPB.t1 VPB.t4 213.084
R59 VPB VPB.t3 192.369
R60 a_205_93.t0 a_205_93.n1 696.434
R61 a_205_93.n0 a_205_93.t2 322.747
R62 a_205_93.n1 a_205_93.t1 269.803
R63 a_205_93.n0 a_205_93.t3 194.213
R64 a_205_93.n1 a_205_93.n0 152
R65 a_393_413.t0 a_393_413.t1 499.582
R66 C_N.n0 C_N.t1 329.902
R67 C_N C_N.n0 153.738
R68 C_N.n0 C_N.t0 132.282
R69 a_27_410.t0 a_27_410.n1 665.061
R70 a_27_410.n1 a_27_410.n0 340.236
R71 a_27_410.n1 a_27_410.t1 312.767
R72 a_27_410.n0 a_27_410.t2 206.19
R73 a_27_410.n0 a_27_410.t3 148.35
R74 X X.t0 359.536
R75 X X.t1 286.675
R76 B.t0 B.t1 397.286
R77 B B.t0 338.192
R78 a_489_297.t0 a_489_297.t1 98.5005
R79 D_N D_N.n0 154.429
R80 D_N.n0 D_N.t1 142.994
R81 D_N.n0 D_N.t0 126.927
C0 C_N VGND 0.031122f
C1 VPB VPWR 0.113906f
C2 A VGND 0.018081f
C3 VPB X 0.010957f
C4 VPWR D_N 0.00402f
C5 D_N X 1.35e-20
C6 VPB VGND 0.012362f
C7 VPB C_N 0.088545f
C8 D_N VGND 0.018273f
C9 C_N D_N 0.081313f
C10 VPWR B 0.107056f
C11 VPB A 0.032658f
C12 B X 7.74e-19
C13 B VGND 0.015175f
C14 VPB D_N 0.037415f
C15 VPWR X 0.088522f
C16 B A 0.082255f
C17 VPWR VGND 0.08158f
C18 C_N VPWR 0.021037f
C19 VPB B 0.094576f
C20 X VGND 0.035904f
C21 VPWR A 0.008054f
C22 A X 0.001365f
C23 VGND VNB 0.518562f
C24 X VNB 0.088401f
C25 A VNB 0.111872f
C26 D_N VNB 0.100883f
C27 B VNB 0.101167f
C28 VPWR VNB 0.406703f
C29 C_N VNB 0.132375f
C30 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4bb_2 VPWR VGND VPB VNB B A C_N D_N X
X0 a_398_413.t0 a_206_93.t2 a_316_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR.t1 a_316_413.t5 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X2 X.t3 a_316_413.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 X.t0 a_316_413.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X4 VGND.t5 C_N.t0 a_27_410.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR.t2 C_N.t1 a_27_410.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND.t4 a_27_410.t2 a_316_413.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X7 VGND.t3 A.t0 a_316_413.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND.t0 a_316_413.t8 X.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_566_297.t0 B.t0 a_494_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_206_93.t1 D_N.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X11 a_316_413.t4 B.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_206_93.t0 D_N.t1 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X13 a_494_297.t1 a_27_410.t3 a_398_413.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X14 a_316_413.t1 a_206_93.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VPWR.t4 A.t1 a_566_297.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
R0 a_206_93.t0 a_206_93.n1 697.085
R1 a_206_93.n0 a_206_93.t2 322.747
R2 a_206_93.n1 a_206_93.t1 270.313
R3 a_206_93.n0 a_206_93.t3 194.213
R4 a_206_93.n1 a_206_93.n0 157.272
R5 a_316_413.t0 a_316_413.n5 835.578
R6 a_316_413.n2 a_316_413.n1 264.435
R7 a_316_413.n3 a_316_413.t5 212.081
R8 a_316_413.n4 a_316_413.t7 212.081
R9 a_316_413.n2 a_316_413.n0 198.929
R10 a_316_413.n5 a_316_413.n4 155.653
R11 a_316_413.n3 a_316_413.t8 139.78
R12 a_316_413.n4 a_316_413.t6 139.78
R13 a_316_413.n5 a_316_413.n2 63.3981
R14 a_316_413.n4 a_316_413.n3 61.346
R15 a_316_413.n1 a_316_413.t3 47.1434
R16 a_316_413.n1 a_316_413.t1 40.0005
R17 a_316_413.n0 a_316_413.t2 38.5719
R18 a_316_413.n0 a_316_413.t4 38.5719
R19 a_398_413.t0 a_398_413.t1 499.582
R20 VPB.t6 VPB.t2 568.225
R21 VPB.t7 VPB.t0 290.031
R22 VPB.t4 VPB.t6 287.072
R23 VPB.t2 VPB.t3 284.113
R24 VPB.t5 VPB.t7 257.478
R25 VPB.t0 VPB.t1 248.599
R26 VPB.t3 VPB.t5 213.084
R27 VPB VPB.t4 189.409
R28 X X.n0 299.197
R29 X X.n1 261.752
R30 X.n0 X.t1 26.5955
R31 X.n0 X.t0 26.5955
R32 X.n1 X.t2 24.9236
R33 X.n1 X.t3 24.9236
R34 VPWR.n14 VPWR.n1 601.679
R35 VPWR.n1 VPWR.t3 327.592
R36 VPWR.n6 VPWR.n4 315.406
R37 VPWR.n5 VPWR.t1 271.224
R38 VPWR.n4 VPWR.t4 96.1553
R39 VPWR.n1 VPWR.t2 63.3219
R40 VPWR.n8 VPWR.n7 34.6358
R41 VPWR.n8 VPWR.n2 34.6358
R42 VPWR.n12 VPWR.n2 34.6358
R43 VPWR.n13 VPWR.n12 34.6358
R44 VPWR.n4 VPWR.t0 26.5955
R45 VPWR.n7 VPWR.n6 24.4711
R46 VPWR.n14 VPWR.n13 22.9652
R47 VPWR.n7 VPWR.n3 9.3005
R48 VPWR.n9 VPWR.n8 9.3005
R49 VPWR.n10 VPWR.n2 9.3005
R50 VPWR.n12 VPWR.n11 9.3005
R51 VPWR.n13 VPWR.n0 9.3005
R52 VPWR.n15 VPWR.n14 7.12063
R53 VPWR.n6 VPWR.n5 6.67589
R54 VPWR.n5 VPWR.n3 0.626956
R55 VPWR.n15 VPWR.n0 0.148519
R56 VPWR.n9 VPWR.n3 0.120292
R57 VPWR.n10 VPWR.n9 0.120292
R58 VPWR.n11 VPWR.n10 0.120292
R59 VPWR.n11 VPWR.n0 0.120292
R60 VPWR VPWR.n15 0.11354
R61 VGND.n13 VGND.t2 237.994
R62 VGND.n1 VGND.n0 228.294
R63 VGND.n4 VGND.n3 200.516
R64 VGND.n7 VGND.n6 198.475
R65 VGND.n5 VGND.t0 166.154
R66 VGND.n6 VGND.t3 52.8576
R67 VGND.n0 VGND.t5 45.7148
R68 VGND.n3 VGND.t7 38.5719
R69 VGND.n3 VGND.t4 38.5719
R70 VGND.n0 VGND.t6 38.5719
R71 VGND.n6 VGND.t1 30.6379
R72 VGND.n14 VGND.n1 30.4946
R73 VGND.n14 VGND.n13 25.977
R74 VGND.n12 VGND.n4 24.4711
R75 VGND.n8 VGND.n4 19.9534
R76 VGND.n8 VGND.n7 18.4476
R77 VGND.n13 VGND.n12 16.5652
R78 VGND.n16 VGND.n1 11.8003
R79 VGND.n9 VGND.n8 9.3005
R80 VGND.n10 VGND.n4 9.3005
R81 VGND.n12 VGND.n11 9.3005
R82 VGND.n13 VGND.n2 9.3005
R83 VGND.n15 VGND.n14 9.3005
R84 VGND.n7 VGND.n5 6.57533
R85 VGND.n9 VGND.n5 0.646345
R86 VGND.n16 VGND.n15 0.141672
R87 VGND VGND.n16 0.120476
R88 VGND.n10 VGND.n9 0.120292
R89 VGND.n11 VGND.n10 0.120292
R90 VGND.n11 VGND.n2 0.120292
R91 VGND.n15 VGND.n2 0.120292
R92 VNB.t6 VNB.t2 2677.02
R93 VNB.t3 VNB.t1 1395.47
R94 VNB.t2 VNB.t4 1295.79
R95 VNB.t5 VNB.t6 1267.31
R96 VNB.t1 VNB.t0 1196.12
R97 VNB.t7 VNB.t3 1196.12
R98 VNB.t4 VNB.t7 1196.12
R99 VNB VNB.t5 1025.24
R100 C_N.n0 C_N.t1 329.902
R101 C_N C_N.n0 153.738
R102 C_N.n0 C_N.t0 132.282
R103 a_27_410.n1 a_27_410.t1 665.061
R104 a_27_410.n1 a_27_410.n0 342.118
R105 a_27_410.t0 a_27_410.n1 310.425
R106 a_27_410.n0 a_27_410.t2 206.19
R107 a_27_410.n0 a_27_410.t3 148.35
R108 A.n0 A.t0 206.19
R109 A A.n0 161.504
R110 A.n0 A.t1 148.35
R111 B.t0 B.t1 397.286
R112 B B.t0 338.192
R113 a_494_297.t0 a_494_297.t1 98.5005
R114 a_566_297.t0 a_566_297.t1 133.679
R115 D_N D_N.n0 154.429
R116 D_N.n0 D_N.t1 142.994
R117 D_N.n0 D_N.t0 126.927
C0 X VGND 0.087597f
C1 D_N VPB 0.037591f
C2 A B 0.082255f
C3 VGND C_N 0.031143f
C4 X VPWR 0.17521f
C5 C_N VPWR 0.021141f
C6 VPB B 0.095698f
C7 A VGND 0.018314f
C8 A VPWR 0.008186f
C9 VGND VPB 0.014432f
C10 VPB VPWR 0.128592f
C11 A X 0.001365f
C12 D_N VGND 0.018248f
C13 D_N VPWR 0.004034f
C14 X VPB 0.003896f
C15 VGND B 0.015175f
C16 VPB C_N 0.088703f
C17 VPWR B 0.107293f
C18 D_N X 1.34e-20
C19 D_N C_N 0.081397f
C20 A VPB 0.033153f
C21 X B 7.74e-19
C22 VGND VPWR 0.103917f
C23 VGND VNB 0.596898f
C24 X VNB 0.020672f
C25 A VNB 0.111376f
C26 D_N VNB 0.101197f
C27 B VNB 0.100059f
C28 VPWR VNB 0.486471f
C29 C_N VNB 0.132365f
C30 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_2 VPB VNB VGND VPWR A Y C_N B
X0 a_281_297.t2 B.t0 a_27_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t3 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t2 A.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t5 a_531_21.t2 Y.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t0 C_N.t0 a_531_21.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t4 A.t1 Y.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t7 A.t2 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND.t1 B.t2 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t1 A.t3 a_27_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297.t3 a_531_21.t3 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y.t1 a_531_21.t4 a_281_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND.t3 C_N.t1 a_531_21.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_27_297.t0 B.t3 a_281_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y.t0 a_531_21.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t0 212.081
R2 B B.n2 152.469
R3 B.n0 B.t2 139.78
R4 B.n1 B.t1 139.78
R5 B.n2 B.n0 32.8641
R6 B.n2 B.n1 28.4823
R7 a_27_297.t0 a_27_297.n1 371.904
R8 a_27_297.n1 a_27_297.t3 276.781
R9 a_27_297.n1 a_27_297.n0 208.507
R10 a_27_297.n0 a_27_297.t1 26.5955
R11 a_27_297.n0 a_27_297.t2 26.5955
R12 a_281_297.n1 a_281_297.n0 354.344
R13 a_281_297.n0 a_281_297.t3 279.796
R14 a_281_297.n0 a_281_297.t0 234.12
R15 a_281_297.n1 a_281_297.t1 26.5955
R16 a_281_297.t2 a_281_297.n1 26.5955
R17 VPB.t5 VPB.t3 580.062
R18 VPB.t1 VPB.t0 580.062
R19 VPB.t0 VPB.t5 248.599
R20 VPB.t2 VPB.t1 248.599
R21 VPB.t4 VPB.t2 248.599
R22 VPB.t6 VPB.t4 248.599
R23 VPB VPB.t6 201.246
R24 VGND.n10 VGND.t1 263.462
R25 VGND.n9 VGND.t0 263.462
R26 VGND.n5 VGND.t3 259.594
R27 VGND.n16 VGND.n1 207.965
R28 VGND.n4 VGND.t5 158.379
R29 VGND.n18 VGND.t6 150.922
R30 VGND.n15 VGND.n2 34.6358
R31 VGND.n17 VGND.n16 32.377
R32 VGND.n8 VGND.n7 30.4887
R33 VGND.n1 VGND.t2 24.9236
R34 VGND.n1 VGND.t4 24.9236
R35 VGND.n18 VGND.n17 24.4711
R36 VGND.n10 VGND.n2 21.6534
R37 VGND.n7 VGND.n4 21.4593
R38 VGND.n19 VGND.n18 9.3005
R39 VGND.n7 VGND.n6 9.3005
R40 VGND.n8 VGND.n3 9.3005
R41 VGND.n12 VGND.n11 9.3005
R42 VGND.n13 VGND.n2 9.3005
R43 VGND.n15 VGND.n14 9.3005
R44 VGND.n17 VGND.n0 9.3005
R45 VGND.n11 VGND.n9 9.0005
R46 VGND.n5 VGND.n4 7.11519
R47 VGND.n16 VGND.n15 2.25932
R48 VGND.n11 VGND.n10 2.2005
R49 VGND.n6 VGND.n5 0.542305
R50 VGND.n9 VGND.n8 0.2005
R51 VGND.n6 VGND.n3 0.120292
R52 VGND.n12 VGND.n3 0.120292
R53 VGND.n13 VGND.n12 0.120292
R54 VGND.n14 VGND.n13 0.120292
R55 VGND.n14 VGND.n0 0.120292
R56 VGND.n19 VGND.n0 0.120292
R57 VGND VGND.n19 0.0213333
R58 Y.n4 Y.n3 336.889
R59 Y Y.n6 186.358
R60 Y.n6 Y.n5 185
R61 Y.n2 Y.n0 135.249
R62 Y.n2 Y.n1 98.982
R63 Y.n4 Y.n2 76.0894
R64 Y.n3 Y.t4 26.5955
R65 Y.n3 Y.t1 26.5955
R66 Y.n6 Y.t6 24.9236
R67 Y.n6 Y.t0 24.9236
R68 Y.n0 Y.t5 24.9236
R69 Y.n0 Y.t7 24.9236
R70 Y.n1 Y.t2 24.9236
R71 Y.n1 Y.t3 24.9236
R72 Y Y.n5 11.8308
R73 Y.n5 Y.n4 3.29747
R74 VNB.t5 VNB.t3 2790.94
R75 VNB.t1 VNB.t0 2790.94
R76 VNB.t0 VNB.t5 1196.12
R77 VNB.t2 VNB.t1 1196.12
R78 VNB.t4 VNB.t2 1196.12
R79 VNB.t6 VNB.t4 1196.12
R80 VNB VNB.t6 968.285
R81 A.n0 A.t0 212.081
R82 A.n1 A.t3 212.081
R83 A A.n2 152.823
R84 A.n0 A.t1 139.78
R85 A.n1 A.t2 139.78
R86 A.n2 A.n0 38.7066
R87 A.n2 A.n1 22.6399
R88 VPWR.n1 VPWR.t0 708.317
R89 VPWR.n1 VPWR.n0 324.24
R90 VPWR.n0 VPWR.t2 26.5955
R91 VPWR.n0 VPWR.t1 26.5955
R92 VPWR VPWR.n1 0.148626
R93 a_531_21.t0 a_531_21.n2 670.135
R94 a_531_21.n2 a_531_21.t1 245.206
R95 a_531_21.n1 a_531_21.t3 212.081
R96 a_531_21.n0 a_531_21.t4 212.081
R97 a_531_21.n2 a_531_21.n1 211.373
R98 a_531_21.n1 a_531_21.t2 139.78
R99 a_531_21.n0 a_531_21.t5 139.78
R100 a_531_21.n1 a_531_21.n0 61.346
R101 C_N C_N.n0 157.487
R102 C_N.n0 C_N.t0 147.814
R103 C_N.n0 C_N.t1 131.748
C0 VPB Y 0.00635f
C1 VGND A 0.058456f
C2 A B 0.069132f
C3 VPWR Y 0.011678f
C4 VPB VPWR 0.127595f
C5 VGND Y 0.465329f
C6 VGND VPB 0.013036f
C7 B Y 0.173598f
C8 VPB B 0.06329f
C9 VGND VPWR 0.091025f
C10 C_N Y 5.12e-19
C11 C_N VPB 0.042561f
C12 A Y 0.061756f
C13 B VPWR 0.023905f
C14 VPB A 0.056279f
C15 VGND B 0.032508f
C16 C_N VPWR 0.034098f
C17 C_N VGND 0.041388f
C18 A VPWR 0.043783f
C19 VGND VNB 0.602664f
C20 C_N VNB 0.138101f
C21 Y VNB 0.023739f
C22 VPWR VNB 0.476696f
C23 B VNB 0.188946f
C24 A VNB 0.207619f
C25 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_4 VPB VNB VGND VPWR A C_N B Y
X0 Y.t15 B.t0 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR.t4 A.t0 a_197_297.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t0 a_27_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t4 A.t1 Y.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_555_297.t3 a_27_47.t3 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_197_297.t2 A.t2 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t2 a_27_47.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_197_297.t7 B.t1 a_555_297.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND.t3 a_27_47.t5 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t11 B.t2 Y.t14 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t7 A.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t0 C_N.t0 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 Y.t8 A.t4 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t4 a_27_47.t6 a_555_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t5 a_27_47.t7 a_555_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t0 C_N.t1 a_27_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X16 a_555_297.t0 a_27_47.t8 Y.t10 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t7 A.t5 Y.t9 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_555_297.t6 B.t3 a_197_297.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_197_297.t6 B.t4 a_555_297.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t10 B.t5 Y.t13 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_555_297.t4 B.t6 a_197_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t2 A.t6 a_197_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 a_197_297.t0 A.t7 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y.t12 B.t7 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X25 Y.t11 a_27_47.t9 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t4 212.081
R2 B.n3 B.t6 212.081
R3 B.n4 B.t1 212.081
R4 B B.n5 163.582
R5 B.n0 B.t2 139.78
R6 B.n1 B.t0 139.78
R7 B.n3 B.t5 139.78
R8 B.n4 B.t7 139.78
R9 B B.n2 79.2697
R10 B.n1 B.n0 61.346
R11 B.n5 B.n3 48.2005
R12 B.n2 B.n1 33.1364
R13 B.n3 B.n2 21.6238
R14 B.n5 B.n4 13.146
R15 VGND.n13 VGND.t3 294.144
R16 VGND.n12 VGND.n11 207.965
R17 VGND.n17 VGND.n9 207.965
R18 VGND.n7 VGND.n6 207.965
R19 VGND.n32 VGND.n3 207.965
R20 VGND.n1 VGND.n0 207.965
R21 VGND.n24 VGND.n4 185
R22 VGND.n26 VGND.n25 185
R23 VGND.n25 VGND.n24 96.0005
R24 VGND.n16 VGND.n10 34.6358
R25 VGND.n19 VGND.n18 34.6358
R26 VGND.n23 VGND.n22 34.6358
R27 VGND.n31 VGND.n30 34.6358
R28 VGND.n33 VGND.n1 33.8829
R29 VGND.n13 VGND.n12 31.1922
R30 VGND.n33 VGND.n32 29.3652
R31 VGND.n25 VGND.t9 24.9236
R32 VGND.n24 VGND.t7 24.9236
R33 VGND.n11 VGND.t8 24.9236
R34 VGND.n11 VGND.t2 24.9236
R35 VGND.n9 VGND.t1 24.9236
R36 VGND.n9 VGND.t11 24.9236
R37 VGND.n6 VGND.t12 24.9236
R38 VGND.n6 VGND.t10 24.9236
R39 VGND.n3 VGND.t6 24.9236
R40 VGND.n3 VGND.t4 24.9236
R41 VGND.n0 VGND.t5 24.9236
R42 VGND.n0 VGND.t0 24.9236
R43 VGND.n22 VGND.n7 21.8358
R44 VGND.n17 VGND.n16 18.824
R45 VGND.n30 VGND.n4 18.6417
R46 VGND.n18 VGND.n17 15.8123
R47 VGND.n19 VGND.n7 12.8005
R48 VGND.n12 VGND.n10 9.78874
R49 VGND.n34 VGND.n33 9.3005
R50 VGND.n31 VGND.n2 9.3005
R51 VGND.n30 VGND.n29 9.3005
R52 VGND.n28 VGND.n27 9.3005
R53 VGND.n14 VGND.n10 9.3005
R54 VGND.n16 VGND.n15 9.3005
R55 VGND.n18 VGND.n8 9.3005
R56 VGND.n20 VGND.n19 9.3005
R57 VGND.n22 VGND.n21 9.3005
R58 VGND.n23 VGND.n5 9.3005
R59 VGND.n35 VGND.n1 8.41204
R60 VGND.n27 VGND.n26 7.4005
R61 VGND.n32 VGND.n31 5.27109
R62 VGND.n27 VGND.n4 3.0005
R63 VGND.n26 VGND.n23 2.07697
R64 VGND.n14 VGND.n13 1.40484
R65 VGND.n35 VGND.n34 0.141672
R66 VGND VGND.n35 0.120476
R67 VGND.n15 VGND.n14 0.120292
R68 VGND.n15 VGND.n8 0.120292
R69 VGND.n20 VGND.n8 0.120292
R70 VGND.n21 VGND.n20 0.120292
R71 VGND.n21 VGND.n5 0.120292
R72 VGND.n28 VGND.n5 0.120292
R73 VGND.n29 VGND.n28 0.120292
R74 VGND.n29 VGND.n2 0.120292
R75 VGND.n34 VGND.n2 0.120292
R76 Y.n2 Y.n0 345.31
R77 Y.n2 Y.n1 300.885
R78 Y.n5 Y.n3 135.249
R79 Y.n5 Y.n4 98.982
R80 Y.n7 Y.n6 98.982
R81 Y.n9 Y.n8 98.982
R82 Y.n11 Y.n10 98.982
R83 Y.n13 Y.n12 98.982
R84 Y.n7 Y.n5 73.2449
R85 Y.n14 Y.n13 56.8057
R86 Y.n9 Y.n7 36.2672
R87 Y.n11 Y.n9 36.2672
R88 Y.n13 Y.n11 36.2672
R89 Y.n14 Y.n2 34.2593
R90 Y.n0 Y.t10 26.5955
R91 Y.n0 Y.t5 26.5955
R92 Y.n1 Y.t1 26.5955
R93 Y.n1 Y.t4 26.5955
R94 Y.n3 Y.t6 24.9236
R95 Y.n3 Y.t7 24.9236
R96 Y.n4 Y.t9 24.9236
R97 Y.n4 Y.t8 24.9236
R98 Y.n6 Y.t13 24.9236
R99 Y.n6 Y.t12 24.9236
R100 Y.n8 Y.t14 24.9236
R101 Y.n8 Y.t15 24.9236
R102 Y.n10 Y.t2 24.9236
R103 Y.n10 Y.t0 24.9236
R104 Y.n12 Y.t3 24.9236
R105 Y.n12 Y.t11 24.9236
R106 Y Y.n14 13.1907
R107 VNB.t7 VNB.t9 2677.02
R108 VNB.t8 VNB.t3 1196.12
R109 VNB.t2 VNB.t8 1196.12
R110 VNB.t1 VNB.t2 1196.12
R111 VNB.t11 VNB.t1 1196.12
R112 VNB.t12 VNB.t11 1196.12
R113 VNB.t10 VNB.t12 1196.12
R114 VNB.t9 VNB.t10 1196.12
R115 VNB.t6 VNB.t7 1196.12
R116 VNB.t4 VNB.t6 1196.12
R117 VNB.t5 VNB.t4 1196.12
R118 VNB.t0 VNB.t5 1196.12
R119 VNB VNB.t0 968.285
R120 A.n1 A.t6 212.081
R121 A.n4 A.t7 212.081
R122 A.n7 A.t0 212.081
R123 A.n6 A.t2 212.081
R124 A A.n8 163.582
R125 A.n3 A.n2 152
R126 A.n5 A.n0 152
R127 A.n1 A.t5 139.78
R128 A.n4 A.t4 139.78
R129 A.n7 A.t1 139.78
R130 A.n6 A.t3 139.78
R131 A.n7 A.n6 61.346
R132 A.n8 A.n5 49.6611
R133 A.n4 A.n3 39.4369
R134 A.n2 A 26.21
R135 A.n3 A.n1 21.9096
R136 A A.n0 18.8957
R137 A.n5 A.n4 10.2247
R138 A A.n0 9.14336
R139 A.n2 A 1.82907
R140 A.n8 A.n7 1.46111
R141 a_197_297.n3 a_197_297.n1 639.12
R142 a_197_297.n3 a_197_297.n2 585
R143 a_197_297.n4 a_197_297.n0 345.31
R144 a_197_297.n5 a_197_297.n4 300.885
R145 a_197_297.n4 a_197_297.n3 88.4254
R146 a_197_297.n2 a_197_297.t5 26.5955
R147 a_197_297.n2 a_197_297.t7 26.5955
R148 a_197_297.n1 a_197_297.t4 26.5955
R149 a_197_297.n1 a_197_297.t6 26.5955
R150 a_197_297.n0 a_197_297.t3 26.5955
R151 a_197_297.n0 a_197_297.t2 26.5955
R152 a_197_297.n5 a_197_297.t1 26.5955
R153 a_197_297.t0 a_197_297.n5 26.5955
R154 VPWR.n2 VPWR.t2 851.365
R155 VPWR.n4 VPWR.n3 606.505
R156 VPWR.n6 VPWR.n1 318.293
R157 VPWR.n1 VPWR.t3 26.5955
R158 VPWR.n1 VPWR.t0 26.5955
R159 VPWR.n3 VPWR.t1 26.5955
R160 VPWR.n3 VPWR.t4 26.5955
R161 VPWR.n6 VPWR.n5 24.4711
R162 VPWR.n5 VPWR.n4 19.9534
R163 VPWR.n5 VPWR.n0 9.3005
R164 VPWR.n7 VPWR.n6 7.34101
R165 VPWR.n4 VPWR.n2 6.8762
R166 VPWR.n2 VPWR.n0 0.688889
R167 VPWR.n7 VPWR.n0 0.145717
R168 VPWR VPWR.n7 0.116379
R169 VPB.t6 VPB.t12 556.386
R170 VPB.t2 VPB.t1 248.599
R171 VPB.t4 VPB.t2 248.599
R172 VPB.t3 VPB.t4 248.599
R173 VPB.t11 VPB.t3 248.599
R174 VPB.t10 VPB.t11 248.599
R175 VPB.t9 VPB.t10 248.599
R176 VPB.t12 VPB.t9 248.599
R177 VPB.t5 VPB.t6 248.599
R178 VPB.t8 VPB.t5 248.599
R179 VPB.t7 VPB.t8 248.599
R180 VPB.t0 VPB.t7 248.599
R181 VPB VPB.t0 201.246
R182 a_27_47.n11 a_27_47.n10 323.801
R183 a_27_47.t1 a_27_47.n11 255.287
R184 a_27_47.n2 a_27_47.t3 212.081
R185 a_27_47.n1 a_27_47.t6 212.081
R186 a_27_47.n7 a_27_47.t8 212.081
R187 a_27_47.n8 a_27_47.t7 212.081
R188 a_27_47.n11 a_27_47.t0 196.149
R189 a_27_47.n4 a_27_47.n3 172.725
R190 a_27_47.n10 a_27_47.n9 152
R191 a_27_47.n6 a_27_47.n0 152
R192 a_27_47.n5 a_27_47.n4 152
R193 a_27_47.n2 a_27_47.t5 139.78
R194 a_27_47.n1 a_27_47.t9 139.78
R195 a_27_47.n7 a_27_47.t4 139.78
R196 a_27_47.n8 a_27_47.t2 139.78
R197 a_27_47.n6 a_27_47.n5 49.6611
R198 a_27_47.n9 a_27_47.n7 48.2005
R199 a_27_47.n3 a_27_47.n1 39.4369
R200 a_27_47.n3 a_27_47.n2 21.9096
R201 a_27_47.n4 a_27_47.n0 20.7243
R202 a_27_47.n10 a_27_47.n0 20.7243
R203 a_27_47.n9 a_27_47.n8 13.146
R204 a_27_47.n5 a_27_47.n1 10.2247
R205 a_27_47.n7 a_27_47.n6 1.46111
R206 a_555_297.n1 a_555_297.t7 877.794
R207 a_555_297.n1 a_555_297.n0 585
R208 a_555_297.t3 a_555_297.n5 371.904
R209 a_555_297.n3 a_555_297.n2 300.885
R210 a_555_297.n5 a_555_297.n4 300.885
R211 a_555_297.n3 a_555_297.n1 49.2725
R212 a_555_297.n5 a_555_297.n3 44.424
R213 a_555_297.n0 a_555_297.t5 26.5955
R214 a_555_297.n0 a_555_297.t4 26.5955
R215 a_555_297.n2 a_555_297.t1 26.5955
R216 a_555_297.n2 a_555_297.t6 26.5955
R217 a_555_297.n4 a_555_297.t2 26.5955
R218 a_555_297.n4 a_555_297.t0 26.5955
R219 C_N.n0 C_N.t1 229.56
R220 C_N C_N.n0 159.619
R221 C_N.n0 C_N.t0 157.26
C0 B Y 0.174302f
C1 A VGND 0.062171f
C2 B VGND 0.050364f
C3 A B 0.029813f
C4 VPB VPWR 0.136599f
C5 VPWR Y 0.05487f
C6 VPB Y 0.032254f
C7 C_N VPWR 0.021656f
C8 VPB C_N 0.038398f
C9 VPWR VGND 0.134334f
C10 A VPWR 0.072992f
C11 C_N Y 8.06e-19
C12 VPB VGND 0.012462f
C13 VPB A 0.12176f
C14 Y VGND 0.885345f
C15 B VPWR 0.030354f
C16 A Y 0.197151f
C17 C_N VGND 0.015201f
C18 VPB B 0.120612f
C19 C_N A 0.050963f
C20 VGND VNB 0.766389f
C21 Y VNB 0.121117f
C22 VPWR VNB 0.626561f
C23 B VNB 0.362678f
C24 A VNB 0.367401f
C25 C_N VNB 0.142994f
C26 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_1 VPB VNB VGND VPWR Y D C B A
X0 Y.t1 B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1 a_191_297.t0 C.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR.t0 A.t0 a_297_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t3 C.t1 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X4 VGND.t2 A.t1 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_297_297.t0 B.t1 a_191_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297.t1 D.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y.t0 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t1 241.536
R1 B B.n0 188.722
R2 B.n0 B.t0 169.237
R3 VGND.n1 VGND.t2 285.038
R4 VGND.n5 VGND.t0 282.663
R5 VGND.n3 VGND.n2 200.127
R6 VGND.n4 VGND.n3 25.977
R7 VGND.n5 VGND.n4 25.977
R8 VGND.n2 VGND.t3 25.8467
R9 VGND.n2 VGND.t1 24.9236
R10 VGND.n6 VGND.n5 9.3005
R11 VGND.n4 VGND.n0 9.3005
R12 VGND.n3 VGND.n1 6.18988
R13 VGND.n1 VGND.n0 0.755914
R14 VGND.n6 VGND.n0 0.120292
R15 VGND VGND.n6 0.0226354
R16 Y Y.n0 593.216
R17 Y.n4 Y.n0 289.288
R18 Y.n3 Y.n2 259.729
R19 Y.n3 Y.n1 189.589
R20 Y.n4 Y.n3 81.9525
R21 Y.n1 Y.t0 42.462
R22 Y.n0 Y.t3 26.5955
R23 Y.n2 Y.t2 24.9236
R24 Y.n2 Y.t1 24.9236
R25 Y.n1 Y.t4 24.9236
R26 Y Y.n4 11.2013
R27 VNB.t0 VNB.t3 1466.67
R28 VNB.t3 VNB.t1 1210.36
R29 VNB.t1 VNB.t2 1196.12
R30 VNB VNB.t0 925.567
R31 C.n0 C.t0 241.536
R32 C.n0 C.t1 169.237
R33 C C.n0 167.065
R34 a_109_297.t0 a_109_297.t1 51.2205
R35 a_191_297.t0 a_191_297.t1 74.8605
R36 VPB.t0 VPB.t1 313.707
R37 VPB.t1 VPB.t2 248.599
R38 VPB.t3 VPB.t0 242.679
R39 VPB VPB.t3 192.369
R40 A.n0 A.t0 230.155
R41 A A.n0 171.446
R42 A.n0 A.t1 157.856
R43 a_297_297.t0 a_297_297.t1 53.1905
R44 VPWR VPWR.t0 349.659
R45 D.n0 D.t0 230.155
R46 D.n0 D.t1 157.856
R47 D D.n0 154.816
C0 A Y 0.017544f
C1 Y VPB 0.012654f
C2 VPB D 0.03755f
C3 VPWR Y 0.056134f
C4 VGND A 0.052553f
C5 VPWR D 0.012791f
C6 VGND VPB 0.004805f
C7 VPWR VGND 0.049214f
C8 B Y 0.040285f
C9 A VPB 0.040967f
C10 VPWR A 0.048251f
C11 VGND B 0.019083f
C12 VPWR VPB 0.052382f
C13 B A 0.110206f
C14 C Y 0.125478f
C15 C D 0.052345f
C16 B VPB 0.0304f
C17 VGND C 0.018387f
C18 VPWR B 0.088682f
C19 C A 0.002684f
C20 C VPB 0.029891f
C21 Y D 0.107589f
C22 VPWR C 0.050897f
C23 VGND Y 0.150668f
C24 VGND D 0.045612f
C25 C B 0.172838f
C26 VGND VNB 0.321875f
C27 VPWR VNB 0.276275f
C28 Y VNB 0.064476f
C29 A VNB 0.174401f
C30 B VNB 0.09682f
C31 C VNB 0.091102f
C32 D VNB 0.158827f
C33 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_2 VNB VPB VGND VPWR B D Y A C
X0 a_281_297.t3 B.t0 a_27_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t9 B.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t0 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297.t1 D.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t2 C.t0 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t0 D.t1 a_475_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t3 D.t2 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t4 A.t1 Y.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t7 A.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VGND.t6 B.t2 Y.t8 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t2 D.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t0 A.t3 a_27_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297.t2 C.t1 a_281_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_281_297.t1 C.t2 a_475_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297.t2 B.t3 a_281_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 Y.t1 C.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t0 212.081
R2 B B.n2 152.875
R3 B.n0 B.t2 139.78
R4 B.n1 B.t1 139.78
R5 B.n2 B.n0 32.8641
R6 B.n2 B.n1 28.4823
R7 a_27_297.n0 a_27_297.t2 371.904
R8 a_27_297.n0 a_27_297.t1 279.267
R9 a_27_297.n1 a_27_297.n0 208.506
R10 a_27_297.n1 a_27_297.t3 26.5955
R11 a_27_297.t0 a_27_297.n1 26.5955
R12 a_281_297.n1 a_281_297.n0 688.359
R13 a_281_297.n0 a_281_297.t0 26.5955
R14 a_281_297.n0 a_281_297.t1 26.5955
R15 a_281_297.t2 a_281_297.n1 26.5955
R16 a_281_297.n1 a_281_297.t3 26.5955
R17 VPB.t6 VPB.t5 580.062
R18 VPB.t1 VPB.t3 248.599
R19 VPB.t4 VPB.t1 248.599
R20 VPB.t5 VPB.t4 248.599
R21 VPB.t7 VPB.t6 248.599
R22 VPB.t0 VPB.t7 248.599
R23 VPB.t2 VPB.t0 248.599
R24 VPB VPB.t2 201.246
R25 VGND.n6 VGND.t3 286.986
R26 VGND.n11 VGND.t6 257.858
R27 VGND.n10 VGND.t0 257.858
R28 VGND.n5 VGND.n4 207.965
R29 VGND.n17 VGND.n1 207.965
R30 VGND.n19 VGND.t5 150.922
R31 VGND.n16 VGND.n2 34.6358
R32 VGND.n18 VGND.n17 32.377
R33 VGND.n9 VGND.n8 30.4887
R34 VGND.n8 VGND.n5 27.8593
R35 VGND.n4 VGND.t1 24.9236
R36 VGND.n4 VGND.t2 24.9236
R37 VGND.n1 VGND.t7 24.9236
R38 VGND.n1 VGND.t4 24.9236
R39 VGND.n19 VGND.n18 24.4711
R40 VGND.n11 VGND.n2 21.6534
R41 VGND.n6 VGND.n5 13.8844
R42 VGND.n20 VGND.n19 9.3005
R43 VGND.n8 VGND.n7 9.3005
R44 VGND.n9 VGND.n3 9.3005
R45 VGND.n13 VGND.n12 9.3005
R46 VGND.n14 VGND.n2 9.3005
R47 VGND.n16 VGND.n15 9.3005
R48 VGND.n18 VGND.n0 9.3005
R49 VGND.n12 VGND.n10 9.0005
R50 VGND.n17 VGND.n16 2.25932
R51 VGND.n12 VGND.n11 2.2005
R52 VGND.n7 VGND.n6 0.61214
R53 VGND.n10 VGND.n9 0.2005
R54 VGND.n7 VGND.n3 0.120292
R55 VGND.n13 VGND.n3 0.120292
R56 VGND.n14 VGND.n13 0.120292
R57 VGND.n15 VGND.n14 0.120292
R58 VGND.n15 VGND.n0 0.120292
R59 VGND.n20 VGND.n0 0.120292
R60 VGND VGND.n20 0.0213333
R61 Y.n8 Y.n7 349.293
R62 Y.n2 Y.n0 135.249
R63 Y.n2 Y.n1 98.982
R64 Y.n4 Y.n3 98.982
R65 Y.n6 Y.n5 98.982
R66 Y.n4 Y.n2 76.0894
R67 Y.n6 Y.n4 36.2672
R68 Y.n7 Y.t3 26.5955
R69 Y.n7 Y.t0 26.5955
R70 Y.n0 Y.t6 24.9236
R71 Y.n0 Y.t7 24.9236
R72 Y.n1 Y.t8 24.9236
R73 Y.n1 Y.t9 24.9236
R74 Y.n3 Y.t4 24.9236
R75 Y.n3 Y.t1 24.9236
R76 Y.n5 Y.t5 24.9236
R77 Y.n5 Y.t2 24.9236
R78 Y.n8 Y.n6 16.7116
R79 Y Y.n8 1.91095
R80 VNB.t6 VNB.t0 2790.94
R81 VNB.t1 VNB.t3 1196.12
R82 VNB.t2 VNB.t1 1196.12
R83 VNB.t0 VNB.t2 1196.12
R84 VNB.t7 VNB.t6 1196.12
R85 VNB.t4 VNB.t7 1196.12
R86 VNB.t5 VNB.t4 1196.12
R87 VNB VNB.t5 968.285
R88 A.n0 A.t0 212.081
R89 A.n1 A.t3 212.081
R90 A A.n2 152.921
R91 A.n0 A.t1 139.78
R92 A.n1 A.t2 139.78
R93 A.n2 A.n0 38.7066
R94 A.n2 A.n1 22.6399
R95 VPWR VPWR.n0 324.387
R96 VPWR.n0 VPWR.t1 26.5955
R97 VPWR.n0 VPWR.t0 26.5955
R98 D.n0 D.t0 212.081
R99 D.n1 D.t1 212.081
R100 D D.n2 174.553
R101 D.n0 D.t2 139.78
R102 D.n1 D.t3 139.78
R103 D.n2 D.n0 33.5944
R104 D.n2 D.n1 27.752
R105 a_475_297.n1 a_475_297.t3 392.906
R106 a_475_297.t1 a_475_297.n1 392.906
R107 a_475_297.n1 a_475_297.n0 187.506
R108 a_475_297.n0 a_475_297.t0 26.5955
R109 a_475_297.n0 a_475_297.t2 26.5955
R110 C.n0 C.t1 212.081
R111 C.n1 C.t2 212.081
R112 C C.n2 180.649
R113 C.n0 C.t0 139.78
R114 C.n1 C.t3 139.78
R115 C.n2 C.n0 30.6732
R116 C.n2 C.n1 30.6732
C0 VPWR VGND 0.090165f
C1 VGND A 0.050759f
C2 VPWR C 0.022213f
C3 Y B 0.098054f
C4 Y VGND 0.610575f
C5 Y C 0.108438f
C6 VGND B 0.030223f
C7 B C 0.031131f
C8 VGND C 0.031089f
C9 D VPB 0.056793f
C10 D VPWR 0.016136f
C11 VPWR VPB 0.092403f
C12 VPB A 0.056022f
C13 D Y 0.154521f
C14 Y VPB 0.016666f
C15 VPWR A 0.04358f
C16 VPB B 0.057664f
C17 D VGND 0.026848f
C18 VPWR Y 0.02023f
C19 VPWR B 0.022495f
C20 VGND VPB 0.011501f
C21 Y A 0.061442f
C22 D C 0.067517f
C23 VPB C 0.060484f
C24 A B 0.069132f
C25 VGND VNB 0.576715f
C26 Y VNB 0.0798f
C27 VPWR VNB 0.440934f
C28 D VNB 0.19659f
C29 C VNB 0.18423f
C30 B VNB 0.181984f
C31 A VNB 0.206594f
C32 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_4 VPB VNB VGND VPWR A B Y D C
X0 VPWR.t3 A.t0 a_27_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_807_297.t7 D.t0 Y.t13 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t7 C.t0 Y.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t4 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t12 D.t1 a_807_297.t6 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297.t3 A.t2 VPWR.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t1 C.t1 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t14 D.t2 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t2 C.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X9 Y.t9 D.t3 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t2 A.t3 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_297.t0 B.t0 a_449_297.t7 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 Y.t6 A.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 VGND.t0 A.t5 Y.t5 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t12 B.t1 Y.t15 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t13 B.t2 Y.t16 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_449_297.t6 B.t3 a_27_297.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_807_297.t0 C.t3 a_449_297.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND.t9 D.t4 Y.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VGND.t8 D.t5 Y.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_807_297.t1 C.t4 a_449_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR.t1 A.t6 a_27_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X22 a_449_297.t1 C.t5 a_807_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y.t17 B.t4 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 Y.t18 B.t5 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_449_297.t0 C.t6 a_807_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_27_297.t6 B.t6 a_449_297.t5 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_807_297.t5 D.t6 Y.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X28 a_449_297.t4 B.t7 a_27_297.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y.t10 D.t7 a_807_297.t4 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_297.t1 A.t7 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VGND.t4 C.t7 Y.t19 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n3 A.t7 212.081
R1 A.n5 A.t0 212.081
R2 A.n7 A.t2 212.081
R3 A.n1 A.t6 212.081
R4 A.n4 A.n0 172.725
R5 A.n9 A.n2 172.725
R6 A.n6 A.n0 152
R7 A.n9 A.n8 152
R8 A.n3 A.t5 139.78
R9 A.n5 A.t1 139.78
R10 A.n7 A.t3 139.78
R11 A.n1 A.t4 139.78
R12 A.n8 A.n6 49.6611
R13 A.n7 A.n2 48.2005
R14 A.n5 A.n4 39.4369
R15 A.n4 A.n3 21.9096
R16 A.n2 A.n1 13.146
R17 A A.n0 11.5815
R18 A.n6 A.n5 10.2247
R19 A A.n9 9.14336
R20 A.n8 A.n7 1.46111
R21 a_27_297.t0 a_27_297.n5 370.401
R22 a_27_297.n5 a_27_297.n4 300.885
R23 a_27_297.n1 a_27_297.t2 276.781
R24 a_27_297.n1 a_27_297.n0 208.507
R25 a_27_297.n3 a_27_297.n2 187.506
R26 a_27_297.n3 a_27_297.n1 65.4262
R27 a_27_297.n5 a_27_297.n3 65.4258
R28 a_27_297.n2 a_27_297.t7 26.5955
R29 a_27_297.n2 a_27_297.t1 26.5955
R30 a_27_297.n0 a_27_297.t4 26.5955
R31 a_27_297.n0 a_27_297.t3 26.5955
R32 a_27_297.n4 a_27_297.t5 26.5955
R33 a_27_297.n4 a_27_297.t6 26.5955
R34 VPWR.n2 VPWR.n0 323.974
R35 VPWR.n2 VPWR.n1 323.86
R36 VPWR.n1 VPWR.t2 26.5955
R37 VPWR.n1 VPWR.t1 26.5955
R38 VPWR.n0 VPWR.t0 26.5955
R39 VPWR.n0 VPWR.t3 26.5955
R40 VPWR VPWR.n2 0.505993
R41 VPB.t0 VPB.t4 556.386
R42 VPB.t10 VPB.t9 248.599
R43 VPB.t11 VPB.t10 248.599
R44 VPB.t12 VPB.t11 248.599
R45 VPB.t1 VPB.t12 248.599
R46 VPB.t3 VPB.t1 248.599
R47 VPB.t2 VPB.t3 248.599
R48 VPB.t4 VPB.t2 248.599
R49 VPB.t13 VPB.t0 248.599
R50 VPB.t14 VPB.t13 248.599
R51 VPB.t15 VPB.t14 248.599
R52 VPB.t5 VPB.t15 248.599
R53 VPB.t8 VPB.t5 248.599
R54 VPB.t7 VPB.t8 248.599
R55 VPB.t6 VPB.t7 248.599
R56 VPB VPB.t6 201.246
R57 D.n2 D.t6 212.081
R58 D.n4 D.t7 212.081
R59 D.n6 D.t0 212.081
R60 D.n1 D.t1 212.081
R61 D.n3 D.n0 172.725
R62 D.n5 D.n0 152
R63 D.n2 D.t5 139.78
R64 D.n4 D.t3 139.78
R65 D.n6 D.t4 139.78
R66 D.n1 D.t2 139.78
R67 D D.n7 78.6602
R68 D.n6 D.n5 46.7399
R69 D.n4 D.n3 35.055
R70 D.n7 D.n1 31.6758
R71 D.n3 D.n2 26.2914
R72 D.n7 D.n6 23.0844
R73 D.n5 D.n4 14.6066
R74 D D.n0 12.191
R75 Y.n17 Y.n15 345.31
R76 Y.n17 Y.n16 300.885
R77 Y.n2 Y.n0 135.249
R78 Y.n2 Y.n1 98.982
R79 Y.n4 Y.n3 98.982
R80 Y.n6 Y.n5 98.982
R81 Y.n8 Y.n7 98.982
R82 Y.n10 Y.n9 98.982
R83 Y.n12 Y.n11 98.982
R84 Y.n14 Y.n13 98.982
R85 Y.n8 Y.n6 73.2449
R86 Y.n18 Y.n17 52.4415
R87 Y.n4 Y.n2 36.2672
R88 Y.n6 Y.n4 36.2672
R89 Y.n10 Y.n8 36.2672
R90 Y.n12 Y.n10 36.2672
R91 Y.n14 Y.n12 36.2672
R92 Y.n15 Y.t13 26.5955
R93 Y.n15 Y.t12 26.5955
R94 Y.n16 Y.t11 26.5955
R95 Y.n16 Y.t10 26.5955
R96 Y.n0 Y.t3 24.9236
R97 Y.n0 Y.t6 24.9236
R98 Y.n1 Y.t5 24.9236
R99 Y.n1 Y.t4 24.9236
R100 Y.n3 Y.t15 24.9236
R101 Y.n3 Y.t17 24.9236
R102 Y.n5 Y.t16 24.9236
R103 Y.n5 Y.t18 24.9236
R104 Y.n7 Y.t0 24.9236
R105 Y.n7 Y.t2 24.9236
R106 Y.n9 Y.t19 24.9236
R107 Y.n9 Y.t1 24.9236
R108 Y.n11 Y.t8 24.9236
R109 Y.n11 Y.t14 24.9236
R110 Y.n13 Y.t7 24.9236
R111 Y.n13 Y.t9 24.9236
R112 Y.n18 Y.n14 14.2227
R113 Y Y.n18 2.37087
R114 a_807_297.n3 a_807_297.t5 371.904
R115 a_807_297.n1 a_807_297.t3 371.01
R116 a_807_297.n3 a_807_297.n2 300.885
R117 a_807_297.n1 a_807_297.n0 300.885
R118 a_807_297.n5 a_807_297.n4 300.885
R119 a_807_297.n4 a_807_297.n1 44.424
R120 a_807_297.n4 a_807_297.n3 44.424
R121 a_807_297.n2 a_807_297.t4 26.5955
R122 a_807_297.n2 a_807_297.t7 26.5955
R123 a_807_297.n0 a_807_297.t2 26.5955
R124 a_807_297.n0 a_807_297.t1 26.5955
R125 a_807_297.t6 a_807_297.n5 26.5955
R126 a_807_297.n5 a_807_297.t0 26.5955
R127 C.n2 C.t3 212.081
R128 C.n1 C.t5 212.081
R129 C.n7 C.t4 212.081
R130 C.n8 C.t6 212.081
R131 C.n4 C.n3 172.725
R132 C C.n9 169.677
R133 C.n5 C.n4 152
R134 C.n6 C.n0 152
R135 C.n2 C.t7 139.78
R136 C.n1 C.t1 139.78
R137 C.n7 C.t0 139.78
R138 C.n8 C.t2 139.78
R139 C.n6 C.n5 49.6611
R140 C.n9 C.n7 48.2005
R141 C.n3 C.n1 39.4369
R142 C.n3 C.n2 21.9096
R143 C.n4 C.n0 20.7243
R144 C.n9 C.n8 13.146
R145 C.n5 C.n1 10.2247
R146 C C.n0 3.04812
R147 C.n7 C.n6 1.46111
R148 VGND.n14 VGND.t8 294.512
R149 VGND.n13 VGND.n12 207.965
R150 VGND.n18 VGND.n10 207.965
R151 VGND.n8 VGND.n7 207.965
R152 VGND.n34 VGND.n4 207.965
R153 VGND.n37 VGND.n36 207.965
R154 VGND.n43 VGND.n1 207.965
R155 VGND.n28 VGND.n27 185
R156 VGND.n26 VGND.n25 185
R157 VGND.n45 VGND.t1 150.922
R158 VGND.n27 VGND.n26 96.0005
R159 VGND.n14 VGND.n13 39.0017
R160 VGND.n17 VGND.n11 34.6358
R161 VGND.n20 VGND.n19 34.6358
R162 VGND.n24 VGND.n23 34.6358
R163 VGND.n33 VGND.n5 34.6358
R164 VGND.n38 VGND.n35 34.6358
R165 VGND.n42 VGND.n2 34.6358
R166 VGND.n44 VGND.n43 32.377
R167 VGND.n18 VGND.n17 27.8593
R168 VGND.n37 VGND.n2 26.3534
R169 VGND.n26 VGND.t5 24.9236
R170 VGND.n27 VGND.t13 24.9236
R171 VGND.n12 VGND.t10 24.9236
R172 VGND.n12 VGND.t9 24.9236
R173 VGND.n10 VGND.t11 24.9236
R174 VGND.n10 VGND.t4 24.9236
R175 VGND.n7 VGND.t6 24.9236
R176 VGND.n7 VGND.t7 24.9236
R177 VGND.n4 VGND.t15 24.9236
R178 VGND.n4 VGND.t12 24.9236
R179 VGND.n36 VGND.t14 24.9236
R180 VGND.n36 VGND.t0 24.9236
R181 VGND.n1 VGND.t3 24.9236
R182 VGND.n1 VGND.t2 24.9236
R183 VGND.n45 VGND.n44 24.4711
R184 VGND.n20 VGND.n8 21.8358
R185 VGND.n35 VGND.n34 20.3299
R186 VGND.n34 VGND.n33 14.3064
R187 VGND.n23 VGND.n8 12.8005
R188 VGND.n25 VGND.n24 11.1123
R189 VGND.n28 VGND.n5 9.60638
R190 VGND.n46 VGND.n45 9.3005
R191 VGND.n15 VGND.n11 9.3005
R192 VGND.n17 VGND.n16 9.3005
R193 VGND.n19 VGND.n9 9.3005
R194 VGND.n21 VGND.n20 9.3005
R195 VGND.n23 VGND.n22 9.3005
R196 VGND.n24 VGND.n6 9.3005
R197 VGND.n30 VGND.n29 9.3005
R198 VGND.n31 VGND.n5 9.3005
R199 VGND.n33 VGND.n32 9.3005
R200 VGND.n35 VGND.n3 9.3005
R201 VGND.n39 VGND.n38 9.3005
R202 VGND.n40 VGND.n2 9.3005
R203 VGND.n42 VGND.n41 9.3005
R204 VGND.n44 VGND.n0 9.3005
R205 VGND.n38 VGND.n37 8.28285
R206 VGND.n19 VGND.n18 6.77697
R207 VGND.n29 VGND.n28 5.4005
R208 VGND.n29 VGND.n25 5.0005
R209 VGND.n15 VGND.n14 2.68138
R210 VGND.n43 VGND.n42 2.25932
R211 VGND.n13 VGND.n11 0.753441
R212 VGND.n16 VGND.n15 0.120292
R213 VGND.n16 VGND.n9 0.120292
R214 VGND.n21 VGND.n9 0.120292
R215 VGND.n22 VGND.n21 0.120292
R216 VGND.n22 VGND.n6 0.120292
R217 VGND.n30 VGND.n6 0.120292
R218 VGND.n31 VGND.n30 0.120292
R219 VGND.n32 VGND.n31 0.120292
R220 VGND.n32 VGND.n3 0.120292
R221 VGND.n39 VGND.n3 0.120292
R222 VGND.n40 VGND.n39 0.120292
R223 VGND.n41 VGND.n40 0.120292
R224 VGND.n41 VGND.n0 0.120292
R225 VGND.n46 VGND.n0 0.120292
R226 VGND VGND.n46 0.0213333
R227 VNB.t13 VNB.t5 2677.02
R228 VNB.t10 VNB.t8 1196.12
R229 VNB.t9 VNB.t10 1196.12
R230 VNB.t11 VNB.t9 1196.12
R231 VNB.t4 VNB.t11 1196.12
R232 VNB.t6 VNB.t4 1196.12
R233 VNB.t7 VNB.t6 1196.12
R234 VNB.t5 VNB.t7 1196.12
R235 VNB.t15 VNB.t13 1196.12
R236 VNB.t12 VNB.t15 1196.12
R237 VNB.t14 VNB.t12 1196.12
R238 VNB.t0 VNB.t14 1196.12
R239 VNB.t3 VNB.t0 1196.12
R240 VNB.t2 VNB.t3 1196.12
R241 VNB.t1 VNB.t2 1196.12
R242 VNB VNB.t1 968.285
R243 B.n3 B.t0 212.081
R244 B.n6 B.t3 212.081
R245 B.n8 B.t6 212.081
R246 B.n1 B.t7 212.081
R247 B.n10 B.n2 172.725
R248 B.n5 B.n4 152
R249 B.n7 B.n0 152
R250 B.n10 B.n9 152
R251 B.n3 B.t2 139.78
R252 B.n6 B.t5 139.78
R253 B.n8 B.t1 139.78
R254 B.n1 B.t4 139.78
R255 B.n9 B.n7 49.6611
R256 B.n8 B.n2 48.2005
R257 B.n6 B.n5 39.4369
R258 B.n5 B.n3 21.9096
R259 B.n4 B.n0 20.7243
R260 B B.n10 18.8957
R261 B.n2 B.n1 13.146
R262 B.n7 B.n6 10.2247
R263 B.n4 B 5.48621
R264 B B.n0 1.82907
R265 B.n9 B.n8 1.46111
R266 a_449_297.n2 a_449_297.n0 345.31
R267 a_449_297.n5 a_449_297.n4 345.308
R268 a_449_297.n2 a_449_297.n1 300.885
R269 a_449_297.n4 a_449_297.n3 300.885
R270 a_449_297.n4 a_449_297.n2 83.577
R271 a_449_297.n0 a_449_297.t5 26.5955
R272 a_449_297.n0 a_449_297.t4 26.5955
R273 a_449_297.n1 a_449_297.t7 26.5955
R274 a_449_297.n1 a_449_297.t6 26.5955
R275 a_449_297.n3 a_449_297.t2 26.5955
R276 a_449_297.n3 a_449_297.t0 26.5955
R277 a_449_297.t3 a_449_297.n5 26.5955
R278 a_449_297.n5 a_449_297.t1 26.5955
C0 A B 0.064024f
C1 Y B 0.228595f
C2 C VGND 0.051297f
C3 D VGND 0.060366f
C4 VGND VPB 0.012049f
C5 C D 0.068777f
C6 VPWR VGND 0.150605f
C7 C VPB 0.120618f
C8 VGND A 0.083785f
C9 C VPWR 0.031063f
C10 Y VGND 1.11928f
C11 D VPB 0.11978f
C12 VGND B 0.051942f
C13 C Y 0.18445f
C14 D VPWR 0.034379f
C15 C B 0.034032f
C16 VPWR VPB 0.140426f
C17 D Y 0.368015f
C18 VPB A 0.119932f
C19 Y VPB 0.01493f
C20 VPWR A 0.08856f
C21 VPWR Y 0.030393f
C22 VPB B 0.122233f
C23 VPWR B 0.032908f
C24 Y A 0.166171f
C25 VGND VNB 0.89449f
C26 Y VNB 0.081809f
C27 VPWR VNB 0.703863f
C28 D VNB 0.380799f
C29 C VNB 0.362819f
C30 B VNB 0.369648f
C31 A VNB 0.391825f
C32 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4b_1 VPB VNB VGND VPWR D_N C Y B A
X0 Y.t3 a_91_199.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1 Y.t0 B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND.t1 C.t0 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_91_199.t0 D_N.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND.t2 A.t0 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t0 A.t1 a_341_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6 a_245_297.t1 C.t1 a_161_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_341_297.t0 B.t1 a_245_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X8 a_91_199.t1 D_N.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X9 a_161_297.t1 a_91_199.t3 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
R0 a_91_199.n1 a_91_199.t1 648.322
R1 a_91_199.t0 a_91_199.n1 338.163
R2 a_91_199.n1 a_91_199.n0 316.959
R3 a_91_199.n0 a_91_199.t3 234.804
R4 a_91_199.n0 a_91_199.t2 162.504
R5 VGND.n8 VGND.t4 284.678
R6 VGND.n2 VGND.n1 200.127
R7 VGND.n4 VGND.n3 116.157
R8 VGND.n3 VGND.t3 57.875
R9 VGND.n7 VGND.n6 34.6358
R10 VGND.n1 VGND.t0 30.462
R11 VGND.n1 VGND.t1 30.462
R12 VGND.n3 VGND.t2 24.6931
R13 VGND.n9 VGND.n8 18.7123
R14 VGND.n4 VGND.n2 10.6873
R15 VGND.n7 VGND.n0 9.3005
R16 VGND.n6 VGND.n5 9.3005
R17 VGND.n6 VGND.n2 5.64756
R18 VGND.n5 VGND.n4 1.15067
R19 VGND.n8 VGND.n7 0.376971
R20 VGND.n5 VGND.n0 0.120292
R21 VGND.n9 VGND.n0 0.120292
R22 VGND VGND.n9 0.0226354
R23 Y Y.t4 382.32
R24 Y.n2 Y.n0 251.127
R25 Y.n2 Y.n1 200.68
R26 Y Y.n2 89.8467
R27 Y.n0 Y.t2 24.9236
R28 Y.n0 Y.t0 24.9236
R29 Y.n1 Y.t1 24.9236
R30 Y.n1 Y.t3 24.9236
R31 VNB VNB.t4 1666.02
R32 VNB.t2 VNB.t3 1381.23
R33 VNB.t1 VNB.t0 1366.99
R34 VNB.t0 VNB.t2 1196.12
R35 VNB.t4 VNB.t1 1196.12
R36 B.n0 B.t1 241.536
R37 B.n0 B.t0 169.237
R38 B B.n0 154.168
R39 C.n0 C.t1 241.536
R40 C.n0 C.t0 169.237
R41 C C.n0 153.756
R42 D_N.n0 D_N.t1 211.01
R43 D_N D_N.n0 154.994
R44 D_N.n0 D_N.t0 132.282
R45 A.n0 A.t1 241.536
R46 A.n0 A.t0 169.237
R47 A A.n0 154.582
R48 a_341_297.t0 a_341_297.t1 53.1905
R49 VPWR VPWR.n0 611.409
R50 VPWR.n0 VPWR.t1 96.1553
R51 VPWR.n0 VPWR.t0 27.9645
R52 VPB VPB.t4 346.262
R53 VPB.t1 VPB.t2 287.072
R54 VPB.t3 VPB.t0 284.113
R55 VPB.t0 VPB.t1 248.599
R56 VPB.t4 VPB.t3 248.599
R57 a_161_297.t0 a_161_297.t1 53.1905
R58 a_245_297.t0 a_245_297.t1 65.0105
C0 VGND A 0.038485f
C1 Y D_N 7.15e-19
C2 VPB C 0.0278f
C3 B A 0.108301f
C4 VPWR VPB 0.077888f
C5 Y C 0.038588f
C6 D_N A 0.090907f
C7 VGND B 0.01441f
C8 Y VPWR 0.053626f
C9 D_N VGND 0.018525f
C10 Y VPB 0.013415f
C11 VGND C 0.013779f
C12 VPWR A 0.016549f
C13 D_N B 3.76e-19
C14 VPWR VGND 0.063428f
C15 C B 0.102789f
C16 VPB A 0.03087f
C17 D_N C 1.64e-19
C18 VPWR B 0.010542f
C19 VGND VPB 0.007986f
C20 Y A 0.003117f
C21 Y VGND 0.252703f
C22 VPWR D_N 0.006724f
C23 VPB B 0.027966f
C24 D_N VPB 0.06112f
C25 VPWR C 0.00875f
C26 Y B 0.040324f
C27 VGND VNB 0.41827f
C28 D_N VNB 0.12553f
C29 VPWR VNB 0.341029f
C30 Y VNB 0.101031f
C31 A VNB 0.095088f
C32 B VNB 0.089124f
C33 C VNB 0.088776f
C34 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4b_2 VNB VPB VGND VPWR A B C Y D_N
X0 VPWR.t2 D_N.t0 a_694_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_27_297.t1 B.t0 a_277_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_474_297.t2 a_694_21.t2 Y.t8 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_277_297.t1 B.t1 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t5 a_694_21.t3 a_474_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t3 C.t0 Y.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND.t6 D_N.t1 a_694_21.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_27_297.t2 A.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t5 A.t1 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t1 B.t2 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t9 C.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_474_297.t3 C.t2 a_277_297.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y.t0 B.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t7 a_694_21.t4 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_277_297.t2 C.t3 a_474_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t7 a_694_21.t5 Y.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t1 A.t2 a_27_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y.t3 A.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 D_N.n0 D_N.t0 334.188
R1 D_N D_N.n0 168.946
R2 D_N.n0 D_N.t1 131.748
R3 a_694_21.n2 a_694_21.t1 720.273
R4 a_694_21.t0 a_694_21.n2 248.66
R5 a_694_21.n2 a_694_21.n1 227.952
R6 a_694_21.n1 a_694_21.t2 212.081
R7 a_694_21.n0 a_694_21.t3 212.081
R8 a_694_21.n1 a_694_21.t5 139.78
R9 a_694_21.n0 a_694_21.t4 139.78
R10 a_694_21.n1 a_694_21.n0 61.346
R11 VPWR.n1 VPWR.t2 678.777
R12 VPWR.n1 VPWR.n0 329.233
R13 VPWR.n0 VPWR.t0 26.5955
R14 VPWR.n0 VPWR.t1 26.5955
R15 VPWR VPWR.n1 0.149648
R16 VPB.t1 VPB.t3 577.104
R17 VPB.t7 VPB.t5 556.386
R18 VPB.t6 VPB.t7 248.599
R19 VPB.t8 VPB.t6 248.599
R20 VPB.t3 VPB.t8 248.599
R21 VPB.t0 VPB.t1 248.599
R22 VPB.t2 VPB.t0 248.599
R23 VPB.t4 VPB.t2 248.599
R24 VPB VPB.t4 192.369
R25 B.n0 B.t0 212.081
R26 B.n1 B.t1 212.081
R27 B B.n2 156.571
R28 B.n0 B.t2 139.78
R29 B.n1 B.t3 139.78
R30 B.n2 B.n1 40.1672
R31 B.n2 B.n0 21.1793
R32 a_277_297.n1 a_277_297.n0 697.17
R33 a_277_297.n0 a_277_297.t3 26.5955
R34 a_277_297.n0 a_277_297.t2 26.5955
R35 a_277_297.t0 a_277_297.n1 26.5955
R36 a_277_297.n1 a_277_297.t1 26.5955
R37 a_27_297.t1 a_27_297.n1 367.259
R38 a_27_297.n1 a_27_297.t3 273.365
R39 a_27_297.n1 a_27_297.n0 208.507
R40 a_27_297.n0 a_27_297.t0 26.5955
R41 a_27_297.n0 a_27_297.t2 26.5955
R42 Y.n8 Y.n0 301.979
R43 Y.n3 Y.n1 135.249
R44 Y.n3 Y.n2 98.982
R45 Y.n5 Y.n4 98.982
R46 Y.n7 Y.n6 98.982
R47 Y.n5 Y.n3 75.7338
R48 Y.n7 Y.n5 36.2672
R49 Y Y.n7 28.906
R50 Y.n0 Y.t8 26.5955
R51 Y.n0 Y.t5 26.5955
R52 Y.n6 Y.t6 24.9236
R53 Y.n6 Y.t7 24.9236
R54 Y.n1 Y.t4 24.9236
R55 Y.n1 Y.t3 24.9236
R56 Y.n2 Y.t1 24.9236
R57 Y.n2 Y.t0 24.9236
R58 Y.n4 Y.t2 24.9236
R59 Y.n4 Y.t9 24.9236
R60 Y.n8 Y 0.4005
R61 Y Y.n8 0.316549
R62 a_474_297.t2 a_474_297.n1 393.075
R63 a_474_297.n1 a_474_297.t0 387.301
R64 a_474_297.n1 a_474_297.n0 187.506
R65 a_474_297.n0 a_474_297.t1 26.5955
R66 a_474_297.n0 a_474_297.t3 26.5955
R67 C.n0 C.t2 212.081
R68 C.n1 C.t3 212.081
R69 C C.n2 156.571
R70 C.n0 C.t0 139.78
R71 C.n1 C.t1 139.78
R72 C.n2 C.n1 40.1672
R73 C.n2 C.n0 21.1793
R74 VGND.n7 VGND.t6 264.7
R75 VGND.n16 VGND.t1 263.462
R76 VGND.n15 VGND.t2 263.462
R77 VGND.n5 VGND.n4 207.965
R78 VGND.n22 VGND.n1 207.965
R79 VGND.n8 VGND.t7 161.185
R80 VGND.n24 VGND.t4 154.988
R81 VGND.n10 VGND.n9 34.6358
R82 VGND.n21 VGND.n2 34.6358
R83 VGND.n14 VGND.n13 31.8711
R84 VGND.n23 VGND.n22 30.8711
R85 VGND.n13 VGND.n5 25.977
R86 VGND.n24 VGND.n23 25.977
R87 VGND.n4 VGND.t8 24.9236
R88 VGND.n4 VGND.t3 24.9236
R89 VGND.n1 VGND.t0 24.9236
R90 VGND.n1 VGND.t5 24.9236
R91 VGND.n16 VGND.n2 20.1476
R92 VGND.n9 VGND.n8 13.5534
R93 VGND.n8 VGND.n7 12.5758
R94 VGND.n25 VGND.n24 9.3005
R95 VGND.n9 VGND.n6 9.3005
R96 VGND.n11 VGND.n10 9.3005
R97 VGND.n13 VGND.n12 9.3005
R98 VGND.n14 VGND.n3 9.3005
R99 VGND.n18 VGND.n17 9.3005
R100 VGND.n19 VGND.n2 9.3005
R101 VGND.n21 VGND.n20 9.3005
R102 VGND.n23 VGND.n0 9.3005
R103 VGND.n10 VGND.n5 8.65932
R104 VGND.n17 VGND.n15 8.5005
R105 VGND.n22 VGND.n21 3.76521
R106 VGND.n17 VGND.n16 2.6005
R107 VGND.n7 VGND.n6 0.792188
R108 VGND.n15 VGND.n14 0.7005
R109 VGND.n11 VGND.n6 0.120292
R110 VGND.n12 VGND.n11 0.120292
R111 VGND.n12 VGND.n3 0.120292
R112 VGND.n18 VGND.n3 0.120292
R113 VGND.n19 VGND.n18 0.120292
R114 VGND.n20 VGND.n19 0.120292
R115 VGND.n20 VGND.n0 0.120292
R116 VGND.n25 VGND.n0 0.120292
R117 VGND VGND.n25 0.0226354
R118 VNB.t1 VNB.t2 2776.7
R119 VNB.t7 VNB.t6 2677.02
R120 VNB.t8 VNB.t7 1196.12
R121 VNB.t3 VNB.t8 1196.12
R122 VNB.t2 VNB.t3 1196.12
R123 VNB.t0 VNB.t1 1196.12
R124 VNB.t5 VNB.t0 1196.12
R125 VNB.t4 VNB.t5 1196.12
R126 VNB VNB.t4 925.567
R127 A.n0 A.t0 212.081
R128 A.n1 A.t2 212.081
R129 A A.n2 152.619
R130 A.n0 A.t1 139.78
R131 A.n1 A.t3 139.78
R132 A.n2 A.n0 38.7066
R133 A.n2 A.n1 22.6399
C0 VGND B 0.031649f
C1 Y B 0.134698f
C2 VPB A 0.056844f
C3 VPB B 0.061511f
C4 C VPWR 0.021029f
C5 VGND C 0.030356f
C6 A B 0.071745f
C7 C Y 0.112979f
C8 D_N VPWR 0.039993f
C9 VGND D_N 0.043568f
C10 D_N Y 0.001445f
C11 VGND VPWR 0.10707f
C12 VPWR Y 0.013832f
C13 C VPB 0.057655f
C14 VGND Y 0.596793f
C15 D_N VPB 0.114753f
C16 C B 0.039237f
C17 VPWR VPB 0.12035f
C18 VGND VPB 0.01388f
C19 Y VPB 0.007074f
C20 VPWR A 0.038692f
C21 VGND A 0.058253f
C22 VPWR B 0.023258f
C23 Y A 0.085441f
C24 VGND VNB 0.6979f
C25 Y VNB 0.024376f
C26 VPWR VNB 0.536012f
C27 D_N VNB 0.176252f
C28 C VNB 0.180624f
C29 B VNB 0.186947f
C30 A VNB 0.210159f
C31 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4b_4 VPB VNB VGND VPWR B D_N A C Y
X0 VGND.t6 B.t0 Y.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t5 B.t1 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t2 D_N.t0 a_1191_21.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_803_297.t7 a_1191_21.t2 Y.t10 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_445_297.t5 B.t2 a_27_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297.t6 A.t0 VPWR.t4 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t11 a_1191_21.t3 a_803_297.t6 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_803_297.t5 a_1191_21.t4 Y.t12 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t7 C.t0 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t3 A.t1 a_27_297.t7 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y.t13 a_1191_21.t5 a_803_297.t4 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y.t8 C.t1 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X12 Y.t14 a_1191_21.t6 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297.t5 A.t2 VPWR.t2 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t0 D_N.t1 a_1191_21.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t16 A.t3 Y.t19 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t0 A.t4 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t10 C.t2 Y.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297.t2 B.t3 a_445_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t15 C.t3 Y.t18 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND.t12 a_1191_21.t7 Y.t15 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t13 a_1191_21.t8 Y.t16 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t1 A.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y.t3 B.t4 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_445_297.t3 B.t5 a_27_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_803_297.t3 C.t4 a_445_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y.t2 B.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 a_27_297.t0 B.t7 a_445_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_445_297.t0 C.t5 a_803_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_803_297.t2 C.t6 a_445_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y.t17 a_1191_21.t9 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR.t1 A.t6 a_27_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_445_297.t1 C.t7 a_803_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 Y.t6 A.t7 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n3 B.t3 212.081
R1 B.n5 B.t5 212.081
R2 B.n7 B.t7 212.081
R3 B.n1 B.t2 212.081
R4 B.n4 B.n0 172.725
R5 B.n9 B.n2 172.725
R6 B.n6 B.n0 152
R7 B.n9 B.n8 152
R8 B.n3 B.t1 139.78
R9 B.n5 B.t6 139.78
R10 B.n7 B.t0 139.78
R11 B.n1 B.t4 139.78
R12 B.n8 B.n6 49.6611
R13 B.n7 B.n2 48.2005
R14 B.n5 B.n4 39.4369
R15 B.n4 B.n3 21.9096
R16 B B.n9 18.8957
R17 B.n2 B.n1 13.146
R18 B.n6 B.n5 10.2247
R19 B B.n0 1.82907
R20 B.n8 B.n7 1.46111
R21 Y Y.n0 593.961
R22 Y.n18 Y.n0 585
R23 Y.n17 Y.n1 337.779
R24 Y.n16 Y.n2 143.427
R25 Y.n6 Y.n4 135.249
R26 Y.n6 Y.n5 98.982
R27 Y.n8 Y.n7 98.982
R28 Y.n10 Y.n9 98.982
R29 Y.n12 Y.n11 98.982
R30 Y.n14 Y.n13 98.982
R31 Y.n15 Y.n3 95.6388
R32 Y.n12 Y.n10 73.2449
R33 Y.n15 Y.n14 48.0005
R34 Y.n8 Y.n6 36.2672
R35 Y.n10 Y.n8 36.2672
R36 Y.n14 Y.n12 36.2672
R37 Y.n0 Y.t12 26.5955
R38 Y.n0 Y.t13 26.5955
R39 Y.n1 Y.t10 26.5955
R40 Y.n1 Y.t11 26.5955
R41 Y.n3 Y.t15 24.9236
R42 Y.n3 Y.t14 24.9236
R43 Y.n4 Y.t19 24.9236
R44 Y.n4 Y.t6 24.9236
R45 Y.n5 Y.t0 24.9236
R46 Y.n5 Y.t1 24.9236
R47 Y.n7 Y.t5 24.9236
R48 Y.n7 Y.t3 24.9236
R49 Y.n9 Y.t4 24.9236
R50 Y.n9 Y.t2 24.9236
R51 Y.n11 Y.t18 24.9236
R52 Y.n11 Y.t8 24.9236
R53 Y.n13 Y.t9 24.9236
R54 Y.n13 Y.t7 24.9236
R55 Y.n2 Y.t16 24.9236
R56 Y.n2 Y.t17 24.9236
R57 Y.n17 Y.n16 23.2234
R58 Y Y.n18 8.37536
R59 Y.n16 Y.n15 3.55606
R60 Y.n18 Y.n17 2.92621
R61 VGND.n15 VGND.t13 286.426
R62 VGND.n12 VGND.n11 207.965
R63 VGND.n21 VGND.n10 207.965
R64 VGND.n8 VGND.n7 207.965
R65 VGND.n37 VGND.n4 207.965
R66 VGND.n40 VGND.n39 207.965
R67 VGND.n46 VGND.n1 207.965
R68 VGND.n31 VGND.n30 185
R69 VGND.n29 VGND.n28 185
R70 VGND.n14 VGND.t2 162.111
R71 VGND.n48 VGND.t7 160.8
R72 VGND.n30 VGND.n29 96.0005
R73 VGND.n17 VGND.n16 34.6358
R74 VGND.n23 VGND.n22 34.6358
R75 VGND.n27 VGND.n26 34.6358
R76 VGND.n36 VGND.n5 34.6358
R77 VGND.n41 VGND.n38 34.6358
R78 VGND.n45 VGND.n2 34.6358
R79 VGND.n20 VGND.n12 33.8829
R80 VGND.n48 VGND.n47 32.377
R81 VGND.n47 VGND.n46 30.8711
R82 VGND.n21 VGND.n20 29.3652
R83 VGND.n16 VGND.n15 27.8593
R84 VGND.n29 VGND.t9 24.9236
R85 VGND.n30 VGND.t5 24.9236
R86 VGND.n11 VGND.t14 24.9236
R87 VGND.n11 VGND.t12 24.9236
R88 VGND.n10 VGND.t11 24.9236
R89 VGND.n10 VGND.t10 24.9236
R90 VGND.n7 VGND.t8 24.9236
R91 VGND.n7 VGND.t15 24.9236
R92 VGND.n4 VGND.t3 24.9236
R93 VGND.n4 VGND.t6 24.9236
R94 VGND.n39 VGND.t4 24.9236
R95 VGND.n39 VGND.t0 24.9236
R96 VGND.n1 VGND.t1 24.9236
R97 VGND.n1 VGND.t16 24.9236
R98 VGND.n40 VGND.n2 24.8476
R99 VGND.n23 VGND.n8 23.3417
R100 VGND.n38 VGND.n37 18.824
R101 VGND.n37 VGND.n36 15.8123
R102 VGND.n15 VGND.n14 13.9879
R103 VGND.n28 VGND.n27 12.6181
R104 VGND.n49 VGND.n48 11.5593
R105 VGND.n26 VGND.n8 11.2946
R106 VGND.n41 VGND.n40 9.78874
R107 VGND.n47 VGND.n0 9.3005
R108 VGND.n45 VGND.n44 9.3005
R109 VGND.n43 VGND.n2 9.3005
R110 VGND.n42 VGND.n41 9.3005
R111 VGND.n38 VGND.n3 9.3005
R112 VGND.n36 VGND.n35 9.3005
R113 VGND.n34 VGND.n5 9.3005
R114 VGND.n33 VGND.n32 9.3005
R115 VGND.n27 VGND.n6 9.3005
R116 VGND.n26 VGND.n25 9.3005
R117 VGND.n24 VGND.n23 9.3005
R118 VGND.n22 VGND.n9 9.3005
R119 VGND.n20 VGND.n19 9.3005
R120 VGND.n18 VGND.n17 9.3005
R121 VGND.n16 VGND.n13 9.3005
R122 VGND.n31 VGND.n5 8.1005
R123 VGND.n32 VGND.n31 5.8005
R124 VGND.n22 VGND.n21 5.27109
R125 VGND.n32 VGND.n28 4.6005
R126 VGND.n46 VGND.n45 3.76521
R127 VGND.n17 VGND.n12 0.753441
R128 VGND.n14 VGND.n13 0.523738
R129 VGND.n18 VGND.n13 0.120292
R130 VGND.n19 VGND.n18 0.120292
R131 VGND.n19 VGND.n9 0.120292
R132 VGND.n24 VGND.n9 0.120292
R133 VGND.n25 VGND.n24 0.120292
R134 VGND.n25 VGND.n6 0.120292
R135 VGND.n33 VGND.n6 0.120292
R136 VGND.n34 VGND.n33 0.120292
R137 VGND.n35 VGND.n34 0.120292
R138 VGND.n35 VGND.n3 0.120292
R139 VGND.n42 VGND.n3 0.120292
R140 VGND.n43 VGND.n42 0.120292
R141 VGND.n44 VGND.n43 0.120292
R142 VGND.n44 VGND.n0 0.120292
R143 VGND.n49 VGND.n0 0.120292
R144 VGND VGND.n49 0.0226354
R145 VNB.t13 VNB.t2 2677.02
R146 VNB.t5 VNB.t9 2677.02
R147 VNB.t14 VNB.t13 1196.12
R148 VNB.t12 VNB.t14 1196.12
R149 VNB.t11 VNB.t12 1196.12
R150 VNB.t10 VNB.t11 1196.12
R151 VNB.t8 VNB.t10 1196.12
R152 VNB.t15 VNB.t8 1196.12
R153 VNB.t9 VNB.t15 1196.12
R154 VNB.t3 VNB.t5 1196.12
R155 VNB.t6 VNB.t3 1196.12
R156 VNB.t4 VNB.t6 1196.12
R157 VNB.t0 VNB.t4 1196.12
R158 VNB.t1 VNB.t0 1196.12
R159 VNB.t16 VNB.t1 1196.12
R160 VNB.t7 VNB.t16 1196.12
R161 VNB VNB.t7 925.567
R162 D_N.n0 D_N.t1 231.718
R163 D_N.n0 D_N.t0 159.417
R164 D_N D_N.n0 152.833
R165 a_1191_21.t0 a_1191_21.n7 267.118
R166 a_1191_21.n0 a_1191_21.t2 212.081
R167 a_1191_21.n4 a_1191_21.t3 212.081
R168 a_1191_21.n2 a_1191_21.t4 212.081
R169 a_1191_21.n1 a_1191_21.t5 212.081
R170 a_1191_21.n7 a_1191_21.n0 190.707
R171 a_1191_21.n6 a_1191_21.n3 172.725
R172 a_1191_21.n7 a_1191_21.t1 169.643
R173 a_1191_21.n6 a_1191_21.n5 152
R174 a_1191_21.n0 a_1191_21.t8 139.78
R175 a_1191_21.n4 a_1191_21.t9 139.78
R176 a_1191_21.n2 a_1191_21.t7 139.78
R177 a_1191_21.n1 a_1191_21.t6 139.78
R178 a_1191_21.n2 a_1191_21.n1 61.346
R179 a_1191_21.n3 a_1191_21.n2 51.1217
R180 a_1191_21.n5 a_1191_21.n4 39.4369
R181 a_1191_21.n7 a_1191_21.n6 25.2957
R182 a_1191_21.n5 a_1191_21.n0 21.9096
R183 a_1191_21.n4 a_1191_21.n3 10.2247
R184 a_803_297.n4 a_803_297.t7 371.904
R185 a_803_297.n1 a_803_297.t1 371.904
R186 a_803_297.n1 a_803_297.n0 300.885
R187 a_803_297.n5 a_803_297.n4 300.885
R188 a_803_297.n3 a_803_297.n2 208.508
R189 a_803_297.n3 a_803_297.n1 44.424
R190 a_803_297.n4 a_803_297.n3 44.424
R191 a_803_297.n0 a_803_297.t0 26.5955
R192 a_803_297.n0 a_803_297.t2 26.5955
R193 a_803_297.n2 a_803_297.t4 26.5955
R194 a_803_297.n2 a_803_297.t3 26.5955
R195 a_803_297.t6 a_803_297.n5 26.5955
R196 a_803_297.n5 a_803_297.t5 26.5955
R197 VPB.t13 VPB.t9 556.386
R198 VPB.t4 VPB.t1 556.386
R199 VPB.t12 VPB.t13 248.599
R200 VPB.t11 VPB.t12 248.599
R201 VPB.t10 VPB.t11 248.599
R202 VPB.t7 VPB.t10 248.599
R203 VPB.t0 VPB.t7 248.599
R204 VPB.t6 VPB.t0 248.599
R205 VPB.t1 VPB.t6 248.599
R206 VPB.t3 VPB.t4 248.599
R207 VPB.t2 VPB.t3 248.599
R208 VPB.t5 VPB.t2 248.599
R209 VPB.t15 VPB.t5 248.599
R210 VPB.t16 VPB.t15 248.599
R211 VPB.t14 VPB.t16 248.599
R212 VPB.t8 VPB.t14 248.599
R213 VPB VPB.t8 192.369
R214 a_27_297.n4 a_27_297.t2 371.904
R215 a_27_297.n5 a_27_297.n4 300.885
R216 a_27_297.n1 a_27_297.t4 273.675
R217 a_27_297.n1 a_27_297.n0 208.507
R218 a_27_297.n3 a_27_297.n2 187.506
R219 a_27_297.n3 a_27_297.n1 65.4262
R220 a_27_297.n4 a_27_297.n3 65.4258
R221 a_27_297.n2 a_27_297.t3 26.5955
R222 a_27_297.n2 a_27_297.t6 26.5955
R223 a_27_297.n0 a_27_297.t7 26.5955
R224 a_27_297.n0 a_27_297.t5 26.5955
R225 a_27_297.n5 a_27_297.t1 26.5955
R226 a_27_297.t0 a_27_297.n5 26.5955
R227 a_445_297.n5 a_445_297.n4 345.31
R228 a_445_297.n2 a_445_297.n0 345.308
R229 a_445_297.n2 a_445_297.n1 300.885
R230 a_445_297.n4 a_445_297.n3 300.885
R231 a_445_297.n4 a_445_297.n2 83.577
R232 a_445_297.n0 a_445_297.t7 26.5955
R233 a_445_297.n0 a_445_297.t0 26.5955
R234 a_445_297.n1 a_445_297.t6 26.5955
R235 a_445_297.n1 a_445_297.t1 26.5955
R236 a_445_297.n3 a_445_297.t4 26.5955
R237 a_445_297.n3 a_445_297.t3 26.5955
R238 a_445_297.n5 a_445_297.t2 26.5955
R239 a_445_297.t5 a_445_297.n5 26.5955
R240 A.n3 A.t0 212.081
R241 A.n5 A.t1 212.081
R242 A.n7 A.t2 212.081
R243 A.n1 A.t6 212.081
R244 A.n4 A.n0 172.725
R245 A.n9 A.n2 172.725
R246 A.n6 A.n0 152
R247 A.n9 A.n8 152
R248 A.n3 A.t4 139.78
R249 A.n5 A.t5 139.78
R250 A.n7 A.t3 139.78
R251 A.n1 A.t7 139.78
R252 A.n8 A.n6 49.6611
R253 A.n7 A.n2 48.2005
R254 A.n5 A.n4 39.4369
R255 A.n4 A.n3 21.9096
R256 A.n2 A.n1 13.146
R257 A A.n0 11.5815
R258 A.n6 A.n5 10.2247
R259 A A.n9 9.14336
R260 A.n8 A.n7 1.46111
R261 VPWR.n6 VPWR.n1 323.192
R262 VPWR.n4 VPWR.n3 318.293
R263 VPWR.n2 VPWR.t0 263.466
R264 VPWR.n1 VPWR.t2 26.5955
R265 VPWR.n1 VPWR.t1 26.5955
R266 VPWR.n3 VPWR.t4 26.5955
R267 VPWR.n3 VPWR.t3 26.5955
R268 VPWR.n6 VPWR.n5 25.977
R269 VPWR.n5 VPWR.n4 18.4476
R270 VPWR.n5 VPWR.n0 9.3005
R271 VPWR.n4 VPWR.n2 7.50979
R272 VPWR.n7 VPWR.n6 7.4049
R273 VPWR.n2 VPWR.n0 0.148605
R274 VPWR.n7 VPWR.n0 0.144904
R275 VPWR VPWR.n7 0.118504
R276 C.n2 C.t4 212.081
R277 C.n1 C.t5 212.081
R278 C.n7 C.t6 212.081
R279 C.n8 C.t7 212.081
R280 C.n4 C.n3 172.725
R281 C C.n9 170.895
R282 C.n5 C.n4 152
R283 C.n6 C.n0 152
R284 C.n2 C.t2 139.78
R285 C.n1 C.t0 139.78
R286 C.n7 C.t3 139.78
R287 C.n8 C.t1 139.78
R288 C.n6 C.n5 49.6611
R289 C.n9 C.n7 48.2005
R290 C.n3 C.n1 39.4369
R291 C.n3 C.n2 21.9096
R292 C.n4 C.n0 20.7243
R293 C.n9 C.n8 13.146
R294 C.n5 C.n1 10.2247
R295 C C.n0 1.82907
R296 C.n7 C.n6 1.46111
C0 Y A 0.166251f
C1 VPWR B 0.032132f
C2 VPB B 0.121375f
C3 Y B 0.204158f
C4 A B 0.064024f
C5 VGND C 0.054186f
C6 VGND D_N 0.048609f
C7 VGND VPWR 0.169623f
C8 VGND VPB 0.015088f
C9 VGND Y 1.08712f
C10 VGND A 0.064884f
C11 C VPWR 0.032374f
C12 C VPB 0.121447f
C13 D_N VPWR 0.047566f
C14 VGND B 0.049943f
C15 C Y 0.219574f
C16 D_N VPB 0.044114f
C17 VPWR VPB 0.174995f
C18 C B 0.033119f
C19 VPWR Y 0.026955f
C20 VPWR A 0.081878f
C21 Y VPB 0.010986f
C22 VPB A 0.119082f
C23 VGND VNB 1.00837f
C24 Y VNB 0.033645f
C25 VPWR VNB 0.821893f
C26 D_N VNB 0.151275f
C27 C VNB 0.366554f
C28 B VNB 0.366269f
C29 A VNB 0.389209f
C30 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4bb_1 VNB VPB VGND VPWR A Y B D_N C_N
X0 Y.t3 B.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND.t3 a_27_410.t2 Y.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t0 C_N.t0 a_27_410.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND.t2 A.t0 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t1 C_N.t1 a_27_410.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_205_93.t1 D_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 VPWR.t2 A.t1 a_573_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_205_93.t0 D_N.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.1226 ps=1.32 w=0.42 l=0.15
X8 a_477_297.t0 a_27_410.t3 a_393_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X9 a_573_297.t0 B.t1 a_477_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X10 a_393_297.t1 a_205_93.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2559 ps=2.52 w=1 l=0.15
X11 Y.t4 a_205_93.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t1 241.536
R1 B.n0 B.t0 169.237
R2 B B.n0 163.055
R3 VGND.n8 VGND.t5 282.817
R4 VGND.n1 VGND.n0 228.294
R5 VGND.n4 VGND.n3 200.127
R6 VGND.n5 VGND.t2 156.573
R7 VGND.n0 VGND.t0 44.2862
R8 VGND.n0 VGND.t1 38.5719
R9 VGND.n9 VGND.n1 30.8711
R10 VGND.n3 VGND.t4 30.462
R11 VGND.n3 VGND.t3 30.462
R12 VGND.n9 VGND.n8 27.4829
R13 VGND.n7 VGND.n4 23.7181
R14 VGND.n8 VGND.n7 16.9417
R15 VGND.n11 VGND.n1 11.4238
R16 VGND.n10 VGND.n9 9.3005
R17 VGND.n8 VGND.n2 9.3005
R18 VGND.n7 VGND.n6 9.3005
R19 VGND.n5 VGND.n4 6.37884
R20 VGND.n6 VGND.n5 0.717338
R21 VGND.n11 VGND.n10 0.141672
R22 VGND VGND.n11 0.120476
R23 VGND.n6 VGND.n2 0.120292
R24 VGND.n10 VGND.n2 0.120292
R25 Y.n1 Y.t0 715.948
R26 Y.n1 Y.n0 195.24
R27 Y.n3 Y.n2 185
R28 Y.n3 Y.n1 73.657
R29 Y.n2 Y.t1 24.9236
R30 Y.n2 Y.t3 24.9236
R31 Y.n0 Y.t2 24.9236
R32 Y.n0 Y.t4 24.9236
R33 Y Y.n3 4.4805
R34 VNB.t1 VNB.t5 2677.02
R35 VNB.t3 VNB.t4 1366.99
R36 VNB.t0 VNB.t1 1253.07
R37 VNB.t4 VNB.t2 1196.12
R38 VNB.t5 VNB.t3 1196.12
R39 VNB VNB.t0 1025.24
R40 a_27_410.t0 a_27_410.n1 663.83
R41 a_27_410.n1 a_27_410.n0 397.623
R42 a_27_410.n1 a_27_410.t1 312.135
R43 a_27_410.n0 a_27_410.t3 241.536
R44 a_27_410.n0 a_27_410.t2 169.237
R45 C_N.n0 C_N.t1 329.902
R46 C_N.n1 C_N.n0 152
R47 C_N.n0 C_N.t0 132.282
R48 C_N.n1 C_N 10.4234
R49 C_N C_N.n1 2.01193
R50 A.n0 A.t1 235.821
R51 A.n0 A.t0 163.52
R52 A A.n0 153.173
R53 VPWR.n1 VPWR.n0 606.069
R54 VPWR.n1 VPWR.t2 344.702
R55 VPWR.n0 VPWR.t0 327.592
R56 VPWR.n0 VPWR.t1 63.3219
R57 VPWR VPWR.n1 0.147188
R58 VPB.t1 VPB.t0 553.428
R59 VPB.t3 VPB.t1 287.072
R60 VPB.t2 VPB.t4 284.113
R61 VPB.t4 VPB.t5 248.599
R62 VPB.t0 VPB.t2 248.599
R63 VPB VPB.t3 189.409
R64 D_N D_N.n0 154.429
R65 D_N.n0 D_N.t1 142.994
R66 D_N.n0 D_N.t0 126.927
R67 a_205_93.n2 a_205_93.n1 636.506
R68 a_205_93.n1 a_205_93.t1 268.209
R69 a_205_93.n0 a_205_93.t2 227.987
R70 a_205_93.n0 a_205_93.t3 155.686
R71 a_205_93.n1 a_205_93.n0 152
R72 a_205_93.n3 a_205_93.n2 54.0789
R73 a_205_93.n2 a_205_93.t0 33.4876
R74 a_573_297.t0 a_573_297.t1 53.1905
R75 a_393_297.t0 a_393_297.t1 53.1905
R76 a_477_297.t0 a_477_297.t1 65.0105
C0 C_N A 6.47e-20
C1 VPB C_N 0.092841f
C2 B A 0.117062f
C3 C_N VPWR 0.020742f
C4 Y C_N 8.35e-19
C5 VPB B 0.030423f
C6 B VPWR 0.093333f
C7 D_N C_N 0.081621f
C8 Y B 0.045178f
C9 VPB A 0.037187f
C10 A VPWR 0.05703f
C11 VGND C_N 0.031388f
C12 Y A 0.003062f
C13 D_N B 7.23e-20
C14 VPB VPWR 0.087631f
C15 Y VPB 0.00728f
C16 VGND B 0.019341f
C17 Y VPWR 0.016454f
C18 D_N VPB 0.039097f
C19 D_N VPWR 0.004144f
C20 VGND A 0.056936f
C21 Y D_N 0.001204f
C22 VGND VPB 0.008641f
C23 VGND VPWR 0.073703f
C24 Y VGND 0.208773f
C25 D_N VGND 0.01804f
C26 C_N B 2.57e-19
C27 VGND VNB 0.487444f
C28 D_N VNB 0.100723f
C29 Y VNB 0.0187f
C30 VPWR VNB 0.391341f
C31 A VNB 0.151061f
C32 B VNB 0.094788f
C33 C_N VNB 0.135087f
C34 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4bb_2 VNB VPB VGND VPWR Y B A D_N C_N
X0 Y.t3 a_27_410.t2 a_336_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t0 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_336_297.t2 a_201_93.t2 a_418_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y.t6 a_201_93.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X4 Y.t4 a_27_410.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t8 B.t0 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_418_297.t1 a_201_93.t4 a_336_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t9 D_N.t0 a_27_410.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR.t3 D_N.t1 a_27_410.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND.t5 A.t1 Y.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t8 B.t1 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_776_297.t3 A.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X12 a_201_93.t1 C_N.t0 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1226 ps=1.32 w=0.42 l=0.15
X13 a_201_93.t0 C_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VPWR.t1 A.t3 a_776_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_776_297.t1 B.t2 a_418_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t4 a_201_93.t5 Y.t7 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_336_297.t0 a_27_410.t4 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 a_418_297.t3 B.t3 a_776_297.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 VGND.t1 a_27_410.t5 Y.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_27_410.t0 a_27_410.n3 664.076
R1 a_27_410.n3 a_27_410.t1 313.127
R2 a_27_410.n3 a_27_410.n2 292.978
R3 a_27_410.n0 a_27_410.t4 212.081
R4 a_27_410.n1 a_27_410.t2 212.081
R5 a_27_410.n0 a_27_410.t5 139.78
R6 a_27_410.n1 a_27_410.t3 139.78
R7 a_27_410.n2 a_27_410.n0 28.0981
R8 a_27_410.n2 a_27_410.n1 26.6803
R9 a_336_297.n1 a_336_297.t3 886.899
R10 a_336_297.t0 a_336_297.n1 866.682
R11 a_336_297.n1 a_336_297.n0 585
R12 a_336_297.n0 a_336_297.t1 26.5955
R13 a_336_297.n0 a_336_297.t2 26.5955
R14 Y Y.n7 599.769
R15 Y.n5 Y.n3 135.249
R16 Y.n2 Y.n0 135.249
R17 Y.n5 Y.n4 98.982
R18 Y.n2 Y.n1 98.982
R19 Y Y.n6 33.5009
R20 Y.n7 Y.t2 26.5955
R21 Y.n7 Y.t3 26.5955
R22 Y.n3 Y.t1 24.9236
R23 Y.n3 Y.t0 24.9236
R24 Y.n4 Y.t9 24.9236
R25 Y.n4 Y.t8 24.9236
R26 Y.n0 Y.t7 24.9236
R27 Y.n0 Y.t6 24.9236
R28 Y.n1 Y.t5 24.9236
R29 Y.n1 Y.t4 24.9236
R30 Y.n6 Y.n2 24.5338
R31 Y.n6 Y.n5 20.2672
R32 VPB.t8 VPB.t6 627.414
R33 VPB.t2 VPB.t9 568.225
R34 VPB.t7 VPB.t8 287.072
R35 VPB.t0 VPB.t1 248.599
R36 VPB.t5 VPB.t0 248.599
R37 VPB.t9 VPB.t5 248.599
R38 VPB.t3 VPB.t2 248.599
R39 VPB.t4 VPB.t3 248.599
R40 VPB.t6 VPB.t4 248.599
R41 VPB VPB.t7 192.369
R42 A.n0 A.t2 212.081
R43 A.n1 A.t3 212.081
R44 A A.n2 157.761
R45 A.n0 A.t1 139.78
R46 A.n1 A.t0 139.78
R47 A.n2 A.n1 32.1338
R48 A.n2 A.n0 29.2126
R49 VGND.n15 VGND.t1 263.462
R50 VGND.n5 VGND.t7 257.858
R51 VGND.n24 VGND.t3 239.821
R52 VGND.n1 VGND.n0 228.294
R53 VGND.n9 VGND.n7 207.965
R54 VGND.n18 VGND.n17 207.965
R55 VGND.n8 VGND.t5 156.958
R56 VGND.n0 VGND.t0 38.5719
R57 VGND.n0 VGND.t9 38.5719
R58 VGND.n9 VGND.n8 37.305
R59 VGND.n11 VGND.n10 34.6358
R60 VGND.n23 VGND.n3 34.6358
R61 VGND.n25 VGND.n1 32.377
R62 VGND.n19 VGND.n16 31.8711
R63 VGND.n25 VGND.n24 30.8711
R64 VGND.n19 VGND.n18 25.977
R65 VGND.n7 VGND.t6 24.9236
R66 VGND.n7 VGND.t8 24.9236
R67 VGND.n17 VGND.t2 24.9236
R68 VGND.n17 VGND.t4 24.9236
R69 VGND.n11 VGND.n5 21.277
R70 VGND.n24 VGND.n23 13.5534
R71 VGND.n27 VGND.n1 9.91792
R72 VGND.n26 VGND.n25 9.3005
R73 VGND.n24 VGND.n2 9.3005
R74 VGND.n23 VGND.n22 9.3005
R75 VGND.n21 VGND.n3 9.3005
R76 VGND.n20 VGND.n19 9.3005
R77 VGND.n16 VGND.n4 9.3005
R78 VGND.n14 VGND.n13 9.3005
R79 VGND.n12 VGND.n11 9.3005
R80 VGND.n10 VGND.n6 9.3005
R81 VGND.n18 VGND.n3 8.65932
R82 VGND.n15 VGND.n14 8.5005
R83 VGND.n10 VGND.n9 2.63579
R84 VGND.n14 VGND.n5 2.3005
R85 VGND.n8 VGND.n6 2.13159
R86 VGND.n16 VGND.n15 0.7005
R87 VGND.n27 VGND.n26 0.141672
R88 VGND VGND.n27 0.121778
R89 VGND.n12 VGND.n6 0.120292
R90 VGND.n13 VGND.n12 0.120292
R91 VGND.n13 VGND.n4 0.120292
R92 VGND.n20 VGND.n4 0.120292
R93 VGND.n21 VGND.n20 0.120292
R94 VGND.n22 VGND.n21 0.120292
R95 VGND.n22 VGND.n2 0.120292
R96 VGND.n26 VGND.n2 0.120292
R97 VNB.t0 VNB.t3 3089.97
R98 VNB.t1 VNB.t7 2733.98
R99 VNB.t6 VNB.t5 1196.12
R100 VNB.t8 VNB.t6 1196.12
R101 VNB.t7 VNB.t8 1196.12
R102 VNB.t2 VNB.t1 1196.12
R103 VNB.t4 VNB.t2 1196.12
R104 VNB.t3 VNB.t4 1196.12
R105 VNB.t9 VNB.t0 1196.12
R106 VNB VNB.t9 1039.48
R107 a_201_93.n3 a_201_93.t1 691.299
R108 a_201_93.t0 a_201_93.n3 264.221
R109 a_201_93.n0 a_201_93.t2 212.081
R110 a_201_93.n1 a_201_93.t4 212.081
R111 a_201_93.n0 a_201_93.t5 139.78
R112 a_201_93.n1 a_201_93.t3 139.78
R113 a_201_93.n3 a_201_93.n2 109.812
R114 a_201_93.n2 a_201_93.n0 45.0371
R115 a_201_93.n2 a_201_93.n1 13.8297
R116 a_418_297.n1 a_418_297.n0 1038.95
R117 a_418_297.n0 a_418_297.t0 26.5955
R118 a_418_297.n0 a_418_297.t3 26.5955
R119 a_418_297.t2 a_418_297.n1 26.5955
R120 a_418_297.n1 a_418_297.t1 26.5955
R121 B.n0 B.t2 212.081
R122 B.n1 B.t3 212.081
R123 B B.n2 163.201
R124 B.n0 B.t1 139.78
R125 B.n1 B.t0 139.78
R126 B.n2 B.n1 32.8641
R127 B.n2 B.n0 28.4823
R128 D_N.n0 D_N.t1 329.902
R129 D_N D_N.n0 153.829
R130 D_N.n0 D_N.t0 132.282
R131 VPWR.n2 VPWR.n1 606.071
R132 VPWR.n2 VPWR.n0 330.416
R133 VPWR.n1 VPWR.t2 327.592
R134 VPWR.n1 VPWR.t3 63.3219
R135 VPWR.n0 VPWR.t0 26.5955
R136 VPWR.n0 VPWR.t1 26.5955
R137 VPWR VPWR.n2 0.148043
R138 a_776_297.n0 a_776_297.t0 867.038
R139 a_776_297.n0 a_776_297.t3 297.284
R140 a_776_297.n1 a_776_297.n0 186.993
R141 a_776_297.n1 a_776_297.t2 26.5955
R142 a_776_297.t1 a_776_297.n1 26.5955
R143 C_N C_N.n0 154.47
R144 C_N.n0 C_N.t0 141.946
R145 C_N.n0 C_N.t1 125.879
C0 C_N D_N 0.084106f
C1 C_N Y 3.39e-19
C2 Y D_N 2.43e-19
C3 C_N VGND 0.017548f
C4 VGND D_N 0.030376f
C5 Y B 0.125788f
C6 Y VGND 0.564951f
C7 Y A 0.055312f
C8 C_N VPWR 0.004164f
C9 VGND B 0.030025f
C10 B A 0.070229f
C11 D_N VPWR 0.020821f
C12 Y VPWR 0.014551f
C13 VGND A 0.059935f
C14 B VPWR 0.017248f
C15 C_N VPB 0.040702f
C16 D_N VPB 0.09413f
C17 VGND VPWR 0.11679f
C18 A VPWR 0.038741f
C19 Y VPB 0.012857f
C20 B VPB 0.057558f
C21 VGND VPB 0.012598f
C22 A VPB 0.056715f
C23 VPWR VPB 0.132033f
C24 VGND VNB 0.729348f
C25 Y VNB 0.037208f
C26 C_N VNB 0.105364f
C27 VPWR VNB 0.560323f
C28 A VNB 0.206969f
C29 B VNB 0.18064f
C30 D_N VNB 0.133196f
C31 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4bb_4 VNB VPB VGND VPWR D_N A B C_N Y
X0 Y.t4 B.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_729_297.t7 k.t2 a_311_297.t7 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t3 B.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t19 A.t0 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_197_47.t1 D_N.t0 VPWR.t5 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 a_311_297.t6 k.t3 a_729_297.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t17 A.t1 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_729_297.t1 B.t2 a_1087_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t10 a_197_47.t2 Y.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t11 a_197_47.t3 Y.t10 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_729_297.t5 k.t4 a_311_297.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_1087_297.t2 B.t3 a_729_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t6 k.t5 Y.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_197_47.t0 D_N.t1 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t7 k.t6 Y.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t5 C_N.t0 k.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X16 a_729_297.t3 B.t4 a_1087_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VGND.t16 A.t2 Y.t18 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t0 A.t3 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_1087_297.t7 A.t4 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X20 Y.t7 k.t7 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t8 k.t8 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t3 A.t5 a_1087_297.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t0 C_N.t1 k.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X24 a_311_297.t0 a_197_47.t4 Y.t11 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t12 a_197_47.t5 a_311_297.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 a_1087_297.t5 A.t6 VPWR.t2 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR.t1 A.t7 a_1087_297.t4 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_311_297.t2 a_197_47.t6 Y.t13 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_1087_297.t0 B.t5 a_729_297.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND.t2 B.t6 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 Y.t14 a_197_47.t7 a_311_297.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 VGND.t1 B.t7 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 Y.t15 a_197_47.t8 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X34 a_311_297.t4 k.t9 a_729_297.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X35 Y.t16 a_197_47.t9 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B.n2 B.t5 212.081
R1 B.n1 B.t2 212.081
R2 B.n7 B.t3 212.081
R3 B.n8 B.t4 212.081
R4 B.n4 B.n3 172.725
R5 B B.n9 164.19
R6 B.n5 B.n4 152
R7 B.n6 B.n0 152
R8 B.n2 B.t7 139.78
R9 B.n1 B.t1 139.78
R10 B.n7 B.t6 139.78
R11 B.n8 B.t0 139.78
R12 B.n6 B.n5 49.6611
R13 B.n3 B.n1 48.2005
R14 B.n9 B.n7 39.4369
R15 B.n9 B.n8 21.9096
R16 B.n4 B.n0 20.7243
R17 B.n3 B.n2 13.146
R18 B.n7 B.n6 10.2247
R19 B B.n0 8.53383
R20 B.n5 B.n1 1.46111
R21 VGND.n48 VGND.t12 286.426
R22 VGND.n15 VGND.n14 207.965
R23 VGND.n20 VGND.n12 207.965
R24 VGND.n23 VGND.n22 207.965
R25 VGND.n36 VGND.n35 207.965
R26 VGND.n42 VGND.n6 207.965
R27 VGND.n4 VGND.n3 207.965
R28 VGND.n1 VGND.n0 207.965
R29 VGND.n33 VGND.n32 185
R30 VGND.n31 VGND.n30 185
R31 VGND.n16 VGND.t0 156.258
R32 VGND.n32 VGND.n31 96.0005
R33 VGND.n16 VGND.n15 37.6466
R34 VGND.n19 VGND.n13 34.6358
R35 VGND.n24 VGND.n21 34.6358
R36 VGND.n29 VGND.n10 34.6358
R37 VGND.n37 VGND.n34 34.6358
R38 VGND.n41 VGND.n7 34.6358
R39 VGND.n44 VGND.n43 34.6358
R40 VGND.n50 VGND.n49 34.6358
R41 VGND.n47 VGND.n4 33.8829
R42 VGND.n50 VGND.n1 33.8829
R43 VGND.n48 VGND.n47 29.3652
R44 VGND.n43 VGND.n42 27.8593
R45 VGND.n20 VGND.n19 26.3534
R46 VGND.n31 VGND.t4 24.9236
R47 VGND.n32 VGND.t7 24.9236
R48 VGND.n14 VGND.t15 24.9236
R49 VGND.n14 VGND.t16 24.9236
R50 VGND.n12 VGND.t17 24.9236
R51 VGND.n12 VGND.t1 24.9236
R52 VGND.n22 VGND.t3 24.9236
R53 VGND.n22 VGND.t2 24.9236
R54 VGND.n35 VGND.t9 24.9236
R55 VGND.n35 VGND.t6 24.9236
R56 VGND.n6 VGND.t8 24.9236
R57 VGND.n6 VGND.t11 24.9236
R58 VGND.n3 VGND.t13 24.9236
R59 VGND.n3 VGND.t10 24.9236
R60 VGND.n0 VGND.t14 24.9236
R61 VGND.n0 VGND.t5 24.9236
R62 VGND.n36 VGND.n7 21.8358
R63 VGND.n24 VGND.n23 20.3299
R64 VGND.n23 VGND.n10 14.3064
R65 VGND.n37 VGND.n36 12.8005
R66 VGND.n34 VGND.n33 11.1123
R67 VGND.n30 VGND.n29 9.60638
R68 VGND.n51 VGND.n50 9.3005
R69 VGND.n49 VGND.n2 9.3005
R70 VGND.n47 VGND.n46 9.3005
R71 VGND.n45 VGND.n44 9.3005
R72 VGND.n43 VGND.n5 9.3005
R73 VGND.n41 VGND.n40 9.3005
R74 VGND.n39 VGND.n7 9.3005
R75 VGND.n38 VGND.n37 9.3005
R76 VGND.n34 VGND.n8 9.3005
R77 VGND.n27 VGND.n9 9.3005
R78 VGND.n29 VGND.n28 9.3005
R79 VGND.n26 VGND.n10 9.3005
R80 VGND.n25 VGND.n24 9.3005
R81 VGND.n21 VGND.n11 9.3005
R82 VGND.n19 VGND.n18 9.3005
R83 VGND.n17 VGND.n13 9.3005
R84 VGND.n52 VGND.n1 8.41204
R85 VGND.n21 VGND.n20 8.28285
R86 VGND.n42 VGND.n41 6.77697
R87 VGND.n30 VGND.n9 5.4005
R88 VGND.n49 VGND.n48 5.27109
R89 VGND.n33 VGND.n9 5.0005
R90 VGND.n15 VGND.n13 2.25932
R91 VGND.n17 VGND.n16 2.14912
R92 VGND.n44 VGND.n4 0.753441
R93 VGND.n52 VGND.n51 0.141672
R94 VGND VGND.n52 0.120476
R95 VGND.n18 VGND.n17 0.120292
R96 VGND.n18 VGND.n11 0.120292
R97 VGND.n25 VGND.n11 0.120292
R98 VGND.n26 VGND.n25 0.120292
R99 VGND.n28 VGND.n26 0.120292
R100 VGND.n28 VGND.n27 0.120292
R101 VGND.n27 VGND.n8 0.120292
R102 VGND.n38 VGND.n8 0.120292
R103 VGND.n39 VGND.n38 0.120292
R104 VGND.n40 VGND.n39 0.120292
R105 VGND.n40 VGND.n5 0.120292
R106 VGND.n45 VGND.n5 0.120292
R107 VGND.n46 VGND.n45 0.120292
R108 VGND.n46 VGND.n2 0.120292
R109 VGND.n51 VGND.n2 0.120292
R110 Y Y.n17 620.311
R111 Y.n16 Y.n15 585
R112 Y.n13 Y.n12 146.982
R113 Y.n2 Y.n0 135.249
R114 Y.n2 Y.n1 98.982
R115 Y.n4 Y.n3 98.982
R116 Y.n6 Y.n5 98.982
R117 Y.n8 Y.n7 98.982
R118 Y.n10 Y.n9 98.982
R119 Y.n13 Y.n11 95.6388
R120 Y.n8 Y.n6 73.2449
R121 Y.n16 Y.n14 45.4626
R122 Y.n14 Y.n10 36.6227
R123 Y.n4 Y.n2 36.2672
R124 Y.n6 Y.n4 36.2672
R125 Y.n10 Y.n8 36.2672
R126 Y.n17 Y.t13 26.5955
R127 Y.n17 Y.t14 26.5955
R128 Y.n15 Y.t11 26.5955
R129 Y.n15 Y.t12 26.5955
R130 Y.n11 Y.t10 24.9236
R131 Y.n11 Y.t16 24.9236
R132 Y.n12 Y.t9 24.9236
R133 Y.n12 Y.t15 24.9236
R134 Y.n0 Y.t0 24.9236
R135 Y.n0 Y.t17 24.9236
R136 Y.n1 Y.t18 24.9236
R137 Y.n1 Y.t19 24.9236
R138 Y.n3 Y.t1 24.9236
R139 Y.n3 Y.t3 24.9236
R140 Y.n5 Y.t2 24.9236
R141 Y.n5 Y.t4 24.9236
R142 Y.n7 Y.t6 24.9236
R143 Y.n7 Y.t8 24.9236
R144 Y.n9 Y.t5 24.9236
R145 Y.n9 Y.t7 24.9236
R146 Y.n14 Y.n13 11.3783
R147 Y Y.n16 1.76602
R148 VNB.t14 VNB.t12 2790.94
R149 VNB.t7 VNB.t4 2677.02
R150 VNB.t15 VNB.t0 1196.12
R151 VNB.t16 VNB.t15 1196.12
R152 VNB.t17 VNB.t16 1196.12
R153 VNB.t1 VNB.t17 1196.12
R154 VNB.t3 VNB.t1 1196.12
R155 VNB.t2 VNB.t3 1196.12
R156 VNB.t4 VNB.t2 1196.12
R157 VNB.t9 VNB.t7 1196.12
R158 VNB.t6 VNB.t9 1196.12
R159 VNB.t8 VNB.t6 1196.12
R160 VNB.t11 VNB.t8 1196.12
R161 VNB.t13 VNB.t11 1196.12
R162 VNB.t10 VNB.t13 1196.12
R163 VNB.t12 VNB.t10 1196.12
R164 VNB.t5 VNB.t14 1196.12
R165 VNB VNB.t5 968.285
R166 k.n11 k.n10 263.529
R167 k.n11 k.t0 233.565
R168 k.n2 k.t9 212.081
R169 k.n1 k.t2 212.081
R170 k.n7 k.t3 212.081
R171 k.n8 k.t4 212.081
R172 k.n4 k.n3 172.725
R173 k.n12 k.n11 166.532
R174 k.n10 k.n9 152
R175 k.n6 k.n0 152
R176 k.n5 k.n4 152
R177 k.n2 k.t6 139.78
R178 k.n1 k.t8 139.78
R179 k.n7 k.t5 139.78
R180 k.n8 k.t7 139.78
R181 k k.n12 64.6541
R182 k.n6 k.n5 49.6611
R183 k.n3 k.n1 48.2005
R184 k.n9 k.n7 39.4369
R185 k.n12 k.t1 36.2466
R186 k.n9 k.n8 21.9096
R187 k.n4 k.n0 20.7243
R188 k.n10 k.n0 20.7243
R189 k.n3 k.n2 13.146
R190 k.n7 k.n6 10.2247
R191 k.n5 k.n1 1.46111
R192 a_311_297.n3 a_311_297.t3 866.682
R193 a_311_297.n3 a_311_297.n2 585
R194 a_311_297.n5 a_311_297.n4 585
R195 a_311_297.n1 a_311_297.t4 371.012
R196 a_311_297.n1 a_311_297.n0 300.885
R197 a_311_297.n4 a_311_297.n1 49.8603
R198 a_311_297.n4 a_311_297.n3 43.0085
R199 a_311_297.n2 a_311_297.t1 26.5955
R200 a_311_297.n2 a_311_297.t2 26.5955
R201 a_311_297.n0 a_311_297.t7 26.5955
R202 a_311_297.n0 a_311_297.t6 26.5955
R203 a_311_297.n5 a_311_297.t5 26.5955
R204 a_311_297.t0 a_311_297.n5 26.5955
R205 a_729_297.n5 a_729_297.n4 346.892
R206 a_729_297.n2 a_729_297.n0 345.308
R207 a_729_297.n2 a_729_297.n1 300.885
R208 a_729_297.n4 a_729_297.n3 300.885
R209 a_729_297.n4 a_729_297.n2 83.577
R210 a_729_297.n0 a_729_297.t2 26.5955
R211 a_729_297.n0 a_729_297.t1 26.5955
R212 a_729_297.n1 a_729_297.t0 26.5955
R213 a_729_297.n1 a_729_297.t3 26.5955
R214 a_729_297.n3 a_729_297.t4 26.5955
R215 a_729_297.n3 a_729_297.t7 26.5955
R216 a_729_297.t6 a_729_297.n5 26.5955
R217 a_729_297.n5 a_729_297.t5 26.5955
R218 VPB.t15 VPB.t10 580.062
R219 VPB.t11 VPB.t2 556.386
R220 VPB.t5 VPB.t6 248.599
R221 VPB.t16 VPB.t5 248.599
R222 VPB.t17 VPB.t16 248.599
R223 VPB.t1 VPB.t17 248.599
R224 VPB.t4 VPB.t1 248.599
R225 VPB.t3 VPB.t4 248.599
R226 VPB.t2 VPB.t3 248.599
R227 VPB.t14 VPB.t11 248.599
R228 VPB.t13 VPB.t14 248.599
R229 VPB.t12 VPB.t13 248.599
R230 VPB.t7 VPB.t12 248.599
R231 VPB.t8 VPB.t7 248.599
R232 VPB.t9 VPB.t8 248.599
R233 VPB.t10 VPB.t9 248.599
R234 VPB.t0 VPB.t15 248.599
R235 VPB VPB.t0 201.246
R236 A.n3 A.t4 212.081
R237 A.n5 A.t5 212.081
R238 A.n7 A.t6 212.081
R239 A.n1 A.t7 212.081
R240 A.n4 A.n0 172.725
R241 A.n9 A.n2 172.725
R242 A.n6 A.n0 152
R243 A.n9 A.n8 152
R244 A.n3 A.t3 139.78
R245 A.n5 A.t1 139.78
R246 A.n7 A.t2 139.78
R247 A.n1 A.t0 139.78
R248 A.n8 A.n6 49.6611
R249 A.n5 A.n4 48.2005
R250 A.n7 A.n2 39.4369
R251 A.n2 A.n1 21.9096
R252 A A.n0 19.5053
R253 A.n4 A.n3 13.146
R254 A.n8 A.n7 10.2247
R255 A.n6 A.n5 1.46111
R256 A A.n9 1.21955
R257 D_N.n0 D_N.t0 229.754
R258 D_N.n0 D_N.t1 157.453
R259 D_N D_N.n0 154.071
R260 VPWR.n33 VPWR.n1 601.292
R261 VPWR.n11 VPWR.n10 323.993
R262 VPWR.n9 VPWR.n8 318.293
R263 VPWR.n14 VPWR.n13 34.6358
R264 VPWR.n15 VPWR.n14 34.6358
R265 VPWR.n15 VPWR.n6 34.6358
R266 VPWR.n19 VPWR.n6 34.6358
R267 VPWR.n20 VPWR.n19 34.6358
R268 VPWR.n21 VPWR.n20 34.6358
R269 VPWR.n21 VPWR.n4 34.6358
R270 VPWR.n25 VPWR.n4 34.6358
R271 VPWR.n26 VPWR.n25 34.6358
R272 VPWR.n27 VPWR.n26 34.6358
R273 VPWR.n27 VPWR.n2 34.6358
R274 VPWR.n31 VPWR.n2 34.6358
R275 VPWR.n32 VPWR.n31 34.6358
R276 VPWR.n13 VPWR.n9 30.4946
R277 VPWR.n1 VPWR.t5 26.5955
R278 VPWR.n1 VPWR.t0 26.5955
R279 VPWR.n8 VPWR.t2 26.5955
R280 VPWR.n8 VPWR.t1 26.5955
R281 VPWR.n10 VPWR.t4 26.5955
R282 VPWR.n10 VPWR.t3 26.5955
R283 VPWR.n33 VPWR.n32 21.4593
R284 VPWR.n13 VPWR.n12 9.3005
R285 VPWR.n14 VPWR.n7 9.3005
R286 VPWR.n16 VPWR.n15 9.3005
R287 VPWR.n17 VPWR.n6 9.3005
R288 VPWR.n19 VPWR.n18 9.3005
R289 VPWR.n20 VPWR.n5 9.3005
R290 VPWR.n22 VPWR.n21 9.3005
R291 VPWR.n23 VPWR.n4 9.3005
R292 VPWR.n25 VPWR.n24 9.3005
R293 VPWR.n26 VPWR.n3 9.3005
R294 VPWR.n28 VPWR.n27 9.3005
R295 VPWR.n29 VPWR.n2 9.3005
R296 VPWR.n31 VPWR.n30 9.3005
R297 VPWR.n32 VPWR.n0 9.3005
R298 VPWR.n34 VPWR.n33 7.1994
R299 VPWR.n11 VPWR.n9 6.47684
R300 VPWR.n12 VPWR.n11 0.58037
R301 VPWR.n34 VPWR.n0 0.147518
R302 VPWR.n12 VPWR.n7 0.120292
R303 VPWR.n16 VPWR.n7 0.120292
R304 VPWR.n17 VPWR.n16 0.120292
R305 VPWR.n18 VPWR.n17 0.120292
R306 VPWR.n18 VPWR.n5 0.120292
R307 VPWR.n22 VPWR.n5 0.120292
R308 VPWR.n23 VPWR.n22 0.120292
R309 VPWR.n24 VPWR.n23 0.120292
R310 VPWR.n24 VPWR.n3 0.120292
R311 VPWR.n28 VPWR.n3 0.120292
R312 VPWR.n29 VPWR.n28 0.120292
R313 VPWR.n30 VPWR.n29 0.120292
R314 VPWR.n30 VPWR.n0 0.120292
R315 VPWR VPWR.n34 0.114555
R316 a_197_47.t1 a_197_47.n7 896.015
R317 a_197_47.n0 a_197_47.t4 212.081
R318 a_197_47.n1 a_197_47.t5 212.081
R319 a_197_47.n3 a_197_47.t6 212.081
R320 a_197_47.n4 a_197_47.t7 212.081
R321 a_197_47.n7 a_197_47.t0 171.192
R322 a_197_47.n6 a_197_47.n5 152
R323 a_197_47.n0 a_197_47.t3 139.78
R324 a_197_47.n1 a_197_47.t9 139.78
R325 a_197_47.n3 a_197_47.t2 139.78
R326 a_197_47.n4 a_197_47.t8 139.78
R327 a_197_47.n6 a_197_47.n2 96.7795
R328 a_197_47.n1 a_197_47.n0 61.346
R329 a_197_47.n5 a_197_47.n3 45.2793
R330 a_197_47.n7 a_197_47.n6 33.8829
R331 a_197_47.n2 a_197_47.n1 30.5591
R332 a_197_47.n3 a_197_47.n2 24.2858
R333 a_197_47.n5 a_197_47.n4 16.0672
R334 a_1087_297.n4 a_1087_297.t1 370.401
R335 a_1087_297.n5 a_1087_297.n4 300.885
R336 a_1087_297.n1 a_1087_297.t7 276.781
R337 a_1087_297.n1 a_1087_297.n0 208.507
R338 a_1087_297.n3 a_1087_297.n2 187.506
R339 a_1087_297.n3 a_1087_297.n1 65.4262
R340 a_1087_297.n4 a_1087_297.n3 65.4258
R341 a_1087_297.n2 a_1087_297.t4 26.5955
R342 a_1087_297.n2 a_1087_297.t0 26.5955
R343 a_1087_297.n0 a_1087_297.t6 26.5955
R344 a_1087_297.n0 a_1087_297.t5 26.5955
R345 a_1087_297.t3 a_1087_297.n5 26.5955
R346 a_1087_297.n5 a_1087_297.t2 26.5955
R347 C_N.n0 C_N.t1 231.017
R348 C_N.n0 C_N.t0 158.716
R349 C_N C_N.n0 157.738
C0 VGND Y 1.0875f
C1 C_N k 0.126555f
C2 VGND VPB 0.01358f
C3 VGND C_N 0.014688f
C4 VGND k 0.159986f
C5 B A 0.064024f
C6 D_N VPWR 0.016553f
C7 B VPWR 0.032923f
C8 VPB D_N 0.040151f
C9 B Y 0.226994f
C10 A VPWR 0.088736f
C11 C_N D_N 0.050963f
C12 VPB B 0.122175f
C13 A Y 0.166162f
C14 D_N k 0.047156f
C15 VPB A 0.12019f
C16 VPWR Y 0.022544f
C17 B k 0.033459f
C18 VGND D_N 0.018179f
C19 VPB VPWR 0.171238f
C20 A k 1.15e-19
C21 VGND B 0.051876f
C22 VPB Y 0.007542f
C23 C_N VPWR 0.015201f
C24 VPWR k 0.186643f
C25 VGND A 0.091482f
C26 Y k 0.376278f
C27 VPB C_N 0.037623f
C28 VGND VPWR 0.177025f
C29 VPB k 0.147127f
C30 VGND VNB 1.02631f
C31 Y VNB 0.032995f
C32 VPWR VNB 0.821363f
C33 A VNB 0.392851f
C34 B VNB 0.369498f
C35 D_N VNB 0.115085f
C36 C_N VNB 0.142861f
C37 VPB VNB 1.84511f
C38 k VNB 0.446549f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2a_1 VNB VPB VPWR VGND X A1_N A2_N B2 B1
X0 a_206_369.t0 A1_N.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369.t1 A2_N.t0 a_205_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND.t1 B2.t0 a_489_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369.t0 B2.t1 a_76_199.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47.t2 a_206_369.t3 a_76_199.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47.t1 B1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR.t3 A2_N.t1 a_206_369.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199.t1 a_206_369.t4 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47.t0 A1_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR.t2 a_76_199.t3 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR.t4 B1.t1 a_585_369.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND.t2 a_76_199.t4 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1_N.n0 A1_N.t0 264.029
R1 A1_N.n0 A1_N.t1 206.19
R2 A1_N A1_N.n0 155.52
R3 VPWR.n4 VPWR.t4 679.928
R4 VPWR.n8 VPWR.n1 642.188
R5 VPWR.n3 VPWR.n2 585
R6 VPWR.n2 VPWR.t1 135.268
R7 VPWR.n2 VPWR.t3 118.549
R8 VPWR.n1 VPWR.t0 96.1553
R9 VPWR.n7 VPWR.n6 34.6358
R10 VPWR.n1 VPWR.t2 32.7439
R11 VPWR.n8 VPWR.n7 22.9652
R12 VPWR.n6 VPWR.n3 12.3976
R13 VPWR.n4 VPWR.n3 10.9214
R14 VPWR.n6 VPWR.n5 9.3005
R15 VPWR.n7 VPWR.n0 9.3005
R16 VPWR.n9 VPWR.n8 7.12063
R17 VPWR.n5 VPWR.n4 0.226183
R18 VPWR.n9 VPWR.n0 0.148519
R19 VPWR.n5 VPWR.n0 0.120292
R20 VPWR VPWR.n9 0.11354
R21 a_206_369.n2 a_206_369.n1 787.759
R22 a_206_369.n1 a_206_369.t1 305.416
R23 a_206_369.n0 a_206_369.t3 292.413
R24 a_206_369.n1 a_206_369.n0 216.998
R25 a_206_369.n0 a_206_369.t4 120.431
R26 a_206_369.n2 a_206_369.t2 93.81
R27 a_206_369.t0 a_206_369.n2 93.81
R28 VPB.t3 VPB.t5 517.913
R29 VPB.t0 VPB.t3 325.546
R30 VPB.t1 VPB.t0 287.072
R31 VPB.t5 VPB.t2 278.193
R32 VPB.t2 VPB.t4 213.084
R33 VPB VPB.t1 189.409
R34 A2_N.n0 A2_N.t1 334.298
R35 A2_N A2_N.n0 190.923
R36 A2_N.n0 A2_N.t0 131.857
R37 a_205_47.t0 a_205_47.t1 90.0005
R38 VNB.t1 VNB.t5 2719.74
R39 VNB.t3 VNB.t0 1366.99
R40 VNB.t0 VNB.t1 1324.27
R41 VNB.t2 VNB.t4 1196.12
R42 VNB.t5 VNB.t2 1196.12
R43 VNB VNB.t3 911.327
R44 B2.n0 B2.t1 264.029
R45 B2.n0 B2.t0 206.19
R46 B2 B2.n0 171.018
R47 a_489_47.n0 a_489_47.t1 476.041
R48 a_489_47.t0 a_489_47.n0 38.5719
R49 a_489_47.n0 a_489_47.t2 38.5719
R50 VGND.n2 VGND.n0 225.345
R51 VGND.n2 VGND.n1 215.535
R52 VGND.n0 VGND.t0 48.5719
R53 VGND.n1 VGND.t3 38.5719
R54 VGND.n1 VGND.t1 38.5719
R55 VGND.n0 VGND.t2 33.0774
R56 VGND VGND.n2 0.151861
R57 a_76_199.n2 a_76_199.n1 588.051
R58 a_76_199.n1 a_76_199.n0 319.154
R59 a_76_199.n1 a_76_199.t2 303.993
R60 a_76_199.n0 a_76_199.t3 241.536
R61 a_76_199.n0 a_76_199.t4 169.237
R62 a_76_199.t0 a_76_199.n2 86.7743
R63 a_76_199.n2 a_76_199.t1 63.3219
R64 a_585_369.t0 a_585_369.t1 98.5005
R65 B1.n0 B1.t1 252.649
R66 B1.n0 B1.t0 194.809
R67 B1 B1.n0 154.042
R68 X X.n0 593.615
R69 X.n1 X.n0 585
R70 X.n1 X.t1 217.732
R71 X.n0 X.t0 26.5955
R72 X X.n1 8.12358
C0 B2 VGND 0.016247f
C1 A1_N VPB 0.062218f
C2 VPWR A2_N 0.009748f
C3 B1 VGND 0.016305f
C4 A2_N VPB 0.053423f
C5 A1_N A2_N 0.09394f
C6 B2 VPWR 0.088044f
C7 B2 VPB 0.055976f
C8 B1 VPWR 0.048982f
C9 VGND X 0.086091f
C10 B1 VPB 0.06625f
C11 VGND VPWR 0.072388f
C12 VGND VPB 0.009258f
C13 VGND A1_N 0.027491f
C14 VGND A2_N 0.064685f
C15 X VPWR 0.061845f
C16 X VPB 0.010949f
C17 X A1_N 0.003606f
C18 B2 B1 0.162675f
C19 VPWR VPB 0.108864f
C20 X A2_N 0.006853f
C21 VPWR A1_N 0.010805f
C22 VGND VNB 0.452597f
C23 B1 VNB 0.181469f
C24 B2 VNB 0.105231f
C25 A2_N VNB 0.125702f
C26 A1_N VNB 0.121561f
C27 VPWR VNB 0.391659f
C28 X VNB 0.094468f
C29 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2a_2 VNB VPB VGND VPWR B1 B2 A2_N X A1_N
X0 a_294_47.t0 A1_N.t0 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X1 VPWR.t4 A2_N.t0 a_295_369.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.2272 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X2 VPWR.t1 B1.t0 a_665_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND.t1 a_84_21.t3 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X.t2 a_84_21.t4 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_581_47.t2 a_295_369.t3 a_84_21.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR.t0 a_84_21.t5 X.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X7 a_665_369.t0 B2.t0 a_84_21.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X8 VGND.t0 B2.t1 a_581_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_295_369.t1 A2_N.t1 a_294_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X10 X.t0 a_84_21.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X11 a_84_21.t1 a_295_369.t4 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.2272 ps=1.35 w=0.64 l=0.15
X12 a_295_369.t0 A1_N.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.335 w=0.64 l=0.15
X13 a_581_47.t1 B1.t1 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 A1_N.n0 A1_N.t1 299.377
R1 A1_N.n0 A1_N.t0 206.19
R2 A1_N A1_N.n0 156.8
R3 VGND.n4 VGND.n1 218.13
R4 VGND.n3 VGND.n2 215.517
R5 VGND.n6 VGND.t2 151.131
R6 VGND.n1 VGND.t3 48.5719
R7 VGND.n2 VGND.t4 38.5719
R8 VGND.n2 VGND.t0 38.5719
R9 VGND.n5 VGND.n4 34.6358
R10 VGND.n1 VGND.t1 33.0774
R11 VGND.n6 VGND.n5 24.4711
R12 VGND.n7 VGND.n6 9.3005
R13 VGND.n5 VGND.n0 9.3005
R14 VGND.n4 VGND.n3 7.5997
R15 VGND.n3 VGND.n0 0.148605
R16 VGND.n7 VGND.n0 0.120292
R17 VGND VGND.n7 0.0252396
R18 a_294_47.t0 a_294_47.t1 90.0005
R19 VNB.t4 VNB.t5 2762.46
R20 VNB.t1 VNB.t3 1366.99
R21 VNB.t3 VNB.t4 1324.27
R22 VNB.t0 VNB.t6 1196.12
R23 VNB.t5 VNB.t0 1196.12
R24 VNB.t2 VNB.t1 1196.12
R25 VNB VNB.t2 1025.24
R26 A2_N.n0 A2_N.t0 369.644
R27 A2_N A2_N.n0 192.357
R28 A2_N.n0 A2_N.t1 131.857
R29 a_295_369.n2 a_295_369.n1 788.78
R30 a_295_369.n1 a_295_369.t1 306.836
R31 a_295_369.n0 a_295_369.t3 295.336
R32 a_295_369.n1 a_295_369.n0 215.536
R33 a_295_369.n0 a_295_369.t4 154.24
R34 a_295_369.n2 a_295_369.t2 61.563
R35 a_295_369.t0 a_295_369.n2 61.563
R36 VPWR.n10 VPWR.n2 600.515
R37 VPWR.n5 VPWR.n4 585
R38 VPWR.n6 VPWR.t1 383.014
R39 VPWR.n12 VPWR.t2 252.894
R40 VPWR.n4 VPWR.t5 113.891
R41 VPWR.n4 VPWR.t4 104.656
R42 VPWR.n2 VPWR.t3 61.563
R43 VPWR.n9 VPWR.n3 34.6358
R44 VPWR.n2 VPWR.t0 30.5947
R45 VPWR.n12 VPWR.n11 24.4711
R46 VPWR.n10 VPWR.n9 24.0946
R47 VPWR.n11 VPWR.n10 20.3299
R48 VPWR.n5 VPWR.n3 11.3805
R49 VPWR.n6 VPWR.n5 11.1689
R50 VPWR.n7 VPWR.n3 9.3005
R51 VPWR.n9 VPWR.n8 9.3005
R52 VPWR.n10 VPWR.n1 9.3005
R53 VPWR.n11 VPWR.n0 9.3005
R54 VPWR.n13 VPWR.n12 9.3005
R55 VPWR.n7 VPWR.n6 0.221987
R56 VPWR.n8 VPWR.n7 0.120292
R57 VPWR.n8 VPWR.n1 0.120292
R58 VPWR.n1 VPWR.n0 0.120292
R59 VPWR.n13 VPWR.n0 0.120292
R60 VPWR VPWR.n13 0.0252396
R61 VPB.t4 VPB.t6 509.034
R62 VPB.t3 VPB.t4 325.546
R63 VPB.t0 VPB.t3 287.072
R64 VPB.t6 VPB.t5 260.437
R65 VPB.t5 VPB.t1 248.599
R66 VPB.t2 VPB.t0 248.599
R67 VPB VPB.t2 213.084
R68 B1.n0 B1.t0 288.416
R69 B1.n0 B1.t1 195.23
R70 B1 B1.n0 154.042
R71 a_665_369.t0 a_665_369.t1 83.1099
R72 a_84_21.n2 a_84_21.n1 326.103
R73 a_84_21.n2 a_84_21.t2 304.502
R74 a_84_21.n3 a_84_21.n2 296.087
R75 a_84_21.n1 a_84_21.t5 212.081
R76 a_84_21.n0 a_84_21.t6 212.081
R77 a_84_21.n1 a_84_21.t3 139.78
R78 a_84_21.n0 a_84_21.t4 139.78
R79 a_84_21.n1 a_84_21.n0 61.346
R80 a_84_21.t0 a_84_21.n3 47.7114
R81 a_84_21.n3 a_84_21.t1 41.5552
R82 X X.n0 593.784
R83 X.n2 X.n0 585
R84 X.n2 X.n1 181.351
R85 X.n0 X.t1 26.5955
R86 X.n0 X.t0 26.5955
R87 X.n1 X.t3 24.9236
R88 X.n1 X.t2 24.9236
R89 X X.n2 8.28285
R90 a_581_47.n0 a_581_47.t1 479.365
R91 a_581_47.t0 a_581_47.n0 38.5719
R92 a_581_47.n0 a_581_47.t2 38.5719
R93 B2.n0 B2.t0 299.377
R94 B2.n0 B2.t1 206.19
R95 B2 B2.n0 170.763
C0 VPWR A1_N 0.017618f
C1 A1_N A2_N 0.09574f
C2 X A1_N 0.003177f
C3 VPWR A2_N 0.015999f
C4 VPWR X 0.149714f
C5 X A2_N 0.006845f
C6 VPWR B2 0.084063f
C7 VGND A1_N 0.027973f
C8 VPWR VGND 0.096397f
C9 A1_N VPB 0.059833f
C10 VPWR VPB 0.100824f
C11 VPWR B1 0.052593f
C12 VGND A2_N 0.064792f
C13 X VGND 0.140484f
C14 A2_N VPB 0.051951f
C15 X VPB 0.003689f
C16 VGND B2 0.016971f
C17 B2 VPB 0.052524f
C18 VGND VPB 0.00924f
C19 B2 B1 0.150852f
C20 VGND B1 0.016331f
C21 B1 VPB 0.066689f
C22 VGND VNB 0.530409f
C23 X VNB 0.023471f
C24 VPWR VNB 0.468225f
C25 B1 VNB 0.181888f
C26 B2 VNB 0.106585f
C27 A2_N VNB 0.12764f
C28 A1_N VNB 0.119854f
C29 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2a_4 VNB VPB VGND VPWR B1 B2 A2_N A1_N X
X0 a_27_47.t4 a_415_21.t6 a_193_297.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR.t2 A2_N.t0 a_415_21.t5 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_415_21.t4 A1_N.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3 a_415_21.t1 A2_N.t1 a_717_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_193_297.t3 a_415_21.t7 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t5 B1.t0 a_109_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t9 a_193_297.t6 X.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t4 a_193_297.t7 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_109_297.t2 B2.t0 a_193_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t2 a_193_297.t8 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_717_47.t3 A1_N.t1 VGND.t5 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_717_47.t0 A2_N.t2 a_415_21.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t7 a_193_297.t9 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_193_297.t1 B2.t1 a_109_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_47.t2 B2.t2 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_27_47.t0 B1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t7 a_193_297.t10 X.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t4 A1_N.t2 a_717_47.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t6 a_193_297.t11 X.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VGND.t0 B2.t3 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_193_297.t4 a_415_21.t8 a_27_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR.t11 a_193_297.t12 X.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t6 a_415_21.t9 a_193_297.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X23 X.t0 a_193_297.t13 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t0 A1_N.t3 a_415_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_109_297.t0 B1.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_415_21.t3 A2_N.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VGND.t1 B1.t3 a_27_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_415_21.n5 a_415_21.n4 585
R1 a_415_21.n6 a_415_21.n5 347.803
R2 a_415_21.n3 a_415_21.n2 275.387
R3 a_415_21.n1 a_415_21.t9 212.081
R4 a_415_21.n0 a_415_21.t7 212.081
R5 a_415_21.n3 a_415_21.n1 195.85
R6 a_415_21.n1 a_415_21.t6 139.78
R7 a_415_21.n0 a_415_21.t8 139.78
R8 a_415_21.n5 a_415_21.n3 84.8748
R9 a_415_21.n1 a_415_21.n0 61.346
R10 a_415_21.n4 a_415_21.t5 26.5955
R11 a_415_21.n4 a_415_21.t4 26.5955
R12 a_415_21.t0 a_415_21.n6 26.5955
R13 a_415_21.n6 a_415_21.t3 26.5955
R14 a_415_21.n2 a_415_21.t2 24.9236
R15 a_415_21.n2 a_415_21.t1 24.9236
R16 a_193_297.n13 a_193_297.n12 655.164
R17 a_193_297.n12 a_193_297.n0 222.315
R18 a_193_297.n11 a_193_297.n1 216.793
R19 a_193_297.n3 a_193_297.t6 212.081
R20 a_193_297.n5 a_193_297.t8 212.081
R21 a_193_297.n7 a_193_297.t12 212.081
R22 a_193_297.n8 a_193_297.t13 212.081
R23 a_193_297.n4 a_193_297.n2 177.601
R24 a_193_297.n10 a_193_297.n9 152
R25 a_193_297.n6 a_193_297.n2 152
R26 a_193_297.n3 a_193_297.t11 139.78
R27 a_193_297.n5 a_193_297.t9 139.78
R28 a_193_297.n7 a_193_297.t10 139.78
R29 a_193_297.n8 a_193_297.t7 139.78
R30 a_193_297.n9 a_193_297.n8 49.6611
R31 a_193_297.n11 a_193_297.n10 42.9594
R32 a_193_297.n7 a_193_297.n6 37.9763
R33 a_193_297.n4 a_193_297.n3 35.055
R34 a_193_297.n0 a_193_297.t2 26.5955
R35 a_193_297.n0 a_193_297.t3 26.5955
R36 a_193_297.t0 a_193_297.n13 26.5955
R37 a_193_297.n13 a_193_297.t1 26.5955
R38 a_193_297.n5 a_193_297.n4 26.2914
R39 a_193_297.n10 a_193_297.n2 25.6005
R40 a_193_297.n1 a_193_297.t5 24.9236
R41 a_193_297.n1 a_193_297.t4 24.9236
R42 a_193_297.n6 a_193_297.n5 23.3702
R43 a_193_297.n9 a_193_297.n7 11.6853
R44 a_193_297.n12 a_193_297.n11 5.66716
R45 a_27_47.t4 a_27_47.n3 316.983
R46 a_27_47.n1 a_27_47.t5 174.512
R47 a_27_47.n1 a_27_47.n0 98.982
R48 a_27_47.n3 a_27_47.n2 88.3446
R49 a_27_47.n3 a_27_47.n1 51.5158
R50 a_27_47.n2 a_27_47.t3 24.9236
R51 a_27_47.n2 a_27_47.t0 24.9236
R52 a_27_47.n0 a_27_47.t1 24.9236
R53 a_27_47.n0 a_27_47.t2 24.9236
R54 VNB.t8 VNB.t0 2677.02
R55 VNB.t11 VNB.t9 1196.12
R56 VNB.t10 VNB.t11 1196.12
R57 VNB.t12 VNB.t10 1196.12
R58 VNB.t1 VNB.t12 1196.12
R59 VNB.t5 VNB.t1 1196.12
R60 VNB.t4 VNB.t5 1196.12
R61 VNB.t0 VNB.t4 1196.12
R62 VNB.t7 VNB.t8 1196.12
R63 VNB.t2 VNB.t7 1196.12
R64 VNB.t3 VNB.t2 1196.12
R65 VNB.t6 VNB.t3 1196.12
R66 VNB.t13 VNB.t6 1196.12
R67 VNB VNB.t13 925.567
R68 A2_N.n0 A2_N.t3 212.081
R69 A2_N.n1 A2_N.t0 212.081
R70 A2_N A2_N.n2 171.201
R71 A2_N.n0 A2_N.t2 139.78
R72 A2_N.n1 A2_N.t1 139.78
R73 A2_N.n2 A2_N.n1 31.4035
R74 A2_N.n2 A2_N.n0 29.9429
R75 VPWR.n28 VPWR.n27 606.505
R76 VPWR.n15 VPWR.n14 606.505
R77 VPWR.n8 VPWR.n7 604.968
R78 VPWR.n25 VPWR.n24 585
R79 VPWR.n23 VPWR.n22 585
R80 VPWR.n35 VPWR.t3 350.533
R81 VPWR.n9 VPWR.t9 349.051
R82 VPWR.n12 VPWR.n6 318.293
R83 VPWR.n24 VPWR.n23 102.441
R84 VPWR.n33 VPWR.n1 34.6358
R85 VPWR.n34 VPWR.n33 34.6358
R86 VPWR.n29 VPWR.n26 34.6358
R87 VPWR.n21 VPWR.n4 34.6358
R88 VPWR.n16 VPWR.n13 34.6358
R89 VPWR.n11 VPWR.n8 30.4946
R90 VPWR.n23 VPWR.t4 26.5955
R91 VPWR.n24 VPWR.t6 26.5955
R92 VPWR.n27 VPWR.t7 26.5955
R93 VPWR.n27 VPWR.t5 26.5955
R94 VPWR.n14 VPWR.t1 26.5955
R95 VPWR.n14 VPWR.t2 26.5955
R96 VPWR.n6 VPWR.t10 26.5955
R97 VPWR.n6 VPWR.t0 26.5955
R98 VPWR.n7 VPWR.t8 26.5955
R99 VPWR.n7 VPWR.t11 26.5955
R100 VPWR.n35 VPWR.n34 25.977
R101 VPWR.n28 VPWR.n1 15.4358
R102 VPWR.n26 VPWR.n25 14.0479
R103 VPWR.n12 VPWR.n11 13.9299
R104 VPWR.n11 VPWR.n10 9.3005
R105 VPWR.n13 VPWR.n5 9.3005
R106 VPWR.n17 VPWR.n16 9.3005
R107 VPWR.n18 VPWR.n4 9.3005
R108 VPWR.n21 VPWR.n20 9.3005
R109 VPWR.n19 VPWR.n3 9.3005
R110 VPWR.n26 VPWR.n2 9.3005
R111 VPWR.n30 VPWR.n29 9.3005
R112 VPWR.n31 VPWR.n1 9.3005
R113 VPWR.n33 VPWR.n32 9.3005
R114 VPWR.n34 VPWR.n0 9.3005
R115 VPWR.n36 VPWR.n35 9.3005
R116 VPWR.n15 VPWR.n4 7.90638
R117 VPWR.n16 VPWR.n15 7.90638
R118 VPWR.n9 VPWR.n8 6.47684
R119 VPWR.n22 VPWR.n3 5.92289
R120 VPWR.n22 VPWR.n21 4.27091
R121 VPWR.n25 VPWR.n3 4.01244
R122 VPWR.n13 VPWR.n12 1.88285
R123 VPWR.n10 VPWR.n9 0.58037
R124 VPWR.n29 VPWR.n28 0.376971
R125 VPWR.n10 VPWR.n5 0.120292
R126 VPWR.n17 VPWR.n5 0.120292
R127 VPWR.n18 VPWR.n17 0.120292
R128 VPWR.n20 VPWR.n18 0.120292
R129 VPWR.n20 VPWR.n19 0.120292
R130 VPWR.n19 VPWR.n2 0.120292
R131 VPWR.n30 VPWR.n2 0.120292
R132 VPWR.n31 VPWR.n30 0.120292
R133 VPWR.n32 VPWR.n31 0.120292
R134 VPWR.n32 VPWR.n0 0.120292
R135 VPWR.n36 VPWR.n0 0.120292
R136 VPWR VPWR.n36 0.0226354
R137 VPB.t8 VPB.t4 556.386
R138 VPB.t12 VPB.t13 248.599
R139 VPB.t11 VPB.t12 248.599
R140 VPB.t10 VPB.t11 248.599
R141 VPB.t0 VPB.t10 248.599
R142 VPB.t1 VPB.t0 248.599
R143 VPB.t2 VPB.t1 248.599
R144 VPB.t4 VPB.t2 248.599
R145 VPB.t9 VPB.t8 248.599
R146 VPB.t6 VPB.t9 248.599
R147 VPB.t5 VPB.t6 248.599
R148 VPB.t7 VPB.t5 248.599
R149 VPB.t3 VPB.t7 248.599
R150 VPB VPB.t3 192.369
R151 A1_N.n2 A1_N.n0 251.79
R152 A1_N.n1 A1_N.t3 241.536
R153 A1_N.n0 A1_N.t0 236.18
R154 A1_N.n1 A1_N.t2 169.237
R155 A1_N.n0 A1_N.t1 163.881
R156 A1_N.n2 A1_N.n1 152
R157 A1_N A1_N.n2 1.95606
R158 a_717_47.n1 a_717_47.n0 338.505
R159 a_717_47.n0 a_717_47.t2 24.9236
R160 a_717_47.n0 a_717_47.t0 24.9236
R161 a_717_47.t1 a_717_47.n1 24.9236
R162 a_717_47.n1 a_717_47.t3 24.9236
R163 B1.n2 B1.n0 244.804
R164 B1.n1 B1.t2 241.536
R165 B1.n0 B1.t0 241.536
R166 B1.n1 B1.t3 169.237
R167 B1.n0 B1.t1 169.237
R168 B1.n2 B1.n1 152
R169 B1 B1.n2 6.28198
R170 a_109_297.n1 a_109_297.n0 935.014
R171 a_109_297.n0 a_109_297.t3 26.5955
R172 a_109_297.n0 a_109_297.t0 26.5955
R173 a_109_297.t1 a_109_297.n1 26.5955
R174 a_109_297.n1 a_109_297.t2 26.5955
R175 X.n2 X.n0 350.113
R176 X.n2 X.n1 196.083
R177 X.n5 X.n3 135.249
R178 X.n5 X.n4 98.982
R179 X X.n5 40.6621
R180 X X.n2 29.2575
R181 X.n1 X.t3 26.5955
R182 X.n1 X.t2 26.5955
R183 X.n0 X.t1 26.5955
R184 X.n0 X.t0 26.5955
R185 X.n3 X.t6 24.9236
R186 X.n3 X.t4 24.9236
R187 X.n4 X.t5 24.9236
R188 X.n4 X.t7 24.9236
R189 VGND.n10 VGND.t6 292.029
R190 VGND.n21 VGND.t5 286.426
R191 VGND.n11 VGND.n9 207.965
R192 VGND.n3 VGND.n2 207.965
R193 VGND.n33 VGND.n1 207.965
R194 VGND.n14 VGND.n13 121.451
R195 VGND.n34 VGND.n33 43.1829
R196 VGND.n11 VGND.n10 35.4566
R197 VGND.n15 VGND.n12 34.6358
R198 VGND.n19 VGND.n7 34.6358
R199 VGND.n20 VGND.n19 34.6358
R200 VGND.n22 VGND.n20 34.6358
R201 VGND.n26 VGND.n5 34.6358
R202 VGND.n27 VGND.n26 34.6358
R203 VGND.n28 VGND.n27 34.6358
R204 VGND.n32 VGND.n31 34.6358
R205 VGND.n31 VGND.n3 27.8593
R206 VGND.n9 VGND.t8 24.9236
R207 VGND.n9 VGND.t7 24.9236
R208 VGND.n13 VGND.t9 24.9236
R209 VGND.n13 VGND.t4 24.9236
R210 VGND.n2 VGND.t2 24.9236
R211 VGND.n2 VGND.t0 24.9236
R212 VGND.n1 VGND.t3 24.9236
R213 VGND.n1 VGND.t1 24.9236
R214 VGND.n15 VGND.n14 23.3417
R215 VGND.n21 VGND.n5 23.3417
R216 VGND.n14 VGND.n7 11.2946
R217 VGND.n22 VGND.n21 11.2946
R218 VGND.n12 VGND.n8 9.3005
R219 VGND.n16 VGND.n15 9.3005
R220 VGND.n17 VGND.n7 9.3005
R221 VGND.n19 VGND.n18 9.3005
R222 VGND.n20 VGND.n6 9.3005
R223 VGND.n23 VGND.n22 9.3005
R224 VGND.n24 VGND.n5 9.3005
R225 VGND.n26 VGND.n25 9.3005
R226 VGND.n27 VGND.n4 9.3005
R227 VGND.n29 VGND.n28 9.3005
R228 VGND.n31 VGND.n30 9.3005
R229 VGND.n32 VGND.n0 9.3005
R230 VGND.n28 VGND.n3 6.77697
R231 VGND.n12 VGND.n11 5.27109
R232 VGND.n10 VGND.n8 1.65809
R233 VGND.n33 VGND.n32 0.753441
R234 VGND.n16 VGND.n8 0.120292
R235 VGND.n17 VGND.n16 0.120292
R236 VGND.n18 VGND.n17 0.120292
R237 VGND.n18 VGND.n6 0.120292
R238 VGND.n23 VGND.n6 0.120292
R239 VGND.n24 VGND.n23 0.120292
R240 VGND.n25 VGND.n24 0.120292
R241 VGND.n25 VGND.n4 0.120292
R242 VGND.n29 VGND.n4 0.120292
R243 VGND.n30 VGND.n29 0.120292
R244 VGND.n30 VGND.n0 0.120292
R245 VGND.n34 VGND.n0 0.120292
R246 VGND VGND.n34 0.0226354
R247 B2.n0 B2.t0 212.081
R248 B2.n1 B2.t1 212.081
R249 B2 B2.n2 153.304
R250 B2.n0 B2.t3 139.78
R251 B2.n1 B2.t2 139.78
R252 B2.n2 B2.n0 30.6732
R253 B2.n2 B2.n1 30.6732
C0 B2 VPWR 0.017715f
C1 A1_N A2_N 0.216681f
C2 B2 VGND 0.028174f
C3 A1_N X 6.19e-19
C4 B2 VPB 0.051071f
C5 A1_N VPWR 0.052809f
C6 A1_N VGND 0.035115f
C7 A2_N X 4.44e-19
C8 A1_N VPB 0.066849f
C9 B2 B1 0.203357f
C10 A2_N VPWR 0.024497f
C11 A2_N VGND 0.01609f
C12 VPWR X 0.310545f
C13 X VGND 0.280222f
C14 X VPB 0.016547f
C15 A2_N VPB 0.051106f
C16 VPWR VGND 0.09406f
C17 VPWR VPB 0.161016f
C18 VGND VPB 0.013541f
C19 VPWR B1 0.067784f
C20 VGND B1 0.030689f
C21 VPB B1 0.066139f
C22 VGND VNB 0.842624f
C23 X VNB 0.058281f
C24 VPWR VNB 0.710313f
C25 A2_N VNB 0.166952f
C26 A1_N VNB 0.193617f
C27 B2 VNB 0.167862f
C28 B1 VNB 0.231381f
C29 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_1 VPB VNB VGND VPWR B1 B2 Y A2_N A1_N
X0 VPWR.t1 A2_N.t0 a_112_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=1.84 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t2 a_112_297.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.42 ps=1.84 w=1 l=0.15
X2 VGND.t1 B2.t0 a_394_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_112_297.t0 A2_N.t1 a_112_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.2405 pd=2.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 a_112_47.t0 A1_N.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17875 ps=1.85 w=0.65 l=0.15
X5 a_112_297.t2 A1_N.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X6 VPWR.t0 B1.t0 a_478_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X7 a_394_47.t2 a_112_297.t4 Y.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_394_47.t0 B1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_478_297.t1 B2.t1 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A2_N.n0 A2_N.t0 241.536
R1 A2_N.n0 A2_N.t1 169.237
R2 A2_N A2_N.n0 163.637
R3 a_112_297.n2 a_112_297.n1 368.839
R4 a_112_297.n1 a_112_297.n0 226.492
R5 a_112_297.n0 a_112_297.t3 212.081
R6 a_112_297.n1 a_112_297.t0 164.242
R7 a_112_297.n0 a_112_297.t4 139.78
R8 a_112_297.t1 a_112_297.n2 26.5955
R9 a_112_297.n2 a_112_297.t2 26.5955
R10 VPWR.n2 VPWR.n1 292.5
R11 VPWR.n4 VPWR.n3 292.5
R12 VPWR.n5 VPWR.t0 259.245
R13 VPWR.n9 VPWR.t3 251.999
R14 VPWR.n3 VPWR.n2 88.6505
R15 VPWR.n3 VPWR.t2 42.3555
R16 VPWR.n2 VPWR.t1 34.4755
R17 VPWR.n8 VPWR.n7 24.7001
R18 VPWR.n9 VPWR.n8 21.8358
R19 VPWR.n7 VPWR.n6 9.3005
R20 VPWR.n8 VPWR.n0 9.3005
R21 VPWR.n10 VPWR.n9 9.3005
R22 VPWR.n5 VPWR.n4 7.17539
R23 VPWR.n4 VPWR.n1 5.93864
R24 VPWR.n6 VPWR.n5 0.239865
R25 VPWR.n6 VPWR.n0 0.120292
R26 VPWR.n10 VPWR.n0 0.120292
R27 VPWR.n7 VPWR.n1 0.0664794
R28 VPWR VPWR.n10 0.0226354
R29 VPB.t2 VPB.t3 585.981
R30 VPB.t0 VPB.t1 248.599
R31 VPB.t3 VPB.t0 248.599
R32 VPB.t4 VPB.t2 248.599
R33 VPB VPB.t4 201.246
R34 Y.n1 Y.n0 585
R35 Y Y.n0 302.55
R36 Y.n1 Y.t1 290.217
R37 Y.n0 Y.t0 26.5955
R38 Y.n0 Y.t2 26.5955
R39 Y Y.n1 6.4005
R40 B2.n0 B2.t1 241.536
R41 B2 B2.n0 172.043
R42 B2.n0 B2.t0 169.237
R43 a_394_47.t0 a_394_47.n0 368.781
R44 a_394_47.n0 a_394_47.t1 24.9236
R45 a_394_47.n0 a_394_47.t2 24.9236
R46 VGND.n1 VGND.n0 215.239
R47 VGND.n1 VGND.t2 154.587
R48 VGND.n0 VGND.t0 24.9236
R49 VGND.n0 VGND.t1 24.9236
R50 VGND VGND.n1 0.0621188
R51 VNB.t3 VNB.t4 2990.29
R52 VNB.t1 VNB.t0 1196.12
R53 VNB.t4 VNB.t1 1196.12
R54 VNB.t2 VNB.t3 1025.24
R55 VNB VNB.t2 968.285
R56 a_112_47.t0 a_112_47.t1 38.7697
R57 A1_N.n0 A1_N.t1 229.56
R58 A1_N A1_N.n0 157.333
R59 A1_N.n0 A1_N.t0 157.26
R60 B1.n0 B1.t0 229.56
R61 B1.n0 B1.t1 157.26
R62 B1 B1.n0 154.012
R63 a_478_297.t0 a_478_297.t1 53.1905
C0 A1_N VPB 0.03925f
C1 Y A2_N 7.8e-19
C2 VPWR B2 0.109959f
C3 VGND A1_N 0.055337f
C4 A2_N VPB 0.031296f
C5 VPWR Y 0.126571f
C6 VPWR VPB 0.084563f
C7 VGND A2_N 0.087547f
C8 Y B2 0.131683f
C9 VPWR B1 0.053617f
C10 B2 VPB 0.029961f
C11 VPWR VGND 0.070693f
C12 Y VPB 0.004898f
C13 B2 B1 0.087918f
C14 VGND B2 0.016554f
C15 Y B1 8.74e-19
C16 B1 VPB 0.03925f
C17 Y VGND 0.028956f
C18 VGND VPB 0.006779f
C19 VGND B1 0.016182f
C20 A1_N A2_N 0.096243f
C21 VPWR A1_N 0.054618f
C22 VPWR A2_N 0.023606f
C23 VGND VNB 0.423292f
C24 Y VNB 0.010059f
C25 VPWR VNB 0.387462f
C26 B1 VNB 0.142474f
C27 B2 VNB 0.094838f
C28 A2_N VNB 0.101393f
C29 A1_N VNB 0.145115f
C30 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_2 VNB VPB VGND VPWR B2 Y A1_N B1 A2_N
X0 a_113_297.t5 A2_N.t0 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_113_47.t2 A2_N.t1 a_113_297.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t2 B1.t0 a_730_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t6 A2_N.t2 a_113_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_730_297.t1 B2.t0 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47.t1 B2.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_471_47.t5 B1.t1 VGND.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t0 B2.t2 a_730_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_113_297.t2 A2_N.t3 a_113_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_113_47.t0 A1_N.t0 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND.t5 A1_N.t1 a_113_47.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t2 B2.t3 a_471_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t4 a_113_297.t6 Y.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X13 a_113_297.t1 A1_N.t2 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 Y.t4 a_113_297.t7 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X15 a_730_297.t2 B1.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X16 Y.t3 a_113_297.t8 a_471_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1755 ps=1.84 w=0.65 l=0.15
X17 a_471_47.t2 a_113_297.t9 Y.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t0 A1_N.t3 a_113_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t4 B1.t3 a_471_47.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
R0 A2_N.n0 A2_N.t0 212.081
R1 A2_N.n1 A2_N.t2 212.081
R2 A2_N A2_N.n2 153.165
R3 A2_N.n0 A2_N.t1 139.78
R4 A2_N.n1 A2_N.t3 139.78
R5 A2_N.n2 A2_N.n0 31.4035
R6 A2_N.n2 A2_N.n1 29.9429
R7 VPWR.n18 VPWR.n2 606.505
R8 VPWR.n6 VPWR.n5 603.864
R9 VPWR.n11 VPWR.n3 585
R10 VPWR.n13 VPWR.n12 585
R11 VPWR.n7 VPWR.t2 360.856
R12 VPWR.n20 VPWR.t3 344.887
R13 VPWR.n12 VPWR.n11 104.41
R14 VPWR.n5 VPWR.t1 33.4905
R15 VPWR.n10 VPWR.n9 32.1073
R16 VPWR.n18 VPWR.n17 27.4829
R17 VPWR.n12 VPWR.t5 26.5955
R18 VPWR.n11 VPWR.t0 26.5955
R19 VPWR.n2 VPWR.t7 26.5955
R20 VPWR.n2 VPWR.t6 26.5955
R21 VPWR.n5 VPWR.t4 26.5955
R22 VPWR.n19 VPWR.n18 22.9652
R23 VPWR.n20 VPWR.n19 21.8358
R24 VPWR.n17 VPWR.n3 19.3297
R25 VPWR.n9 VPWR.n6 16.1887
R26 VPWR.n9 VPWR.n8 9.3005
R27 VPWR.n10 VPWR.n4 9.3005
R28 VPWR.n15 VPWR.n14 9.3005
R29 VPWR.n17 VPWR.n16 9.3005
R30 VPWR.n18 VPWR.n1 9.3005
R31 VPWR.n19 VPWR.n0 9.3005
R32 VPWR.n21 VPWR.n20 9.3005
R33 VPWR.n14 VPWR.n13 8.02438
R34 VPWR.n7 VPWR.n6 7.46771
R35 VPWR.n14 VPWR.n3 2.10199
R36 VPWR.n13 VPWR.n10 0.764679
R37 VPWR.n8 VPWR.n7 0.177017
R38 VPWR.n8 VPWR.n4 0.120292
R39 VPWR.n15 VPWR.n4 0.120292
R40 VPWR.n16 VPWR.n15 0.120292
R41 VPWR.n16 VPWR.n1 0.120292
R42 VPWR.n1 VPWR.n0 0.120292
R43 VPWR.n21 VPWR.n0 0.120292
R44 VPWR VPWR.n21 0.0213333
R45 a_113_297.n6 a_113_297.n5 585
R46 a_113_297.n5 a_113_297.n4 347.803
R47 a_113_297.n3 a_113_297.n0 269.558
R48 a_113_297.n1 a_113_297.t6 212.081
R49 a_113_297.n2 a_113_297.t7 212.081
R50 a_113_297.n3 a_113_297.n2 182.673
R51 a_113_297.n1 a_113_297.t9 139.78
R52 a_113_297.n2 a_113_297.t8 139.78
R53 a_113_297.n5 a_113_297.n3 81.9774
R54 a_113_297.n2 a_113_297.n1 61.346
R55 a_113_297.n4 a_113_297.t4 26.5955
R56 a_113_297.n4 a_113_297.t1 26.5955
R57 a_113_297.n6 a_113_297.t0 26.5955
R58 a_113_297.t5 a_113_297.n6 26.5955
R59 a_113_297.n0 a_113_297.t3 24.9236
R60 a_113_297.n0 a_113_297.t2 24.9236
R61 VPB.t1 VPB.t6 562.306
R62 VPB.t7 VPB.t2 269.315
R63 VPB.t3 VPB.t4 248.599
R64 VPB.t0 VPB.t3 248.599
R65 VPB.t2 VPB.t0 248.599
R66 VPB.t6 VPB.t7 248.599
R67 VPB.t9 VPB.t1 248.599
R68 VPB.t8 VPB.t9 248.599
R69 VPB.t5 VPB.t8 248.599
R70 VPB VPB.t5 201.246
R71 a_113_47.n1 a_113_47.n0 338.505
R72 a_113_47.n0 a_113_47.t1 24.9236
R73 a_113_47.n0 a_113_47.t0 24.9236
R74 a_113_47.n1 a_113_47.t3 24.9236
R75 a_113_47.t2 a_113_47.n1 24.9236
R76 VNB.t9 VNB.t6 2705.5
R77 VNB.t5 VNB.t2 1295.79
R78 VNB.t0 VNB.t1 1196.12
R79 VNB.t3 VNB.t0 1196.12
R80 VNB.t2 VNB.t3 1196.12
R81 VNB.t6 VNB.t5 1196.12
R82 VNB.t8 VNB.t9 1196.12
R83 VNB.t7 VNB.t8 1196.12
R84 VNB.t4 VNB.t7 1196.12
R85 VNB VNB.t4 968.285
R86 B1.n2 B1.n0 244.804
R87 B1.n1 B1.t0 241.536
R88 B1.n0 B1.t2 241.536
R89 B1.n1 B1.t1 169.237
R90 B1.n0 B1.t3 169.237
R91 B1.n2 B1.n1 152
R92 B1 B1.n2 7.34865
R93 a_730_297.n1 a_730_297.n0 935.015
R94 a_730_297.n0 a_730_297.t3 26.5955
R95 a_730_297.n0 a_730_297.t1 26.5955
R96 a_730_297.n1 a_730_297.t0 26.5955
R97 a_730_297.t2 a_730_297.n1 26.5955
R98 B2.n0 B2.t0 212.081
R99 B2.n1 B2.t2 212.081
R100 B2 B2.n2 158.72
R101 B2.n0 B2.t3 139.78
R102 B2.n1 B2.t1 139.78
R103 B2.n2 B2.n0 30.6732
R104 B2.n2 B2.n1 30.6732
R105 Y.n2 Y.n1 657.12
R106 Y Y.n3 208.458
R107 Y.n2 Y.n0 196.244
R108 Y.n1 Y.t1 26.5955
R109 Y.n1 Y.t0 26.5955
R110 Y.n0 Y.t5 26.5955
R111 Y.n0 Y.t4 26.5955
R112 Y.n3 Y.t2 24.9236
R113 Y.n3 Y.t3 24.9236
R114 Y Y.n2 9.23946
R115 VGND.n12 VGND.t5 286.426
R116 VGND.n7 VGND.n6 219.756
R117 VGND.n5 VGND.n4 207.965
R118 VGND.n19 VGND.t0 157.993
R119 VGND.n10 VGND.n3 34.6358
R120 VGND.n11 VGND.n10 34.6358
R121 VGND.n13 VGND.n11 34.6358
R122 VGND.n17 VGND.n1 34.6358
R123 VGND.n18 VGND.n17 34.6358
R124 VGND.n19 VGND.n18 30.8711
R125 VGND.n12 VGND.n1 26.3534
R126 VGND.n5 VGND.n3 25.224
R127 VGND.n6 VGND.t3 24.9236
R128 VGND.n6 VGND.t2 24.9236
R129 VGND.n4 VGND.t1 24.9236
R130 VGND.n4 VGND.t4 24.9236
R131 VGND.n7 VGND.n5 16.2661
R132 VGND.n20 VGND.n19 13.0652
R133 VGND.n8 VGND.n3 9.3005
R134 VGND.n10 VGND.n9 9.3005
R135 VGND.n11 VGND.n2 9.3005
R136 VGND.n14 VGND.n13 9.3005
R137 VGND.n15 VGND.n1 9.3005
R138 VGND.n17 VGND.n16 9.3005
R139 VGND.n18 VGND.n0 9.3005
R140 VGND.n13 VGND.n12 8.28285
R141 VGND.n8 VGND.n7 0.893984
R142 VGND.n9 VGND.n8 0.120292
R143 VGND.n9 VGND.n2 0.120292
R144 VGND.n14 VGND.n2 0.120292
R145 VGND.n15 VGND.n14 0.120292
R146 VGND.n16 VGND.n15 0.120292
R147 VGND.n16 VGND.n0 0.120292
R148 VGND.n20 VGND.n0 0.120292
R149 VGND VGND.n20 0.0213333
R150 a_471_47.n1 a_471_47.t3 311.62
R151 a_471_47.n2 a_471_47.t5 174.512
R152 a_471_47.n3 a_471_47.n2 98.982
R153 a_471_47.n1 a_471_47.n0 88.8348
R154 a_471_47.n2 a_471_47.n1 49.9695
R155 a_471_47.n0 a_471_47.t4 31.3851
R156 a_471_47.n0 a_471_47.t2 24.9236
R157 a_471_47.n3 a_471_47.t0 24.9236
R158 a_471_47.t1 a_471_47.n3 24.9236
R159 A1_N.n2 A1_N.n0 244.804
R160 A1_N.n1 A1_N.t2 236.18
R161 A1_N.n0 A1_N.t3 236.18
R162 A1_N.n1 A1_N.t0 163.881
R163 A1_N.n0 A1_N.t1 163.881
R164 A1_N.n2 A1_N.n1 152
R165 A1_N A1_N.n2 7.34865
C0 B2 Y 0.014468f
C1 Y VPB 0.005407f
C2 VPWR A1_N 0.082986f
C3 VPB A2_N 0.051079f
C4 VPWR Y 0.164208f
C5 VPWR A2_N 0.035863f
C6 Y A1_N 5.18e-19
C7 A1_N A2_N 0.213033f
C8 Y A2_N 9.39e-20
C9 B1 VGND 0.034644f
C10 B2 VGND 0.023446f
C11 VGND VPB 0.007942f
C12 B1 B2 0.203357f
C13 B1 VPB 0.074012f
C14 VPWR VGND 0.112313f
C15 VGND A1_N 0.058727f
C16 B1 VPWR 0.070185f
C17 B2 VPB 0.051071f
C18 Y VGND 0.012757f
C19 VGND A2_N 0.020843f
C20 B2 VPWR 0.015998f
C21 B1 Y 0.133324f
C22 VPWR VPB 0.120694f
C23 VPB A1_N 0.077469f
C24 VGND VNB 0.663699f
C25 Y VNB 0.012258f
C26 VPWR VNB 0.56065f
C27 B2 VNB 0.167862f
C28 B1 VNB 0.236335f
C29 A2_N VNB 0.167001f
C30 A1_N VNB 0.250905f
C31 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_4 VPB VNB VGND VPWR A2_N A1_N B2 Y B1
X0 a_1241_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_113_47.t6 A2_N.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_807_47.t3 a_113_47.t12 Y.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_113_47.t7 A2_N.t1 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t10 A2_N.t2 a_113_47.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t6 a_113_47.t13 a_807_47.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_1241_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y B2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t5 a_113_47.t14 a_807_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_27_47.t2 A2_N.t3 a_113_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t2 A1_N.t0 a_113_47.t8 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.135 ps=1.27 w=1 l=0.15
X12 a_113_47.t1 A2_N.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 a_27_47.t0 A2_N.t5 a_113_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_27_47.t4 A1_N.t1 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_1241_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47.t5 A1_N.t2 VGND.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_113_47.t11 A1_N.t3 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y B2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y.t2 a_113_47.t15 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t7 a_113_47.t16 Y.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_113_47.t4 A2_N.t6 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X22 a_1241_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND.t2 A1_N.t4 a_27_47.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 Y.t0 a_113_47.t17 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.38 ps=1.76 w=1 l=0.15
X25 VGND.t3 A1_N.t5 a_27_47.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR B1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR.t4 A1_N.t6 a_113_47.t9 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_113_47.t10 A1_N.t7 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR.t1 A2_N.t7 a_113_47.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_807_47.t0 a_113_47.t18 Y.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.247 pd=1.41 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B1.n10 B1.n8 212.081
R1 B1.n12 B1.n6 212.081
R2 B1.n14 B1.n4 212.081
R3 B1.n3 B1.n1 212.081
R4 B1.n11 B1.n0 172.725
R5 B1.n13 B1.n0 152
R6 B1.n10 B1.n9 139.78
R7 B1.n12 B1.n7 139.78
R8 B1.n14 B1.n5 139.78
R9 B1.n3 B1.n2 139.78
R10 B1 B1.n15 86.2792
R11 B1.n14 B1.n13 46.7399
R12 B1.n12 B1.n11 35.055
R13 B1.n15 B1.n3 31.6758
R14 B1.n11 B1.n10 26.2914
R15 B1.n15 B1.n14 23.0844
R16 B1.n13 B1.n12 14.6066
R17 B1 B1.n0 4.57193
R18 VPWR.n22 VPWR.t0 344.887
R19 VPWR.n10 VPWR.n9 324.276
R20 VPWR.n20 VPWR.n2 318.293
R21 VPWR.n4 VPWR.n3 318.293
R22 VPWR.n14 VPWR.n6 318.293
R23 VPWR.n8 VPWR.n7 134.257
R24 VPWR.n7 VPWR.t2 68.0259
R25 VPWR.n7 VPWR.t8 68.0256
R26 VPWR.n13 VPWR.n12 34.6358
R27 VPWR.n15 VPWR.n4 33.5064
R28 VPWR.n20 VPWR.n19 27.4829
R29 VPWR.n2 VPWR.t3 26.5955
R30 VPWR.n2 VPWR.t10 26.5955
R31 VPWR.n3 VPWR.t5 26.5955
R32 VPWR.n3 VPWR.t1 26.5955
R33 VPWR.n6 VPWR.t9 26.5955
R34 VPWR.n6 VPWR.t4 26.5955
R35 VPWR.n9 VPWR.t6 26.5955
R36 VPWR.n9 VPWR.t7 26.5955
R37 VPWR.n21 VPWR.n20 22.9652
R38 VPWR.n22 VPWR.n21 21.4593
R39 VPWR.n19 VPWR.n4 16.9417
R40 VPWR.n15 VPWR.n14 10.9181
R41 VPWR.n12 VPWR.n11 9.3005
R42 VPWR.n13 VPWR.n5 9.3005
R43 VPWR.n16 VPWR.n15 9.3005
R44 VPWR.n17 VPWR.n4 9.3005
R45 VPWR.n19 VPWR.n18 9.3005
R46 VPWR.n20 VPWR.n1 9.3005
R47 VPWR.n21 VPWR.n0 9.3005
R48 VPWR.n23 VPWR.n22 9.3005
R49 VPWR.n10 VPWR.n8 5.46011
R50 VPWR.n12 VPWR.n8 4.89462
R51 VPWR.n14 VPWR.n13 4.89462
R52 VPWR.n11 VPWR.n10 0.592895
R53 VPWR.n11 VPWR.n5 0.120292
R54 VPWR.n16 VPWR.n5 0.120292
R55 VPWR.n17 VPWR.n16 0.120292
R56 VPWR.n18 VPWR.n17 0.120292
R57 VPWR.n18 VPWR.n1 0.120292
R58 VPWR.n1 VPWR.n0 0.120292
R59 VPWR.n23 VPWR.n0 0.120292
R60 VPWR VPWR.n23 0.0252396
R61 VPB.t2 VPB.t8 538.63
R62 VPB.t7 VPB.t6 248.599
R63 VPB.t8 VPB.t7 248.599
R64 VPB.t9 VPB.t2 248.599
R65 VPB.t4 VPB.t9 248.599
R66 VPB.t5 VPB.t4 248.599
R67 VPB.t1 VPB.t5 248.599
R68 VPB.t3 VPB.t1 248.599
R69 VPB.t10 VPB.t3 248.599
R70 VPB.t0 VPB.t10 248.599
R71 VPB VPB.t0 210.125
R72 A2_N.n3 A2_N.t7 212.081
R73 A2_N.n5 A2_N.t0 212.081
R74 A2_N.n7 A2_N.t2 212.081
R75 A2_N.n1 A2_N.t6 212.081
R76 A2_N.n4 A2_N.n0 172.725
R77 A2_N.n9 A2_N.n2 172.725
R78 A2_N.n6 A2_N.n0 152
R79 A2_N.n9 A2_N.n8 152
R80 A2_N.n3 A2_N.t5 139.78
R81 A2_N.n5 A2_N.t1 139.78
R82 A2_N.n7 A2_N.t3 139.78
R83 A2_N.n1 A2_N.t4 139.78
R84 A2_N.n8 A2_N.n6 49.6611
R85 A2_N.n7 A2_N.n2 46.7399
R86 A2_N.n5 A2_N.n4 40.8975
R87 A2_N.n4 A2_N.n3 20.449
R88 A2_N.n2 A2_N.n1 14.6066
R89 A2_N A2_N.n0 13.1053
R90 A2_N.n6 A2_N.n5 8.76414
R91 A2_N A2_N.n9 7.61955
R92 A2_N.n8 A2_N.n7 2.92171
R93 a_113_47.n2 a_113_47.n0 226.355
R94 a_113_47.n16 a_113_47.t17 216.463
R95 a_113_47.n8 a_113_47.n7 212.081
R96 a_113_47.n6 a_113_47.t15 212.081
R97 a_113_47.n15 a_113_47.t16 212.081
R98 a_113_47.n4 a_113_47.n3 208.508
R99 a_113_47.n20 a_113_47.n19 208.507
R100 a_113_47.n22 a_113_47.n21 208.507
R101 a_113_47.n24 a_113_47.n23 208.506
R102 a_113_47.n2 a_113_47.n1 185
R103 a_113_47.n11 a_113_47.n10 172.725
R104 a_113_47.n18 a_113_47.n17 152
R105 a_113_47.n13 a_113_47.n5 152
R106 a_113_47.n12 a_113_47.n11 152
R107 a_113_47.n8 a_113_47.t18 144.162
R108 a_113_47.n16 a_113_47.t14 139.78
R109 a_113_47.n14 a_113_47.t12 139.78
R110 a_113_47.n9 a_113_47.t13 139.78
R111 a_113_47.n4 a_113_47.n2 97.9987
R112 a_113_47.n20 a_113_47.n18 87.7182
R113 a_113_47.n13 a_113_47.n12 49.6611
R114 a_113_47.n22 a_113_47.n20 44.424
R115 a_113_47.n23 a_113_47.n4 44.424
R116 a_113_47.n23 a_113_47.n22 44.424
R117 a_113_47.n17 a_113_47.n15 43.8187
R118 a_113_47.n10 a_113_47.n9 39.4369
R119 a_113_47.n19 a_113_47.t8 26.5955
R120 a_113_47.n19 a_113_47.t11 26.5955
R121 a_113_47.n21 a_113_47.t9 26.5955
R122 a_113_47.n21 a_113_47.t10 26.5955
R123 a_113_47.n3 a_113_47.t5 26.5955
R124 a_113_47.n3 a_113_47.t4 26.5955
R125 a_113_47.n24 a_113_47.t3 26.5955
R126 a_113_47.t6 a_113_47.n24 26.5955
R127 a_113_47.n1 a_113_47.t2 24.9236
R128 a_113_47.n1 a_113_47.t1 24.9236
R129 a_113_47.n0 a_113_47.t0 24.9236
R130 a_113_47.n0 a_113_47.t7 24.9236
R131 a_113_47.n11 a_113_47.n5 20.7243
R132 a_113_47.n18 a_113_47.n5 20.7243
R133 a_113_47.n10 a_113_47.n8 17.5278
R134 a_113_47.n17 a_113_47.n16 13.146
R135 a_113_47.n12 a_113_47.n6 5.84292
R136 a_113_47.n9 a_113_47.n6 4.38232
R137 a_113_47.n15 a_113_47.n14 4.38232
R138 a_113_47.n14 a_113_47.n13 1.46111
R139 Y.n1 Y.n0 252.931
R140 Y.n1 Y.t2 235.102
R141 Y.n4 Y.n2 226.355
R142 Y.n4 Y.n3 185
R143 Y Y.n5 92.3076
R144 Y.n5 Y.n4 57.3719
R145 Y.n5 Y.n1 27.1064
R146 Y.n0 Y.t1 26.5955
R147 Y.n0 Y.t0 26.5955
R148 Y.n2 Y.t3 24.9236
R149 Y.n2 Y.t5 24.9236
R150 Y.n3 Y.t4 24.9236
R151 Y.n3 Y.t6 24.9236
R152 a_807_47.n0 a_807_47.t1 266.642
R153 a_807_47.n1 a_807_47.n0 185
R154 a_807_47.n0 a_807_47.t0 174.833
R155 a_807_47.n1 a_807_47.t2 24.9236
R156 a_807_47.t3 a_807_47.n1 24.9236
R157 VNB.t9 VNB.t6 2677.02
R158 VNB.t7 VNB.t5 1196.12
R159 VNB.t8 VNB.t7 1196.12
R160 VNB.t6 VNB.t8 1196.12
R161 VNB.t11 VNB.t9 1196.12
R162 VNB.t4 VNB.t11 1196.12
R163 VNB.t10 VNB.t4 1196.12
R164 VNB.t0 VNB.t10 1196.12
R165 VNB.t3 VNB.t0 1196.12
R166 VNB.t2 VNB.t3 1196.12
R167 VNB.t1 VNB.t2 1196.12
R168 VNB VNB.t1 1011
R169 B2.n9 B2.n7 212.081
R170 B2.n11 B2.n5 212.081
R171 B2.n15 B2.n13 212.081
R172 B2.n3 B2.n1 212.081
R173 B2.n10 B2.n0 172.725
R174 B2.n17 B2.n4 172.725
R175 B2.n12 B2.n0 152
R176 B2.n17 B2.n16 152
R177 B2.n9 B2.n8 139.78
R178 B2.n11 B2.n6 139.78
R179 B2.n15 B2.n14 139.78
R180 B2.n3 B2.n2 139.78
R181 B2.n16 B2.n12 49.6611
R182 B2.n15 B2.n4 48.2005
R183 B2.n11 B2.n10 39.4369
R184 B2.n10 B2.n9 21.9096
R185 B2 B2.n0 16.1529
R186 B2.n4 B2.n3 13.146
R187 B2.n12 B2.n11 10.2247
R188 B2 B2.n17 4.57193
R189 B2.n16 B2.n15 1.46111
R190 VGND.n2 VGND.n1 220.102
R191 VGND.n2 VGND.n0 219.156
R192 VGND.n1 VGND.t1 24.9236
R193 VGND.n1 VGND.t3 24.9236
R194 VGND.n0 VGND.t0 24.9236
R195 VGND.n0 VGND.t2 24.9236
R196 VGND VGND.n2 1.08714
R197 a_27_47.n4 a_27_47.t1 306.731
R198 a_27_47.n5 a_27_47.n4 185
R199 a_27_47.n1 a_27_47.t5 174.512
R200 a_27_47.n1 a_27_47.n0 98.982
R201 a_27_47.n3 a_27_47.n2 88.3446
R202 a_27_47.n4 a_27_47.n3 53.5212
R203 a_27_47.n3 a_27_47.n1 48.9326
R204 a_27_47.n2 a_27_47.t6 24.9236
R205 a_27_47.n2 a_27_47.t0 24.9236
R206 a_27_47.n0 a_27_47.t7 24.9236
R207 a_27_47.n0 a_27_47.t4 24.9236
R208 a_27_47.t3 a_27_47.n5 24.9236
R209 a_27_47.n5 a_27_47.t2 24.9236
R210 A1_N.n3 A1_N.t0 212.081
R211 A1_N.n5 A1_N.t3 212.081
R212 A1_N.n7 A1_N.t6 212.081
R213 A1_N.n1 A1_N.t7 212.081
R214 A1_N.n4 A1_N.n0 172.725
R215 A1_N.n9 A1_N.n2 172.725
R216 A1_N.n6 A1_N.n0 152
R217 A1_N.n9 A1_N.n8 152
R218 A1_N.n3 A1_N.t2 139.78
R219 A1_N.n5 A1_N.t5 139.78
R220 A1_N.n7 A1_N.t1 139.78
R221 A1_N.n1 A1_N.t4 139.78
R222 A1_N.n8 A1_N.n6 49.6611
R223 A1_N.n7 A1_N.n2 48.2005
R224 A1_N.n5 A1_N.n4 39.4369
R225 A1_N.n4 A1_N.n3 21.9096
R226 A1_N A1_N.n9 17.9815
R227 A1_N.n2 A1_N.n1 13.146
R228 A1_N.n6 A1_N.n5 10.2247
R229 A1_N A1_N.n0 2.74336
R230 A1_N.n8 A1_N.n7 1.46111
C0 A2_N Y 1.31e-19
C1 A1_N Y 6.7e-19
C2 B2 B1 0.068777f
C3 a_1241_297# VPWR 0.641453f
C4 B2 VPWR 0.036901f
C5 a_1241_297# Y 0.26408f
C6 VPB VGND 0.015096f
C7 B2 Y 0.180922f
C8 B1 VPWR 0.084948f
C9 A2_N VGND 0.035782f
C10 VGND A1_N 0.049612f
C11 B1 Y 7.54e-19
C12 VPB A2_N 0.119261f
C13 a_1241_297# VGND 0.010123f
C14 VPWR Y 0.387841f
C15 VPB A1_N 0.120425f
C16 VGND B2 0.059771f
C17 A2_N A1_N 0.064024f
C18 a_1241_297# VPB 0.024807f
C19 VGND B1 0.060712f
C20 VPB B2 0.120606f
C21 VGND VPWR 0.199679f
C22 VPB B1 0.124186f
C23 VGND Y 0.030451f
C24 VPB VPWR 0.203244f
C25 a_1241_297# B2 0.064299f
C26 A2_N VPWR 0.087232f
C27 VPB Y 0.024371f
C28 A1_N VPWR 0.074066f
C29 a_1241_297# B1 0.231076f
C30 VGND VNB 1.08735f
C31 Y VNB 0.023331f
C32 VPWR VNB 0.911503f
C33 B1 VNB 0.395164f
C34 B2 VNB 0.362816f
C35 A1_N VNB 0.363082f
C36 A2_N VNB 0.380578f
C37 VPB VNB 2.0223f
C38 a_1241_297# VNB 0.034305f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR.t1 A1.t0 a_382_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47.t0 B1.t0 a_79_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47.t1 A1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t2 A2.t0 a_297_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR.t0 a_79_21.t3 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21.t2 B1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297.t0 A2.t1 a_79_21.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND.t0 a_79_21.t4 X.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t0 226.392
R1 A1 A1.n0 167.862
R2 A1.n0 A1.t1 158.275
R3 a_382_297.t0 a_382_297.t1 60.0855
R4 VPWR.n2 VPWR.n0 585
R5 VPWR.n1 VPWR.n0 585
R6 VPWR.n5 VPWR.t1 344.36
R7 VPWR.n4 VPWR.n3 275.348
R8 VPWR.n3 VPWR.n2 34.3087
R9 VPWR.n3 VPWR.n1 34.3087
R10 VPWR.n2 VPWR.t0 28.5655
R11 VPWR.n1 VPWR.t2 27.5805
R12 VPWR.n5 VPWR.n4 10.3977
R13 VPWR.n4 VPWR.n0 6.13008
R14 VPWR VPWR.n5 0.245228
R15 VPB.t0 VPB.t3 476.481
R16 VPB.t3 VPB.t1 319.627
R17 VPB.t1 VPB.t2 269.315
R18 VPB VPB.t0 204.207
R19 B1.n0 B1.t1 239.986
R20 B1 B1.n0 168.975
R21 B1.n0 B1.t0 167.685
R22 a_79_21.n2 a_79_21.n1 255.995
R23 a_79_21.n0 a_79_21.t3 231.017
R24 a_79_21.n1 a_79_21.t1 162.386
R25 a_79_21.n0 a_79_21.t4 158.716
R26 a_79_21.n1 a_79_21.n0 152
R27 a_79_21.n2 a_79_21.t2 41.3705
R28 a_79_21.t0 a_79_21.n2 35.4605
R29 a_297_47.n0 a_297_47.t1 364.741
R30 a_297_47.t0 a_297_47.n0 32.3082
R31 a_297_47.n0 a_297_47.t2 24.9236
R32 VNB.t0 VNB.t1 2677.02
R33 VNB.t1 VNB.t3 1310.03
R34 VNB.t3 VNB.t2 1196.12
R35 VNB VNB.t0 925.567
R36 VGND.n1 VGND.t0 297.233
R37 VGND.n1 VGND.n0 214.512
R38 VGND.n0 VGND.t1 24.9236
R39 VGND.n0 VGND.t2 24.9236
R40 VGND VGND.n1 0.182274
R41 A2.n0 A2.t1 241.536
R42 A2.n0 A2.t0 169.237
R43 A2 A2.n0 157.179
R44 X.n1 X.n0 585
R45 X X.n0 304.337
R46 X.n1 X.t1 172.978
R47 X.n0 X.t0 26.5955
R48 X X.n1 7.54336
C0 X VPWR 0.095752f
C1 X B1 3.56e-19
C2 VPWR VPB 0.062388f
C3 VPB B1 0.032789f
C4 X VGND 0.073624f
C5 VGND VPB 0.004903f
C6 VPWR B1 0.021269f
C7 VPB A2 0.033371f
C8 VPWR VGND 0.058833f
C9 VGND B1 0.018231f
C10 VPWR A2 0.083453f
C11 B1 A2 0.06645f
C12 VPB A1 0.041226f
C13 VGND A2 0.017086f
C14 VPWR A1 0.044921f
C15 VGND A1 0.015749f
C16 A2 A1 0.102437f
C17 X VPB 0.011001f
C18 VGND VNB 0.351611f
C19 VPWR VNB 0.304004f
C20 X VNB 0.09354f
C21 A1 VNB 0.152087f
C22 A2 VNB 0.098105f
C23 B1 VNB 0.101193f
C24 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21a_2 VNB VPB VGND VPWR X B1 A2 A1
X0 VPWR.t2 A1.t0 a_470_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21.t1 B1.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND.t1 a_79_21.t3 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 VGND.t2 A2.t0 a_384_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297.t1 A2.t1 a_79_21.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR.t0 a_79_21.t4 X.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15
X6 a_384_47.t2 B1.t1 a_79_21.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_384_47.t0 A1.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X.t0 a_79_21.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 X.t3 a_79_21.t6 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t0 230.155
R1 A1.n0 A1.t1 157.856
R2 A1 A1.n0 154.111
R3 a_470_297.t0 a_470_297.t1 63.0405
R4 VPWR.n9 VPWR.n8 585
R5 VPWR.n7 VPWR.n6 585
R6 VPWR.n11 VPWR.t1 415.579
R7 VPWR.n2 VPWR.t2 409.036
R8 VPWR.n8 VPWR.n7 102.441
R9 VPWR.n6 VPWR.n2 31.2874
R10 VPWR.n7 VPWR.t3 27.5805
R11 VPWR.n8 VPWR.t0 27.5805
R12 VPWR.n11 VPWR.n10 25.977
R13 VPWR.n10 VPWR.n9 22.607
R14 VPWR.n5 VPWR.n1 9.49727
R15 VPWR.n5 VPWR.n4 9.3005
R16 VPWR.n3 VPWR.n1 9.3005
R17 VPWR.n10 VPWR.n0 9.3005
R18 VPWR.n12 VPWR.n11 9.3005
R19 VPWR.n9 VPWR.n1 0.826306
R20 VPWR.n4 VPWR.n2 0.554787
R21 VPWR.n6 VPWR.n5 0.413403
R22 VPWR.n4 VPWR.n3 0.120292
R23 VPWR.n3 VPWR.n0 0.120292
R24 VPWR.n12 VPWR.n0 0.120292
R25 VPWR VPWR.n12 0.0213333
R26 VPB.t0 VPB.t4 562.306
R27 VPB.t3 VPB.t2 278.193
R28 VPB.t4 VPB.t3 254.518
R29 VPB.t1 VPB.t0 251.559
R30 VPB VPB.t1 189.409
R31 B1.n0 B1.t0 232.214
R32 B1 B1.n0 160.899
R33 B1.n0 B1.t1 159.915
R34 a_79_21.n3 a_79_21.n2 384.279
R35 a_79_21.n1 a_79_21.t4 208.868
R36 a_79_21.n0 a_79_21.t5 208.868
R37 a_79_21.n2 a_79_21.n1 183.082
R38 a_79_21.n2 a_79_21.t2 162.88
R39 a_79_21.n1 a_79_21.t3 139.78
R40 a_79_21.n0 a_79_21.t6 139.78
R41 a_79_21.n1 a_79_21.n0 60.2505
R42 a_79_21.t0 a_79_21.n3 27.5805
R43 a_79_21.n3 a_79_21.t1 27.5805
R44 X X.n0 594.144
R45 X.n2 X.n0 585
R46 X.n2 X.n1 257.62
R47 X.n0 X.t1 27.5805
R48 X.n0 X.t0 26.5955
R49 X.n1 X.t2 25.8467
R50 X.n1 X.t3 24.9236
R51 X X.n2 16.4576
R52 VGND.n3 VGND.t1 281.25
R53 VGND.n2 VGND.n1 205.72
R54 VGND.n5 VGND.t0 156.495
R55 VGND.n1 VGND.t3 29.539
R56 VGND.n1 VGND.t2 29.539
R57 VGND.n5 VGND.n4 25.977
R58 VGND.n4 VGND.n3 19.2005
R59 VGND.n6 VGND.n5 9.3005
R60 VGND.n4 VGND.n0 9.3005
R61 VGND.n3 VGND.n2 7.14895
R62 VGND.n2 VGND.n0 0.225736
R63 VGND.n6 VGND.n0 0.120292
R64 VGND VGND.n6 0.0213333
R65 VNB.t1 VNB.t4 2705.5
R66 VNB.t2 VNB.t3 1338.51
R67 VNB.t4 VNB.t2 1224.6
R68 VNB.t0 VNB.t1 1210.36
R69 VNB VNB.t0 911.327
R70 A2.n0 A2.t1 236.18
R71 A2 A2.n0 181.291
R72 A2.n0 A2.t0 163.881
R73 a_384_47.t0 a_384_47.n0 449.534
R74 a_384_47.n0 a_384_47.t1 25.8467
R75 a_384_47.n0 a_384_47.t2 25.8467
C0 A1 VPWR 0.048873f
C1 A1 VPB 0.040155f
C2 A1 B1 4.59e-19
C3 VPWR VPB 0.078997f
C4 A1 VGND 0.017567f
C5 VPWR X 0.13299f
C6 A1 A2 0.090246f
C7 VPWR B1 0.024191f
C8 X VPB 0.00507f
C9 VPWR VGND 0.07997f
C10 VPB B1 0.039443f
C11 VGND VPB 0.006428f
C12 X B1 3.33e-19
C13 VPWR A2 0.059208f
C14 X VGND 0.105923f
C15 VPB A2 0.033772f
C16 VGND B1 0.019516f
C17 B1 A2 0.099478f
C18 VGND A2 0.019566f
C19 VGND VNB 0.43148f
C20 X VNB 0.027585f
C21 VPWR VNB 0.383466f
C22 A1 VNB 0.150768f
C23 A2 VNB 0.101916f
C24 B1 VNB 0.1061f
C25 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND.t2 A2.t0 a_29_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y.t3 B1.t0 a_29_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR.t3 B1.t1 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR.t1 A1.t0 a_112_297.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47.t3 A2.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y.t1 A2.t2 a_112_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND.t0 A1.t1 a_29_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297.t2 A1.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297.t0 A2.t3 Y.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47.t0 B1.t2 Y.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y.t4 B1.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47.t5 A1.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
R0 A2.n0 A2.t3 212.081
R1 A2.n1 A2.t2 212.081
R2 A2.n0 A2.t0 139.78
R3 A2.n1 A2.t1 139.78
R4 A2 A2.n2 71.2431
R5 A2.n2 A2.n0 35.2128
R6 A2.n2 A2.n1 21.2357
R7 a_29_47.t0 a_29_47.n3 266.411
R8 a_29_47.n1 a_29_47.t2 176.514
R9 a_29_47.n1 a_29_47.n0 98.0123
R10 a_29_47.n3 a_29_47.n2 89.3175
R11 a_29_47.n3 a_29_47.n1 56.8835
R12 a_29_47.n2 a_29_47.t1 25.8467
R13 a_29_47.n2 a_29_47.t5 25.8467
R14 a_29_47.n0 a_29_47.t4 25.8467
R15 a_29_47.n0 a_29_47.t3 25.8467
R16 VGND.n2 VGND.n1 213.952
R17 VGND.n2 VGND.n0 213.636
R18 VGND.n0 VGND.t3 36.9236
R19 VGND.n0 VGND.t2 35.0774
R20 VGND.n1 VGND.t1 25.8467
R21 VGND.n1 VGND.t0 25.8467
R22 VGND VGND.n2 0.381594
R23 VNB.t4 VNB.t5 1537.86
R24 VNB.t1 VNB.t0 1224.6
R25 VNB.t5 VNB.t1 1224.6
R26 VNB.t3 VNB.t4 1224.6
R27 VNB.t2 VNB.t3 1224.6
R28 VNB VNB.t2 982.524
R29 B1.n2 B1.t1 265.101
R30 B1.n0 B1.t3 263.493
R31 B1 B1.n2 175.415
R32 B1.n1 B1.t2 160.667
R33 B1.n0 B1.t0 128.534
R34 B1.n1 B1.n0 83.4688
R35 B1.n2 B1.n1 32.1338
R36 Y.n3 Y.n0 596.712
R37 Y.n2 Y.n0 585
R38 Y.n5 Y.n4 585
R39 Y.n2 Y.n1 238.03
R40 Y Y.n3 30.5783
R41 Y.n4 Y.t0 27.5805
R42 Y.n4 Y.t1 27.5805
R43 Y.n0 Y.t5 27.5805
R44 Y.n0 Y.t4 27.5805
R45 Y.n1 Y.t2 25.8467
R46 Y.n1 Y.t3 25.8467
R47 Y Y.n5 22.2123
R48 Y Y.n2 9.44812
R49 Y.n3 Y 4.90263
R50 Y.n5 Y 2.63579
R51 VPWR.n3 VPWR.n2 599.74
R52 VPWR.n4 VPWR.t3 402.134
R53 VPWR.n9 VPWR.t0 338.553
R54 VPWR.n7 VPWR.n1 34.6358
R55 VPWR.n8 VPWR.n7 34.6358
R56 VPWR.n2 VPWR.t2 32.5055
R57 VPWR.n2 VPWR.t1 30.5355
R58 VPWR.n3 VPWR.n1 22.5887
R59 VPWR.n9 VPWR.n8 19.2005
R60 VPWR.n5 VPWR.n1 9.3005
R61 VPWR.n7 VPWR.n6 9.3005
R62 VPWR.n8 VPWR.n0 9.3005
R63 VPWR.n10 VPWR.n9 9.3005
R64 VPWR.n4 VPWR.n3 6.49172
R65 VPWR.n5 VPWR.n4 0.677932
R66 VPWR.n6 VPWR.n5 0.120292
R67 VPWR.n6 VPWR.n0 0.120292
R68 VPWR.n10 VPWR.n0 0.120292
R69 VPWR VPWR.n10 0.0239375
R70 VPB.t2 VPB.t1 295.95
R71 VPB.t1 VPB.t4 278.193
R72 VPB.t4 VPB.t5 254.518
R73 VPB.t3 VPB.t2 254.518
R74 VPB.t0 VPB.t3 254.518
R75 VPB VPB.t0 204.207
R76 A1 A1.n0 251.453
R77 A1.n0 A1.t0 236.18
R78 A1.n1 A1.t2 234.392
R79 A1.n0 A1.t3 163.881
R80 A1.n2 A1.n1 152
R81 A1.n1 A1.t1 150.442
R82 A1.n2 A1 11.055
R83 A1 A1.n2 2.13383
R84 a_112_297.n1 a_112_297.n0 943.162
R85 a_112_297.n0 a_112_297.t0 37.4305
R86 a_112_297.n0 a_112_297.t3 31.5205
R87 a_112_297.t1 a_112_297.n1 27.5805
R88 a_112_297.n1 a_112_297.t2 27.5805
C0 VGND VPB 0.005313f
C1 VGND Y 0.010009f
C2 VGND A1 0.03345f
C3 A2 VPWR 0.018401f
C4 A2 VPB 0.05711f
C5 B1 VPWR 0.073571f
C6 A2 Y 0.014024f
C7 B1 VPB 0.069214f
C8 A2 A1 0.221218f
C9 B1 Y 0.112227f
C10 VPWR VPB 0.077635f
C11 B1 A1 0.058994f
C12 VPWR Y 0.194637f
C13 Y VPB 0.005213f
C14 VPWR A1 0.082322f
C15 VGND A2 0.029375f
C16 VPB A1 0.079187f
C17 Y A1 0.135839f
C18 VGND B1 0.0228f
C19 VGND VPWR 0.06541f
C20 VGND VNB 0.387326f
C21 Y VNB 0.020784f
C22 VPWR VNB 0.378429f
C23 B1 VNB 0.254047f
C24 A2 VNB 0.179711f
C25 A1 VNB 0.254318f
C26 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y.t2 A2.t0 a_109_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR.t1 B1.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47.t2 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y.t0 B1.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND.t0 A1.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t0 240.484
R1 A2.n0 A2.t1 168.185
R2 A2.n1 A2.n0 159.952
R3 A2 A2.n1 7.87742
R4 A2.n1 A2 2.90959
R5 a_109_297.t0 a_109_297.t1 41.3705
R6 Y.n0 Y 593.34
R7 Y.n1 Y.n0 585
R8 Y Y.t0 305.245
R9 Y.n0 Y.t2 56.9025
R10 Y.n0 Y.t1 46.4362
R11 Y Y.n1 8.33989
R12 Y.n1 Y 4.84898
R13 VPB.t2 VPB.t1 319.627
R14 VPB.t0 VPB.t2 213.084
R15 VPB VPB.t0 189.409
R16 B1.n0 B1.t1 254.256
R17 B1.n0 B1.t0 181.956
R18 B1 B1.n0 154.667
R19 VPWR.n0 VPWR.t1 361.24
R20 VPWR.n0 VPWR.t0 251.102
R21 VPWR VPWR.n0 0.142966
R22 VGND VGND.n0 204.819
R23 VGND.n0 VGND.t0 36.0005
R24 VGND.n0 VGND.t1 24.9236
R25 a_27_47.t0 a_27_47.n0 471.692
R26 a_27_47.n0 a_27_47.t1 24.9236
R27 a_27_47.n0 a_27_47.t2 24.9236
R28 VNB.t0 VNB.t2 1366.99
R29 VNB.t2 VNB.t1 1196.12
R30 VNB VNB.t0 911.327
R31 A1.n0 A1.t0 234.483
R32 A1.n0 A1.t1 162.184
R33 A1 A1.n0 158.788
C0 A2 B1 0.047196f
C1 VPWR Y 0.105149f
C2 VPWR VGND 0.038082f
C3 VPWR VPB 0.056004f
C4 Y VGND 0.028878f
C5 Y VPB 0.00672f
C6 VPWR A1 0.049725f
C7 VPWR A2 0.10874f
C8 VGND VPB 0.004618f
C9 Y A1 8.9e-19
C10 VPWR B1 0.043328f
C11 Y A2 0.123701f
C12 VGND A1 0.016299f
C13 VPB A1 0.032652f
C14 VGND A2 0.01829f
C15 Y B1 0.081114f
C16 VPB A2 0.030454f
C17 VGND B1 0.016035f
C18 VPB B1 0.074099f
C19 A1 A2 0.098638f
C20 VGND VNB 0.253652f
C21 Y VNB 0.054462f
C22 VPWR VNB 0.271009f
C23 B1 VNB 0.151859f
C24 A2 VNB 0.096175f
C25 A1 VNB 0.138363f
C26 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_0 VNB VPB VGND VPWR B1 A1 Y A2
X0 a_120_369.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0768 pd=0.88 as=0.1696 ps=1.81 w=0.64 l=0.15
X1 VGND.t1 A1.t1 a_32_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X2 Y.t0 A2.t0 a_120_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0896 pd=0.92 as=0.0768 ps=0.88 w=0.64 l=0.15
X3 a_32_47.t0 A2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR.t1 B1.t0 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X5 Y.t1 B1.t1 a_32_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A1.n0 A1.t0 257.56
R1 A1.n0 A1.t1 197.018
R2 A1 A1.n0 68.9673
R3 VPWR.n0 VPWR.t0 382.204
R4 VPWR.n0 VPWR.t1 380.885
R5 VPWR VPWR.n0 0.166667
R6 a_120_369.t0 a_120_369.t1 73.8755
R7 VPB.t1 VPB.t2 254.518
R8 VPB.t0 VPB.t1 230.841
R9 VPB VPB.t0 224.923
R10 a_32_47.n0 a_32_47.t1 486.89
R11 a_32_47.n0 a_32_47.t2 40.0005
R12 a_32_47.t0 a_32_47.n0 40.0005
R13 VGND VGND.n0 204.85
R14 VGND.n0 VGND.t0 40.0005
R15 VGND.n0 VGND.t1 40.0005
R16 VNB.t0 VNB.t2 1224.6
R17 VNB.t1 VNB.t0 1224.6
R18 VNB VNB.t1 1011
R19 A2.n0 A2.t0 280.363
R20 A2.n0 A2.t1 219.31
R21 A2 A2.n0 164.534
R22 Y Y.n0 593.216
R23 Y.n1 Y.n0 585
R24 Y.n1 Y.t1 312.966
R25 Y.n0 Y.t2 43.0943
R26 Y.n0 Y.t0 43.0943
R27 Y Y.n1 5.15871
R28 B1.n0 B1.t1 309.517
R29 B1.n0 B1.t0 171.344
R30 B1 B1.n0 154.91
C0 Y A1 0.009573f
C1 VGND Y 0.043922f
C2 A2 B1 0.082922f
C3 A2 VPWR 0.025473f
C4 VPB A1 0.077136f
C5 A2 Y 0.059496f
C6 B1 VPWR 0.041323f
C7 VGND VPB 0.006029f
C8 B1 Y 0.089469f
C9 VGND A1 0.019176f
C10 VPWR Y 0.129332f
C11 A2 VPB 0.053524f
C12 A2 A1 0.119838f
C13 B1 VPB 0.071952f
C14 VGND A2 0.016172f
C15 VPWR VPB 0.057722f
C16 VGND B1 0.013944f
C17 Y VPB 0.011815f
C18 VPWR A1 0.051245f
C19 VGND VPWR 0.036805f
C20 VGND VNB 0.254196f
C21 Y VNB 0.069992f
C22 VPWR VNB 0.259532f
C23 B1 VNB 0.169823f
C24 A2 VNB 0.108932f
C25 A1 VNB 0.209504f
C26 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21a_4 VNB VPB VPWR VGND A2 A1 X B1
X0 X.t4 a_80_21.t6 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_475_47.t5 A1.t0 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X.t0 a_80_21.t7 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND.t2 a_80_21.t8 X.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_762_297.t0 A1.t1 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X5 a_475_47.t2 B1.t0 a_80_21.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND.t5 A2.t0 a_475_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND.t1 a_80_21.t9 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR.t2 a_80_21.t10 X.t7 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 X.t1 a_80_21.t11 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 a_80_21.t3 A2.t1 a_762_297.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_80_21.t1 B1.t1 a_475_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X12 a_80_21.t4 B1.t2 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X13 a_475_47.t0 A2.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X14 X.t6 a_80_21.t12 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR.t4 A1.t2 a_934_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X16 a_934_297.t0 A2.t3 a_80_21.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 VPWR.t7 B1.t3 a_80_21.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR.t0 a_80_21.t13 X.t5 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND.t7 A1.t3 a_475_47.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
R0 a_80_21.n18 a_80_21.n17 374.195
R1 a_80_21.n17 a_80_21.n0 297.127
R2 a_80_21.n16 a_80_21.n1 235.567
R3 a_80_21.n14 a_80_21.t13 225.226
R4 a_80_21.n12 a_80_21.t12 212.081
R5 a_80_21.n3 a_80_21.t10 212.081
R6 a_80_21.n5 a_80_21.t7 212.081
R7 a_80_21.n8 a_80_21.n4 164.8
R8 a_80_21.n4 a_80_21.t11 163.15
R9 a_80_21.n8 a_80_21.n7 152
R10 a_80_21.n10 a_80_21.n9 152
R11 a_80_21.n12 a_80_21.n2 152
R12 a_80_21.n15 a_80_21.n14 152
R13 a_80_21.n6 a_80_21.t9 139.78
R14 a_80_21.n11 a_80_21.t6 139.78
R15 a_80_21.n13 a_80_21.t8 139.78
R16 a_80_21.n17 a_80_21.n16 56.6999
R17 a_80_21.n12 a_80_21.n11 46.7399
R18 a_80_21.n7 a_80_21.n3 36.5157
R19 a_80_21.n14 a_80_21.n13 33.5944
R20 a_80_21.n0 a_80_21.t5 27.5805
R21 a_80_21.n0 a_80_21.t4 27.5805
R22 a_80_21.t2 a_80_21.n18 27.5805
R23 a_80_21.n18 a_80_21.t3 27.5805
R24 a_80_21.n1 a_80_21.t0 25.8467
R25 a_80_21.n1 a_80_21.t1 25.8467
R26 a_80_21.n5 a_80_21.n4 23.3702
R27 a_80_21.n13 a_80_21.n12 16.0672
R28 a_80_21.n6 a_80_21.n5 16.0672
R29 a_80_21.n10 a_80_21.n3 13.146
R30 a_80_21.n15 a_80_21.n2 12.8005
R31 a_80_21.n9 a_80_21.n2 12.8005
R32 a_80_21.n9 a_80_21.n8 12.8005
R33 a_80_21.n7 a_80_21.n6 10.2247
R34 a_80_21.n16 a_80_21.n15 8.28285
R35 a_80_21.n11 a_80_21.n10 2.92171
R36 VGND.n13 VGND.t2 281.25
R37 VGND.n19 VGND.t0 281.25
R38 VGND.n8 VGND.n5 204.392
R39 VGND.n17 VGND.n2 198.964
R40 VGND.n7 VGND.n6 198.554
R41 VGND.n6 VGND.t7 38.7697
R42 VGND.n11 VGND.n4 34.6358
R43 VGND.n12 VGND.n11 34.6358
R44 VGND.n13 VGND.n12 28.9887
R45 VGND.n6 VGND.t4 27.6928
R46 VGND.n5 VGND.t6 25.8467
R47 VGND.n5 VGND.t5 25.8467
R48 VGND.n2 VGND.t3 25.8467
R49 VGND.n2 VGND.t1 25.8467
R50 VGND.n7 VGND.n4 24.4711
R51 VGND.n17 VGND.n1 24.4711
R52 VGND.n18 VGND.n17 19.9534
R53 VGND.n19 VGND.n18 19.9534
R54 VGND.n13 VGND.n1 15.4358
R55 VGND.n20 VGND.n19 9.3005
R56 VGND.n9 VGND.n4 9.3005
R57 VGND.n11 VGND.n10 9.3005
R58 VGND.n12 VGND.n3 9.3005
R59 VGND.n14 VGND.n13 9.3005
R60 VGND.n15 VGND.n1 9.3005
R61 VGND.n17 VGND.n16 9.3005
R62 VGND.n18 VGND.n0 9.3005
R63 VGND.n8 VGND.n7 6.36102
R64 VGND.n9 VGND.n8 0.631783
R65 VGND.n10 VGND.n9 0.120292
R66 VGND.n10 VGND.n3 0.120292
R67 VGND.n14 VGND.n3 0.120292
R68 VGND.n15 VGND.n14 0.120292
R69 VGND.n16 VGND.n15 0.120292
R70 VGND.n16 VGND.n0 0.120292
R71 VGND.n20 VGND.n0 0.120292
R72 VGND VGND.n20 0.0213333
R73 X.n2 X.n0 366.902
R74 X.n2 X.n1 315.207
R75 X.n5 X.n3 242.938
R76 X.n5 X.n4 185
R77 X X.n2 92.1048
R78 X X.n5 29.6107
R79 X.n0 X.t5 27.5805
R80 X.n0 X.t6 27.5805
R81 X.n1 X.t7 27.5805
R82 X.n1 X.t0 27.5805
R83 X.n4 X.t2 25.8467
R84 X.n4 X.t1 25.8467
R85 X.n3 X.t3 25.8467
R86 X.n3 X.t4 25.8467
R87 VNB.t2 VNB.t7 2705.5
R88 VNB.t9 VNB.t4 1452.43
R89 VNB.t6 VNB.t9 1452.43
R90 VNB.t5 VNB.t8 1224.6
R91 VNB.t4 VNB.t5 1224.6
R92 VNB.t7 VNB.t6 1224.6
R93 VNB.t3 VNB.t2 1224.6
R94 VNB.t1 VNB.t3 1224.6
R95 VNB.t0 VNB.t1 1224.6
R96 VNB VNB.t0 925.567
R97 A1 A1.n0 251.714
R98 A1.n1 A1.t2 236.18
R99 A1.n0 A1.t1 233.288
R100 A1.n1 A1.t0 163.881
R101 A1 A1.n1 161.859
R102 A1.n0 A1.t3 160.988
R103 a_475_47.n2 a_475_47.t3 315.834
R104 a_475_47.n1 a_475_47.t5 275.599
R105 a_475_47.n1 a_475_47.n0 185
R106 a_475_47.n3 a_475_47.n2 89.5048
R107 a_475_47.n2 a_475_47.n1 64.5337
R108 a_475_47.n3 a_475_47.t2 40.6159
R109 a_475_47.n0 a_475_47.t1 25.8467
R110 a_475_47.n0 a_475_47.t0 25.8467
R111 a_475_47.t4 a_475_47.n3 25.8467
R112 VPWR.n13 VPWR.n12 598.898
R113 VPWR.n10 VPWR.n9 585
R114 VPWR.n8 VPWR.n7 585
R115 VPWR.n6 VPWR.t4 342.918
R116 VPWR.n21 VPWR.t3 338.507
R117 VPWR.n19 VPWR.n1 310.928
R118 VPWR.n9 VPWR.n8 66.9805
R119 VPWR.n18 VPWR.n2 34.6358
R120 VPWR.n14 VPWR.n11 34.6358
R121 VPWR.n12 VPWR.t0 31.5205
R122 VPWR.n21 VPWR.n20 30.4946
R123 VPWR.n7 VPWR.n6 28.45
R124 VPWR.n8 VPWR.t5 27.5805
R125 VPWR.n9 VPWR.t7 27.5805
R126 VPWR.n1 VPWR.t1 27.5805
R127 VPWR.n1 VPWR.t2 27.5805
R128 VPWR.n12 VPWR.t6 27.5805
R129 VPWR.n20 VPWR.n19 9.41227
R130 VPWR.n5 VPWR.n4 9.3005
R131 VPWR.n11 VPWR.n3 9.3005
R132 VPWR.n15 VPWR.n14 9.3005
R133 VPWR.n16 VPWR.n2 9.3005
R134 VPWR.n18 VPWR.n17 9.3005
R135 VPWR.n20 VPWR.n0 9.3005
R136 VPWR.n22 VPWR.n21 6.61781
R137 VPWR.n10 VPWR.n4 6.52125
R138 VPWR.n11 VPWR.n10 5.86776
R139 VPWR.n13 VPWR.n2 4.89462
R140 VPWR.n14 VPWR.n13 3.38874
R141 VPWR.n7 VPWR.n4 1.69107
R142 VPWR.n19 VPWR.n18 0.376971
R143 VPWR.n6 VPWR.n5 0.223724
R144 VPWR.n22 VPWR.n0 0.154914
R145 VPWR.n5 VPWR.n3 0.120292
R146 VPWR.n15 VPWR.n3 0.120292
R147 VPWR.n16 VPWR.n15 0.120292
R148 VPWR.n17 VPWR.n16 0.120292
R149 VPWR.n17 VPWR.n0 0.120292
R150 VPWR VPWR.n22 0.107063
R151 VPB.t9 VPB.t6 455.764
R152 VPB VPB.t3 381.776
R153 VPB.t0 VPB.t8 266.356
R154 VPB.t4 VPB.t5 254.518
R155 VPB.t7 VPB.t4 254.518
R156 VPB.t6 VPB.t7 254.518
R157 VPB.t8 VPB.t9 254.518
R158 VPB.t1 VPB.t0 254.518
R159 VPB.t2 VPB.t1 254.518
R160 VPB.t3 VPB.t2 254.518
R161 a_762_297.t0 a_762_297.t1 55.1605
R162 B1.n3 B1.t2 228.877
R163 B1.n1 B1.t3 212.081
R164 B1.n0 B1.t0 162.419
R165 B1 B1.n3 158.637
R166 B1 B1.n0 153.423
R167 B1.n2 B1.t1 139.78
R168 B1.n2 B1.n1 36.5157
R169 B1.n3 B1.n2 9.49444
R170 B1.n1 B1.n0 3.65202
R171 A2.n0 A2.t3 212.081
R172 A2.n1 A2.t1 212.081
R173 A2.n0 A2.t0 139.78
R174 A2.n1 A2.t2 139.78
R175 A2 A2.n2 68.4298
R176 A2.n2 A2.n1 31.1903
R177 A2.n2 A2.n0 23.8138
R178 a_934_297.t0 a_934_297.t1 55.1605
C0 VPWR X 0.320138f
C1 VPB A2 0.055963f
C2 B1 A1 0.076697f
C3 VPWR VGND 0.112219f
C4 X VGND 0.14134f
C5 A1 A2 0.20474f
C6 VPB VPWR 0.122982f
C7 B1 VPWR 0.030977f
C8 VPB X 0.021402f
C9 VPB VGND 0.009535f
C10 A1 VPWR 0.09105f
C11 B1 X 6.82e-19
C12 B1 VGND 0.021643f
C13 A2 VPWR 0.026983f
C14 A1 VGND 0.036414f
C15 A2 VGND 0.033295f
C16 VPB B1 0.06822f
C17 VPB A1 0.080302f
C18 VGND VNB 0.642083f
C19 X VNB 0.05864f
C20 VPWR VNB 0.557258f
C21 A2 VNB 0.179165f
C22 A1 VNB 0.256876f
C23 B1 VNB 0.193817f
C24 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ba_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_2 VNB VPB VGND VPWR A2 A1 B1_N X
X0 VGND.t2 B1_N.t0 a_27_93.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND.t1 A2.t0 a_478_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X2 a_478_47.t1 a_27_93.t2 a_174_21.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_478_47.t2 A1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X.t2 a_174_21.t3 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5 VPWR.t2 a_174_21.t4 X.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 X.t3 a_174_21.t5 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 VPWR.t4 A1.t1 a_574_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND.t0 a_174_21.t6 X.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t3 B1_N.t1 a_27_93.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 a_574_297.t0 A2.t1 a_174_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X11 a_174_21.t2 a_27_93.t3 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.395 ps=1.79 w=1 l=0.15
R0 B1_N B1_N.n0 154.012
R1 B1_N.n0 B1_N.t1 148.35
R2 B1_N.n0 B1_N.t0 132.282
R3 a_27_93.t0 a_27_93.n1 648.322
R4 a_27_93.n1 a_27_93.n0 394.529
R5 a_27_93.n1 a_27_93.t1 288.954
R6 a_27_93.n0 a_27_93.t3 212.081
R7 a_27_93.n0 a_27_93.t2 139.78
R8 VGND.n3 VGND.t0 281.589
R9 VGND.n6 VGND.n5 231.934
R10 VGND.n2 VGND.n1 215.212
R11 VGND.n5 VGND.t4 41.6488
R12 VGND.n5 VGND.t2 38.5719
R13 VGND.n6 VGND.n4 28.2358
R14 VGND.n1 VGND.t3 24.9236
R15 VGND.n1 VGND.t1 24.9236
R16 VGND.n4 VGND.n3 19.577
R17 VGND.n4 VGND.n0 9.3005
R18 VGND.n7 VGND.n6 7.4049
R19 VGND.n3 VGND.n2 7.02737
R20 VGND.n2 VGND.n0 0.212293
R21 VGND.n7 VGND.n0 0.144904
R22 VGND VGND.n7 0.118504
R23 VNB.t0 VNB.t2 2705.5
R24 VNB.t2 VNB.t1 1352.75
R25 VNB.t3 VNB.t5 1352.75
R26 VNB.t1 VNB.t4 1196.12
R27 VNB.t5 VNB.t0 1196.12
R28 VNB VNB.t3 925.567
R29 A2.n0 A2.t1 241.536
R30 A2 A2.n0 169.677
R31 A2.n0 A2.t0 169.237
R32 a_478_47.n0 a_478_47.t2 371.981
R33 a_478_47.n0 a_478_47.t1 35.0774
R34 a_478_47.t0 a_478_47.n0 24.9236
R35 a_174_21.n3 a_174_21.n2 253.478
R36 a_174_21.n0 a_174_21.t4 212.81
R37 a_174_21.n1 a_174_21.t5 212.081
R38 a_174_21.n2 a_174_21.n0 203.82
R39 a_174_21.n1 a_174_21.t3 141.242
R40 a_174_21.n0 a_174_21.t6 139.78
R41 a_174_21.n2 a_174_21.t1 135.516
R42 a_174_21.n0 a_174_21.n1 60.6157
R43 a_174_21.n3 a_174_21.t2 38.4155
R44 a_174_21.t0 a_174_21.n3 26.5955
R45 A1.n0 A1.t1 234.804
R46 A1.n0 A1.t0 162.504
R47 A1 A1.n0 154.327
R48 X X.n0 668.782
R49 X X.n1 185.218
R50 X.n0 X.t0 26.5955
R51 X.n0 X.t3 26.5955
R52 X.n1 X.t1 24.9236
R53 X.n1 X.t2 24.9236
R54 VPWR.n10 VPWR.n1 600.812
R55 VPWR.n8 VPWR.n7 585
R56 VPWR.n6 VPWR.n5 585
R57 VPWR.n4 VPWR.t4 345.462
R58 VPWR.n1 VPWR.t3 96.1553
R59 VPWR.n7 VPWR.n6 90.6205
R60 VPWR.n6 VPWR.t0 34.4755
R61 VPWR.n7 VPWR.t2 30.5355
R62 VPWR.n1 VPWR.t1 25.6105
R63 VPWR.n9 VPWR.n8 24.0068
R64 VPWR.n10 VPWR.n9 18.0711
R65 VPWR.n5 VPWR.n2 9.70717
R66 VPWR.n3 VPWR.n2 9.3005
R67 VPWR.n9 VPWR.n0 9.3005
R68 VPWR.n5 VPWR.n4 7.26622
R69 VPWR.n11 VPWR.n10 7.14087
R70 VPWR.n4 VPWR.n3 0.251847
R71 VPWR.n11 VPWR.n0 0.148262
R72 VPWR.n3 VPWR.n0 0.120292
R73 VPWR VPWR.n11 0.115103
R74 VPWR.n8 VPWR.n2 0.107167
R75 VPB.t3 VPB.t1 556.386
R76 VPB.t4 VPB.t2 287.072
R77 VPB.t1 VPB.t0 284.113
R78 VPB.t2 VPB.t3 248.599
R79 VPB.t0 VPB.t5 213.084
R80 VPB VPB.t4 192.369
R81 a_574_297.t0 a_574_297.t1 41.3705
C0 VPB A1 0.039065f
C1 VPWR B1_N 0.010054f
C2 A2 A1 0.08184f
C3 VPB VPWR 0.089281f
C4 VPWR X 0.014526f
C5 A2 VPWR 0.0222f
C6 VPB B1_N 0.038629f
C7 B1_N X 0.059031f
C8 VGND A1 0.01629f
C9 VPB X 0.00312f
C10 VPB A2 0.025723f
C11 VGND VPWR 0.076383f
C12 VGND B1_N 0.034972f
C13 VPB VGND 0.007751f
C14 VGND X 0.111699f
C15 A2 VGND 0.015205f
C16 A1 VPWR 0.053552f
C17 VGND VNB 0.453428f
C18 X VNB 0.005337f
C19 B1_N VNB 0.12157f
C20 VPWR VNB 0.395412f
C21 A1 VNB 0.145852f
C22 A2 VNB 0.089905f
C23 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ba_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_1 VNB VPB VGND VPWR B1_N A1 A2 X
X0 a_222_93.t1 B1_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR.t2 A1.t0 a_544_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND.t3 a_79_199.t3 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93.t0 B1_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND.t2 A2.t0 a_448_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47.t2 a_222_93.t2 a_79_199.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199.t1 a_222_93.t3 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297.t0 A2.t1 a_79_199.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47.t1 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t1 a_79_199.t4 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
R0 B1_N B1_N.n0 154.715
R1 B1_N.n0 B1_N.t1 144.548
R2 B1_N.n0 B1_N.t0 128.482
R3 VGND.n2 VGND.n0 238.963
R4 VGND.n2 VGND.n1 219.91
R5 VGND.n0 VGND.t1 47.1434
R6 VGND.n0 VGND.t3 35.4291
R7 VGND.n1 VGND.t0 24.9236
R8 VGND.n1 VGND.t2 24.9236
R9 VGND VGND.n2 0.180332
R10 a_222_93.t0 a_222_93.n1 703.663
R11 a_222_93.n1 a_222_93.t1 276.654
R12 a_222_93.n1 a_222_93.n0 232.333
R13 a_222_93.n0 a_222_93.t3 212.081
R14 a_222_93.n0 a_222_93.t2 139.78
R15 VNB.t1 VNB.t3 3218.12
R16 VNB.t4 VNB.t1 1381.23
R17 VNB.t3 VNB.t2 1366.99
R18 VNB.t2 VNB.t0 1196.12
R19 VNB VNB.t4 1153.4
R20 A1.n0 A1.t0 234.804
R21 A1 A1.n0 167.238
R22 A1.n0 A1.t1 162.504
R23 a_544_297.t0 a_544_297.t1 41.3705
R24 VPWR.n2 VPWR.t3 808.141
R25 VPWR.n7 VPWR.n1 613.71
R26 VPWR.n3 VPWR.t2 251.738
R27 VPWR.n1 VPWR.t0 114.918
R28 VPWR.n6 VPWR.n5 34.6358
R29 VPWR.n1 VPWR.t1 33.4905
R30 VPWR.n7 VPWR.n6 10.9181
R31 VPWR.n5 VPWR.n2 10.5417
R32 VPWR.n5 VPWR.n4 9.3005
R33 VPWR.n6 VPWR.n0 9.3005
R34 VPWR.n3 VPWR.n2 7.41335
R35 VPWR.n8 VPWR.n7 7.4049
R36 VPWR.n4 VPWR.n3 0.308712
R37 VPWR.n8 VPWR.n0 0.144904
R38 VPWR.n4 VPWR.n0 0.120292
R39 VPWR VPWR.n8 0.118504
R40 VPB.t0 VPB.t4 668.847
R41 VPB.t1 VPB.t0 334.425
R42 VPB.t4 VPB.t2 284.113
R43 VPB.t2 VPB.t3 213.084
R44 VPB VPB.t1 192.369
R45 a_79_199.n1 a_79_199.t2 283.509
R46 a_79_199.n1 a_79_199.n0 266.269
R47 a_79_199.n0 a_79_199.t4 235.821
R48 a_79_199.n2 a_79_199.n1 195.048
R49 a_79_199.n0 a_79_199.t3 163.52
R50 a_79_199.n2 a_79_199.t1 38.4155
R51 a_79_199.t0 a_79_199.n2 26.5955
R52 X X.n0 592.529
R53 X.n1 X.n0 289.336
R54 X.n1 X.t1 261.212
R55 X.n0 X.t0 26.5955
R56 X X.n1 11.6023
R57 A2.n0 A2.t1 241.536
R58 A2.n0 A2.t0 169.237
R59 A2 A2.n0 160.534
R60 a_448_47.n0 a_448_47.t1 275.274
R61 a_448_47.n0 a_448_47.t2 36.0005
R62 a_448_47.t0 a_448_47.n0 24.9236
C0 VPWR B1_N 0.004485f
C1 VPWR VGND 0.074192f
C2 VPB VPWR 0.109668f
C3 B1_N VGND 0.016051f
C4 A2 VPWR 0.022715f
C5 VPB B1_N 0.041907f
C6 VPB VGND 0.011612f
C7 A1 VPWR 0.050783f
C8 A2 VGND 0.015713f
C9 X VPWR 0.072913f
C10 VPB A2 0.02588f
C11 A1 VGND 0.017036f
C12 X B1_N 0.001139f
C13 VPB A1 0.038356f
C14 X VGND 0.060887f
C15 A2 A1 0.079314f
C16 VPB X 0.013182f
C17 VGND VNB 0.468282f
C18 B1_N VNB 0.105165f
C19 VPWR VNB 0.400387f
C20 X VNB 0.086477f
C21 A1 VNB 0.13607f
C22 A2 VNB 0.09044f
C23 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_4 VNB VPB VPWR VGND B1 Y A1 A2
X0 VPWR.t6 B1.t0 Y.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297.t4 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297.t5 A2.t0 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR.t1 A1.t1 a_115_297.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND.t7 A2.t1 a_32_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y.t2 B1.t1 a_32_47.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND.t3 A1.t2 a_32_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 Y.t5 B1.t2 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47.t10 B1.t3 Y.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y.t8 B1.t4 a_32_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y.t0 A2.t2 a_115_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47.t6 A2.t3 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47.t8 B1.t5 Y.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47.t5 A2.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297.t6 A2.t5 Y.t10 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47.t2 A1.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR.t4 B1.t6 Y.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47.t1 A1.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND.t4 A2.t6 a_32_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y.t3 B1.t7 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR.t2 A1.t5 a_115_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y.t11 A2.t7 a_115_297.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND.t0 A1.t6 a_32_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297.t1 A1.t7 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
R0 B1.n6 B1.t0 212.081
R1 B1.n2 B1.t6 212.081
R2 B1.n1 B1.t2 212.081
R3 B1.n7 B1.t7 212.081
R4 B1.n4 B1.n3 168.738
R5 B1 B1.n8 162.585
R6 B1.n5 B1.n4 152
R7 B1.n6 B1.n0 152
R8 B1.n6 B1.t5 139.78
R9 B1.n2 B1.t3 139.78
R10 B1.n1 B1.t1 139.78
R11 B1.n7 B1.t4 139.78
R12 B1.n6 B1.n5 49.6611
R13 B1.n8 B1.n6 49.6611
R14 B1.n3 B1.n1 36.5157
R15 B1.n3 B1.n2 26.2914
R16 B1.n4 B1.n0 16.739
R17 B1.n5 B1.n1 13.146
R18 B1.n8 B1.n7 13.146
R19 B1 B1.n0 6.15435
R20 Y.n3 Y.n1 649.754
R21 Y.n3 Y.n2 585
R22 Y.n6 Y.n0 296.077
R23 Y.n5 Y.n4 295.69
R24 Y.n9 Y.n7 232.862
R25 Y.n9 Y.n8 185
R26 Y.n5 Y.n3 100.864
R27 Y Y.n6 40.8361
R28 Y.n0 Y.t4 27.5805
R29 Y.n0 Y.t5 27.5805
R30 Y.n1 Y.t10 27.5805
R31 Y.n1 Y.t0 27.5805
R32 Y.n2 Y.t1 27.5805
R33 Y.n2 Y.t11 27.5805
R34 Y.n4 Y.t6 27.5805
R35 Y.n4 Y.t3 27.5805
R36 Y.n7 Y.t7 25.8467
R37 Y.n7 Y.t8 25.8467
R38 Y.n8 Y.t9 25.8467
R39 Y.n8 Y.t2 25.8467
R40 Y Y.n9 21.6845
R41 Y.n6 Y.n5 17.2999
R42 VPWR.n6 VPWR.n5 601.457
R43 VPWR.n21 VPWR.n2 599.74
R44 VPWR.n9 VPWR.n8 599.74
R45 VPWR.n7 VPWR.t4 343.728
R46 VPWR.n23 VPWR.t7 340.916
R47 VPWR.n15 VPWR.n14 34.6358
R48 VPWR.n16 VPWR.n15 34.6358
R49 VPWR.n16 VPWR.n3 34.6358
R50 VPWR.n20 VPWR.n3 34.6358
R51 VPWR.n10 VPWR.n6 34.6358
R52 VPWR.n5 VPWR.t3 31.5205
R53 VPWR.n5 VPWR.t1 31.5205
R54 VPWR.n2 VPWR.t0 27.5805
R55 VPWR.n2 VPWR.t2 27.5805
R56 VPWR.n8 VPWR.t5 27.5805
R57 VPWR.n8 VPWR.t6 27.5805
R58 VPWR.n21 VPWR.n20 22.5887
R59 VPWR.n22 VPWR.n21 21.8358
R60 VPWR.n23 VPWR.n22 21.4593
R61 VPWR.n14 VPWR.n6 13.5534
R62 VPWR.n9 VPWR.n7 9.54996
R63 VPWR.n11 VPWR.n10 9.3005
R64 VPWR.n12 VPWR.n6 9.3005
R65 VPWR.n14 VPWR.n13 9.3005
R66 VPWR.n15 VPWR.n4 9.3005
R67 VPWR.n17 VPWR.n16 9.3005
R68 VPWR.n18 VPWR.n3 9.3005
R69 VPWR.n20 VPWR.n19 9.3005
R70 VPWR.n21 VPWR.n1 9.3005
R71 VPWR.n22 VPWR.n0 9.3005
R72 VPWR.n24 VPWR.n23 9.3005
R73 VPWR.n10 VPWR.n9 6.77697
R74 VPWR.n11 VPWR.n7 1.16488
R75 VPWR.n12 VPWR.n11 0.120292
R76 VPWR.n13 VPWR.n12 0.120292
R77 VPWR.n13 VPWR.n4 0.120292
R78 VPWR.n17 VPWR.n4 0.120292
R79 VPWR.n18 VPWR.n17 0.120292
R80 VPWR.n19 VPWR.n18 0.120292
R81 VPWR.n19 VPWR.n1 0.120292
R82 VPWR.n1 VPWR.n0 0.120292
R83 VPWR.n24 VPWR.n0 0.120292
R84 VPWR VPWR.n24 0.0226354
R85 VPB.t1 VPB.t5 278.193
R86 VPB.t7 VPB.t6 254.518
R87 VPB.t8 VPB.t7 254.518
R88 VPB.t5 VPB.t8 254.518
R89 VPB.t4 VPB.t1 254.518
R90 VPB.t10 VPB.t4 254.518
R91 VPB.t9 VPB.t10 254.518
R92 VPB.t3 VPB.t9 254.518
R93 VPB.t0 VPB.t3 254.518
R94 VPB.t2 VPB.t0 254.518
R95 VPB.t11 VPB.t2 254.518
R96 VPB VPB.t11 210.125
R97 A1.n1 A1.n0 326.01
R98 A1.n0 A1.t1 236.18
R99 A1.n4 A1.t0 212.081
R100 A1.n6 A1.t5 212.081
R101 A1.n2 A1.t7 212.081
R102 A1.n0 A1.t3 163.881
R103 A1.n5 A1.n1 152
R104 A1.n8 A1.n7 152
R105 A1.n4 A1.t6 139.78
R106 A1.n6 A1.t4 139.78
R107 A1.n2 A1.t2 139.78
R108 A1.n8 A1.n3 87.6153
R109 A1.n6 A1.n3 51.6904
R110 A1.n7 A1.n5 49.6611
R111 A1.n3 A1.n2 10.1344
R112 A1.n5 A1.n4 7.30353
R113 A1.n7 A1.n6 5.84292
R114 A1 A1.n1 4.6811
R115 A1 A1.n8 1.81543
R116 a_115_297.n4 a_115_297.n0 670.314
R117 a_115_297.n3 a_115_297.n1 642.938
R118 a_115_297.n3 a_115_297.n2 585
R119 a_115_297.n5 a_115_297.n4 585
R120 a_115_297.n4 a_115_297.n3 57.9373
R121 a_115_297.n0 a_115_297.t2 27.5805
R122 a_115_297.n0 a_115_297.t1 27.5805
R123 a_115_297.n2 a_115_297.t7 27.5805
R124 a_115_297.n2 a_115_297.t6 27.5805
R125 a_115_297.n1 a_115_297.t3 27.5805
R126 a_115_297.n1 a_115_297.t5 27.5805
R127 a_115_297.n5 a_115_297.t0 27.5805
R128 a_115_297.t4 a_115_297.n5 27.5805
R129 A2.n1 A2.t0 212.081
R130 A2.n3 A2.t7 212.081
R131 A2.n5 A2.t5 212.081
R132 A2.n6 A2.t2 212.081
R133 A2.n2 A2.n0 170.619
R134 A2.n4 A2.n0 152
R135 A2.n8 A2.n7 152
R136 A2.n1 A2.t1 139.78
R137 A2.n3 A2.t3 139.78
R138 A2.n5 A2.t6 139.78
R139 A2.n6 A2.t4 139.78
R140 A2.n5 A2.n4 54.0429
R141 A2.n7 A2.n6 54.0429
R142 A2.n3 A2.n2 49.6611
R143 A2.n8 A2.n0 20.015
R144 A2.n2 A2.n1 13.146
R145 A2.n4 A2.n3 8.76414
R146 A2.n7 A2.n5 8.76414
R147 A2 A2.n8 8.14595
R148 a_32_47.t10 a_32_47.n9 327.147
R149 a_32_47.n1 a_32_47.t3 264.545
R150 a_32_47.n5 a_32_47.n4 185
R151 a_32_47.n3 a_32_47.n2 185
R152 a_32_47.n1 a_32_47.n0 185
R153 a_32_47.n7 a_32_47.n6 185
R154 a_32_47.n9 a_32_47.n8 185
R155 a_32_47.n9 a_32_47.n7 62.1113
R156 a_32_47.n7 a_32_47.n5 57.5055
R157 a_32_47.n5 a_32_47.n3 53.6981
R158 a_32_47.n3 a_32_47.n1 53.6981
R159 a_32_47.n8 a_32_47.t11 25.8467
R160 a_32_47.n8 a_32_47.t8 25.8467
R161 a_32_47.n6 a_32_47.t9 25.8467
R162 a_32_47.n6 a_32_47.t2 25.8467
R163 a_32_47.n0 a_32_47.t0 25.8467
R164 a_32_47.n0 a_32_47.t1 25.8467
R165 a_32_47.n2 a_32_47.t4 25.8467
R166 a_32_47.n2 a_32_47.t5 25.8467
R167 a_32_47.n4 a_32_47.t7 25.8467
R168 a_32_47.n4 a_32_47.t6 25.8467
R169 VGND.n6 VGND.n3 203.915
R170 VGND.n5 VGND.n4 198.964
R171 VGND.n9 VGND.n2 198.964
R172 VGND.n12 VGND.n11 198.964
R173 VGND.n3 VGND.t2 33.2313
R174 VGND.n3 VGND.t7 25.8467
R175 VGND.n4 VGND.t6 25.8467
R176 VGND.n4 VGND.t4 25.8467
R177 VGND.n2 VGND.t5 25.8467
R178 VGND.n2 VGND.t0 25.8467
R179 VGND.n11 VGND.t1 25.8467
R180 VGND.n11 VGND.t3 25.8467
R181 VGND.n9 VGND.n1 24.8476
R182 VGND.n12 VGND.n10 20.3299
R183 VGND.n10 VGND.n9 19.577
R184 VGND.n5 VGND.n1 15.0593
R185 VGND.n7 VGND.n1 9.3005
R186 VGND.n9 VGND.n8 9.3005
R187 VGND.n10 VGND.n0 9.3005
R188 VGND.n13 VGND.n12 7.25484
R189 VGND.n6 VGND.n5 6.8128
R190 VGND.n7 VGND.n6 0.684746
R191 VGND.n13 VGND.n0 0.146813
R192 VGND.n8 VGND.n7 0.120292
R193 VGND.n8 VGND.n0 0.120292
R194 VGND VGND.n13 0.116571
R195 VNB.t7 VNB.t2 1338.51
R196 VNB.t11 VNB.t10 1224.6
R197 VNB.t8 VNB.t11 1224.6
R198 VNB.t9 VNB.t8 1224.6
R199 VNB.t2 VNB.t9 1224.6
R200 VNB.t6 VNB.t7 1224.6
R201 VNB.t4 VNB.t6 1224.6
R202 VNB.t5 VNB.t4 1224.6
R203 VNB.t0 VNB.t5 1224.6
R204 VNB.t1 VNB.t0 1224.6
R205 VNB.t3 VNB.t1 1224.6
R206 VNB VNB.t3 1011
C0 B1 VPWR 0.053036f
C1 A2 Y 0.024846f
C2 B1 Y 0.36131f
C3 A2 VGND 0.065981f
C4 VPB A1 0.151717f
C5 VPWR Y 0.34787f
C6 B1 VGND 0.031015f
C7 VPWR VGND 0.117721f
C8 Y VGND 0.043236f
C9 VPB A2 0.118886f
C10 VPB B1 0.123824f
C11 A1 A2 0.290574f
C12 A1 B1 0.076799f
C13 VPB VPWR 0.130182f
C14 A1 VPWR 0.106383f
C15 VPB Y 0.019834f
C16 VPB VGND 0.009998f
C17 A1 Y 0.19145f
C18 A1 VGND 0.073118f
C19 A2 VPWR 0.034747f
C20 VGND VNB 0.669095f
C21 Y VNB 0.069548f
C22 VPWR VNB 0.596421f
C23 B1 VNB 0.380316f
C24 A2 VNB 0.355607f
C25 A1 VNB 0.444055f
C26 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21bai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21bai_2 VNB VPB VGND VPWR B1_N Y A2 A1
X0 a_397_297.t2 A2.t0 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t4 B1_N.t0 a_28_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 Y.t2 A2.t1 a_397_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND.t1 A2.t2 a_229_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND.t4 A1.t0 a_229_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_28_297.t1 B1_N.t1 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 Y.t0 a_28_297.t2 a_229_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR.t2 a_28_297.t3 Y.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_297.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_229_47.t2 a_28_297.t4 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t4 a_28_297.t5 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X11 a_229_47.t0 A2.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_229_47.t4 A1.t2 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR.t3 A1.t3 a_397_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A2.n0 A2.t0 212.081
R1 A2.n1 A2.t1 212.081
R2 A2 A2.n2 157.44
R3 A2.n0 A2.t3 139.78
R4 A2.n1 A2.t2 139.78
R5 A2.n2 A2.n0 30.6732
R6 A2.n2 A2.n1 30.6732
R7 Y.n2 Y.n1 348.635
R8 Y.n2 Y.n0 235.773
R9 Y Y.n3 218.894
R10 Y.n1 Y.t3 26.5955
R11 Y.n1 Y.t2 26.5955
R12 Y.n0 Y.t5 26.5955
R13 Y.n0 Y.t4 26.5955
R14 Y.n3 Y.t1 24.9236
R15 Y.n3 Y.t0 24.9236
R16 Y Y.n2 4.26717
R17 a_397_297.n0 a_397_297.t1 403.692
R18 a_397_297.n0 a_397_297.t0 301.301
R19 a_397_297.n1 a_397_297.n0 184.905
R20 a_397_297.n1 a_397_297.t3 26.5955
R21 a_397_297.t2 a_397_297.n1 26.5955
R22 VPB.t6 VPB.t1 556.386
R23 VPB.t3 VPB.t5 287.072
R24 VPB.t4 VPB.t0 248.599
R25 VPB.t2 VPB.t4 248.599
R26 VPB.t1 VPB.t2 248.599
R27 VPB.t5 VPB.t6 248.599
R28 VPB VPB.t3 195.327
R29 B1_N B1_N.n0 160.145
R30 B1_N.n0 B1_N.t0 140.101
R31 B1_N.n0 B1_N.t1 124.035
R32 a_28_297.t0 a_28_297.n3 710.439
R33 a_28_297.n3 a_28_297.t1 250.365
R34 a_28_297.n2 a_28_297.t5 242.754
R35 a_28_297.n1 a_28_297.t3 212.081
R36 a_28_297.n0 a_28_297.t4 201.125
R37 a_28_297.n3 a_28_297.n2 181.365
R38 a_28_297.n0 a_28_297.t2 139.78
R39 a_28_297.n2 a_28_297.n1 30.6732
R40 a_28_297.n1 a_28_297.n0 14.6066
R41 VPWR.n4 VPWR.t2 344.889
R42 VPWR.n3 VPWR.n2 316.553
R43 VPWR.n6 VPWR.n1 313.75
R44 VPWR.n1 VPWR.t4 96.1553
R45 VPWR.n2 VPWR.t0 26.5955
R46 VPWR.n2 VPWR.t3 26.5955
R47 VPWR.n1 VPWR.t1 25.6105
R48 VPWR.n5 VPWR.n4 24.0946
R49 VPWR.n6 VPWR.n5 17.6946
R50 VPWR.n5 VPWR.n0 9.3005
R51 VPWR.n7 VPWR.n6 7.37348
R52 VPWR.n4 VPWR.n3 7.26177
R53 VPWR.n3 VPWR.n0 0.167133
R54 VPWR.n7 VPWR.n0 0.145304
R55 VPWR VPWR.n7 0.118099
R56 a_229_47.t3 a_229_47.n3 185.225
R57 a_229_47.n1 a_229_47.t4 171.256
R58 a_229_47.n1 a_229_47.n0 98.982
R59 a_229_47.n3 a_229_47.n2 88.3446
R60 a_229_47.n3 a_229_47.n1 48.9326
R61 a_229_47.n2 a_229_47.t1 24.9236
R62 a_229_47.n2 a_229_47.t2 24.9236
R63 a_229_47.n0 a_229_47.t5 24.9236
R64 a_229_47.n0 a_229_47.t0 24.9236
R65 VGND.n12 VGND.t2 266.866
R66 VGND.n3 VGND.n2 217.615
R67 VGND.n5 VGND.n4 207.965
R68 VGND.n6 VGND.n5 34.6358
R69 VGND.n6 VGND.n1 34.6358
R70 VGND.n10 VGND.n1 34.6358
R71 VGND.n11 VGND.n10 34.6358
R72 VGND.n12 VGND.n11 32.0005
R73 VGND.n4 VGND.t0 24.9236
R74 VGND.n4 VGND.t1 24.9236
R75 VGND.n2 VGND.t3 24.9236
R76 VGND.n2 VGND.t4 24.9236
R77 VGND.n13 VGND.n12 11.9358
R78 VGND.n7 VGND.n6 9.3005
R79 VGND.n8 VGND.n1 9.3005
R80 VGND.n10 VGND.n9 9.3005
R81 VGND.n11 VGND.n0 9.3005
R82 VGND.n5 VGND.n3 7.15882
R83 VGND.n7 VGND.n3 0.589543
R84 VGND.n8 VGND.n7 0.120292
R85 VGND.n9 VGND.n8 0.120292
R86 VGND.n9 VGND.n0 0.120292
R87 VGND.n13 VGND.n0 0.120292
R88 VGND VGND.n13 0.0226354
R89 VNB.t4 VNB.t3 2862.14
R90 VNB.t6 VNB.t5 1196.12
R91 VNB.t0 VNB.t6 1196.12
R92 VNB.t1 VNB.t0 1196.12
R93 VNB.t2 VNB.t1 1196.12
R94 VNB.t3 VNB.t2 1196.12
R95 VNB VNB.t4 939.807
R96 A1.n0 A1.t1 212.081
R97 A1.n1 A1.t3 212.081
R98 A1 A1.n2 155.84
R99 A1.n0 A1.t2 139.78
R100 A1.n1 A1.t0 139.78
R101 A1.n2 A1.n1 38.7066
R102 A1.n2 A1.n0 22.6399
C0 Y VGND 0.0115f
C1 VPWR VGND 0.081288f
C2 VPB A2 0.057933f
C3 VPB B1_N 0.043887f
C4 VPB A1 0.058332f
C5 VPB Y 0.016573f
C6 VPB VPWR 0.110807f
C7 A2 A1 0.071165f
C8 VPB VGND 0.010723f
C9 A2 Y 0.102058f
C10 B1_N Y 0.001034f
C11 A2 VPWR 0.020263f
C12 A1 Y 9.56e-19
C13 VPWR B1_N 0.010231f
C14 A2 VGND 0.030584f
C15 B1_N VGND 0.037965f
C16 A1 VPWR 0.043335f
C17 VPWR Y 0.172769f
C18 A1 VGND 0.030808f
C19 VGND VNB 0.523474f
C20 Y VNB 0.015429f
C21 B1_N VNB 0.149047f
C22 VPWR VNB 0.415751f
C23 A1 VNB 0.207848f
C24 A2 VNB 0.173371f
C25 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21bai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21bai_1 VPB VNB VPWR VGND A1 B1_N Y A2
X0 a_388_297.t1 A2.t0 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352.t1 B1_N.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47.t2 a_105_352.t2 Y.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47.t1 A1.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t1 A1.t1 a_388_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND.t1 A2.t1 a_297_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR.t0 B1_N.t1 a_105_352.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y.t1 a_105_352.t3 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
R0 A2.n0 A2.t0 241.536
R1 A2 A2.n0 171.81
R2 A2.n0 A2.t1 169.237
R3 Y Y.n0 591.893
R4 Y.n1 Y.t0 299.318
R5 Y.n1 Y.n0 289.192
R6 Y.n0 Y.t1 33.4905
R7 Y.n0 Y.t2 26.5955
R8 Y Y.n1 13.1191
R9 a_388_297.t0 a_388_297.t1 50.2355
R10 VPB VPB.t3 423.209
R11 VPB.t3 VPB.t1 325.546
R12 VPB.t1 VPB.t2 269.315
R13 VPB.t2 VPB.t0 239.72
R14 B1_N.n0 B1_N.t1 300.983
R15 B1_N B1_N.n0 165.153
R16 B1_N.n0 B1_N.t0 132.282
R17 VGND.n1 VGND.t0 261.486
R18 VGND.n1 VGND.n0 215.381
R19 VGND.n0 VGND.t2 24.9236
R20 VGND.n0 VGND.t1 24.9236
R21 VGND VGND.n1 0.065416
R22 a_105_352.t0 a_105_352.n1 691.898
R23 a_105_352.n1 a_105_352.t1 250.345
R24 a_105_352.n1 a_105_352.n0 222.109
R25 a_105_352.n0 a_105_352.t3 212.081
R26 a_105_352.n0 a_105_352.t2 139.78
R27 VNB.t0 VNB.t3 2677.02
R28 VNB.t3 VNB.t1 1310.03
R29 VNB.t1 VNB.t2 1196.12
R30 VNB VNB.t0 925.567
R31 a_297_47.n0 a_297_47.t1 287.736
R32 a_297_47.n0 a_297_47.t2 31.3851
R33 a_297_47.t0 a_297_47.n0 25.8467
R34 A1.n0 A1.t1 234.804
R35 A1.n0 A1.t0 162.504
R36 A1 A1.n0 155.963
R37 VPWR.n1 VPWR.n0 331.12
R38 VPWR.n1 VPWR.t1 249.058
R39 VPWR.n0 VPWR.t0 101.528
R40 VPWR.n0 VPWR.t2 43.3144
R41 VPWR VPWR.n1 0.348665
C0 B1_N VGND 0.055241f
C1 A2 Y 0.052594f
C2 A1 VPWR 0.053335f
C3 A2 VGND 0.015186f
C4 A1 Y 0.004082f
C5 A1 VGND 0.014794f
C6 VPWR Y 0.153593f
C7 VPB B1_N 0.143535f
C8 VPWR VGND 0.057787f
C9 VPB A2 0.026254f
C10 Y VGND 0.03965f
C11 VPB A1 0.034048f
C12 A2 A1 0.07506f
C13 VPB VPWR 0.075403f
C14 B1_N VPWR 0.070917f
C15 VPB Y 0.006653f
C16 A2 VPWR 0.024707f
C17 VPB VGND 0.007193f
C18 B1_N Y 0.004901f
C19 VGND VNB 0.383651f
C20 Y VNB 0.018294f
C21 VPWR VNB 0.326522f
C22 A1 VNB 0.1335f
C23 A2 VNB 0.090367f
C24 B1_N VNB 0.231947f
C25 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ba_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_4 VNB VPB VGND VPWR B1_N X A2 A1
X0 VPWR.t4 B1_N.t0 a_27_297.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.38 ps=2.76 w=1 l=0.15
X1 VPWR.t0 A1.t0 a_743_297.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_743_297.t2 A1.t1 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_575_47.t3 a_27_297.t2 a_187_21.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_743_297.t0 A2.t0 a_187_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t2 a_27_297.t3 a_187_21.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_187_21.t1 A2.t1 a_743_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_187_21.t2 a_27_297.t4 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_187_21.t4 a_27_297.t5 a_575_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VGND.t0 B1_N.t1 a_27_297.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.91 w=0.65 l=0.15
X10 VGND.t6 A2.t2 a_575_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t5 a_187_21.t6 X.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t8 A1.t2 a_575_47.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t2 a_187_21.t7 X.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 X.t2 a_187_21.t8 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t7 a_187_21.t9 X.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_575_47.t4 A1.t3 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_575_47.t1 A2.t3 VGND.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 X.t0 a_187_21.t10 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X.t6 a_187_21.t11 VGND.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 X.t5 a_187_21.t12 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t3 a_187_21.t13 X.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B1_N.n0 B1_N.t0 241.536
R1 B1_N.n0 B1_N.t1 169.237
R2 B1_N B1_N.n0 156.851
R3 a_27_297.n3 a_27_297.n2 381.623
R4 a_27_297.n2 a_27_297.t4 252.977
R5 a_27_297.t0 a_27_297.n3 226.135
R6 a_27_297.n1 a_27_297.t3 212.081
R7 a_27_297.n0 a_27_297.t2 201.125
R8 a_27_297.n3 a_27_297.t1 191.101
R9 a_27_297.n0 a_27_297.t5 139.78
R10 a_27_297.n2 a_27_297.n1 20.449
R11 a_27_297.n1 a_27_297.n0 14.6066
R12 VPWR.n8 VPWR.t2 845.178
R13 VPWR.n16 VPWR.n1 601.292
R14 VPWR.n14 VPWR.n3 601.292
R15 VPWR.n5 VPWR.n4 601.292
R16 VPWR.n7 VPWR.n6 316.76
R17 VPWR.n1 VPWR.t8 26.5955
R18 VPWR.n1 VPWR.t4 26.5955
R19 VPWR.n3 VPWR.t6 26.5955
R20 VPWR.n3 VPWR.t7 26.5955
R21 VPWR.n4 VPWR.t3 26.5955
R22 VPWR.n4 VPWR.t5 26.5955
R23 VPWR.n6 VPWR.t1 26.5955
R24 VPWR.n6 VPWR.t0 26.5955
R25 VPWR.n9 VPWR.n5 25.977
R26 VPWR.n15 VPWR.n14 24.4711
R27 VPWR.n14 VPWR.n13 19.9534
R28 VPWR.n13 VPWR.n5 18.4476
R29 VPWR.n9 VPWR.n8 15.8123
R30 VPWR.n16 VPWR.n15 13.9299
R31 VPWR.n10 VPWR.n9 9.3005
R32 VPWR.n11 VPWR.n5 9.3005
R33 VPWR.n13 VPWR.n12 9.3005
R34 VPWR.n14 VPWR.n2 9.3005
R35 VPWR.n15 VPWR.n0 9.3005
R36 VPWR.n8 VPWR.n7 7.58106
R37 VPWR.n17 VPWR.n16 7.52093
R38 VPWR.n10 VPWR.n7 0.167193
R39 VPWR.n17 VPWR.n0 0.143429
R40 VPWR.n11 VPWR.n10 0.120292
R41 VPWR.n12 VPWR.n11 0.120292
R42 VPWR.n12 VPWR.n2 0.120292
R43 VPWR.n2 VPWR.n0 0.120292
R44 VPWR VPWR.n17 0.119998
R45 VPB.t5 VPB.t1 556.386
R46 VPB VPB.t6 263.397
R47 VPB.t2 VPB.t3 248.599
R48 VPB.t0 VPB.t2 248.599
R49 VPB.t1 VPB.t0 248.599
R50 VPB.t4 VPB.t5 248.599
R51 VPB.t7 VPB.t4 248.599
R52 VPB.t8 VPB.t7 248.599
R53 VPB.t9 VPB.t8 248.599
R54 VPB.t10 VPB.t9 248.599
R55 VPB.t6 VPB.t10 248.599
R56 A1.n0 A1.t1 212.081
R57 A1.n1 A1.t0 212.081
R58 A1 A1.n2 152.779
R59 A1.n0 A1.t3 139.78
R60 A1.n1 A1.t2 139.78
R61 A1.n2 A1.n1 38.7066
R62 A1.n2 A1.n0 22.6399
R63 a_743_297.n1 a_743_297.t1 907.087
R64 a_743_297.t2 a_743_297.n1 301.301
R65 a_743_297.n1 a_743_297.n0 184.905
R66 a_743_297.n0 a_743_297.t3 26.5955
R67 a_743_297.n0 a_743_297.t0 26.5955
R68 a_187_21.n10 a_187_21.n0 338.336
R69 a_187_21.n11 a_187_21.n10 335.945
R70 a_187_21.n4 a_187_21.t6 212.081
R71 a_187_21.n5 a_187_21.t8 212.081
R72 a_187_21.n2 a_187_21.t9 212.081
R73 a_187_21.n1 a_187_21.t10 212.081
R74 a_187_21.n9 a_187_21.n8 185
R75 a_187_21.n7 a_187_21.n3 173.761
R76 a_187_21.n7 a_187_21.n6 152
R77 a_187_21.n4 a_187_21.t13 139.78
R78 a_187_21.n5 a_187_21.t12 139.78
R79 a_187_21.n2 a_187_21.t7 139.78
R80 a_187_21.n1 a_187_21.t11 139.78
R81 a_187_21.n9 a_187_21.n7 101.632
R82 a_187_21.n10 a_187_21.n9 69.9424
R83 a_187_21.n2 a_187_21.n1 61.346
R84 a_187_21.n3 a_187_21.n2 54.0429
R85 a_187_21.n6 a_187_21.n5 42.3581
R86 a_187_21.n0 a_187_21.t0 26.5955
R87 a_187_21.n0 a_187_21.t1 26.5955
R88 a_187_21.t3 a_187_21.n11 26.5955
R89 a_187_21.n11 a_187_21.t2 26.5955
R90 a_187_21.n8 a_187_21.t5 24.9236
R91 a_187_21.n8 a_187_21.t4 24.9236
R92 a_187_21.n6 a_187_21.n4 18.9884
R93 a_187_21.n5 a_187_21.n3 7.30353
R94 a_575_47.n2 a_575_47.t2 316.983
R95 a_575_47.n1 a_575_47.t4 171.256
R96 a_575_47.n1 a_575_47.n0 98.982
R97 a_575_47.n3 a_575_47.n2 88.3446
R98 a_575_47.n2 a_575_47.n1 48.9326
R99 a_575_47.n0 a_575_47.t5 24.9236
R100 a_575_47.n0 a_575_47.t1 24.9236
R101 a_575_47.n3 a_575_47.t0 24.9236
R102 a_575_47.t3 a_575_47.n3 24.9236
R103 VNB.t5 VNB.t2 2677.02
R104 VNB VNB.t4 1267.31
R105 VNB.t10 VNB.t9 1196.12
R106 VNB.t1 VNB.t10 1196.12
R107 VNB.t0 VNB.t1 1196.12
R108 VNB.t3 VNB.t0 1196.12
R109 VNB.t2 VNB.t3 1196.12
R110 VNB.t6 VNB.t5 1196.12
R111 VNB.t8 VNB.t6 1196.12
R112 VNB.t7 VNB.t8 1196.12
R113 VNB.t4 VNB.t7 1196.12
R114 A2.n0 A2.t0 212.081
R115 A2.n1 A2.t1 212.081
R116 A2 A2.n2 152.678
R117 A2.n0 A2.t3 139.78
R118 A2.n1 A2.t2 139.78
R119 A2.n2 A2.n0 30.6732
R120 A2.n2 A2.n1 30.6732
R121 VGND.n4 VGND.t3 286.426
R122 VGND.n10 VGND.n9 219.685
R123 VGND.n8 VGND.n7 207.965
R124 VGND.n19 VGND.n3 207.965
R125 VGND.n1 VGND.n0 121.453
R126 VGND.n13 VGND.n6 34.6358
R127 VGND.n14 VGND.n13 34.6358
R128 VGND.n15 VGND.n14 34.6358
R129 VGND.n21 VGND.n20 34.6358
R130 VGND.n19 VGND.n18 32.377
R131 VGND.n18 VGND.n4 30.8711
R132 VGND.n8 VGND.n6 26.3534
R133 VGND.n21 VGND.n1 26.3534
R134 VGND.n9 VGND.t7 24.9236
R135 VGND.n9 VGND.t8 24.9236
R136 VGND.n7 VGND.t5 24.9236
R137 VGND.n7 VGND.t6 24.9236
R138 VGND.n3 VGND.t4 24.9236
R139 VGND.n3 VGND.t2 24.9236
R140 VGND.n0 VGND.t1 24.9236
R141 VGND.n0 VGND.t0 24.9236
R142 VGND.n23 VGND.n1 15.9414
R143 VGND.n10 VGND.n8 15.1733
R144 VGND.n11 VGND.n6 9.3005
R145 VGND.n13 VGND.n12 9.3005
R146 VGND.n14 VGND.n5 9.3005
R147 VGND.n16 VGND.n15 9.3005
R148 VGND.n18 VGND.n17 9.3005
R149 VGND.n20 VGND.n2 9.3005
R150 VGND.n22 VGND.n21 9.3005
R151 VGND.n15 VGND.n4 3.76521
R152 VGND.n20 VGND.n19 2.25932
R153 VGND.n11 VGND.n10 0.857451
R154 VGND.n23 VGND.n22 0.141672
R155 VGND VGND.n23 0.121778
R156 VGND.n12 VGND.n11 0.120292
R157 VGND.n12 VGND.n5 0.120292
R158 VGND.n16 VGND.n5 0.120292
R159 VGND.n17 VGND.n16 0.120292
R160 VGND.n17 VGND.n2 0.120292
R161 VGND.n22 VGND.n2 0.120292
R162 X.n2 X.n0 614.785
R163 X.n2 X.n1 586.441
R164 X X.n6 186.358
R165 X.n6 X.n5 185
R166 X.n4 X.n3 98.3961
R167 X.n5 X.n4 34.5864
R168 X.n1 X.t1 26.5955
R169 X.n1 X.t0 26.5955
R170 X.n0 X.t3 26.5955
R171 X.n0 X.t2 26.5955
R172 X.n6 X.t4 24.9236
R173 X.n6 X.t5 24.9236
R174 X.n3 X.t7 24.9236
R175 X.n3 X.t6 24.9236
R176 X.n4 X.n2 24.3205
R177 X X.n5 11.8308
C0 X VGND 0.26017f
C1 VPWR B1_N 0.020565f
C2 X VPB 0.005674f
C3 VGND VPB 0.010368f
C4 X B1_N 0.053065f
C5 VGND B1_N 0.034605f
C6 VPB B1_N 0.032459f
C7 A2 A1 0.071165f
C8 A2 VPWR 0.019235f
C9 A1 VPWR 0.038443f
C10 A2 VGND 0.028567f
C11 A2 VPB 0.057831f
C12 A1 VGND 0.029007f
C13 VPWR X 0.0315f
C14 A1 VPB 0.061266f
C15 VPWR VGND 0.117298f
C16 VPWR VPB 0.122933f
C17 VGND VNB 0.679566f
C18 X VNB 0.009062f
C19 VPWR VNB 0.555182f
C20 A1 VNB 0.209776f
C21 A2 VNB 0.172798f
C22 B1_N VNB 0.118957f
C23 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21bai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21bai_4 VNB VPB VGND VPWR A2 A1 B1_N Y
X0 Y.t11 a_33_297.t2 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47.t9 a_33_297.t3 Y.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t5 a_33_297.t4 Y.t10 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297.t0 B1_N.t0 VGND.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y.t9 a_33_297.t5 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t0 A2.t0 a_561_297.t5 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y.t6 a_33_297.t6 a_225_47.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y.t5 a_33_297.t7 a_225_47.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND.t6 A2.t1 a_225_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t3 A2.t2 a_225_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_225_47.t6 a_33_297.t8 Y.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_225_47.t1 A1.t0 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_225_47.t3 A2.t3 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_225_47.t4 A2.t4 VGND.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t1 A1.t1 a_561_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_561_297.t0 A1.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR.t2 B1_N.t1 a_33_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X17 a_561_297.t4 A2.t5 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t2 A2.t6 a_561_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t1 A1.t3 a_225_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_561_297.t2 A2.t7 Y.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR.t3 a_33_297.t9 Y.t8 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 a_33_297.t1 a_33_297.n13 269.899
R1 a_33_297.n11 a_33_297.t5 225.226
R2 a_33_297.n3 a_33_297.t9 212.081
R3 a_33_297.n1 a_33_297.t2 212.081
R4 a_33_297.n10 a_33_297.t4 212.081
R5 a_33_297.n2 a_33_297.t8 201.125
R6 a_33_297.n6 a_33_297.n5 172.725
R7 a_33_297.n13 a_33_297.t0 154.901
R8 a_33_297.n12 a_33_297.n11 152
R9 a_33_297.n9 a_33_297.n0 152
R10 a_33_297.n7 a_33_297.n6 152
R11 a_33_297.n8 a_33_297.t6 139.78
R12 a_33_297.n4 a_33_297.t3 139.78
R13 a_33_297.n2 a_33_297.t7 139.78
R14 a_33_297.n11 a_33_297.n10 48.2005
R15 a_33_297.n8 a_33_297.n7 36.5157
R16 a_33_297.n5 a_33_297.n4 24.8308
R17 a_33_297.n5 a_33_297.n3 21.9096
R18 a_33_297.n6 a_33_297.n0 20.7243
R19 a_33_297.n12 a_33_297.n0 20.7243
R20 a_33_297.n3 a_33_297.n2 14.6066
R21 a_33_297.n4 a_33_297.n1 14.6066
R22 a_33_297.n13 a_33_297.n12 13.41
R23 a_33_297.n9 a_33_297.n8 13.146
R24 a_33_297.n7 a_33_297.n1 10.2247
R25 a_33_297.n10 a_33_297.n9 1.46111
R26 VPWR.n4 VPWR.t3 344.889
R27 VPWR.n6 VPWR.n5 326.454
R28 VPWR.n11 VPWR.n1 323.192
R29 VPWR.n9 VPWR.n3 318.293
R30 VPWR.n9 VPWR.n8 28.2358
R31 VPWR.n1 VPWR.t4 26.5955
R32 VPWR.n1 VPWR.t2 26.5955
R33 VPWR.n3 VPWR.t6 26.5955
R34 VPWR.n3 VPWR.t5 26.5955
R35 VPWR.n5 VPWR.t0 26.5955
R36 VPWR.n5 VPWR.t1 26.5955
R37 VPWR.n10 VPWR.n9 22.2123
R38 VPWR.n11 VPWR.n10 22.2123
R39 VPWR.n8 VPWR.n4 16.1887
R40 VPWR.n8 VPWR.n7 9.3005
R41 VPWR.n9 VPWR.n2 9.3005
R42 VPWR.n10 VPWR.n0 9.3005
R43 VPWR.n6 VPWR.n4 7.58767
R44 VPWR.n12 VPWR.n11 7.54776
R45 VPWR.n7 VPWR.n6 0.148358
R46 VPWR.n12 VPWR.n0 0.143088
R47 VPWR VPWR.n12 0.120344
R48 VPWR.n7 VPWR.n2 0.120292
R49 VPWR.n2 VPWR.n0 0.120292
R50 Y.n2 Y.n0 343.096
R51 Y.n2 Y.n1 301.14
R52 Y.n5 Y.n3 255.446
R53 Y.n9 Y.n7 243.353
R54 Y.n5 Y.n4 208.507
R55 Y.n9 Y.n8 185
R56 Y Y.n9 29.7249
R57 Y.n3 Y.t10 26.5955
R58 Y.n3 Y.t9 26.5955
R59 Y.n4 Y.t8 26.5955
R60 Y.n4 Y.t11 26.5955
R61 Y.n0 Y.t1 26.5955
R62 Y.n0 Y.t2 26.5955
R63 Y.n1 Y.t3 26.5955
R64 Y.n1 Y.t0 26.5955
R65 Y.n6 Y.n5 24.9898
R66 Y.n8 Y.t4 24.9236
R67 Y.n8 Y.t5 24.9236
R68 Y.n7 Y.t7 24.9236
R69 Y.n7 Y.t6 24.9236
R70 Y.n6 Y.n2 23.4672
R71 Y Y.n6 2.5605
R72 VPB.t7 VPB.t0 556.386
R73 VPB.t2 VPB.t1 248.599
R74 VPB.t3 VPB.t2 248.599
R75 VPB.t4 VPB.t3 248.599
R76 VPB.t5 VPB.t4 248.599
R77 VPB.t0 VPB.t5 248.599
R78 VPB.t10 VPB.t7 248.599
R79 VPB.t9 VPB.t10 248.599
R80 VPB.t8 VPB.t9 248.599
R81 VPB.t6 VPB.t8 248.599
R82 VPB VPB.t6 221.964
R83 a_225_47.t8 a_225_47.n7 326.709
R84 a_225_47.n7 a_225_47.n6 185
R85 a_225_47.n1 a_225_47.t1 173.059
R86 a_225_47.n1 a_225_47.n0 98.982
R87 a_225_47.n3 a_225_47.n2 98.982
R88 a_225_47.n5 a_225_47.n4 88.3446
R89 a_225_47.n7 a_225_47.n5 65.1609
R90 a_225_47.n5 a_225_47.n3 48.9326
R91 a_225_47.n3 a_225_47.n1 36.2672
R92 a_225_47.n6 a_225_47.t7 24.9236
R93 a_225_47.n6 a_225_47.t9 24.9236
R94 a_225_47.n4 a_225_47.t5 24.9236
R95 a_225_47.n4 a_225_47.t6 24.9236
R96 a_225_47.n0 a_225_47.t0 24.9236
R97 a_225_47.n0 a_225_47.t4 24.9236
R98 a_225_47.n2 a_225_47.t2 24.9236
R99 a_225_47.n2 a_225_47.t3 24.9236
R100 VNB.t5 VNB.t9 2677.02
R101 VNB.t0 VNB.t1 1196.12
R102 VNB.t4 VNB.t0 1196.12
R103 VNB.t2 VNB.t4 1196.12
R104 VNB.t3 VNB.t2 1196.12
R105 VNB.t6 VNB.t3 1196.12
R106 VNB.t7 VNB.t6 1196.12
R107 VNB.t8 VNB.t7 1196.12
R108 VNB.t10 VNB.t8 1196.12
R109 VNB.t9 VNB.t10 1196.12
R110 VNB VNB.t5 1067.96
R111 B1_N.n0 B1_N.t1 232.738
R112 B1_N B1_N.n0 166.934
R113 B1_N.n0 B1_N.t0 160.438
R114 VGND.n8 VGND.n7 219.567
R115 VGND.n9 VGND.n6 207.965
R116 VGND.n4 VGND.n3 207.965
R117 VGND.n22 VGND.t0 157.993
R118 VGND.n11 VGND.n10 34.6358
R119 VGND.n15 VGND.n14 34.6358
R120 VGND.n16 VGND.n15 34.6358
R121 VGND.n16 VGND.n1 34.6358
R122 VGND.n20 VGND.n1 34.6358
R123 VGND.n21 VGND.n20 34.6358
R124 VGND.n22 VGND.n21 28.6123
R125 VGND.n14 VGND.n4 27.1064
R126 VGND.n7 VGND.t2 24.9236
R127 VGND.n7 VGND.t1 24.9236
R128 VGND.n6 VGND.t5 24.9236
R129 VGND.n6 VGND.t3 24.9236
R130 VGND.n3 VGND.t4 24.9236
R131 VGND.n3 VGND.t6 24.9236
R132 VGND.n10 VGND.n9 21.0829
R133 VGND.n9 VGND.n8 20.2741
R134 VGND.n23 VGND.n22 15.324
R135 VGND.n10 VGND.n5 9.3005
R136 VGND.n12 VGND.n11 9.3005
R137 VGND.n14 VGND.n13 9.3005
R138 VGND.n15 VGND.n2 9.3005
R139 VGND.n17 VGND.n16 9.3005
R140 VGND.n18 VGND.n1 9.3005
R141 VGND.n20 VGND.n19 9.3005
R142 VGND.n21 VGND.n0 9.3005
R143 VGND.n11 VGND.n4 7.52991
R144 VGND.n8 VGND.n5 1.02717
R145 VGND.n12 VGND.n5 0.120292
R146 VGND.n13 VGND.n12 0.120292
R147 VGND.n13 VGND.n2 0.120292
R148 VGND.n17 VGND.n2 0.120292
R149 VGND.n18 VGND.n17 0.120292
R150 VGND.n19 VGND.n18 0.120292
R151 VGND.n19 VGND.n0 0.120292
R152 VGND.n23 VGND.n0 0.120292
R153 VGND VGND.n23 0.0226354
R154 A2.n3 A2.t5 212.081
R155 A2.n5 A2.t6 212.081
R156 A2.n7 A2.t7 212.081
R157 A2.n1 A2.t0 212.081
R158 A2.n4 A2.n0 173.761
R159 A2.n9 A2.n2 173.761
R160 A2.n6 A2.n0 152
R161 A2.n9 A2.n8 152
R162 A2.n3 A2.t4 139.78
R163 A2.n5 A2.t2 139.78
R164 A2.n7 A2.t3 139.78
R165 A2.n1 A2.t1 139.78
R166 A2.n8 A2.n6 49.6611
R167 A2.n7 A2.n2 48.2005
R168 A2.n5 A2.n4 39.4369
R169 A2.n4 A2.n3 21.9096
R170 A2 A2.n9 16.3205
R171 A2.n2 A2.n1 13.146
R172 A2.n6 A2.n5 10.2247
R173 A2 A2.n0 5.4405
R174 A2.n8 A2.n7 1.46111
R175 a_561_297.n1 a_561_297.t5 371.01
R176 a_561_297.n1 a_561_297.n0 300.885
R177 a_561_297.n2 a_561_297.t0 300.527
R178 a_561_297.n3 a_561_297.n2 187.506
R179 a_561_297.n2 a_561_297.n1 65.4262
R180 a_561_297.n0 a_561_297.t3 26.5955
R181 a_561_297.n0 a_561_297.t2 26.5955
R182 a_561_297.n3 a_561_297.t1 26.5955
R183 a_561_297.t4 a_561_297.n3 26.5955
R184 A1.n6 A1.n4 212.081
R185 A1.n3 A1.n1 212.081
R186 A1.n10 A1.t2 212.081
R187 A1.n12 A1.t1 212.081
R188 A1.n8 A1.n7 172.725
R189 A1 A1.n13 171.81
R190 A1.n9 A1.n8 152
R191 A1.n11 A1.n0 152
R192 A1.n6 A1.n5 139.78
R193 A1.n3 A1.n2 139.78
R194 A1.n10 A1.t0 139.78
R195 A1.n12 A1.t3 139.78
R196 A1.n13 A1.n11 49.6611
R197 A1.n10 A1.n9 46.7399
R198 A1.n7 A1.n3 35.055
R199 A1.n7 A1.n6 26.2914
R200 A1.n8 A1.n0 20.7243
R201 A1.n9 A1.n3 14.6066
R202 A1.n13 A1.n12 8.76414
R203 A1.n11 A1.n10 2.92171
R204 A1 A1.n0 0.914786
C0 Y VGND 0.025861f
C1 VPB B1_N 0.036636f
C2 VPB A2 0.120104f
C3 VPB VPWR 0.144968f
C4 VPB A1 0.147882f
C5 B1_N VPWR 0.017721f
C6 VPB Y 0.023337f
C7 A2 VPWR 0.034611f
C8 VPB VGND 0.011588f
C9 B1_N Y 3.37e-19
C10 A2 A1 0.068563f
C11 A1 VPWR 0.110511f
C12 B1_N VGND 0.042692f
C13 A2 Y 0.186533f
C14 VPWR Y 0.374864f
C15 A2 VGND 0.053334f
C16 A1 Y 0.00215f
C17 VPWR VGND 0.134064f
C18 A1 VGND 0.065156f
C19 VGND VNB 0.802067f
C20 Y VNB 0.016124f
C21 VPWR VNB 0.630025f
C22 A1 VNB 0.441025f
C23 A2 VNB 0.352617f
C24 B1_N VNB 0.144077f
C25 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199.t3 B1.t0 a_215_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR.t1 A1.t0 a_493_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297.t0 A2.t0 a_78_199.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR.t0 a_78_199.t4 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND.t0 A2.t1 a_215_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199.t2 B2.t0 a_292_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47.t1 A1.t1 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47.t2 B2.t1 a_78_199.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297.t1 B1.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND.t1 a_78_199.t5 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n0 B1.t1 1578.82
R1 B1.n0 B1.t0 157.453
R2 B1 B1.n0 157.376
R3 a_215_47.n0 a_215_47.t3 323.712
R4 a_215_47.n0 a_215_47.t1 183.446
R5 a_215_47.n1 a_215_47.n0 89.3175
R6 a_215_47.n1 a_215_47.t2 39.6928
R7 a_215_47.t0 a_215_47.n1 24.9236
R8 a_78_199.n3 a_78_199.n2 278.697
R9 a_78_199.n2 a_78_199.n0 255.142
R10 a_78_199.n1 a_78_199.t4 230.363
R11 a_78_199.n1 a_78_199.t5 158.064
R12 a_78_199.n2 a_78_199.n1 152
R13 a_78_199.t1 a_78_199.n3 65.9955
R14 a_78_199.n3 a_78_199.t2 26.5955
R15 a_78_199.n0 a_78_199.t0 24.9236
R16 a_78_199.n0 a_78_199.t3 24.9236
R17 VNB.t3 VNB.t4 2677.02
R18 VNB.t2 VNB.t0 1423.95
R19 VNB.t0 VNB.t1 1196.12
R20 VNB.t4 VNB.t2 1196.12
R21 VNB VNB.t3 925.567
R22 A1.n0 A1.t0 235.471
R23 A1.n0 A1.t1 163.172
R24 A1 A1.n0 156.481
R25 a_493_297.t0 a_493_297.t1 41.3705
R26 VPWR.n6 VPWR.n5 292.5
R27 VPWR.n4 VPWR.n3 292.5
R28 VPWR.n2 VPWR.t1 251.44
R29 VPWR.n5 VPWR.n4 89.6355
R30 VPWR.n5 VPWR.t0 30.5355
R31 VPWR.n3 VPWR.n2 30.1305
R32 VPWR.n4 VPWR.t2 26.5955
R33 VPWR.n1 VPWR.n0 9.3005
R34 VPWR.n7 VPWR.n6 7.76924
R35 VPWR.n6 VPWR.n1 5.91878
R36 VPWR.n3 VPWR.n1 0.344586
R37 VPWR.n2 VPWR.n0 0.217659
R38 VPWR.n7 VPWR.n0 0.145522
R39 VPWR VPWR.n7 0.117878
R40 VPB.t0 VPB.t4 529.751
R41 VPB.t3 VPB.t1 366.978
R42 VPB.t4 VPB.t3 227.882
R43 VPB.t1 VPB.t2 213.084
R44 VPB VPB.t0 204.207
R45 A2.n0 A2.t0 239.505
R46 A2 A2.n0 184.407
R47 A2.n0 A2.t1 167.204
R48 X X.n0 593
R49 X.n1 X.n0 288.666
R50 X.n1 X.t1 264.45
R51 X.n0 X.t0 26.5955
R52 X X.n1 15.2134
R53 VGND.n1 VGND.t1 297.262
R54 VGND.n1 VGND.n0 213.156
R55 VGND.n0 VGND.t2 24.9236
R56 VGND.n0 VGND.t0 24.9236
R57 VGND VGND.n1 0.152279
R58 B2.n0 B2.t0 241.536
R59 B2.n0 B2.t1 169.237
R60 B2 B2.n0 166.337
R61 a_292_297.t0 a_292_297.t1 46.2955
C0 VGND B1 0.011856f
C1 VPWR B2 0.010367f
C2 A2 A1 0.087859f
C3 VPWR A2 0.120404f
C4 VGND B2 0.010267f
C5 X VPWR 0.091108f
C6 VGND A2 0.015286f
C7 VPWR A1 0.05704f
C8 X VGND 0.047175f
C9 VGND A1 0.014626f
C10 VPWR VGND 0.066763f
C11 VPB B1 0.038762f
C12 VPB B2 0.028066f
C13 VPB A2 0.034104f
C14 B1 B2 0.081466f
C15 X VPB 0.010691f
C16 VPB A1 0.031899f
C17 B1 A2 3.91e-19
C18 VPWR VPB 0.074428f
C19 X B1 6.11e-19
C20 B2 A2 0.06759f
C21 X B2 1.65e-19
C22 VGND VPB 0.005957f
C23 VPWR B1 0.022722f
C24 VGND VNB 0.402531f
C25 VPWR VNB 0.35911f
C26 X VNB 0.088397f
C27 A1 VNB 0.132282f
C28 A2 VNB 0.097054f
C29 B2 VNB 0.091305f
C30 B1 VNB 0.109674f
C31 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_2 VNB VPB VGND VPWR A1 A2 B2 B1 X
X0 a_301_47.t1 B2.t0 a_81_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t0 A2.t0 a_301_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297.t1 B1.t0 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR.t2 a_81_21.t4 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47.t2 A1.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t3 a_81_21.t5 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 X.t2 a_81_21.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X.t0 a_81_21.t7 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR.t0 A1.t1 a_579_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21.t2 B1.t1 a_301_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297.t1 A2.t1 a_81_21.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21.t0 B2.t1 a_383_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
R0 B2.n0 B2.t1 241.536
R1 B2.n0 B2.t0 169.237
R2 B2 B2.n0 166.337
R3 a_81_21.n5 a_81_21.n4 278.94
R4 a_81_21.n4 a_81_21.n0 253.78
R5 a_81_21.n3 a_81_21.t4 212.081
R6 a_81_21.n1 a_81_21.t7 212.081
R7 a_81_21.n4 a_81_21.n3 184.864
R8 a_81_21.n1 a_81_21.t6 141.242
R9 a_81_21.n2 a_81_21.t5 139.78
R10 a_81_21.n5 a_81_21.t3 65.9955
R11 a_81_21.n2 a_81_21.n1 59.8853
R12 a_81_21.t0 a_81_21.n5 26.5955
R13 a_81_21.n0 a_81_21.t1 24.9236
R14 a_81_21.n0 a_81_21.t2 24.9236
R15 a_81_21.n3 a_81_21.n2 1.46111
R16 a_301_47.n0 a_301_47.t3 323.87
R17 a_301_47.n0 a_301_47.t2 199.306
R18 a_301_47.n1 a_301_47.n0 92.501
R19 a_301_47.n1 a_301_47.t1 40.6159
R20 a_301_47.t0 a_301_47.n1 29.539
R21 VNB.t4 VNB.t5 2677.02
R22 VNB.t1 VNB.t0 1509.39
R23 VNB.t0 VNB.t2 1196.12
R24 VNB.t5 VNB.t1 1196.12
R25 VNB.t3 VNB.t4 1196.12
R26 VNB VNB.t3 996.764
R27 A2.n0 A2.t1 239.505
R28 A2 A2.n0 183.944
R29 A2.n0 A2.t0 167.204
R30 VGND.n3 VGND.t3 295.099
R31 VGND.n2 VGND.n1 213.127
R32 VGND.n5 VGND.t2 160.222
R33 VGND.n5 VGND.n4 31.624
R34 VGND.n4 VGND.n3 25.224
R35 VGND.n1 VGND.t1 24.9236
R36 VGND.n1 VGND.t0 24.9236
R37 VGND.n6 VGND.n5 12.3123
R38 VGND.n4 VGND.n0 9.3005
R39 VGND.n3 VGND.n2 7.44449
R40 VGND.n2 VGND.n0 0.15805
R41 VGND.n6 VGND.n0 0.120292
R42 VGND VGND.n6 0.0265417
R43 B1.n0 B1.t0 230.793
R44 B1.n0 B1.t1 158.494
R45 B1 B1.n0 157.376
R46 VPWR.n2 VPWR.t0 346.481
R47 VPWR.n3 VPWR.n1 292.5
R48 VPWR.n5 VPWR.n4 292.5
R49 VPWR.n11 VPWR.t1 252.511
R50 VPWR.n4 VPWR.n3 92.5905
R51 VPWR.n3 VPWR.t2 34.4755
R52 VPWR.n5 VPWR.n2 30.5063
R53 VPWR.n4 VPWR.t3 26.5955
R54 VPWR.n10 VPWR.n9 25.0985
R55 VPWR.n11 VPWR.n10 24.4711
R56 VPWR.n7 VPWR.n6 9.3005
R57 VPWR.n9 VPWR.n8 9.3005
R58 VPWR.n10 VPWR.n0 9.3005
R59 VPWR.n12 VPWR.n11 9.3005
R60 VPWR.n6 VPWR.n1 6.19405
R61 VPWR.n6 VPWR.n5 0.275769
R62 VPWR.n7 VPWR.n2 0.218365
R63 VPWR.n9 VPWR.n1 0.138134
R64 VPWR.n8 VPWR.n7 0.120292
R65 VPWR.n8 VPWR.n0 0.120292
R66 VPWR.n12 VPWR.n0 0.120292
R67 VPWR VPWR.n12 0.0265417
R68 a_383_297.t0 a_383_297.t1 41.3705
R69 VPB.t4 VPB.t5 550.467
R70 VPB.t2 VPB.t0 366.978
R71 VPB.t3 VPB.t4 248.599
R72 VPB.t0 VPB.t1 213.084
R73 VPB.t5 VPB.t2 213.084
R74 VPB VPB.t3 213.084
R75 X X.n0 595.419
R76 X.n2 X.n0 287.526
R77 X.n2 X.n1 255.974
R78 X.n0 X.t1 26.5955
R79 X.n0 X.t0 26.5955
R80 X.n1 X.t3 24.9236
R81 X.n1 X.t2 24.9236
R82 X X.n2 19.7731
R83 A1.n0 A1.t1 235.471
R84 A1.n0 A1.t0 163.172
R85 A1 A1.n0 153.66
R86 a_579_297.t0 a_579_297.t1 41.3705
C0 VPWR X 0.155514f
C1 VPWR VPB 0.088063f
C2 X VPB 0.003521f
C3 VPWR B1 0.022598f
C4 VPWR VGND 0.088636f
C5 VPWR B2 0.011063f
C6 X B1 6.07e-19
C7 VGND VPB 0.00728f
C8 X VGND 0.077934f
C9 VPB B1 0.037367f
C10 VPWR A2 0.09588f
C11 VPB B2 0.027613f
C12 X B2 2.02e-19
C13 VGND B1 0.011669f
C14 VPWR A1 0.05728f
C15 VGND B2 0.01041f
C16 B1 B2 0.085052f
C17 VPB A2 0.03391f
C18 VGND A2 0.015886f
C19 B1 A2 4.07e-19
C20 VPB A1 0.036054f
C21 VGND A1 0.015816f
C22 B2 A2 0.066724f
C23 A2 A1 0.111848f
C24 VGND VNB 0.477071f
C25 X VNB 0.021756f
C26 VPWR VNB 0.424953f
C27 A1 VNB 0.14472f
C28 A2 VNB 0.097645f
C29 B2 VNB 0.091641f
C30 B1 VNB 0.107405f
C31 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_4 VNB VPB VGND VPWR A1 B1 B2 A2 X
X0 VPWR.t1 B1.t0 a_566_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_484_47.t1 B1.t1 a_96_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X.t3 a_96_21.t8 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t4 a_96_21.t9 X.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4 X.t6 a_96_21.t10 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_566_297.t2 B2.t0 a_96_21.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t6 a_96_21.t11 X.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t2 a_96_21.t12 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND.t4 a_96_21.t13 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_96_21.t6 B2.t1 a_566_297.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t3 A1.t0 a_918_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 a_484_47.t6 A1.t1 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_566_297.t0 B1.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X13 a_484_47.t7 B2.t2 a_96_21.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_96_21.t3 A2.t0 a_918_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_918_297.t2 A2.t1 a_96_21.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_484_47.t4 A2.t2 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_918_297.t0 A1.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_96_21.t0 B1.t3 a_484_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 VGND.t1 A2.t3 a_484_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_96_21.t4 B2.t3 a_484_47.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t0 A1.t3 a_484_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X22 X.t4 a_96_21.t14 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND.t3 a_96_21.t15 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B1.n1 B1.t2 241.536
R1 B1.n0 B1.t0 241.536
R2 B1.n2 B1.n0 238.481
R3 B1.n1 B1.t3 169.237
R4 B1.n0 B1.t1 169.237
R5 B1.n2 B1.n1 152
R6 B1 B1.n2 6.87457
R7 a_566_297.n1 a_566_297.n0 1223.84
R8 a_566_297.n0 a_566_297.t1 26.5955
R9 a_566_297.n0 a_566_297.t2 26.5955
R10 a_566_297.n1 a_566_297.t3 26.5955
R11 a_566_297.t0 a_566_297.n1 26.5955
R12 VPWR.n8 VPWR.n7 601.292
R13 VPWR.n14 VPWR.n3 585
R14 VPWR.n16 VPWR.n15 585
R15 VPWR.n24 VPWR.t7 343.351
R16 VPWR.n22 VPWR.n2 316.757
R17 VPWR.n6 VPWR.t3 269.519
R18 VPWR.n15 VPWR.n14 102.441
R19 VPWR.n7 VPWR.t2 42.3555
R20 VPWR.n9 VPWR.n5 34.6358
R21 VPWR.n13 VPWR.n5 34.6358
R22 VPWR.n23 VPWR.n22 27.8593
R23 VPWR.n15 VPWR.t0 26.5955
R24 VPWR.n14 VPWR.t4 26.5955
R25 VPWR.n2 VPWR.t5 26.5955
R26 VPWR.n2 VPWR.t6 26.5955
R27 VPWR.n7 VPWR.t1 26.5955
R28 VPWR.n16 VPWR.n13 26.4476
R29 VPWR.n21 VPWR.n3 24.1887
R30 VPWR.n22 VPWR.n21 22.5887
R31 VPWR.n24 VPWR.n23 16.5652
R32 VPWR.n9 VPWR.n8 14.3064
R33 VPWR.n10 VPWR.n9 9.3005
R34 VPWR.n11 VPWR.n5 9.3005
R35 VPWR.n13 VPWR.n12 9.3005
R36 VPWR.n17 VPWR.n4 9.3005
R37 VPWR.n19 VPWR.n18 9.3005
R38 VPWR.n21 VPWR.n20 9.3005
R39 VPWR.n22 VPWR.n1 9.3005
R40 VPWR.n23 VPWR.n0 9.3005
R41 VPWR.n25 VPWR.n24 9.3005
R42 VPWR.n18 VPWR.n17 8.65932
R43 VPWR.n8 VPWR.n6 7.41157
R44 VPWR.n18 VPWR.n3 0.847559
R45 VPWR.n17 VPWR.n16 0.282853
R46 VPWR.n10 VPWR.n6 0.176425
R47 VPWR.n11 VPWR.n10 0.120292
R48 VPWR.n12 VPWR.n11 0.120292
R49 VPWR.n12 VPWR.n4 0.120292
R50 VPWR.n19 VPWR.n4 0.120292
R51 VPWR.n20 VPWR.n19 0.120292
R52 VPWR.n20 VPWR.n1 0.120292
R53 VPWR.n1 VPWR.n0 0.120292
R54 VPWR.n25 VPWR.n0 0.120292
R55 VPWR VPWR.n25 0.0226354
R56 VPB.t7 VPB.t0 556.386
R57 VPB.t1 VPB.t2 295.95
R58 VPB.t3 VPB.t6 248.599
R59 VPB.t4 VPB.t3 248.599
R60 VPB.t2 VPB.t4 248.599
R61 VPB.t5 VPB.t1 248.599
R62 VPB.t11 VPB.t5 248.599
R63 VPB.t0 VPB.t11 248.599
R64 VPB.t8 VPB.t7 248.599
R65 VPB.t9 VPB.t8 248.599
R66 VPB.t10 VPB.t9 248.599
R67 VPB VPB.t10 242.679
R68 a_96_21.n17 a_96_21.n16 708.106
R69 a_96_21.n16 a_96_21.n15 585
R70 a_96_21.n13 a_96_21.n11 226.355
R71 a_96_21.n1 a_96_21.t9 212.081
R72 a_96_21.n8 a_96_21.t10 212.081
R73 a_96_21.n2 a_96_21.t11 212.081
R74 a_96_21.n3 a_96_21.t14 212.081
R75 a_96_21.n13 a_96_21.n12 185
R76 a_96_21.n5 a_96_21.n4 173.761
R77 a_96_21.n6 a_96_21.n5 152
R78 a_96_21.n7 a_96_21.n0 152
R79 a_96_21.n10 a_96_21.n9 152
R80 a_96_21.n1 a_96_21.t13 139.78
R81 a_96_21.n8 a_96_21.t8 139.78
R82 a_96_21.n2 a_96_21.t15 139.78
R83 a_96_21.n3 a_96_21.t12 139.78
R84 a_96_21.n16 a_96_21.n14 109.216
R85 a_96_21.n14 a_96_21.n13 56.1408
R86 a_96_21.n7 a_96_21.n6 49.6611
R87 a_96_21.n9 a_96_21.n8 48.2005
R88 a_96_21.n4 a_96_21.n2 39.4369
R89 a_96_21.n15 a_96_21.t5 26.5955
R90 a_96_21.n15 a_96_21.t6 26.5955
R91 a_96_21.t2 a_96_21.n17 26.5955
R92 a_96_21.n17 a_96_21.t3 26.5955
R93 a_96_21.n12 a_96_21.t7 24.9236
R94 a_96_21.n12 a_96_21.t0 24.9236
R95 a_96_21.n11 a_96_21.t1 24.9236
R96 a_96_21.n11 a_96_21.t4 24.9236
R97 a_96_21.n4 a_96_21.n3 21.9096
R98 a_96_21.n10 a_96_21.n0 21.7605
R99 a_96_21.n5 a_96_21.n0 21.7605
R100 a_96_21.n9 a_96_21.n1 13.146
R101 a_96_21.n14 a_96_21.n10 11.2005
R102 a_96_21.n6 a_96_21.n2 10.2247
R103 a_96_21.n8 a_96_21.n7 1.46111
R104 a_484_47.n1 a_484_47.t0 312.334
R105 a_484_47.n1 a_484_47.n0 185
R106 a_484_47.n3 a_484_47.t6 174.512
R107 a_484_47.n3 a_484_47.n2 98.982
R108 a_484_47.n5 a_484_47.n4 89.3175
R109 a_484_47.n4 a_484_47.n1 51.265
R110 a_484_47.n4 a_484_47.n3 48.4528
R111 a_484_47.t1 a_484_47.n5 33.2313
R112 a_484_47.n5 a_484_47.t2 31.3851
R113 a_484_47.n0 a_484_47.t5 24.9236
R114 a_484_47.n0 a_484_47.t7 24.9236
R115 a_484_47.n2 a_484_47.t3 24.9236
R116 a_484_47.n2 a_484_47.t4 24.9236
R117 VNB.t6 VNB.t0 2677.02
R118 VNB.t1 VNB.t2 1423.95
R119 VNB.t3 VNB.t10 1196.12
R120 VNB.t4 VNB.t3 1196.12
R121 VNB.t2 VNB.t4 1196.12
R122 VNB.t9 VNB.t1 1196.12
R123 VNB.t11 VNB.t9 1196.12
R124 VNB.t0 VNB.t11 1196.12
R125 VNB.t8 VNB.t6 1196.12
R126 VNB.t5 VNB.t8 1196.12
R127 VNB.t7 VNB.t5 1196.12
R128 VNB VNB.t7 1167.64
R129 VGND.n19 VGND.t4 286.426
R130 VGND.n25 VGND.t5 280.822
R131 VGND.n9 VGND.n8 219.65
R132 VGND.n7 VGND.n6 207.965
R133 VGND.n2 VGND.n1 207.965
R134 VGND.n12 VGND.n11 34.6358
R135 VGND.n13 VGND.n12 34.6358
R136 VGND.n13 VGND.n4 34.6358
R137 VGND.n17 VGND.n4 34.6358
R138 VGND.n18 VGND.n17 34.6358
R139 VGND.n24 VGND.n23 34.6358
R140 VGND.n20 VGND.n2 32.0005
R141 VGND.n20 VGND.n19 31.2476
R142 VGND.n11 VGND.n7 26.7299
R143 VGND.n25 VGND.n24 25.977
R144 VGND.n8 VGND.t7 24.9236
R145 VGND.n8 VGND.t1 24.9236
R146 VGND.n6 VGND.t2 24.9236
R147 VGND.n6 VGND.t0 24.9236
R148 VGND.n1 VGND.t6 24.9236
R149 VGND.n1 VGND.t3 24.9236
R150 VGND.n26 VGND.n25 17.9593
R151 VGND.n9 VGND.n7 14.809
R152 VGND.n11 VGND.n10 9.3005
R153 VGND.n12 VGND.n5 9.3005
R154 VGND.n14 VGND.n13 9.3005
R155 VGND.n15 VGND.n4 9.3005
R156 VGND.n17 VGND.n16 9.3005
R157 VGND.n18 VGND.n3 9.3005
R158 VGND.n21 VGND.n20 9.3005
R159 VGND.n23 VGND.n22 9.3005
R160 VGND.n24 VGND.n0 9.3005
R161 VGND.n19 VGND.n18 3.38874
R162 VGND.n23 VGND.n2 2.63579
R163 VGND.n10 VGND.n9 0.845273
R164 VGND.n10 VGND.n5 0.120292
R165 VGND.n14 VGND.n5 0.120292
R166 VGND.n15 VGND.n14 0.120292
R167 VGND.n16 VGND.n15 0.120292
R168 VGND.n16 VGND.n3 0.120292
R169 VGND.n21 VGND.n3 0.120292
R170 VGND.n22 VGND.n21 0.120292
R171 VGND.n22 VGND.n0 0.120292
R172 VGND.n26 VGND.n0 0.120292
R173 VGND VGND.n26 0.0226354
R174 X.n2 X.n0 253.444
R175 X.n2 X.n1 209.02
R176 X.n5 X.n3 135.249
R177 X.n5 X.n4 98.982
R178 X X.n2 39.4176
R179 X X.n5 29.3806
R180 X.n0 X.t7 26.5955
R181 X.n0 X.t6 26.5955
R182 X.n1 X.t5 26.5955
R183 X.n1 X.t4 26.5955
R184 X.n3 X.t1 24.9236
R185 X.n3 X.t3 24.9236
R186 X.n4 X.t0 24.9236
R187 X.n4 X.t2 24.9236
R188 B2.n0 B2.t0 212.081
R189 B2.n1 B2.t1 212.081
R190 B2 B2.n2 153.268
R191 B2.n0 B2.t3 139.78
R192 B2.n1 B2.t2 139.78
R193 B2.n2 B2.n0 30.6732
R194 B2.n2 B2.n1 30.6732
R195 A1.n2 A1.n0 260.188
R196 A1.n1 A1.t0 241.536
R197 A1.n0 A1.t2 241.536
R198 A1.n1 A1.t1 169.237
R199 A1.n0 A1.t3 169.237
R200 A1.n2 A1.n1 152
R201 A1 A1.n2 23.6805
R202 a_918_297.n1 a_918_297.n0 935.015
R203 a_918_297.n0 a_918_297.t3 26.5955
R204 a_918_297.n0 a_918_297.t0 26.5955
R205 a_918_297.t1 a_918_297.n1 26.5955
R206 a_918_297.n1 a_918_297.t2 26.5955
R207 A2.n0 A2.t1 212.081
R208 A2.n1 A2.t0 212.081
R209 A2 A2.n2 157.12
R210 A2.n0 A2.t3 139.78
R211 A2.n1 A2.t2 139.78
R212 A2.n2 A2.n0 30.6732
R213 A2.n2 A2.n1 30.6732
C0 VPB B1 0.066215f
C1 B2 VGND 0.016122f
C2 B1 A1 0.092645f
C3 VPB VGND 0.009561f
C4 VPB B2 0.050999f
C5 A1 VGND 0.033334f
C6 B1 X 5.7e-19
C7 VPB A1 0.071126f
C8 A2 VGND 0.02453f
C9 B1 VPWR 0.044326f
C10 X VGND 0.26292f
C11 B2 X 3.6e-19
C12 VPB A2 0.050973f
C13 VPWR VGND 0.128603f
C14 A1 A2 0.209888f
C15 B2 VPWR 0.016799f
C16 VPB X 0.014393f
C17 VPB VPWR 0.141425f
C18 A1 VPWR 0.077937f
C19 A2 VPWR 0.016891f
C20 VPWR X 0.336901f
C21 B1 VGND 0.022322f
C22 B1 B2 0.212706f
C23 VGND VNB 0.73852f
C24 X VNB 0.060903f
C25 VPWR VNB 0.645667f
C26 A2 VNB 0.166288f
C27 A1 VNB 0.227657f
C28 B2 VNB 0.166404f
C29 B1 VNB 0.194216f
C30 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22ai_1 VPB VNB VGND VPWR A1 A2 B1 B2 Y
X0 VGND.t1 A2.t0 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1 a_27_47.t2 B2.t0 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.092625 ps=0.935 w=0.65 l=0.15
X2 VPWR.t1 A1.t0 a_307_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297.t1 A2.t1 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2325 ps=1.465 w=1 l=0.15
X4 a_27_47.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t0 B2.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2325 pd=1.465 as=0.1125 ps=1.225 w=1 l=0.15
X6 a_109_297.t1 B1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.26 ps=2.52 w=1 l=0.15
X7 Y.t2 B1.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t1 241.536
R1 A2 A2.n0 190.323
R2 A2.n0 A2.t0 169.237
R3 a_27_47.n1 a_27_47.t1 323.514
R4 a_27_47.t0 a_27_47.n1 200.645
R5 a_27_47.n1 a_27_47.n0 92.501
R6 a_27_47.n0 a_27_47.t2 36.9236
R7 a_27_47.n0 a_27_47.t3 28.6159
R8 VGND VGND.n0 213.067
R9 VGND.n0 VGND.t0 24.9236
R10 VGND.n0 VGND.t1 24.9236
R11 VNB.t2 VNB.t3 1438.19
R12 VNB.t1 VNB.t2 1238.83
R13 VNB.t3 VNB.t0 1196.12
R14 VNB VNB.t1 925.567
R15 B2.n0 B2.t1 239.986
R16 B2 B2.n0 178.625
R17 B2.n0 B2.t0 167.685
R18 Y Y.n0 589.481
R19 Y.n2 Y.n0 585
R20 Y.n2 Y.n1 284.214
R21 Y.n0 Y.t3 65.0105
R22 Y.n1 Y.t1 27.6928
R23 Y.n0 Y.t0 26.5955
R24 Y.n1 Y.t2 24.9236
R25 Y Y.n2 4.2245
R26 A1.n0 A1.t0 236.18
R27 A1.n0 A1.t1 163.881
R28 A1 A1.n0 156.161
R29 a_307_297.t0 a_307_297.t1 41.3705
R30 VPWR.n0 VPWR.t0 884.386
R31 VPWR.n0 VPWR.t1 252.41
R32 VPWR VPWR.n0 0.070077
R33 VPB.t0 VPB.t3 364.019
R34 VPB.t1 VPB.t0 221.964
R35 VPB.t3 VPB.t2 213.084
R36 VPB VPB.t1 192.369
R37 a_109_297.t0 a_109_297.t1 44.3255
R38 B1.n0 B1.t0 230.155
R39 B1 B1.n0 173.067
R40 B1.n0 B1.t1 157.856
C0 Y B1 0.132195f
C1 VPWR B2 0.011443f
C2 VGND VPB 0.004703f
C3 VGND B1 0.01416f
C4 Y B2 0.120033f
C5 VPWR A2 0.119219f
C6 Y A2 0.063042f
C7 VPWR A1 0.056942f
C8 VGND B2 0.010519f
C9 VPB B1 0.042669f
C10 VGND A2 0.015811f
C11 Y A1 5.15e-19
C12 VPB B2 0.030207f
C13 VGND A1 0.014673f
C14 VPB A2 0.030858f
C15 B1 B2 0.057563f
C16 VPB A1 0.031536f
C17 B2 A2 0.090951f
C18 VPWR Y 0.101555f
C19 B2 A1 4.27e-19
C20 VPWR VGND 0.045923f
C21 A2 A1 0.089045f
C22 Y VGND 0.00968f
C23 VPWR VPB 0.061209f
C24 Y VPB 0.00499f
C25 VPWR B1 0.045146f
C26 VGND VNB 0.297636f
C27 Y VNB 0.014366f
C28 VPWR VNB 0.298221f
C29 A1 VNB 0.131261f
C30 A2 VNB 0.097299f
C31 B2 VNB 0.093928f
C32 B1 VNB 0.184404f
C33 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22ai_2 VPB VNB VGND VPWR A1 A2 Y B2 B1
X0 Y.t2 B2.t0 a_27_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t4 B2.t1 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t3 B1.t0 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297.t3 A1.t0 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47.t0 A2.t0 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t2 A1.t1 a_475_297.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47.t7 A1.t2 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47.t4 B1.t1 Y.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t6 B1.t2 a_27_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47.t2 B2.t2 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.26975 pd=1.48 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t2 A1.t3 a_27_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t0 B1.t3 a_27_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297.t1 A2.t1 Y.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y.t0 A2.t2 a_475_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297.t0 B2.t3 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t0 A2.t3 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26975 ps=1.48 w=0.65 l=0.15
R0 B2.n0 B2.t3 212.081
R1 B2.n1 B2.t0 212.081
R2 B2.n0 B2.t2 139.78
R3 B2.n1 B2.t1 139.78
R4 B2 B2.n2 71.2476
R5 B2.n2 B2.n1 33.5655
R6 B2.n2 B2.n0 21.5936
R7 a_27_297.t0 a_27_297.n1 392.906
R8 a_27_297.n1 a_27_297.t2 300.269
R9 a_27_297.n1 a_27_297.n0 187.506
R10 a_27_297.n0 a_27_297.t1 26.5955
R11 a_27_297.n0 a_27_297.t3 26.5955
R12 Y.n2 Y.n0 334.918
R13 Y Y.n1 324.252
R14 Y.n5 Y.n3 237.513
R15 Y.n5 Y.n4 185
R16 Y Y.n5 68.7712
R17 Y.n1 Y.t1 26.5955
R18 Y.n1 Y.t2 26.5955
R19 Y.n0 Y.t7 26.5955
R20 Y.n0 Y.t0 26.5955
R21 Y.n4 Y.t3 24.9236
R22 Y.n4 Y.t4 24.9236
R23 Y.n3 Y.t5 24.9236
R24 Y.n3 Y.t6 24.9236
R25 Y.n2 Y 7.46717
R26 Y Y.n2 4.70254
R27 VPB.t2 VPB.t0 580.062
R28 VPB.t1 VPB.t7 248.599
R29 VPB.t5 VPB.t1 248.599
R30 VPB.t0 VPB.t5 248.599
R31 VPB.t3 VPB.t2 248.599
R32 VPB.t6 VPB.t3 248.599
R33 VPB.t4 VPB.t6 248.599
R34 VPB VPB.t4 201.246
R35 a_27_47.n6 a_27_47.t5 189.614
R36 a_27_47.n5 a_27_47.n4 185
R37 a_27_47.n3 a_27_47.n2 185
R38 a_27_47.n7 a_27_47.n6 185
R39 a_27_47.n1 a_27_47.t7 174.512
R40 a_27_47.n4 a_27_47.n3 102.463
R41 a_27_47.n1 a_27_47.n0 98.982
R42 a_27_47.n2 a_27_47.n1 67.5142
R43 a_27_47.n6 a_27_47.n5 63.2476
R44 a_27_47.n5 a_27_47.n2 41.7887
R45 a_27_47.n3 a_27_47.t1 25.8467
R46 a_27_47.n4 a_27_47.t2 24.9236
R47 a_27_47.n0 a_27_47.t6 24.9236
R48 a_27_47.n0 a_27_47.t0 24.9236
R49 a_27_47.t3 a_27_47.n7 24.9236
R50 a_27_47.n7 a_27_47.t4 24.9236
R51 VNB.t2 VNB.t1 2790.94
R52 VNB.t6 VNB.t7 1196.12
R53 VNB.t0 VNB.t6 1196.12
R54 VNB.t1 VNB.t0 1196.12
R55 VNB.t3 VNB.t2 1196.12
R56 VNB.t4 VNB.t3 1196.12
R57 VNB.t5 VNB.t4 1196.12
R58 VNB VNB.t5 968.285
R59 B1.n0 B1.t0 212.081
R60 B1.n1 B1.t3 212.081
R61 B1.n0 B1.t1 139.78
R62 B1.n1 B1.t2 139.78
R63 B1 B1.n2 71.0407
R64 B1.n2 B1.n0 34.3636
R65 B1.n2 B1.n1 20.7784
R66 VPWR.n2 VPWR.n0 325.031
R67 VPWR.n2 VPWR.n1 324.24
R68 VPWR.n1 VPWR.t1 26.5955
R69 VPWR.n1 VPWR.t0 26.5955
R70 VPWR.n0 VPWR.t3 26.5955
R71 VPWR.n0 VPWR.t2 26.5955
R72 VPWR VPWR.n2 0.148694
R73 A1.n0 A1.t0 212.081
R74 A1.n1 A1.t1 212.081
R75 A1.n0 A1.t2 139.78
R76 A1.n1 A1.t3 139.78
R77 A1 A1.n2 71.0478
R78 A1.n2 A1.n1 34.2066
R79 A1.n2 A1.n0 20.9353
R80 a_475_297.n0 a_475_297.t0 392.906
R81 a_475_297.n0 a_475_297.t3 300.267
R82 a_475_297.n1 a_475_297.n0 187.506
R83 a_475_297.t2 a_475_297.n1 26.5955
R84 a_475_297.n1 a_475_297.t1 26.5955
R85 A2.n0 A2.t1 212.081
R86 A2.n1 A2.t2 212.081
R87 A2.n0 A2.t0 139.78
R88 A2.n1 A2.t3 139.78
R89 A2 A2.n2 71.2744
R90 A2.n2 A2.n0 33.7298
R91 A2.n2 A2.n1 21.4293
R92 VGND.n2 VGND.n1 219.055
R93 VGND.n2 VGND.n0 216.274
R94 VGND.n1 VGND.t3 24.9236
R95 VGND.n1 VGND.t2 24.9236
R96 VGND.n0 VGND.t1 24.9236
R97 VGND.n0 VGND.t0 24.9236
R98 VGND VGND.n2 1.1645
C0 VPWR VGND 0.088529f
C1 VPB VPWR 0.100418f
C2 Y VGND 0.022889f
C3 VPB Y 0.019705f
C4 B1 VPWR 0.043776f
C5 VPB VGND 0.011072f
C6 B1 Y 0.052485f
C7 B1 VGND 0.019505f
C8 VPB B1 0.060643f
C9 B2 A2 0.018598f
C10 B2 VPWR 0.018617f
C11 A2 A1 0.068184f
C12 A2 VPWR 0.018799f
C13 B2 Y 0.174078f
C14 B2 VGND 0.019466f
C15 VPB B2 0.062102f
C16 A2 Y 0.089289f
C17 A1 VPWR 0.039696f
C18 A2 VGND 0.030408f
C19 B1 B2 0.068122f
C20 VPB A2 0.061811f
C21 A1 Y 0.001363f
C22 A1 VGND 0.027354f
C23 VPB A1 0.061545f
C24 VPWR Y 0.0265f
C25 VGND VNB 0.530218f
C26 Y VNB 0.028982f
C27 VPWR VNB 0.445348f
C28 A1 VNB 0.214995f
C29 A2 VNB 0.188367f
C30 B2 VNB 0.189319f
C31 B1 VNB 0.217195f
C32 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22ai_4 VNB VPB VGND VPWR A1 A2 B2 Y B1
X0 a_33_47.t15 B2.t0 Y.t9 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t3 A1.t0 a_33_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t4 A2.t0 a_33_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_33_47.t10 B1.t0 Y.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_797_297.t3 B2.t1 Y.t13 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t3 A2.t1 a_115_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_797_297.t7 B1.t1 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t12 B2.t2 a_797_297.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_115_297.t2 A2.t2 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR.t6 B1.t2 a_797_297.t6 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_33_47.t5 A1.t1 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t1 A1.t2 a_33_47.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_33_47.t7 A2.t3 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_33_47.t8 A2.t4 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t5 A2.t5 a_115_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_33_47.t3 A1.t3 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_797_297.t5 B1.t3 VPWR.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.32 w=1 l=0.15
X17 a_115_297.t7 A1.t4 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR.t2 A1.t5 a_115_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t4 B1.t4 a_797_297.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t7 A2.t6 a_33_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_33_47.t0 B1.t5 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_797_297.t1 B2.t3 Y.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t1 A1.t6 a_115_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.135 ps=1.27 w=1 l=0.15
X24 Y.t8 B2.t4 a_33_47.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 Y.t10 B2.t5 a_797_297.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y.t1 B1.t6 a_33_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.104 ps=0.97 w=0.65 l=0.15
X27 Y.t15 B2.t6 a_33_47.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_115_297.t0 A2.t7 Y.t6 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y.t2 B1.t7 a_33_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_33_47.t12 B2.t7 Y.t14 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_115_297.t4 A1.t7 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
R0 B2.n0 B2.t3 212.081
R1 B2.n3 B2.t5 212.081
R2 B2.n6 B2.t1 212.081
R3 B2.n4 B2.t2 212.081
R4 B2.n5 B2.n2 173.761
R5 B2 B2.n1 162.881
R6 B2.n9 B2.n8 152
R7 B2.n7 B2.n2 152
R8 B2.n0 B2.t6 139.78
R9 B2.n3 B2.t0 139.78
R10 B2.n6 B2.t4 139.78
R11 B2.n4 B2.t7 139.78
R12 B2.n8 B2.n7 49.6611
R13 B2.n6 B2.n5 46.0096
R14 B2.n3 B2.n1 41.6278
R15 B2.n9 B2.n2 21.7605
R16 B2.n1 B2.n0 19.7187
R17 B2.n5 B2.n4 15.3369
R18 B2 B2.n9 10.8805
R19 B2.n8 B2.n3 8.03383
R20 B2.n7 B2.n6 3.65202
R21 Y.n13 Y.n11 638.836
R22 Y.n2 Y.n0 638.836
R23 Y.n2 Y.n1 585
R24 Y.n13 Y.n12 585
R25 Y.n4 Y.n3 185
R26 Y.n6 Y.n5 185
R27 Y.n8 Y.n7 185
R28 Y.n10 Y.n9 185
R29 Y.n4 Y.n2 181.218
R30 Y.n14 Y.n10 148.911
R31 Y.n6 Y.n4 61.4405
R32 Y.n8 Y.n6 61.4405
R33 Y.n10 Y.n8 61.4405
R34 Y.n12 Y.t6 26.5955
R35 Y.n12 Y.t3 26.5955
R36 Y.n11 Y.t4 26.5955
R37 Y.n11 Y.t5 26.5955
R38 Y.n1 Y.t11 26.5955
R39 Y.n1 Y.t10 26.5955
R40 Y.n0 Y.t13 26.5955
R41 Y.n0 Y.t12 26.5955
R42 Y.n9 Y.t0 24.9236
R43 Y.n9 Y.t1 24.9236
R44 Y.n7 Y.t14 24.9236
R45 Y.n7 Y.t2 24.9236
R46 Y.n5 Y.t9 24.9236
R47 Y.n5 Y.t8 24.9236
R48 Y.n3 Y.t7 24.9236
R49 Y.n3 Y.t15 24.9236
R50 Y Y.n13 3.57697
R51 Y Y.n14 2.25932
R52 Y.n14 Y 1.12991
R53 a_33_47.n1 a_33_47.t10 312.334
R54 a_33_47.n1 a_33_47.n0 185
R55 a_33_47.n11 a_33_47.n10 185
R56 a_33_47.n13 a_33_47.n12 185
R57 a_33_47.n3 a_33_47.t11 174.512
R58 a_33_47.n3 a_33_47.n2 98.982
R59 a_33_47.n5 a_33_47.n4 98.982
R60 a_33_47.n7 a_33_47.n6 98.982
R61 a_33_47.n9 a_33_47.n8 89.0112
R62 a_33_47.n11 a_33_47.n9 51.9746
R63 a_33_47.n9 a_33_47.n7 49.4146
R64 a_33_47.n12 a_33_47.n1 48.8732
R65 a_33_47.n12 a_33_47.n11 48.8732
R66 a_33_47.n5 a_33_47.n3 38.7884
R67 a_33_47.n7 a_33_47.n5 36.2672
R68 a_33_47.n8 a_33_47.t1 34.1543
R69 a_33_47.n10 a_33_47.t2 24.9236
R70 a_33_47.n10 a_33_47.t0 24.9236
R71 a_33_47.n0 a_33_47.t13 24.9236
R72 a_33_47.n0 a_33_47.t15 24.9236
R73 a_33_47.n8 a_33_47.t3 24.9236
R74 a_33_47.n6 a_33_47.t9 24.9236
R75 a_33_47.n6 a_33_47.t8 24.9236
R76 a_33_47.n4 a_33_47.t6 24.9236
R77 a_33_47.n4 a_33_47.t7 24.9236
R78 a_33_47.n2 a_33_47.t4 24.9236
R79 a_33_47.n2 a_33_47.t5 24.9236
R80 a_33_47.t14 a_33_47.n13 24.9236
R81 a_33_47.n13 a_33_47.t12 24.9236
R82 VNB.t3 VNB.t1 1338.51
R83 VNB.t13 VNB.t10 1196.12
R84 VNB.t15 VNB.t13 1196.12
R85 VNB.t14 VNB.t15 1196.12
R86 VNB.t12 VNB.t14 1196.12
R87 VNB.t2 VNB.t12 1196.12
R88 VNB.t0 VNB.t2 1196.12
R89 VNB.t1 VNB.t0 1196.12
R90 VNB.t9 VNB.t3 1196.12
R91 VNB.t8 VNB.t9 1196.12
R92 VNB.t6 VNB.t8 1196.12
R93 VNB.t7 VNB.t6 1196.12
R94 VNB.t4 VNB.t7 1196.12
R95 VNB.t5 VNB.t4 1196.12
R96 VNB.t11 VNB.t5 1196.12
R97 VNB VNB.t11 1011
R98 A1.n1 A1.n0 324.981
R99 A1.n0 A1.t6 241.536
R100 A1.n2 A1.t4 212.081
R101 A1.n5 A1.t5 212.081
R102 A1.n3 A1.t7 212.081
R103 A1.n0 A1.t3 169.237
R104 A1.n7 A1.n6 152
R105 A1.n2 A1.t0 139.78
R106 A1.n5 A1.t1 139.78
R107 A1.n3 A1.t2 139.78
R108 A1.n4 A1 80.2728
R109 A1.n6 A1.n5 48.2005
R110 A1.n4 A1.n3 33.2102
R111 A1.n5 A1.n4 21.5682
R112 A1.n6 A1.n2 13.146
R113 A1 A1.n1 5.4405
R114 A1 A1.n7 2.6571
R115 A1.n7 A1.n1 0.725028
R116 VGND.n7 VGND.n6 219.762
R117 VGND.n5 VGND.n4 207.965
R118 VGND.n11 VGND.n3 207.965
R119 VGND.n1 VGND.n0 207.965
R120 VGND.n10 VGND.n9 34.6358
R121 VGND.n12 VGND.n1 33.1299
R122 VGND.n12 VGND.n11 30.1181
R123 VGND.n6 VGND.t0 24.9236
R124 VGND.n6 VGND.t7 24.9236
R125 VGND.n4 VGND.t6 24.9236
R126 VGND.n4 VGND.t4 24.9236
R127 VGND.n3 VGND.t5 24.9236
R128 VGND.n3 VGND.t3 24.9236
R129 VGND.n0 VGND.t2 24.9236
R130 VGND.n0 VGND.t1 24.9236
R131 VGND.n9 VGND.n5 24.0946
R132 VGND.n7 VGND.n5 17.3598
R133 VGND.n9 VGND.n8 9.3005
R134 VGND.n10 VGND.n2 9.3005
R135 VGND.n13 VGND.n12 9.3005
R136 VGND.n14 VGND.n1 9.16498
R137 VGND.n11 VGND.n10 4.51815
R138 VGND.n8 VGND.n7 0.929644
R139 VGND.n14 VGND.n13 0.141672
R140 VGND VGND.n14 0.121778
R141 VGND.n8 VGND.n2 0.120292
R142 VGND.n13 VGND.n2 0.120292
R143 A2.n3 A2.t7 212.081
R144 A2.n5 A2.t1 212.081
R145 A2.n7 A2.t2 212.081
R146 A2.n1 A2.t5 212.081
R147 A2.n4 A2.n0 173.761
R148 A2.n9 A2.n2 173.761
R149 A2.n6 A2.n0 152
R150 A2.n9 A2.n8 152
R151 A2.n3 A2.t6 139.78
R152 A2.n5 A2.t4 139.78
R153 A2.n7 A2.t0 139.78
R154 A2.n1 A2.t3 139.78
R155 A2.n8 A2.n6 49.6611
R156 A2.n5 A2.n4 48.2005
R157 A2.n7 A2.n2 39.4369
R158 A2.n2 A2.n1 21.9096
R159 A2.n4 A2.n3 13.146
R160 A2 A2.n9 12.4805
R161 A2.n8 A2.n7 10.2247
R162 A2 A2.n0 9.2805
R163 A2.n6 A2.n5 1.46111
R164 B1 B1.n0 311.2
R165 B1.n0 B1.t4 238.59
R166 B1.n3 B1.t1 212.081
R167 B1.n2 B1.t2 212.081
R168 B1.n1 B1.t3 212.081
R169 B1.n0 B1.t0 166.291
R170 B1.n3 B1.t7 139.78
R171 B1.n2 B1.t5 139.78
R172 B1.n1 B1.t6 139.78
R173 B1 B1.n4 67.5321
R174 B1.n2 B1.n1 61.346
R175 B1.n4 B1.n2 29.1988
R176 B1.n4 B1.n3 25.3111
R177 a_797_297.n3 a_797_297.n1 668.523
R178 a_797_297.n4 a_797_297.n0 638.979
R179 a_797_297.n5 a_797_297.n4 585
R180 a_797_297.n3 a_797_297.n2 288.212
R181 a_797_297.n4 a_797_297.n3 61.8028
R182 a_797_297.n2 a_797_297.t2 26.5955
R183 a_797_297.n2 a_797_297.t7 26.5955
R184 a_797_297.n1 a_797_297.t6 26.5955
R185 a_797_297.n1 a_797_297.t5 26.5955
R186 a_797_297.n0 a_797_297.t4 26.5955
R187 a_797_297.n0 a_797_297.t1 26.5955
R188 a_797_297.n5 a_797_297.t0 26.5955
R189 a_797_297.t3 a_797_297.n5 26.5955
R190 VPB.t5 VPB.t13 278.193
R191 VPB.t9 VPB.t12 248.599
R192 VPB.t8 VPB.t9 248.599
R193 VPB.t11 VPB.t8 248.599
R194 VPB.t10 VPB.t11 248.599
R195 VPB.t15 VPB.t10 248.599
R196 VPB.t14 VPB.t15 248.599
R197 VPB.t13 VPB.t14 248.599
R198 VPB.t0 VPB.t5 248.599
R199 VPB.t3 VPB.t0 248.599
R200 VPB.t2 VPB.t3 248.599
R201 VPB.t1 VPB.t2 248.599
R202 VPB.t7 VPB.t1 248.599
R203 VPB.t6 VPB.t7 248.599
R204 VPB.t4 VPB.t6 248.599
R205 VPB VPB.t4 210.125
R206 a_115_297.n4 a_115_297.n0 638.836
R207 a_115_297.n5 a_115_297.n4 585
R208 a_115_297.n3 a_115_297.n2 288.212
R209 a_115_297.n3 a_115_297.n1 257.983
R210 a_115_297.n4 a_115_297.n3 61.8028
R211 a_115_297.n2 a_115_297.t1 26.5955
R212 a_115_297.n2 a_115_297.t7 26.5955
R213 a_115_297.n1 a_115_297.t6 26.5955
R214 a_115_297.n1 a_115_297.t4 26.5955
R215 a_115_297.n0 a_115_297.t5 26.5955
R216 a_115_297.n0 a_115_297.t0 26.5955
R217 a_115_297.t3 a_115_297.n5 26.5955
R218 a_115_297.n5 a_115_297.t2 26.5955
R219 VPWR.n9 VPWR.t4 850.336
R220 VPWR.n6 VPWR.n5 609.437
R221 VPWR.n10 VPWR.n8 607.4
R222 VPWR.n22 VPWR.n2 606.505
R223 VPWR.n24 VPWR.t0 252.511
R224 VPWR.n16 VPWR.n15 34.6358
R225 VPWR.n17 VPWR.n16 34.6358
R226 VPWR.n17 VPWR.n3 34.6358
R227 VPWR.n21 VPWR.n3 34.6358
R228 VPWR.n12 VPWR.n11 34.6358
R229 VPWR.n5 VPWR.t1 34.4755
R230 VPWR.n5 VPWR.t5 28.5655
R231 VPWR.n22 VPWR.n21 26.7299
R232 VPWR.n2 VPWR.t3 26.5955
R233 VPWR.n2 VPWR.t2 26.5955
R234 VPWR.n8 VPWR.t7 26.5955
R235 VPWR.n8 VPWR.t6 26.5955
R236 VPWR.n23 VPWR.n22 23.7181
R237 VPWR.n24 VPWR.n23 20.7064
R238 VPWR.n10 VPWR.n9 20.0223
R239 VPWR.n12 VPWR.n6 9.41227
R240 VPWR.n11 VPWR.n7 9.3005
R241 VPWR.n13 VPWR.n12 9.3005
R242 VPWR.n15 VPWR.n14 9.3005
R243 VPWR.n16 VPWR.n4 9.3005
R244 VPWR.n18 VPWR.n17 9.3005
R245 VPWR.n19 VPWR.n3 9.3005
R246 VPWR.n21 VPWR.n20 9.3005
R247 VPWR.n22 VPWR.n1 9.3005
R248 VPWR.n23 VPWR.n0 9.3005
R249 VPWR.n25 VPWR.n24 9.3005
R250 VPWR.n15 VPWR.n6 8.65932
R251 VPWR.n11 VPWR.n10 4.14168
R252 VPWR.n9 VPWR.n7 0.149563
R253 VPWR.n13 VPWR.n7 0.120292
R254 VPWR.n14 VPWR.n13 0.120292
R255 VPWR.n14 VPWR.n4 0.120292
R256 VPWR.n18 VPWR.n4 0.120292
R257 VPWR.n19 VPWR.n18 0.120292
R258 VPWR.n20 VPWR.n19 0.120292
R259 VPWR.n20 VPWR.n1 0.120292
R260 VPWR.n1 VPWR.n0 0.120292
R261 VPWR.n25 VPWR.n0 0.120292
R262 VPWR VPWR.n25 0.0226354
C0 VGND A1 0.060596f
C1 VGND VPWR 0.141786f
C2 VPB Y 0.013714f
C3 A1 A2 0.291492f
C4 B1 B2 0.300687f
C5 A2 VPWR 0.032168f
C6 VPB VGND 0.008742f
C7 A1 B1 0.049228f
C8 B1 VPWR 0.068294f
C9 VPB A2 0.114794f
C10 B2 VPWR 0.034174f
C11 VPB B1 0.128129f
C12 A1 VPWR 0.110538f
C13 VPB B2 0.114723f
C14 Y VGND 0.041926f
C15 VPB A1 0.130485f
C16 VPB VPWR 0.14836f
C17 Y A2 0.034931f
C18 VGND A2 0.052363f
C19 Y B1 0.413514f
C20 VGND B1 0.036078f
C21 Y B2 0.156323f
C22 Y A1 0.194596f
C23 VGND B2 0.033543f
C24 Y VPWR 0.12838f
C25 VGND VNB 0.798187f
C26 Y VNB 0.07909f
C27 VPWR VNB 0.713952f
C28 B2 VNB 0.35175f
C29 B1 VNB 0.387614f
C30 A2 VNB 0.351925f
C31 A1 VNB 0.401914f
C32 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31a_1 X A1 A2 A3 B1 VPB VNB VGND VPWR
X0 a_103_199.t1 B1.t0 a_253_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR.t1 a_103_199.t3 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297.t0 A2.t0 a_253_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199.t0 A3.t0 a_337_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297.t1 A1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR.t0 B1.t1 a_103_199.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND.t2 a_103_199.t4 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47.t1 A1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47.t3 A3.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND.t0 A2.t1 a_253_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B1.n0 B1.t1 238.155
R1 B1.n0 B1.t0 165.856
R2 B1 B1.n0 156.849
R3 a_253_47.n1 a_253_47.n0 450.795
R4 a_253_47.t0 a_253_47.n1 30.462
R5 a_253_47.n1 a_253_47.t3 30.462
R6 a_253_47.n0 a_253_47.t2 24.9236
R7 a_253_47.n0 a_253_47.t1 24.9236
R8 a_103_199.n1 a_103_199.n0 373.822
R9 a_103_199.n2 a_103_199.n1 284.533
R10 a_103_199.n0 a_103_199.t3 241.536
R11 a_103_199.n1 a_103_199.t1 231.631
R12 a_103_199.n0 a_103_199.t4 169.237
R13 a_103_199.t0 a_103_199.n2 56.1455
R14 a_103_199.n2 a_103_199.t2 27.5805
R15 VNB.t2 VNB.t1 1537.86
R16 VNB VNB.t2 1438.19
R17 VNB.t4 VNB.t0 1366.99
R18 VNB.t3 VNB.t4 1366.99
R19 VNB.t1 VNB.t3 1196.12
R20 X.n0 X 590.091
R21 X.n1 X.n0 585
R22 X.n3 X 186.892
R23 X.n4 X.n3 185
R24 X.n0 X.t1 42.3555
R25 X.n3 X.t0 39.6928
R26 X X.n5 11.5618
R27 X.n4 X 8.0005
R28 X.n1 X 4.8005
R29 X.n2 X.n1 3.63686
R30 X.n5 X 2.47792
R31 X X.n2 2.06502
R32 X X.n4 1.89141
R33 X.n5 X 1.74595
R34 X.n2 X 1.45505
R35 VPWR.n1 VPWR.t0 362.846
R36 VPWR.n1 VPWR.n0 318.649
R37 VPWR.n0 VPWR.t2 38.4155
R38 VPWR.n0 VPWR.t1 38.4155
R39 VPWR VPWR.n1 0.180156
R40 VPB.t0 VPB.t1 340.344
R41 VPB.t3 VPB.t4 319.627
R42 VPB VPB.t3 298.911
R43 VPB.t2 VPB.t0 284.113
R44 VPB.t4 VPB.t2 248.599
R45 A2.n0 A2.t0 241.536
R46 A2.n0 A2.t1 169.237
R47 A2.n1 A2.n0 152
R48 A2 A2.n1 16.3009
R49 A2.n1 A2 2.87397
R50 a_253_297.t0 a_253_297.t1 53.1905
R51 a_337_297.t0 a_337_297.t1 65.0105
R52 A3.n0 A3.t0 241.536
R53 A3.n0 A3.t1 169.237
R54 A3 A3.n0 153.19
R55 A1.n0 A1.t0 241.536
R56 A1.n0 A1.t1 169.237
R57 A1 A1.n0 154.971
R58 VGND.n2 VGND.n1 191.714
R59 VGND.n2 VGND.n0 108.688
R60 VGND.n0 VGND.t1 36.0005
R61 VGND.n0 VGND.t2 36.0005
R62 VGND.n1 VGND.t3 30.462
R63 VGND.n1 VGND.t0 30.462
R64 VGND VGND.n2 0.567674
C0 VPWR VGND 0.06508f
C1 B1 VPB 0.034421f
C2 A2 A3 0.136697f
C3 X VPB 0.01546f
C4 X A1 7.36e-19
C5 VPWR VPB 0.072655f
C6 VPWR A1 0.011487f
C7 VGND VPB 0.006333f
C8 B1 A3 0.073596f
C9 X A2 2.55e-19
C10 VGND A1 0.04324f
C11 VPWR A2 0.00974f
C12 X A3 1.42e-19
C13 VPWR A3 0.011038f
C14 VGND A2 0.013332f
C15 B1 X 8.93e-20
C16 VGND A3 0.013887f
C17 B1 VPWR 0.018978f
C18 VPB A1 0.027104f
C19 B1 VGND 0.015441f
C20 X VPWR 0.120185f
C21 VPB A2 0.028397f
C22 X VGND 0.109334f
C23 VPB A3 0.031009f
C24 A1 A2 0.080246f
C25 VGND VNB 0.39103f
C26 VPWR VNB 0.349144f
C27 X VNB 0.097222f
C28 B1 VNB 0.121351f
C29 A3 VNB 0.089564f
C30 A2 VNB 0.08849f
C31 A1 VNB 0.090241f
C32 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_108_21.t1 B1.t0 a_346_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_346_47.t2 A3.t0 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X.t2 a_108_21.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.26325 ps=2.11 w=0.65 l=0.15
X3 a_108_21.t0 A3.t1 a_430_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297.t0 A2.t0 a_346_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t1 a_108_21.t4 X.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297.t0 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND.t2 A2.t1 a_346_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X.t0 a_108_21.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR.t3 B1.t1 a_108_21.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.2125 ps=1.425 w=1 l=0.15
X10 VGND.t0 a_108_21.t6 X.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11375 ps=1 w=0.65 l=0.15
X11 a_346_47.t1 A1.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
R0 B1.n0 B1.t1 238.155
R1 B1.n0 B1.t0 165.856
R2 B1 B1.n0 156.849
R3 a_346_47.n1 a_346_47.n0 450.795
R4 a_346_47.n0 a_346_47.t3 30.462
R5 a_346_47.n0 a_346_47.t2 30.462
R6 a_346_47.t0 a_346_47.n1 24.9236
R7 a_346_47.n1 a_346_47.t1 24.9236
R8 a_108_21.n2 a_108_21.n1 373.822
R9 a_108_21.n3 a_108_21.n2 284.533
R10 a_108_21.n2 a_108_21.t1 231.31
R11 a_108_21.n1 a_108_21.t4 212.081
R12 a_108_21.n0 a_108_21.t5 212.081
R13 a_108_21.n1 a_108_21.t6 139.78
R14 a_108_21.n0 a_108_21.t3 139.78
R15 a_108_21.n1 a_108_21.n0 73.0308
R16 a_108_21.t0 a_108_21.n3 56.1455
R17 a_108_21.n3 a_108_21.t2 27.5805
R18 VNB.t0 VNB.t3 1537.86
R19 VNB.t1 VNB.t0 1423.95
R20 VNB.t4 VNB.t5 1366.99
R21 VNB.t2 VNB.t4 1366.99
R22 VNB VNB.t1 1324.27
R23 VNB.t3 VNB.t2 1196.12
R24 A3.n0 A3.t1 241.536
R25 A3.n0 A3.t0 169.237
R26 A3 A3.n0 153.19
R27 VGND.n4 VGND.n3 191.365
R28 VGND.n8 VGND.t1 164.429
R29 VGND.n2 VGND.n1 105.097
R30 VGND.n1 VGND.t3 36.0005
R31 VGND.n1 VGND.t0 36.0005
R32 VGND.n7 VGND.n6 34.6358
R33 VGND.n3 VGND.t4 30.462
R34 VGND.n3 VGND.t2 30.462
R35 VGND.n8 VGND.n7 23.3417
R36 VGND.n9 VGND.n8 9.3005
R37 VGND.n6 VGND.n5 9.3005
R38 VGND.n7 VGND.n0 9.3005
R39 VGND.n4 VGND.n2 6.84797
R40 VGND.n5 VGND.n4 0.860247
R41 VGND.n6 VGND.n2 0.753441
R42 VGND.n5 VGND.n0 0.120292
R43 VGND.n9 VGND.n0 0.120292
R44 VGND VGND.n9 0.0213333
R45 X.n0 X 590.091
R46 X.n1 X.n0 585
R47 X.n3 X 186.892
R48 X.n4 X.n3 185
R49 X.n0 X.t3 42.3555
R50 X.n3 X.t1 39.6928
R51 X.n0 X.t0 26.5955
R52 X.n3 X.t2 24.9236
R53 X.n6 X 23.2732
R54 X X.n5 11.5618
R55 X X.n6 10.736
R56 X.n4 X 8.0005
R57 X.n1 X 4.8005
R58 X.n2 X.n1 3.63686
R59 X.n6 X 3.30373
R60 X.n5 X 2.47792
R61 X X.n2 2.06502
R62 X X.n4 1.89141
R63 X.n5 X 1.74595
R64 X.n2 X 1.45505
R65 a_430_297.t0 a_430_297.t1 65.0105
R66 VPB.t4 VPB.t5 340.344
R67 VPB.t1 VPB.t3 319.627
R68 VPB.t0 VPB.t1 295.95
R69 VPB.t2 VPB.t4 284.113
R70 VPB VPB.t0 275.235
R71 VPB.t3 VPB.t2 248.599
R72 A2.n0 A2.t0 241.536
R73 A2.n0 A2.t1 169.237
R74 A2.n1 A2.n0 152
R75 A2 A2.n1 16.3009
R76 A2.n1 A2 2.87397
R77 a_346_297.t0 a_346_297.t1 53.1905
R78 VPWR.n3 VPWR.t3 361.447
R79 VPWR.n2 VPWR.n1 312.981
R80 VPWR.n7 VPWR.t0 275.002
R81 VPWR.n1 VPWR.t2 38.4155
R82 VPWR.n1 VPWR.t1 38.4155
R83 VPWR.n6 VPWR.n5 34.6358
R84 VPWR.n7 VPWR.n6 23.3417
R85 VPWR.n3 VPWR.n2 17.3761
R86 VPWR.n5 VPWR.n4 9.3005
R87 VPWR.n6 VPWR.n0 9.3005
R88 VPWR.n8 VPWR.n7 9.3005
R89 VPWR.n5 VPWR.n2 1.12991
R90 VPWR.n4 VPWR.n3 0.160392
R91 VPWR.n4 VPWR.n0 0.120292
R92 VPWR.n8 VPWR.n0 0.120292
R93 VPWR VPWR.n8 0.0213333
R94 A1.n0 A1.t0 241.536
R95 A1.n0 A1.t1 169.237
R96 A1 A1.n0 154.971
C0 VPB A3 0.030998f
C1 A1 A2 0.080246f
C2 VPB B1 0.034363f
C3 A2 A3 0.136697f
C4 VPB VPWR 0.090218f
C5 A1 VPWR 0.011533f
C6 VPB X 0.006936f
C7 A3 B1 0.073596f
C8 VPB VGND 0.007017f
C9 A1 X 7.36e-19
C10 A2 VPWR 0.009742f
C11 A3 VPWR 0.011087f
C12 A2 X 2.55e-19
C13 A1 VGND 0.043406f
C14 B1 VPWR 0.019038f
C15 A3 X 1.42e-19
C16 A2 VGND 0.013332f
C17 A3 VGND 0.014017f
C18 B1 X 8.93e-20
C19 VPWR X 0.238902f
C20 B1 VGND 0.015575f
C21 VPWR VGND 0.077728f
C22 VPB A1 0.027104f
C23 X VGND 0.197649f
C24 VPB A2 0.028397f
C25 VGND VNB 0.465904f
C26 X VNB 0.030618f
C27 VPWR VNB 0.421343f
C28 B1 VNB 0.121321f
C29 A3 VNB 0.089564f
C30 A2 VNB 0.08849f
C31 A1 VNB 0.090241f
C32 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31a_4 VGND VPWR VPB VNB X A2 A1 A3 B1
X0 VPWR.t6 A1.t0 a_926_297.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t8 A1.t1 a_496_47.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_926_297.t2 A1.t2 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t0 A3.t0 a_496_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VGND.t2 a_102_21.t6 X.t7 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t9 A2.t0 a_496_47.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_926_297.t0 A2.t1 a_672_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_102_21.t5 B1.t0 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X8 a_496_47.t1 A2.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X.t6 a_102_21.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X10 a_102_21.t4 B1.t1 a_496_47.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11 VPWR.t1 a_102_21.t8 X.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X.t5 a_102_21.t9 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 X.t2 a_102_21.t10 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X14 VPWR.t3 a_102_21.t11 X.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X15 a_672_297.t3 A3.t1 a_102_21.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_496_47.t2 B1.t2 a_102_21.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_102_21.t2 A3.t2 a_672_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X18 VGND.t1 a_102_21.t12 X.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X.t0 a_102_21.t13 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 a_496_47.t3 A3.t3 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR.t4 B1.t3 a_102_21.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.145 ps=1.29 w=1 l=0.15
X22 a_496_47.t4 A1.t3 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_672_297.t0 A2.t3 a_926_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A1.n0 A1.t2 221.72
R1 A1.n1 A1.t0 221.72
R2 A1 A1.n2 156.197
R3 A1.n0 A1.t1 149.421
R4 A1.n1 A1.t3 149.421
R5 A1.n2 A1.n1 58.9116
R6 A1.n2 A1.n0 16.0672
R7 a_926_297.n1 a_926_297.n0 1223.76
R8 a_926_297.n0 a_926_297.t1 26.5955
R9 a_926_297.n0 a_926_297.t2 26.5955
R10 a_926_297.n1 a_926_297.t3 26.5955
R11 a_926_297.t0 a_926_297.n1 26.5955
R12 VPWR.n7 VPWR.t4 862.803
R13 VPWR.n6 VPWR.n5 605.035
R14 VPWR.n15 VPWR.t0 333.079
R15 VPWR.n13 VPWR.n2 309.726
R16 VPWR.n4 VPWR.n3 216.142
R17 VPWR.n2 VPWR.t2 29.5505
R18 VPWR.n2 VPWR.t3 29.5505
R19 VPWR.n14 VPWR.n13 28.2358
R20 VPWR.n3 VPWR.t7 26.5955
R21 VPWR.n3 VPWR.t1 26.5955
R22 VPWR.n5 VPWR.t5 26.5955
R23 VPWR.n5 VPWR.t6 26.5955
R24 VPWR.n12 VPWR.n4 23.3417
R25 VPWR.n8 VPWR.n4 21.0829
R26 VPWR.n8 VPWR.n7 18.824
R27 VPWR.n13 VPWR.n12 16.1887
R28 VPWR.n15 VPWR.n14 13.5534
R29 VPWR.n9 VPWR.n8 9.3005
R30 VPWR.n10 VPWR.n4 9.3005
R31 VPWR.n12 VPWR.n11 9.3005
R32 VPWR.n13 VPWR.n1 9.3005
R33 VPWR.n14 VPWR.n0 9.3005
R34 VPWR.n16 VPWR.n15 9.3005
R35 VPWR.n7 VPWR.n6 7.23807
R36 VPWR.n9 VPWR.n6 0.155689
R37 VPWR.n10 VPWR.n9 0.120292
R38 VPWR.n11 VPWR.n10 0.120292
R39 VPWR.n11 VPWR.n1 0.120292
R40 VPWR.n1 VPWR.n0 0.120292
R41 VPWR.n16 VPWR.n0 0.120292
R42 VPWR VPWR.n16 0.0278438
R43 VPB.t8 VPB.t3 580.062
R44 VPB VPB.t4 272.274
R45 VPB.t7 VPB.t6 266.356
R46 VPB.t11 VPB.t8 260.437
R47 VPB.t9 VPB.t1 248.599
R48 VPB.t10 VPB.t9 248.599
R49 VPB.t0 VPB.t10 248.599
R50 VPB.t2 VPB.t0 248.599
R51 VPB.t3 VPB.t2 248.599
R52 VPB.t5 VPB.t11 248.599
R53 VPB.t6 VPB.t5 248.599
R54 VPB.t4 VPB.t7 248.599
R55 a_496_47.n4 a_496_47.t6 328.925
R56 a_496_47.n2 a_496_47.t1 254.749
R57 a_496_47.n3 a_496_47.n0 190.648
R58 a_496_47.n2 a_496_47.n1 190.648
R59 a_496_47.n5 a_496_47.n4 185
R60 a_496_47.n4 a_496_47.n3 49.5971
R61 a_496_47.n3 a_496_47.n2 43.0085
R62 a_496_47.t0 a_496_47.n5 30.462
R63 a_496_47.n5 a_496_47.t2 26.7697
R64 a_496_47.n0 a_496_47.t7 24.9236
R65 a_496_47.n0 a_496_47.t3 24.9236
R66 a_496_47.n1 a_496_47.t5 24.9236
R67 a_496_47.n1 a_496_47.t4 24.9236
R68 VGND.n24 VGND.t4 268.077
R69 VGND.n7 VGND.n6 203.972
R70 VGND.n9 VGND.n8 198.964
R71 VGND.n12 VGND.n11 198.964
R72 VGND.n22 VGND.n2 198.964
R73 VGND.n18 VGND.t2 150.618
R74 VGND.n16 VGND.n4 34.6358
R75 VGND.n17 VGND.n16 34.6358
R76 VGND.n23 VGND.n22 28.2358
R77 VGND.n2 VGND.t3 27.6928
R78 VGND.n2 VGND.t1 27.6928
R79 VGND.n6 VGND.t5 24.9236
R80 VGND.n6 VGND.t8 24.9236
R81 VGND.n8 VGND.t7 24.9236
R82 VGND.n8 VGND.t9 24.9236
R83 VGND.n11 VGND.t6 24.9236
R84 VGND.n11 VGND.t0 24.9236
R85 VGND.n18 VGND.n1 24.4711
R86 VGND.n12 VGND.n4 23.3417
R87 VGND.n12 VGND.n10 21.0829
R88 VGND.n18 VGND.n17 21.0829
R89 VGND.n10 VGND.n9 17.3181
R90 VGND.n24 VGND.n23 16.2963
R91 VGND.n22 VGND.n1 16.1887
R92 VGND.n25 VGND.n24 12.2465
R93 VGND.n23 VGND.n0 9.3005
R94 VGND.n22 VGND.n21 9.3005
R95 VGND.n20 VGND.n1 9.3005
R96 VGND.n19 VGND.n18 9.3005
R97 VGND.n10 VGND.n5 9.3005
R98 VGND.n13 VGND.n12 9.3005
R99 VGND.n14 VGND.n4 9.3005
R100 VGND.n16 VGND.n15 9.3005
R101 VGND.n17 VGND.n3 9.3005
R102 VGND.n9 VGND.n7 6.69995
R103 VGND.n7 VGND.n5 0.699886
R104 VGND.n13 VGND.n5 0.120292
R105 VGND.n14 VGND.n13 0.120292
R106 VGND.n15 VGND.n14 0.120292
R107 VGND.n15 VGND.n3 0.120292
R108 VGND.n19 VGND.n3 0.120292
R109 VGND.n20 VGND.n19 0.120292
R110 VGND.n21 VGND.n20 0.120292
R111 VGND.n21 VGND.n0 0.120292
R112 VGND.n25 VGND.n0 0.120292
R113 VGND VGND.n25 0.0278438
R114 VNB.t2 VNB.t10 2733.98
R115 VNB.t6 VNB.t0 1310.03
R116 VNB VNB.t4 1310.03
R117 VNB.t1 VNB.t3 1281.55
R118 VNB.t9 VNB.t5 1196.12
R119 VNB.t8 VNB.t9 1196.12
R120 VNB.t11 VNB.t8 1196.12
R121 VNB.t7 VNB.t11 1196.12
R122 VNB.t0 VNB.t7 1196.12
R123 VNB.t10 VNB.t6 1196.12
R124 VNB.t3 VNB.t2 1196.12
R125 VNB.t4 VNB.t1 1196.12
R126 A3.n0 A3.t1 221.72
R127 A3.n1 A3.t2 221.72
R128 A3 A3.n2 156.407
R129 A3.n0 A3.t3 149.421
R130 A3.n1 A3.t0 149.421
R131 A3.n2 A3.n1 38.382
R132 A3.n2 A3.n0 36.5968
R133 a_102_21.n10 a_102_21.n9 378.815
R134 a_102_21.n11 a_102_21.n10 293.06
R135 a_102_21.n8 a_102_21.n0 224.424
R136 a_102_21.n4 a_102_21.t8 221.72
R137 a_102_21.n5 a_102_21.t10 221.72
R138 a_102_21.n2 a_102_21.t11 221.72
R139 a_102_21.n1 a_102_21.t13 221.72
R140 a_102_21.n7 a_102_21.n6 152
R141 a_102_21.n4 a_102_21.t6 149.421
R142 a_102_21.n5 a_102_21.t7 149.421
R143 a_102_21.n2 a_102_21.t12 149.421
R144 a_102_21.n1 a_102_21.t9 149.421
R145 a_102_21.n7 a_102_21.n3 86.1555
R146 a_102_21.n2 a_102_21.n1 74.9783
R147 a_102_21.n6 a_102_21.n5 58.9116
R148 a_102_21.n3 a_102_21.n2 44.8609
R149 a_102_21.n10 a_102_21.n8 41.5825
R150 a_102_21.n8 a_102_21.n7 40.3069
R151 a_102_21.n11 a_102_21.t5 30.5355
R152 a_102_21.n9 a_102_21.t3 26.5955
R153 a_102_21.n9 a_102_21.t2 26.5955
R154 a_102_21.t1 a_102_21.n11 26.5955
R155 a_102_21.n5 a_102_21.n3 25.861
R156 a_102_21.n0 a_102_21.t0 24.9236
R157 a_102_21.n0 a_102_21.t4 24.9236
R158 a_102_21.n6 a_102_21.n4 16.0672
R159 X.n8 X.n5 356.098
R160 X.n8 X.n6 312.658
R161 X.n3 X.n2 232.304
R162 X.n1 X.n0 185
R163 X X.n3 88.146
R164 X.n9 X.n4 73.3096
R165 X.n5 X.t3 26.5955
R166 X.n5 X.t2 26.5955
R167 X.n6 X.t1 26.5955
R168 X.n6 X.t0 26.5955
R169 X.n0 X.t4 24.9236
R170 X.n0 X.t5 24.9236
R171 X.n2 X.t7 24.9236
R172 X.n2 X.t6 24.9236
R173 X X.n9 6.88453
R174 X.n8 X.n7 5.95399
R175 X.n9 X 4.65505
R176 X.n7 X 3.49141
R177 X.n4 X.n1 3.33963
R178 X X.n8 2.47445
R179 X.n4 X 1.16414
R180 X.n3 X.n1 1.11354
R181 X.n7 X 0.893523
R182 X.n9 X 0.430752
R183 A2.n0 A2.t1 241.536
R184 A2.n2 A2.t3 241.439
R185 A2.n0 A2.t0 169.237
R186 A2.n2 A2.t2 169.138
R187 A2.n1 A2.n0 152
R188 A2.n3 A2.n2 152
R189 A2.n1 A2 11.3316
R190 A2 A2.n1 7.97427
R191 A2 A2.n3 5.1026
R192 A2.n3 A2 0.985115
R193 a_672_297.n0 a_672_297.t2 920.986
R194 a_672_297.n0 a_672_297.t0 749.322
R195 a_672_297.n1 a_672_297.n0 288.212
R196 a_672_297.t1 a_672_297.n1 26.5955
R197 a_672_297.n1 a_672_297.t3 26.5955
R198 B1.n0 B1.t0 300.269
R199 B1.n0 B1.t3 221.72
R200 B1.n2 B1.t2 172.627
R201 B1.n3 B1.n2 152
R202 B1.n1 B1.t1 149.421
R203 B1.n2 B1.n1 51.7709
R204 B1.n1 B1.n0 17.8524
R205 B1.n4 B1 8.3205
R206 B1 B1.n4 8.3032
R207 B1.n3 B1 1.9032
R208 B1.n4 B1.n3 1.55726
C0 VGND VPB 0.008895f
C1 X B1 2.08e-19
C2 VPWR A3 0.023946f
C3 A1 VGND 0.027449f
C4 A1 VPB 0.051503f
C5 VGND B1 0.025447f
C6 VPWR A2 0.028239f
C7 VPB B1 0.090073f
C8 VGND A3 0.030304f
C9 VPB A3 0.057616f
C10 VGND A2 0.035866f
C11 B1 A3 0.06365f
C12 VPB A2 0.073668f
C13 A1 A2 0.212472f
C14 B1 A2 0.002794f
C15 A3 A2 0.08625f
C16 VPWR X 0.396699f
C17 VPWR VGND 0.087393f
C18 VPWR VPB 0.133978f
C19 A1 VPWR 0.021889f
C20 X VGND 0.28516f
C21 VPWR B1 0.05007f
C22 X VPB 0.015061f
C23 VGND VNB 0.727012f
C24 X VNB 0.06309f
C25 VPWR VNB 0.607096f
C26 A1 VNB 0.167317f
C27 A2 VNB 0.24143f
C28 A3 VNB 0.168689f
C29 B1 VNB 0.228809f
C30 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31ai_1 VPB VNB A1 A2 A3 Y B1 VPWR VGND
X0 Y.t2 B1.t0 a_109_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1 Y.t0 A3.t0 a_193_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297.t0 A2.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t0 A2.t1 a_109_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t0 B1.t1 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X5 a_109_47.t1 A3.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_297.t1 A1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47.t2 A1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n0 B1.t1 212.081
R1 B1 B1.n0 193.615
R2 B1.n0 B1.t0 165.341
R3 a_109_47.n1 a_109_47.n0 237.103
R4 a_109_47.n0 a_109_47.t3 84.9236
R5 a_109_47.n0 a_109_47.t1 27.6928
R6 a_109_47.t0 a_109_47.n1 24.9236
R7 a_109_47.n1 a_109_47.t2 24.9236
R8 Y.n2 Y 595.419
R9 Y.n3 Y.n2 585
R10 Y.n0 Y.t2 128.5
R11 Y.n2 Y.t0 127.066
R12 Y.n2 Y.t1 27.5805
R13 Y Y.n1 16.6703
R14 Y.n3 Y 11.3121
R15 Y Y.n3 8.93073
R16 Y.n1 Y.n0 6.57041
R17 Y.n1 Y 3.57259
R18 Y.n0 Y 2.49254
R19 Y.n1 Y 1.35979
R20 VNB.t1 VNB.t3 2164.4
R21 VNB.t0 VNB.t1 1196.12
R22 VNB.t2 VNB.t0 1196.12
R23 VNB VNB.t2 911.327
R24 A3.n0 A3.t0 232.472
R25 A3.n0 A3.t1 160.173
R26 A3 A3.n0 153.482
R27 a_193_297.t0 a_193_297.t1 53.1905
R28 VPB.t1 VPB.t2 553.428
R29 VPB.t0 VPB.t1 248.599
R30 VPB.t3 VPB.t0 248.599
R31 VPB VPB.t3 189.409
R32 A2.n0 A2.t0 241.536
R33 A2.n0 A2.t1 169.237
R34 A2.n1 A2.n0 152
R35 A2 A2.n1 8.19825
R36 A2.n1 A2 1.58252
R37 a_109_297.t0 a_109_297.t1 53.1905
R38 VGND.n1 VGND.n0 217.203
R39 VGND.n1 VGND.t2 169.786
R40 VGND.n0 VGND.t1 24.9236
R41 VGND.n0 VGND.t0 24.9236
R42 VGND VGND.n1 0.512003
R43 VPWR.n0 VPWR.t0 257.87
R44 VPWR.n0 VPWR.t1 249.114
R45 VPWR VPWR.n0 0.0633232
R46 A1.n0 A1.t0 230.363
R47 A1.n0 A1.t1 158.064
R48 A1 A1.n0 157.376
C0 B1 VPWR 0.059285f
C1 A2 A3 0.136905f
C2 B1 Y 0.099222f
C3 VPWR Y 0.127902f
C4 B1 VGND 0.009398f
C5 B1 VPB 0.054005f
C6 VPWR VGND 0.059246f
C7 VPWR VPB 0.075586f
C8 Y VGND 0.097538f
C9 Y VPB 0.004596f
C10 VPWR A1 0.058076f
C11 VPWR A2 0.146446f
C12 B1 A3 0.027405f
C13 VGND VPB 0.005833f
C14 Y A1 3.1e-19
C15 VGND A1 0.041685f
C16 Y A2 0.004498f
C17 VPWR A3 0.047373f
C18 VPB A1 0.037546f
C19 VGND A2 0.016981f
C20 Y A3 0.113883f
C21 VPB A2 0.030204f
C22 VGND A3 0.017789f
C23 VPB A3 0.040048f
C24 A1 A2 0.088074f
C25 VGND VNB 0.373865f
C26 Y VNB 0.05192f
C27 VPWR VNB 0.360149f
C28 B1 VNB 0.172832f
C29 A3 VNB 0.106588f
C30 A2 VNB 0.093658f
C31 A1 VNB 0.142767f
C32 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31ai_2 VGND VPWR VPB VNB Y A3 A2 A1 B1
X0 a_281_297.t3 A3.t0 Y.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1 a_281_297.t1 A2.t0 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t1 A2.t1 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297.t0 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47.t5 A1.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t5 A1.t2 a_27_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_27_47.t4 A3.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR.t0 B1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t1 A1.t3 a_27_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_27_47.t7 B1.t1 Y.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X10 a_27_47.t1 A2.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.19825 ps=1.26 w=0.65 l=0.15
X11 VGND.t2 A3.t2 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 Y.t1 B1.t2 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t2 A3.t3 a_281_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t4 B1.t3 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X15 a_27_297.t1 A2.t3 a_281_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A3.n0 A3.t3 221.72
R1 A3.n2 A3.t0 221.72
R2 A3.n3 A3.t2 161.917
R3 A3.n1 A3 158.163
R4 A3.n4 A3.n3 152
R5 A3.n0 A3.t1 149.421
R6 A3.n2 A3.n1 58.9116
R7 A3.n1 A3.n0 16.0672
R8 A3 A3.n4 11.8524
R9 A3.n4 A3 9.95606
R10 A3.n3 A3.n2 1.78569
R11 Y.n0 Y 594.115
R12 Y.n5 Y.n4 585
R13 Y.n6 Y.n5 585
R14 Y.n1 Y.n0 585
R15 Y.n3 Y.n2 206.056
R16 Y Y.n8 185.388
R17 Y.n3 Y.n1 42.2793
R18 Y.n8 Y.t1 39.6928
R19 Y.n8 Y.t5 32.3082
R20 Y.n5 Y.t4 26.5955
R21 Y.n0 Y.t3 26.5955
R22 Y.n2 Y.t0 26.5955
R23 Y.n2 Y.t2 26.5955
R24 Y.n7 Y.n6 19.7652
R25 Y.n7 Y.n3 12.8005
R26 Y.n4 Y 12.0476
R27 Y Y.n7 5.23686
R28 Y.n1 Y 4.07323
R29 Y.n4 Y 0.753441
R30 Y.n6 Y 0.753441
R31 a_281_297.n1 a_281_297.n0 1298
R32 a_281_297.n0 a_281_297.t0 26.5955
R33 a_281_297.n0 a_281_297.t1 26.5955
R34 a_281_297.t2 a_281_297.n1 26.5955
R35 a_281_297.n1 a_281_297.t3 26.5955
R36 VPB.t1 VPB.t5 568.225
R37 VPB.t0 VPB.t6 319.627
R38 VPB.t4 VPB.t0 248.599
R39 VPB.t5 VPB.t4 248.599
R40 VPB.t2 VPB.t1 248.599
R41 VPB.t3 VPB.t2 248.599
R42 VPB.t7 VPB.t3 248.599
R43 VPB VPB.t7 201.246
R44 A2.n2 A2.t3 221.72
R45 A2.n3 A2.t0 221.72
R46 A2.n1 A2.t2 180.661
R47 A2.n1 A2.n0 152
R48 A2.n5 A2.n4 152
R49 A2.n3 A2.t1 149.421
R50 A2.n4 A2.n3 43.7375
R51 A2.n4 A2.n2 31.2412
R52 A2.n2 A2.n1 29.4561
R53 A2.n5 A2.n0 16.119
R54 A2.n0 A2 3.55606
R55 A2 A2.n5 2.13383
R56 a_27_297.n0 a_27_297.t1 364.635
R57 a_27_297.n0 a_27_297.t3 270.283
R58 a_27_297.n1 a_27_297.n0 206.055
R59 a_27_297.t2 a_27_297.n1 26.5955
R60 a_27_297.n1 a_27_297.t0 26.5955
R61 a_27_47.n4 a_27_47.t7 312.055
R62 a_27_47.n1 a_27_47.t6 173.317
R63 a_27_47.n1 a_27_47.n0 99.5638
R64 a_27_47.n3 a_27_47.n2 99.5638
R65 a_27_47.n5 a_27_47.n4 89.3175
R66 a_27_47.n3 a_27_47.n1 67.0123
R67 a_27_47.n4 a_27_47.n3 60.6938
R68 a_27_47.n2 a_27_47.t3 39.6928
R69 a_27_47.n2 a_27_47.t1 32.3082
R70 a_27_47.n0 a_27_47.t2 24.9236
R71 a_27_47.n0 a_27_47.t5 24.9236
R72 a_27_47.t0 a_27_47.n5 24.9236
R73 a_27_47.n5 a_27_47.t4 24.9236
R74 VGND.n1 VGND.n0 207.213
R75 VGND.n5 VGND.n4 204.025
R76 VGND.n9 VGND.n8 185
R77 VGND.n7 VGND.n6 185
R78 VGND.n8 VGND.n7 62.7697
R79 VGND.n4 VGND.t3 39.6928
R80 VGND.n10 VGND.n1 33.8829
R81 VGND.n7 VGND.t0 24.9236
R82 VGND.n8 VGND.t1 24.9236
R83 VGND.n4 VGND.t2 24.9236
R84 VGND.n0 VGND.t4 24.9236
R85 VGND.n0 VGND.t5 24.9236
R86 VGND.n10 VGND.n9 24.6922
R87 VGND.n6 VGND.n5 16.7157
R88 VGND.n11 VGND.n10 9.3005
R89 VGND.n3 VGND.n2 9.3005
R90 VGND.n12 VGND.n1 8.41204
R91 VGND.n6 VGND.n3 5.48621
R92 VGND.n9 VGND.n3 1.42272
R93 VGND.n5 VGND.n2 0.618089
R94 VGND.n12 VGND.n11 0.141672
R95 VGND VGND.n12 0.120476
R96 VGND.n11 VGND.n2 0.120292
R97 VNB.t2 VNB.t1 2164.4
R98 VNB.t0 VNB.t7 1537.86
R99 VNB.t1 VNB.t3 1537.86
R100 VNB.t3 VNB.t4 1423.95
R101 VNB.t4 VNB.t0 1196.12
R102 VNB.t5 VNB.t2 1196.12
R103 VNB.t6 VNB.t5 1196.12
R104 VNB VNB.t6 968.285
R105 A1.n0 A1.t0 221.72
R106 A1.n2 A1.t3 221.72
R107 A1.n2 A1.n1 153.786
R108 A1.n4 A1.n3 152
R109 A1.n0 A1.t1 149.421
R110 A1.n2 A1.t2 149.421
R111 A1.n3 A1.n2 58.9116
R112 A1.n3 A1.n0 16.0672
R113 A1.n1 A1 15.6449
R114 A1 A1.n4 11.8524
R115 A1.n4 A1 9.95606
R116 A1.n1 A1 6.16346
R117 VPWR.n2 VPWR.n0 327.945
R118 VPWR.n2 VPWR.n1 316.202
R119 VPWR.n1 VPWR.t0 42.3555
R120 VPWR.n1 VPWR.t3 34.4755
R121 VPWR.n0 VPWR.t2 26.5955
R122 VPWR.n0 VPWR.t1 26.5955
R123 VPWR VPWR.n2 0.149281
R124 B1.n1 B1.t3 212.081
R125 B1.n0 B1.t0 212.081
R126 B1 B1.n1 193.507
R127 B1.n1 B1.t1 139.78
R128 B1.n0 B1.t2 139.78
R129 B1.n1 B1.n0 78.8732
C0 VPB B1 0.080569f
C1 VPB VPWR 0.09313f
C2 VPB A2 0.075182f
C3 VPB Y 0.024814f
C4 A1 VPWR 0.032669f
C5 A1 A2 0.077584f
C6 A1 Y 2.19e-19
C7 A3 VGND 0.03168f
C8 B1 VGND 0.022648f
C9 A3 B1 0.053228f
C10 VPWR VGND 0.089341f
C11 A3 VPWR 0.020628f
C12 A2 VGND 0.031806f
C13 VPB A1 0.062544f
C14 A2 A3 0.052603f
C15 Y VGND 0.01598f
C16 B1 VPWR 0.041228f
C17 A3 Y 0.113339f
C18 B1 Y 0.160721f
C19 A2 VPWR 0.022144f
C20 VPWR Y 0.258059f
C21 A2 Y 5.06e-19
C22 VPB VGND 0.009256f
C23 VPB A3 0.062789f
C24 A1 VGND 0.030858f
C25 VGND VNB 0.522607f
C26 Y VNB 0.055751f
C27 VPWR VNB 0.440807f
C28 B1 VNB 0.26682f
C29 A3 VNB 0.186976f
C30 A2 VNB 0.213289f
C31 A1 VNB 0.222131f
C32 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31ai_4 VGND VPWR VPB VNB A1 Y B1 A3 A2
X0 Y.t9 A3.t0 a_449_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t7 A1.t0 a_27_297.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_449_297.t4 A3.t1 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y.t7 A3.t2 a_449_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t9 A1.t1 a_31_47.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297.t4 A1.t2 VPWR.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t10 B1.t0 a_31_47.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_449_297.t2 A3.t3 Y.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2628 ps=2.57 w=1 l=0.15
X8 Y.t11 B1.t1 a_31_47.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_31_47.t10 A1.t3 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297.t7 A2.t0 a_449_297.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.2605 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t7 A1.t4 a_31_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_31_47.t8 A1.t5 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t0 B1.t2 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_31_47.t14 A2.t1 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_31_47.t15 A2.t2 VGND.t11 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_449_297.t0 A2.t3 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR.t1 B1.t3 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t2 B1.t4 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t5 A1.t6 a_27_297.t3 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 VGND.t0 A2.t4 a_31_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR.t3 B1.t5 Y.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND.t1 A2.t5 a_31_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VGND.t5 A3.t4 a_31_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.222625 pd=1.335 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_31_47.t6 A3.t5 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.222625 ps=1.335 w=0.65 l=0.15
X25 a_27_297.t1 A2.t6 a_449_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND.t3 A3.t6 a_31_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 a_31_47.t4 A3.t7 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X28 a_449_297.t6 A2.t7 a_27_297.t6 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_31_47.t2 B1.t6 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_27_297.t2 A1.t7 VPWR.t4 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_31_47.t3 B1.t7 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A3.n0 A3.t0 221.72
R1 A3.n13 A3.t1 221.72
R2 A3.n1 A3.t2 221.72
R3 A3.n7 A3.t3 221.72
R4 A3.n3 A3.t4 165.488
R5 A3.n15 A3.n14 152
R6 A3.n11 A3.n10 152
R7 A3.n9 A3.n8 152
R8 A3.n6 A3.n5 152
R9 A3.n4 A3.n3 152
R10 A3.n0 A3.t7 149.421
R11 A3.n2 A3.t5 149.421
R12 A3.n12 A3.t6 149.421
R13 A3.n14 A3.n0 61.5894
R14 A3.n6 A3.n3 60.6968
R15 A3.n8 A3.n7 41.9524
R16 A3.n11 A3.n1 27.6709
R17 A3.n12 A3.n11 25.8857
R18 A3.n13 A3.n12 21.4227
R19 A3.n2 A3.n1 21.4227
R20 A3 A3.n15 21.2369
R21 A3.n5 A3.n4 19.7823
R22 A3.n9 A3 19.4914
R23 A3.n7 A3.n6 18.7449
R24 A3.n10 A3 14.255
R25 A3.n14 A3.n13 13.3894
R26 A3.n10 A3 12.5096
R27 A3.n8 A3.n2 11.6042
R28 A3 A3.n9 7.27323
R29 A3.n4 A3 6.4005
R30 A3.n15 A3 5.52777
R31 A3.n5 A3 0.291409
R32 a_449_297.n4 a_449_297.n3 644.321
R33 a_449_297.n5 a_449_297.n4 585
R34 a_449_297.n2 a_449_297.n0 310.421
R35 a_449_297.n2 a_449_297.n1 292.5
R36 a_449_297.n4 a_449_297.n2 57.9519
R37 a_449_297.n3 a_449_297.t1 26.5955
R38 a_449_297.n3 a_449_297.t6 26.5955
R39 a_449_297.n1 a_449_297.t3 26.5955
R40 a_449_297.n1 a_449_297.t2 26.5955
R41 a_449_297.n0 a_449_297.t5 26.5955
R42 a_449_297.n0 a_449_297.t4 26.5955
R43 a_449_297.n5 a_449_297.t7 26.5955
R44 a_449_297.t0 a_449_297.n5 26.5955
R45 Y.n12 Y.t6 765.871
R46 Y.n6 Y.n5 585
R47 Y.n7 Y.n6 585
R48 Y.n14 Y.n13 585
R49 Y.n2 Y.n0 229.8
R50 Y.n15 Y.n11 206
R51 Y.n9 Y.n4 206
R52 Y.n2 Y.n1 185
R53 Y.n13 Y.t8 26.5955
R54 Y.n13 Y.t7 26.5955
R55 Y.n11 Y.t3 26.5955
R56 Y.n11 Y.t9 26.5955
R57 Y.n4 Y.t1 26.5955
R58 Y.n4 Y.t2 26.5955
R59 Y.n6 Y.t0 26.5955
R60 Y.n1 Y.t4 24.9236
R61 Y.n1 Y.t10 24.9236
R62 Y.n0 Y.t5 24.9236
R63 Y.n0 Y.t11 24.9236
R64 Y.n10 Y 23.5248
R65 Y Y.n8 20.7365
R66 Y.n10 Y 19.7125
R67 Y.n9 Y 17.9205
R68 Y.n12 Y 17.6645
R69 Y Y.n3 15.2221
R70 Y Y.n15 13.8245
R71 Y.n14 Y 13.8245
R72 Y.n5 Y 11.004
R73 Y.n15 Y 9.7285
R74 Y Y.n14 9.7285
R75 Y.n3 Y 8.3032
R76 Y Y.n9 5.6325
R77 Y Y.n12 5.6325
R78 Y.n8 Y 5.61454
R79 Y.n8 Y.n7 5.38997
R80 Y.n5 Y 4.26717
R81 Y.n7 Y 4.26717
R82 Y.n3 Y.n2 4.0005
R83 Y.n3 Y 4.0005
R84 Y Y.n10 3.8405
R85 VPB.t12 VPB.t6 565.265
R86 VPB.t3 VPB.t2 248.599
R87 VPB.t4 VPB.t3 248.599
R88 VPB.t5 VPB.t4 248.599
R89 VPB.t9 VPB.t5 248.599
R90 VPB.t8 VPB.t9 248.599
R91 VPB.t7 VPB.t8 248.599
R92 VPB.t6 VPB.t7 248.599
R93 VPB.t0 VPB.t12 248.599
R94 VPB.t1 VPB.t0 248.599
R95 VPB.t11 VPB.t1 248.599
R96 VPB.t15 VPB.t11 248.599
R97 VPB.t10 VPB.t15 248.599
R98 VPB.t13 VPB.t10 248.599
R99 VPB.t14 VPB.t13 248.599
R100 VPB VPB.t14 204.207
R101 A1.n1 A1.t7 221.72
R102 A1.n2 A1.t0 221.72
R103 A1.n7 A1.t2 221.72
R104 A1.n8 A1.t6 221.72
R105 A1 A1.n3 154.941
R106 A1.n4 A1.n0 152
R107 A1.n6 A1.n5 152
R108 A1.n10 A1.n9 152
R109 A1.n1 A1.t5 149.421
R110 A1.n2 A1.t1 149.421
R111 A1.n7 A1.t3 149.421
R112 A1.n8 A1.t4 149.421
R113 A1.n6 A1.n0 60.6968
R114 A1.n9 A1.n7 56.2338
R115 A1.n3 A1.n2 50.8783
R116 A1.n3 A1.n1 24.1005
R117 A1.n9 A1.n8 18.7449
R118 A1 A1.n10 15.3951
R119 A1.n5 A1 11.2437
R120 A1.n2 A1.n0 9.81902
R121 A1.n4 A1 8.82212
R122 A1 A1.n4 7.09239
R123 A1.n5 A1 4.67077
R124 A1.n7 A1.n6 4.46346
R125 A1.n10 A1 0.519419
R126 a_27_297.n4 a_27_297.t7 832.289
R127 a_27_297.n5 a_27_297.n4 295.772
R128 a_27_297.n2 a_27_297.t3 249.304
R129 a_27_297.n2 a_27_297.n1 201.392
R130 a_27_297.n3 a_27_297.n0 190.411
R131 a_27_297.n4 a_27_297.n3 36.5751
R132 a_27_297.n3 a_27_297.n2 32.7419
R133 a_27_297.n0 a_27_297.t6 26.5955
R134 a_27_297.n0 a_27_297.t2 26.5955
R135 a_27_297.n1 a_27_297.t5 26.5955
R136 a_27_297.n1 a_27_297.t4 26.5955
R137 a_27_297.t0 a_27_297.n5 26.5955
R138 a_27_297.n5 a_27_297.t1 26.5955
R139 VPWR.n29 VPWR.n1 607.212
R140 VPWR.n27 VPWR.n2 607.212
R141 VPWR.n11 VPWR.n8 315.13
R142 VPWR.n10 VPWR.n9 309.726
R143 VPWR.n14 VPWR.n7 34.6358
R144 VPWR.n15 VPWR.n14 34.6358
R145 VPWR.n16 VPWR.n15 34.6358
R146 VPWR.n16 VPWR.n5 34.6358
R147 VPWR.n20 VPWR.n5 34.6358
R148 VPWR.n21 VPWR.n20 34.6358
R149 VPWR.n22 VPWR.n21 34.6358
R150 VPWR.n22 VPWR.n3 34.6358
R151 VPWR.n26 VPWR.n3 34.6358
R152 VPWR.n29 VPWR.n28 33.8829
R153 VPWR.n28 VPWR.n27 29.3652
R154 VPWR.n10 VPWR.n7 27.1064
R155 VPWR.n1 VPWR.t6 26.5955
R156 VPWR.n1 VPWR.t5 26.5955
R157 VPWR.n2 VPWR.t4 26.5955
R158 VPWR.n2 VPWR.t7 26.5955
R159 VPWR.n9 VPWR.t2 26.5955
R160 VPWR.n9 VPWR.t3 26.5955
R161 VPWR.n8 VPWR.t0 26.5955
R162 VPWR.n8 VPWR.t1 26.5955
R163 VPWR.n12 VPWR.n7 9.3005
R164 VPWR.n14 VPWR.n13 9.3005
R165 VPWR.n15 VPWR.n6 9.3005
R166 VPWR.n17 VPWR.n16 9.3005
R167 VPWR.n18 VPWR.n5 9.3005
R168 VPWR.n20 VPWR.n19 9.3005
R169 VPWR.n21 VPWR.n4 9.3005
R170 VPWR.n23 VPWR.n22 9.3005
R171 VPWR.n24 VPWR.n3 9.3005
R172 VPWR.n26 VPWR.n25 9.3005
R173 VPWR.n28 VPWR.n0 9.3005
R174 VPWR.n30 VPWR.n29 8.41204
R175 VPWR.n11 VPWR.n10 6.20499
R176 VPWR.n27 VPWR.n26 5.27109
R177 VPWR.n12 VPWR.n11 0.653912
R178 VPWR.n30 VPWR.n0 0.141672
R179 VPWR VPWR.n30 0.121778
R180 VPWR.n13 VPWR.n12 0.120292
R181 VPWR.n13 VPWR.n6 0.120292
R182 VPWR.n17 VPWR.n6 0.120292
R183 VPWR.n18 VPWR.n17 0.120292
R184 VPWR.n19 VPWR.n18 0.120292
R185 VPWR.n19 VPWR.n4 0.120292
R186 VPWR.n23 VPWR.n4 0.120292
R187 VPWR.n24 VPWR.n23 0.120292
R188 VPWR.n25 VPWR.n24 0.120292
R189 VPWR.n25 VPWR.n0 0.120292
R190 a_31_47.n7 a_31_47.n2 196.672
R191 a_31_47.n4 a_31_47.n3 185
R192 a_31_47.n6 a_31_47.n5 185
R193 a_31_47.n4 a_31_47.t3 180.133
R194 a_31_47.n1 a_31_47.t9 175.868
R195 a_31_47.n9 a_31_47.n8 99.5638
R196 a_31_47.n11 a_31_47.n10 99.5638
R197 a_31_47.n1 a_31_47.n0 99.5638
R198 a_31_47.n13 a_31_47.n12 99.5638
R199 a_31_47.n7 a_31_47.n6 83.9534
R200 a_31_47.n9 a_31_47.n7 82.0711
R201 a_31_47.n6 a_31_47.n4 55.2732
R202 a_31_47.n11 a_31_47.n9 38.4005
R203 a_31_47.n12 a_31_47.n1 38.4005
R204 a_31_47.n12 a_31_47.n11 38.4005
R205 a_31_47.n2 a_31_47.t5 24.9236
R206 a_31_47.n2 a_31_47.t6 24.9236
R207 a_31_47.n5 a_31_47.t12 24.9236
R208 a_31_47.n5 a_31_47.t4 24.9236
R209 a_31_47.n3 a_31_47.t13 24.9236
R210 a_31_47.n3 a_31_47.t2 24.9236
R211 a_31_47.n8 a_31_47.t7 24.9236
R212 a_31_47.n8 a_31_47.t15 24.9236
R213 a_31_47.n10 a_31_47.t1 24.9236
R214 a_31_47.n10 a_31_47.t14 24.9236
R215 a_31_47.n0 a_31_47.t11 24.9236
R216 a_31_47.n0 a_31_47.t10 24.9236
R217 a_31_47.t0 a_31_47.n13 24.9236
R218 a_31_47.n13 a_31_47.t8 24.9236
R219 VGND.n20 VGND.n7 207.213
R220 VGND.n5 VGND.n4 207.213
R221 VGND.n27 VGND.n3 207.213
R222 VGND.n1 VGND.n0 207.213
R223 VGND.n10 VGND.n9 190.28
R224 VGND.n14 VGND.n13 185
R225 VGND.n12 VGND.n11 185
R226 VGND.n13 VGND.n12 62.7697
R227 VGND.n13 VGND.t5 38.7697
R228 VGND.n9 VGND.t2 36.0005
R229 VGND.n9 VGND.t3 36.0005
R230 VGND.n19 VGND.n8 34.6358
R231 VGND.n22 VGND.n21 34.6358
R232 VGND.n26 VGND.n25 34.6358
R233 VGND.n28 VGND.n1 33.8829
R234 VGND.n28 VGND.n27 29.3652
R235 VGND.n12 VGND.t4 24.9236
R236 VGND.n7 VGND.t11 24.9236
R237 VGND.n7 VGND.t1 24.9236
R238 VGND.n4 VGND.t10 24.9236
R239 VGND.n4 VGND.t0 24.9236
R240 VGND.n3 VGND.t6 24.9236
R241 VGND.n3 VGND.t9 24.9236
R242 VGND.n0 VGND.t8 24.9236
R243 VGND.n0 VGND.t7 24.9236
R244 VGND.n11 VGND.n10 23.5636
R245 VGND.n25 VGND.n5 23.3417
R246 VGND.n20 VGND.n19 17.3181
R247 VGND.n21 VGND.n20 17.3181
R248 VGND.n22 VGND.n5 11.2946
R249 VGND.n29 VGND.n28 9.3005
R250 VGND.n26 VGND.n2 9.3005
R251 VGND.n25 VGND.n24 9.3005
R252 VGND.n23 VGND.n22 9.3005
R253 VGND.n21 VGND.n6 9.3005
R254 VGND.n19 VGND.n18 9.3005
R255 VGND.n17 VGND.n8 9.3005
R256 VGND.n16 VGND.n15 9.3005
R257 VGND.n14 VGND.n8 9.24494
R258 VGND.n30 VGND.n1 8.41204
R259 VGND.n27 VGND.n26 5.27109
R260 VGND.n15 VGND.n14 4.7751
R261 VGND.n15 VGND.n11 2.13383
R262 VGND.n16 VGND.n10 1.51263
R263 VGND.n30 VGND.n29 0.141672
R264 VGND VGND.n30 0.121778
R265 VGND.n17 VGND.n16 0.120292
R266 VGND.n18 VGND.n17 0.120292
R267 VGND.n18 VGND.n6 0.120292
R268 VGND.n23 VGND.n6 0.120292
R269 VGND.n24 VGND.n23 0.120292
R270 VGND.n24 VGND.n2 0.120292
R271 VGND.n29 VGND.n2 0.120292
R272 VNB.t7 VNB.t6 2377.99
R273 VNB.t5 VNB.t4 1537.86
R274 VNB.t13 VNB.t3 1196.12
R275 VNB.t2 VNB.t13 1196.12
R276 VNB.t12 VNB.t2 1196.12
R277 VNB.t4 VNB.t12 1196.12
R278 VNB.t6 VNB.t5 1196.12
R279 VNB.t15 VNB.t7 1196.12
R280 VNB.t1 VNB.t15 1196.12
R281 VNB.t14 VNB.t1 1196.12
R282 VNB.t0 VNB.t14 1196.12
R283 VNB.t8 VNB.t0 1196.12
R284 VNB.t11 VNB.t8 1196.12
R285 VNB.t10 VNB.t11 1196.12
R286 VNB.t9 VNB.t10 1196.12
R287 VNB VNB.t9 982.524
R288 B1.n1 B1.t2 221.72
R289 B1.n5 B1.t3 221.72
R290 B1.n7 B1.t4 221.72
R291 B1.n6 B1.t5 221.72
R292 B1.n3 B1.n2 152
R293 B1.n4 B1.n0 152
R294 B1.n9 B1.n8 152
R295 B1.n1 B1.t7 149.421
R296 B1.n5 B1.t1 149.421
R297 B1.n7 B1.t6 149.421
R298 B1.n6 B1.t0 149.421
R299 B1.n7 B1.n6 74.9783
R300 B1.n4 B1.n3 60.6968
R301 B1.n8 B1.n5 49.0931
R302 B1.n8 B1.n7 25.8857
R303 B1.n9 B1.n0 19.7823
R304 B1.n2 B1 15.4187
R305 B1.n5 B1.n4 11.6042
R306 B1.n2 B1 11.346
R307 B1 B1.n0 4.36414
R308 B1.n3 B1.n1 2.67828
R309 B1 B1.n9 2.61868
R310 A2.n1 A2.t0 221.72
R311 A2.n2 A2.t3 221.72
R312 A2.n8 A2.t6 221.72
R313 A2.n9 A2.t7 221.72
R314 A2.n4 A2.n3 152
R315 A2.n5 A2.n0 152
R316 A2.n7 A2.n6 152
R317 A2.n11 A2.n10 152
R318 A2.n1 A2.t2 149.421
R319 A2.n2 A2.t5 149.421
R320 A2.n8 A2.t1 149.421
R321 A2.n9 A2.t4 149.421
R322 A2.n7 A2.n0 60.6968
R323 A2.n10 A2.n8 58.9116
R324 A2.n3 A2.n2 48.2005
R325 A2.n3 A2.n1 26.7783
R326 A2.n10 A2.n9 16.0672
R327 A2.n2 A2.n0 12.4968
R328 A2.n5 A2.n4 11.7627
R329 A2.n6 A2 10.7248
R330 A2 A2.n11 9.34104
R331 A2.n11 A2 6.57347
R332 A2.n6 A2 5.18969
R333 A2.n4 A2 3.11401
R334 A2.n8 A2.n7 1.78569
R335 A2 A2.n5 1.03834
C0 Y A1 3.34e-19
C1 VPWR A2 0.030113f
C2 VPB A1 0.124631f
C3 A2 A3 0.058653f
C4 Y A2 0.003818f
C5 VGND A1 0.060402f
C6 VPWR A3 0.030497f
C7 VPB A2 0.127479f
C8 A2 B1 5.04e-20
C9 VPWR Y 0.388444f
C10 VPWR VPB 0.14494f
C11 VGND A2 0.050456f
C12 VPWR B1 0.080946f
C13 Y A3 0.246233f
C14 VPB A3 0.146714f
C15 A3 B1 0.053857f
C16 VPWR VGND 0.150466f
C17 Y VPB 0.031782f
C18 Y B1 0.308241f
C19 VGND A3 0.071616f
C20 VPB B1 0.122991f
C21 Y VGND 0.027144f
C22 VGND VPB 0.009713f
C23 VGND B1 0.035568f
C24 A1 A2 0.083775f
C25 VPWR A1 0.061805f
C26 VGND VNB 0.841426f
C27 Y VNB 0.062783f
C28 VPWR VNB 0.705525f
C29 B1 VNB 0.398183f
C30 A3 VNB 0.419748f
C31 A2 VNB 0.357083f
C32 A1 VNB 0.398845f
C33 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32a_1 VPB VNB VPWR VGND X A1 A2 A3 B2 B1
X0 a_77_199.t1 B2.t0 a_227_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1 a_323_297.t1 A2.t0 a_227_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297.t1 A1.t0 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47.t4 B1.t0 a_77_199.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4 VGND.t3 a_77_199.t4 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR.t1 B1.t1 a_539_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47.t0 A3.t0 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 VPWR.t2 a_77_199.t5 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199.t0 A3.t1 a_323_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND.t2 A2.t1 a_227_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 a_227_47.t2 A1.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_539_297.t1 B2.t1 a_77_199.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
R0 B2.n0 B2.t1 236.18
R1 B2.n0 B2.t0 163.881
R2 B2.n1 B2.n0 152
R3 B2.n1 B2 10.2766
R4 B2 B2.n1 1.9836
R5 a_227_47.n1 a_227_47.t4 315.522
R6 a_227_47.n1 a_227_47.n0 159.321
R7 a_227_47.n2 a_227_47.n1 89.3175
R8 a_227_47.t0 a_227_47.n2 40.6159
R9 a_227_47.n0 a_227_47.t2 31.3851
R10 a_227_47.n2 a_227_47.t3 31.3851
R11 a_227_47.n0 a_227_47.t1 29.539
R12 a_77_199.n2 a_77_199.n0 335.647
R13 a_77_199.n2 a_77_199.n1 308.558
R14 a_77_199.n3 a_77_199.n2 289.24
R15 a_77_199.n0 a_77_199.t5 236.18
R16 a_77_199.n0 a_77_199.t4 163.881
R17 a_77_199.n1 a_77_199.t3 42.462
R18 a_77_199.n3 a_77_199.t2 39.4005
R19 a_77_199.t0 a_77_199.n3 37.4305
R20 a_77_199.n1 a_77_199.t1 33.2313
R21 VNB.t3 VNB.t5 1594.82
R22 VNB.t0 VNB.t3 1537.86
R23 VNB.t1 VNB.t0 1537.86
R24 VNB VNB.t4 1423.95
R25 VNB.t2 VNB.t1 1366.99
R26 VNB.t4 VNB.t2 1196.12
R27 A2.n0 A2.t0 236.18
R28 A2.n0 A2.t1 163.881
R29 A2.n1 A2.n0 152
R30 A2 A2.n1 10.8484
R31 A2.n1 A2 2.04108
R32 a_227_297.t0 a_227_297.t1 65.0105
R33 a_323_297.t0 a_323_297.t1 76.8305
R34 VPB.t4 VPB.t1 331.464
R35 VPB.t0 VPB.t4 319.627
R36 VPB.t2 VPB.t0 319.627
R37 VPB VPB.t5 295.95
R38 VPB.t3 VPB.t2 284.113
R39 VPB.t5 VPB.t3 248.599
R40 A1.n0 A1.t0 236.18
R41 A1.n0 A1.t1 163.881
R42 A1 A1.n0 154.816
R43 VPWR.n1 VPWR.n0 318.534
R44 VPWR.n1 VPWR.t1 254.321
R45 VPWR.n0 VPWR.t0 26.5955
R46 VPWR.n0 VPWR.t2 26.5955
R47 VPWR VPWR.n1 0.168791
R48 B1.n0 B1.t1 229.184
R49 B1.n0 B1.t0 156.883
R50 B1 B1.n0 154.56
R51 X.t1 X 769.845
R52 X.n1 X.t1 717.313
R53 X.n0 X.t0 130.138
R54 X.n1 X.n0 64.0315
R55 X.n0 X 3.7234
R56 X X.n1 0.831669
R57 VGND.n2 VGND.n0 218.712
R58 VGND.n2 VGND.n1 205.607
R59 VGND.n1 VGND.t1 36.0005
R60 VGND.n1 VGND.t2 36.0005
R61 VGND.n0 VGND.t0 24.9236
R62 VGND.n0 VGND.t3 24.9236
R63 VGND VGND.n2 0.565628
R64 a_539_297.t0 a_539_297.t1 80.7705
R65 A3.n0 A3.t1 236.18
R66 A3.n0 A3.t0 163.881
R67 A3.n1 A3.n0 152
R68 A3.n1 A3 13.266
R69 A3 A3.n1 2.5605
C0 A1 VPWR 0.018718f
C1 A2 A3 0.106179f
C2 VPB A2 0.033537f
C3 VPWR B1 0.046731f
C4 A2 B2 4.92e-19
C5 VPB A3 0.033035f
C6 A1 A2 0.075092f
C7 VPWR X 0.102456f
C8 A3 B2 0.102249f
C9 VPB B2 0.033813f
C10 VPB A1 0.029013f
C11 A2 X 2.33e-19
C12 VPB B1 0.041119f
C13 A3 X 1.25e-19
C14 B2 B1 0.04397f
C15 VPB X 0.015707f
C16 VPWR VGND 0.072113f
C17 B2 X 7.64e-20
C18 A1 X 0.001481f
C19 VGND A2 0.016397f
C20 VGND A3 0.013109f
C21 VPB VGND 0.006316f
C22 VGND B2 0.010524f
C23 A1 VGND 0.019687f
C24 VPWR A2 0.013495f
C25 VGND B1 0.010652f
C26 VPWR A3 0.008806f
C27 VPB VPWR 0.083235f
C28 VGND X 0.103165f
C29 VPWR B2 0.012246f
C30 VGND VNB 0.437857f
C31 VPWR VNB 0.404492f
C32 X VNB 0.100953f
C33 B1 VNB 0.150231f
C34 B2 VNB 0.097709f
C35 A3 VNB 0.096505f
C36 A2 VNB 0.096218f
C37 A1 VNB 0.094556f
C38 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32a_2 VNB VPB VGND VPWR B1 B2 A3 A2 A1 X
X0 a_429_297.t1 A2.t0 a_345_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t3 A2.t1 a_345_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t3 a_79_21.t4 X.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t0 a_79_21.t5 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_345_47.t1 A3.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X5 a_345_297.t0 A1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297.t1 B2.t0 a_79_21.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t0 B1.t0 a_629_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21.t3 B2.t1 a_345_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_345_47.t0 B1.t1 a_79_21.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1235 ps=1.03 w=0.65 l=0.15
X10 a_79_21.t1 A3.t1 a_429_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X.t2 a_79_21.t6 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X.t0 a_79_21.t7 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47.t4 A1.t1 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
R0 A2.n0 A2.t0 241.536
R1 A2.n0 A2.t1 169.237
R2 A2 A2.n0 153.653
R3 a_345_297.t0 a_345_297.t1 53.1905
R4 a_429_297.t0 a_429_297.t1 84.7105
R5 VPB.t0 VPB.t3 449.844
R6 VPB.t6 VPB.t4 343.303
R7 VPB.t5 VPB.t2 313.707
R8 VPB.t4 VPB.t5 248.599
R9 VPB.t3 VPB.t6 248.599
R10 VPB.t1 VPB.t0 248.599
R11 VPB VPB.t1 189.409
R12 a_345_47.t0 a_345_47.n2 186.209
R13 a_345_47.n2 a_345_47.n0 154.05
R14 a_345_47.n2 a_345_47.n1 89.3175
R15 a_345_47.n1 a_345_47.t2 24.9236
R16 a_345_47.n1 a_345_47.t1 24.9236
R17 a_345_47.n0 a_345_47.t3 24.9236
R18 a_345_47.n0 a_345_47.t4 24.9236
R19 VGND.n2 VGND.n1 205.26
R20 VGND.n6 VGND.t1 154.599
R21 VGND.n4 VGND.n3 110.424
R22 VGND.n3 VGND.t4 58.1543
R23 VGND.n3 VGND.t0 54.462
R24 VGND.n1 VGND.t2 39.6928
R25 VGND.n1 VGND.t3 39.6928
R26 VGND.n5 VGND.n4 30.4946
R27 VGND.n6 VGND.n5 25.977
R28 VGND.n7 VGND.n6 9.3005
R29 VGND.n5 VGND.n0 9.3005
R30 VGND.n4 VGND.n2 6.3043
R31 VGND.n2 VGND.n0 0.320723
R32 VGND.n7 VGND.n0 0.120292
R33 VGND VGND.n7 0.0213333
R34 VNB.t1 VNB.t6 2164.4
R35 VNB.t5 VNB.t3 1651.78
R36 VNB.t4 VNB.t0 1509.39
R37 VNB.t3 VNB.t4 1196.12
R38 VNB.t6 VNB.t5 1196.12
R39 VNB.t2 VNB.t1 1196.12
R40 VNB VNB.t2 911.327
R41 a_79_21.n3 a_79_21.n1 315.142
R42 a_79_21.n4 a_79_21.n3 300.805
R43 a_79_21.n3 a_79_21.n2 278.541
R44 a_79_21.n1 a_79_21.t4 212.081
R45 a_79_21.n0 a_79_21.t6 212.081
R46 a_79_21.n1 a_79_21.t5 139.78
R47 a_79_21.n0 a_79_21.t7 139.78
R48 a_79_21.n1 a_79_21.n0 61.346
R49 a_79_21.n2 a_79_21.t3 39.6928
R50 a_79_21.n2 a_79_21.t0 30.462
R51 a_79_21.n4 a_79_21.t2 26.5955
R52 a_79_21.t1 a_79_21.n4 26.5955
R53 X X.n0 593.34
R54 X.n4 X.n0 585
R55 X.n3 X.n0 585
R56 X.n1 X 186.745
R57 X.n2 X.n1 185
R58 X.n0 X.t3 26.5955
R59 X.n0 X.t2 26.5955
R60 X.n1 X.t1 24.9236
R61 X.n1 X.t0 24.9236
R62 X.n2 X 11.4429
R63 X.n4 X 8.33989
R64 X.n3 X 8.33989
R65 X X.n4 4.84898
R66 X X.n3 4.84898
R67 X X.n2 1.74595
R68 VPWR.n7 VPWR.n6 585
R69 VPWR.n5 VPWR.n4 585
R70 VPWR.n9 VPWR.t2 249.362
R71 VPWR.n3 VPWR.t0 249.056
R72 VPWR.n6 VPWR.n5 66.9805
R73 VPWR.n5 VPWR.t1 26.5955
R74 VPWR.n6 VPWR.t3 26.5955
R75 VPWR.n8 VPWR.n7 26.0711
R76 VPWR.n9 VPWR.n8 25.977
R77 VPWR.n4 VPWR.n3 15.5986
R78 VPWR.n2 VPWR.n1 9.3005
R79 VPWR.n8 VPWR.n0 9.3005
R80 VPWR.n10 VPWR.n9 9.3005
R81 VPWR.n4 VPWR.n1 5.45932
R82 VPWR.n7 VPWR.n1 0.941676
R83 VPWR.n3 VPWR.n2 0.149666
R84 VPWR.n2 VPWR.n0 0.120292
R85 VPWR.n10 VPWR.n0 0.120292
R86 VPWR VPWR.n10 0.0213333
R87 A3.n0 A3.t1 237.736
R88 A3.n0 A3.t0 165.435
R89 A3 A3.n0 154.065
R90 A1.n0 A1.t0 240.484
R91 A1.n0 A1.t1 168.185
R92 A1 A1.n0 155.201
R93 B2.n0 B2.t0 241.536
R94 B2.n0 B2.t1 169.237
R95 B2 B2.n0 155.304
R96 a_629_297.t0 a_629_297.t1 74.8605
R97 B1.n0 B1.t0 232.212
R98 B1.n0 B1.t1 159.911
R99 B1 B1.n0 153.536
C0 B1 VPWR 0.060063f
C1 VGND VPB 0.007592f
C2 VGND A1 0.021511f
C3 VGND A2 0.011828f
C4 VPB A1 0.031149f
C5 VPB A2 0.028871f
C6 X VGND 0.140264f
C7 VGND A3 0.014884f
C8 X VPB 0.004427f
C9 A1 A2 0.096219f
C10 VPB A3 0.031318f
C11 VGND B2 0.008947f
C12 X A1 9.65e-19
C13 VPB B2 0.028285f
C14 X A2 5.03e-19
C15 A2 A3 0.086246f
C16 VGND B1 0.011469f
C17 VPB B1 0.043332f
C18 X A3 2.29e-19
C19 VGND VPWR 0.0996f
C20 VPB VPWR 0.098316f
C21 X B2 8.55e-20
C22 A3 B2 0.09813f
C23 A1 VPWR 0.014586f
C24 A2 VPWR 0.00904f
C25 X VPWR 0.16003f
C26 B2 B1 0.038848f
C27 A3 VPWR 0.011162f
C28 B2 VPWR 0.011762f
C29 VGND VNB 0.511332f
C30 X VNB 0.025586f
C31 VPWR VNB 0.478925f
C32 B1 VNB 0.150793f
C33 B2 VNB 0.091004f
C34 A3 VNB 0.094014f
C35 A2 VNB 0.089842f
C36 A1 VNB 0.092057f
C37 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32a_4 VNB VPB VGND VPWR A2 A3 B2 X A1 B1
X0 a_27_47.t2 B2.t0 a_549_297.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_297.t2 A2.t0 a_277_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_297.t0 A2.t1 a_27_297.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_549_297.t3 B2.t1 a_739_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47.t4 A3.t0 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297.t0 A1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_739_297.t1 B2.t2 a_549_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X7 a_739_297.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47.t7 A1.t1 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47.t6 A2.t2 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_549_297.t0 B2.t3 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X11 a_277_297.t2 A3.t1 a_549_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR.t3 B1.t1 a_739_297.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_27_47.t5 B1.t2 a_549_297.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_549_297.t5 A3.t2 a_277_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t5 A3.t3 a_27_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X16 VGND.t1 A2.t3 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_549_297.t7 B1.t3 a_27_47.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t2 A1.t2 a_27_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND.t0 A1.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B2.n0 B2.t2 221.72
R1 B2.n1 B2.t1 221.72
R2 B2 B2.n2 171.52
R3 B2.n0 B2.t3 149.421
R4 B2.n1 B2.t0 149.421
R5 B2.n2 B2.n0 40.1672
R6 B2.n2 B2.n1 40.1672
R7 a_549_297.n1 a_549_297.n0 717.558
R8 a_549_297.n24 a_549_297.n23 694.245
R9 a_549_297.n20 a_549_297.t0 258.846
R10 a_549_297.n1 a_549_297.t6 258.846
R11 a_549_297.n12 a_549_297.n10 221.72
R12 a_549_297.n9 a_549_297.n7 221.72
R13 a_549_297.n16 a_549_297.n5 221.72
R14 a_549_297.n18 a_549_297.n3 221.72
R15 a_549_297.n19 a_549_297.n18 188.596
R16 a_549_297.n22 a_549_297.n21 185
R17 a_549_297.n14 a_549_297.n13 183.625
R18 a_549_297.n17 a_549_297.n2 152
R19 a_549_297.n15 a_549_297.n14 152
R20 a_549_297.n12 a_549_297.n11 149.421
R21 a_549_297.n9 a_549_297.n8 149.421
R22 a_549_297.n16 a_549_297.n6 149.421
R23 a_549_297.n18 a_549_297.n4 149.421
R24 a_549_297.n22 a_549_297.n20 64.7534
R25 a_549_297.n23 a_549_297.n1 43.6711
R26 a_549_297.n20 a_549_297.n19 41.4519
R27 a_549_297.n13 a_549_297.n12 37.4894
R28 a_549_297.n13 a_549_297.n9 37.4894
R29 a_549_297.n15 a_549_297.n9 37.4894
R30 a_549_297.n16 a_549_297.n15 37.4894
R31 a_549_297.n17 a_549_297.n16 37.4894
R32 a_549_297.n18 a_549_297.n17 37.4894
R33 a_549_297.n24 a_549_297.t3 32.5055
R34 a_549_297.n14 a_549_297.n2 31.624
R35 a_549_297.n19 a_549_297.n2 30.6135
R36 a_549_297.n0 a_549_297.t4 26.5955
R37 a_549_297.n0 a_549_297.t5 26.5955
R38 a_549_297.t2 a_549_297.n24 26.5955
R39 a_549_297.n21 a_549_297.t1 24.9236
R40 a_549_297.n21 a_549_297.t7 24.9236
R41 a_549_297.n23 a_549_297.n22 3.01226
R42 a_27_47.n1 a_27_47.t0 261.134
R43 a_27_47.n7 a_27_47.n6 238.03
R44 a_27_47.n4 a_27_47.t4 209.923
R45 a_27_47.n3 a_27_47.n2 185
R46 a_27_47.n1 a_27_47.n0 185
R47 a_27_47.n6 a_27_47.n5 185
R48 a_27_47.n6 a_27_47.n4 85.1388
R49 a_27_47.n4 a_27_47.n3 51.7125
R50 a_27_47.n3 a_27_47.n1 44.0325
R51 a_27_47.t2 a_27_47.n7 30.462
R52 a_27_47.n2 a_27_47.t6 28.6159
R53 a_27_47.n5 a_27_47.t8 24.9236
R54 a_27_47.n5 a_27_47.t5 24.9236
R55 a_27_47.n0 a_27_47.t3 24.9236
R56 a_27_47.n0 a_27_47.t7 24.9236
R57 a_27_47.n2 a_27_47.t9 24.9236
R58 a_27_47.n7 a_27_47.t1 24.9236
R59 VNB.t4 VNB.t5 4100.97
R60 VNB.t2 VNB.t1 1281.55
R61 VNB.t6 VNB.t9 1253.07
R62 VNB.t8 VNB.t2 1196.12
R63 VNB.t5 VNB.t8 1196.12
R64 VNB.t9 VNB.t4 1196.12
R65 VNB.t3 VNB.t6 1196.12
R66 VNB.t7 VNB.t3 1196.12
R67 VNB.t0 VNB.t7 1196.12
R68 VNB VNB.t0 911.327
R69 VGND.n4 VGND.n3 189.856
R70 VGND.n2 VGND.n1 185
R71 VGND.n9 VGND.n8 185
R72 VGND.n10 VGND.n9 34.5993
R73 VGND.n8 VGND.t4 24.9236
R74 VGND.n8 VGND.t0 24.9236
R75 VGND.n1 VGND.t3 24.9236
R76 VGND.n1 VGND.t1 24.9236
R77 VGND.n3 VGND.t2 24.9236
R78 VGND.n3 VGND.t5 24.9236
R79 VGND.n7 VGND.n6 10.706
R80 VGND.n7 VGND.n0 9.3005
R81 VGND.n6 VGND.n5 9.3005
R82 VGND.n6 VGND.n2 8.61141
R83 VGND.n4 VGND.n2 6.73577
R84 VGND.n5 VGND.n4 1.49284
R85 VGND.n9 VGND.n7 0.233227
R86 VGND.n5 VGND.n0 0.120292
R87 VGND.n10 VGND.n0 0.120292
R88 VGND VGND.n10 0.0213333
R89 VPWR.n2 VPWR.n0 623.186
R90 VPWR.n2 VPWR.n1 327.955
R91 VPWR.n1 VPWR.t1 26.5955
R92 VPWR.n1 VPWR.t2 26.5955
R93 VPWR.n0 VPWR.t0 26.5955
R94 VPWR.n0 VPWR.t3 26.5955
R95 VPWR VPWR.n2 0.144411
R96 VPB.t5 VPB.t9 556.386
R97 VPB.t2 VPB.t6 556.386
R98 VPB.t4 VPB.t3 266.356
R99 VPB.t0 VPB.t4 248.599
R100 VPB.t9 VPB.t0 248.599
R101 VPB.t6 VPB.t5 248.599
R102 VPB.t8 VPB.t2 248.599
R103 VPB.t1 VPB.t8 248.599
R104 VPB.t7 VPB.t1 248.599
R105 VPB VPB.t7 189.409
R106 A2.n0 A2.t0 221.72
R107 A2.n1 A2.t1 221.72
R108 A2 A2.n2 152.321
R109 A2.n0 A2.t2 149.421
R110 A2.n1 A2.t3 149.421
R111 A2.n2 A2.n1 40.1672
R112 A2.n2 A2.n0 34.8116
R113 a_277_297.n1 a_277_297.n0 655.25
R114 a_277_297.n0 a_277_297.t2 283.173
R115 a_277_297.n0 a_277_297.t3 215.875
R116 a_277_297.n1 a_277_297.t1 26.5955
R117 a_277_297.t0 a_277_297.n1 26.5955
R118 a_27_297.t2 a_27_297.n1 376.757
R119 a_27_297.n1 a_27_297.t3 279.163
R120 a_27_297.n1 a_27_297.n0 189.28
R121 a_27_297.n0 a_27_297.t1 26.5955
R122 a_27_297.n0 a_27_297.t0 26.5955
R123 a_739_297.n1 a_739_297.n0 289.24
R124 a_739_297.n0 a_739_297.t1 276.409
R125 a_739_297.n0 a_739_297.t3 276.147
R126 a_739_297.t2 a_739_297.n1 26.5955
R127 a_739_297.n1 a_739_297.t0 26.5955
R128 A3.n0 A3.t1 296.699
R129 A3.n0 A3.t2 221.72
R130 A3 A3.n2 168
R131 A3.n2 A3.t3 165.488
R132 A3.n1 A3.t0 149.421
R133 A3.n2 A3.n1 58.9116
R134 A3.n1 A3.n0 14.282
R135 A1.n0 A1.t0 221.72
R136 A1.n1 A1.t2 221.72
R137 A1.n2 A1.n1 152.893
R138 A1.n0 A1.t1 149.421
R139 A1.n1 A1.t3 149.421
R140 A1.n1 A1.n0 74.9783
R141 A1 A1.n2 20.1605
R142 A1.n2 A1 9.2805
R143 B1.n0 B1.t0 221.72
R144 B1.n1 B1.t1 221.72
R145 B1 B1.n2 164.481
R146 B1.n0 B1.t3 149.421
R147 B1.n1 B1.t2 149.421
R148 B1.n2 B1.n0 68.7301
R149 B1.n2 B1.n1 6.24865
C0 VPB VGND 0.01783f
C1 A1 VGND 0.030583f
C2 A2 VGND 0.027956f
C3 B1 B2 0.050987f
C4 VPB VPWR 0.186784f
C5 A1 VPWR 0.031822f
C6 A3 VGND 0.03069f
C7 A2 VPWR 0.016547f
C8 B2 X 2.55e-19
C9 B1 VGND 0.015494f
C10 A3 VPWR 0.018179f
C11 B2 VGND 0.016391f
C12 B1 VPWR 0.025064f
C13 X VGND 0.301753f
C14 VPB A1 0.068761f
C15 B2 VPWR 0.015723f
C16 VPB A2 0.057294f
C17 A1 A2 0.065715f
C18 VPWR X 0.378772f
C19 VPB A3 0.085515f
C20 VPWR VGND 0.160905f
C21 VPB B1 0.0592f
C22 A2 A3 0.049084f
C23 VPB B2 0.0593f
C24 VPB X 0.022773f
C25 A3 B1 0.015771f
C26 VGND VNB 0.923963f
C27 X VNB 0.066502f
C28 VPWR VNB 0.786602f
C29 B2 VNB 0.18112f
C30 B1 VNB 0.186113f
C31 A3 VNB 0.22961f
C32 A2 VNB 0.171836f
C33 A1 VNB 0.232509f
C34 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32ai_1 VPB VNB VGND VPWR A1 A2 B1 Y B2 A3
X0 VGND.t2 A3.t0 a_27_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.219375 pd=1.325 as=0.10075 ps=0.96 w=0.65 l=0.15
X1 a_27_47.t3 A2.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.219375 ps=1.325 w=0.65 l=0.15
X2 Y.t1 B2.t0 a_109_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.105 ps=1.21 w=1 l=0.15
X3 a_333_297.t1 A3.t1 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.49 as=0.305 ps=1.61 w=1 l=0.15
X4 VGND.t0 A1.t0 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47.t0 B2.t1 Y.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.105625 ps=0.975 w=0.65 l=0.15
X6 VPWR.t0 A1.t1 a_461_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_297.t1 B1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8 a_461_297.t0 A2.t1 a_333_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.49 w=1 l=0.15
X9 Y.t0 B1.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A3.n0 A3.t1 235.821
R1 A3.n0 A3.t0 215.421
R2 A3 A3.n0 154.429
R3 a_27_47.n1 a_27_47.t1 316.851
R4 a_27_47.n1 a_27_47.n0 283.25
R5 a_27_47.n2 a_27_47.n1 89.3175
R6 a_27_47.t0 a_27_47.n2 29.539
R7 a_27_47.n2 a_27_47.t4 27.6928
R8 a_27_47.n0 a_27_47.t2 24.9236
R9 a_27_47.n0 a_27_47.t3 24.9236
R10 VGND.n3 VGND.n2 185
R11 VGND.n1 VGND.n0 185
R12 VGND.n4 VGND.t0 140.243
R13 VGND.n2 VGND.n1 62.7697
R14 VGND.n1 VGND.t2 36.9236
R15 VGND.n2 VGND.t1 24.9236
R16 VGND.n5 VGND.n0 8.99046
R17 VGND.n4 VGND.n3 7.86735
R18 VGND.n3 VGND.n0 7.63559
R19 VGND.n5 VGND.n4 0.763298
R20 VGND VGND.n5 0.353068
R21 VNB.t4 VNB.t3 2349.51
R22 VNB.t1 VNB.t0 1352.75
R23 VNB.t0 VNB.t4 1310.03
R24 VNB.t3 VNB.t2 1196.12
R25 VNB VNB.t1 911.327
R26 A2.n0 A2.t1 236.18
R27 A2.n0 A2.t0 163.881
R28 A2.n1 A2.n0 152
R29 A2.n1 A2 12.3666
R30 A2 A2.n1 2.38694
R31 B2.n0 B2.t0 233.869
R32 B2.n0 B2.t1 162.549
R33 B2 B2.n0 154.375
R34 a_109_297.t0 a_109_297.t1 41.3705
R35 Y.n2 Y.n0 260.579
R36 Y Y.n1 148.886
R37 Y.n1 Y.t3 60.0855
R38 Y.n1 Y.t1 60.0855
R39 Y.n0 Y.t2 35.0774
R40 Y.n0 Y.t0 24.9236
R41 Y.n2 Y 8.56521
R42 Y Y.n2 0.0946176
R43 VPB.t1 VPB.t3 449.844
R44 VPB.t3 VPB.t0 378.817
R45 VPB.t0 VPB.t4 248.599
R46 VPB.t2 VPB.t1 213.084
R47 VPB VPB.t2 189.409
R48 a_333_297.t0 a_333_297.t1 96.5305
R49 A1.n0 A1.t1 236.18
R50 A1.n0 A1.t0 163.881
R51 A1 A1.n0 158.595
R52 a_461_297.t0 a_461_297.t1 53.1905
R53 VPWR.n0 VPWR.t1 255.544
R54 VPWR.n0 VPWR.t0 245.023
R55 VPWR VPWR.n0 0.0550601
R56 B1.n0 B1.t0 230.363
R57 B1.n0 B1.t1 158.064
R58 B1 B1.n0 154.607
C0 VPB A2 0.035981f
C1 VPB B1 0.036383f
C2 VPB VGND 0.00559f
C3 VPB A1 0.034198f
C4 VGND A2 0.020709f
C5 VPB B2 0.035039f
C6 A2 A1 0.074868f
C7 B1 VGND 0.012893f
C8 VPB VPWR 0.086152f
C9 B2 A2 3e-19
C10 VGND A1 0.063864f
C11 B1 B2 0.058292f
C12 A2 VPWR 0.094677f
C13 VPB A3 0.037151f
C14 B2 VGND 0.01122f
C15 B1 VPWR 0.050169f
C16 VPB Y 0.005999f
C17 A3 A2 0.081117f
C18 VGND VPWR 0.066422f
C19 A2 Y 0.038364f
C20 A1 VPWR 0.064733f
C21 B2 VPWR 0.009831f
C22 B1 Y 0.073988f
C23 VGND A3 0.01787f
C24 VGND Y 0.011045f
C25 A1 Y 1.1e-19
C26 B2 A3 0.099991f
C27 B2 Y 0.115881f
C28 A3 VPWR 0.013001f
C29 VPWR Y 0.215002f
C30 A3 Y 0.023748f
C31 VGND VNB 0.40808f
C32 Y VNB 0.016066f
C33 VPWR VNB 0.400137f
C34 A1 VNB 0.138892f
C35 A2 VNB 0.105715f
C36 A3 VNB 0.100696f
C37 B2 VNB 0.098855f
C38 B1 VNB 0.159818f
C39 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32ai_2 VPB VNB VGND VPWR A1 A2 Y B1 B2 A3
X0 VGND.t5 A1.t0 a_27_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_27_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X2 a_475_297.t3 A2.t0 a_729_297.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_729_297.t1 A1.t1 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR.t1 A1.t2 a_729_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47.t5 A2.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_297.t3 B1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_729_297.t2 A2.t2 a_475_297.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t3 B1.t1 a_27_297.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t2 A2.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297.t0 B2.t0 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47.t3 B2.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_47.t8 B1.t2 Y.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_475_297.t1 A3.t1 Y.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t4 A3.t2 a_475_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y.t6 B1.t3 a_27_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47.t6 A1.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t1 A3.t3 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t0 B2.t2 a_27_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y.t2 B2.t3 a_27_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t2 223.766
R1 A1.n1 A1.t1 212.081
R2 A1.n3 A1.n2 152
R3 A1.n1 A1.t0 151.465
R4 A1.n0 A1.t3 139.78
R5 A1.n2 A1.n0 29.2126
R6 A1.n2 A1.n1 20.449
R7 A1 A1.n3 17.4085
R8 A1.n3 A1 6.1445
R9 a_27_47.n4 a_27_47.t6 190.526
R10 a_27_47.n3 a_27_47.n2 185
R11 a_27_47.n1 a_27_47.n0 185
R12 a_27_47.n1 a_27_47.t9 180.929
R13 a_27_47.n9 a_27_47.n8 98.5806
R14 a_27_47.n8 a_27_47.n3 93.3712
R15 a_27_47.n7 a_27_47.n6 92.5005
R16 a_27_47.n5 a_27_47.n4 92.5005
R17 a_27_47.n6 a_27_47.n5 62.7697
R18 a_27_47.n3 a_27_47.n1 46.7483
R19 a_27_47.n5 a_27_47.t7 43.3851
R20 a_27_47.n8 a_27_47.n7 42.9971
R21 a_27_47.n6 a_27_47.t5 39.6928
R22 a_27_47.n0 a_27_47.t4 24.9236
R23 a_27_47.n0 a_27_47.t3 24.9236
R24 a_27_47.n2 a_27_47.t1 24.9236
R25 a_27_47.n2 a_27_47.t8 24.9236
R26 a_27_47.n9 a_27_47.t2 24.9236
R27 a_27_47.t0 a_27_47.n9 24.9236
R28 a_27_47.n7 a_27_47.n4 6.69588
R29 VGND.n6 VGND.n3 207.213
R30 VGND.n5 VGND.n4 206.079
R31 VGND.n1 VGND.n0 199.739
R32 VGND.n0 VGND.t1 103.385
R33 VGND.n0 VGND.t0 42.462
R34 VGND.n8 VGND.n7 34.6358
R35 VGND.n4 VGND.t4 24.9236
R36 VGND.n4 VGND.t5 24.9236
R37 VGND.n3 VGND.t3 24.9236
R38 VGND.n3 VGND.t2 24.9236
R39 VGND.n6 VGND.n5 21.7681
R40 VGND.n7 VGND.n6 20.3299
R41 VGND.n10 VGND.n1 14.3776
R42 VGND.n7 VGND.n2 9.3005
R43 VGND.n9 VGND.n8 9.3005
R44 VGND.n8 VGND.n1 3.01226
R45 VGND VGND.n10 0.597808
R46 VGND.n5 VGND.n2 0.284459
R47 VGND.n10 VGND.n9 0.147181
R48 VGND.n9 VGND.n2 0.120292
R49 VNB.t5 VNB.t7 2677.02
R50 VNB.t1 VNB.t0 2677.02
R51 VNB.t7 VNB.t6 1196.12
R52 VNB.t2 VNB.t5 1196.12
R53 VNB.t0 VNB.t2 1196.12
R54 VNB.t8 VNB.t1 1196.12
R55 VNB.t4 VNB.t8 1196.12
R56 VNB.t3 VNB.t4 1196.12
R57 VNB.t9 VNB.t3 1196.12
R58 VNB VNB.t9 925.567
R59 A3.n1 A3.t3 351.568
R60 A3.n0 A3.t1 220.845
R61 A3.n1 A3.t2 212.081
R62 A3 A3.n2 175.041
R63 A3.n0 A3.t0 139.78
R64 A3.n2 A3.n0 27.752
R65 A3.n2 A3.n1 24.8308
R66 A2.n0 A2.t0 220.845
R67 A2.n1 A2.t2 212.081
R68 A2.n3 A2.n2 152
R69 A2.n1 A2.t3 148.544
R70 A2.n0 A2.t1 139.78
R71 A2.n3 A2 28.1605
R72 A2.n2 A2.n0 27.752
R73 A2.n2 A2.n1 24.8308
R74 A2 A2.n3 18.9445
R75 a_729_297.n1 a_729_297.n0 583.202
R76 a_729_297.n0 a_729_297.t3 26.5955
R77 a_729_297.n0 a_729_297.t2 26.5955
R78 a_729_297.t0 a_729_297.n1 26.5955
R79 a_729_297.n1 a_729_297.t1 26.5955
R80 a_475_297.n0 a_475_297.t3 380.048
R81 a_475_297.n0 a_475_297.t0 380.046
R82 a_475_297.n1 a_475_297.n0 206
R83 a_475_297.t2 a_475_297.n1 26.5955
R84 a_475_297.n1 a_475_297.t1 26.5955
R85 VPB.t1 VPB.t3 591.9
R86 VPB.t9 VPB.t6 568.225
R87 VPB.t6 VPB.t5 248.599
R88 VPB.t8 VPB.t9 248.599
R89 VPB.t4 VPB.t8 248.599
R90 VPB.t3 VPB.t4 248.599
R91 VPB.t7 VPB.t1 248.599
R92 VPB.t0 VPB.t7 248.599
R93 VPB.t2 VPB.t0 248.599
R94 VPB VPB.t2 192.369
R95 VPWR.n1 VPWR.n0 607.212
R96 VPWR.n5 VPWR.t2 348.036
R97 VPWR.n6 VPWR.t1 265.752
R98 VPWR.n18 VPWR.n1 35.4627
R99 VPWR.n9 VPWR.n8 34.6358
R100 VPWR.n10 VPWR.n9 34.6358
R101 VPWR.n10 VPWR.n3 34.6358
R102 VPWR.n14 VPWR.n3 34.6358
R103 VPWR.n15 VPWR.n14 34.6358
R104 VPWR.n16 VPWR.n15 34.6358
R105 VPWR.n0 VPWR.t0 26.5955
R106 VPWR.n0 VPWR.t3 26.5955
R107 VPWR.n8 VPWR.n5 18.824
R108 VPWR.n8 VPWR.n7 9.3005
R109 VPWR.n9 VPWR.n4 9.3005
R110 VPWR.n11 VPWR.n10 9.3005
R111 VPWR.n12 VPWR.n3 9.3005
R112 VPWR.n14 VPWR.n13 9.3005
R113 VPWR.n15 VPWR.n2 9.3005
R114 VPWR.n17 VPWR.n16 9.3005
R115 VPWR.n6 VPWR.n5 7.4042
R116 VPWR.n16 VPWR.n1 6.77697
R117 VPWR.n7 VPWR.n6 0.698357
R118 VPWR VPWR.n18 0.237687
R119 VPWR.n18 VPWR.n17 0.146169
R120 VPWR.n7 VPWR.n4 0.120292
R121 VPWR.n11 VPWR.n4 0.120292
R122 VPWR.n12 VPWR.n11 0.120292
R123 VPWR.n13 VPWR.n12 0.120292
R124 VPWR.n13 VPWR.n2 0.120292
R125 VPWR.n17 VPWR.n2 0.120292
R126 B1.n0 B1.t0 212.081
R127 B1.n1 B1.t1 212.081
R128 B1.n3 B1.n2 152
R129 B1.n0 B1.t2 139.78
R130 B1.n1 B1.t3 139.78
R131 B1.n2 B1.n0 30.6732
R132 B1.n2 B1.n1 30.6732
R133 B1.n3 B1 23.0405
R134 B1 B1.n3 0.5125
R135 a_27_297.n0 a_27_297.t3 376.531
R136 a_27_297.n0 a_27_297.t1 293.906
R137 a_27_297.n1 a_27_297.n0 288.212
R138 a_27_297.t2 a_27_297.n1 26.5955
R139 a_27_297.n1 a_27_297.t0 26.5955
R140 B2.n0 B2.t0 212.081
R141 B2.n1 B2.t2 212.081
R142 B2 B2.n2 155.584
R143 B2.n0 B2.t1 139.78
R144 B2.n1 B2.t3 139.78
R145 B2.n2 B2.n0 30.6732
R146 B2.n2 B2.n1 30.6732
R147 Y.n5 Y.n3 376.418
R148 Y.n5 Y.n4 344.416
R149 Y.n2 Y.n0 228.008
R150 Y.n2 Y.n1 185
R151 Y Y.n2 37.5873
R152 Y.n4 Y.t5 26.5955
R153 Y.n4 Y.t4 26.5955
R154 Y.n3 Y.t1 26.5955
R155 Y.n3 Y.t0 26.5955
R156 Y.n0 Y.t3 24.9236
R157 Y.n0 Y.t2 24.9236
R158 Y.n1 Y.t7 24.9236
R159 Y.n1 Y.t6 24.9236
R160 Y Y.n5 5.85813
C0 VPB B2 0.056675f
C1 VPB B1 0.058139f
C2 Y VPB 0.02167f
C3 B2 B1 0.074816f
C4 VPB A3 0.082884f
C5 Y B2 0.0949f
C6 VPWR VPB 0.140615f
C7 VPB A2 0.06195f
C8 VGND VPB 0.014058f
C9 VPWR B2 0.017581f
C10 Y B1 0.178547f
C11 A1 VPB 0.070658f
C12 B1 A3 0.03697f
C13 Y A3 0.113372f
C14 VPWR B1 0.025372f
C15 VGND B2 0.017667f
C16 Y VPWR 0.034088f
C17 VPWR A3 0.019636f
C18 VGND B1 0.016258f
C19 Y A2 7.69e-19
C20 Y VGND 0.02392f
C21 A3 A2 0.073419f
C22 VGND A3 0.028466f
C23 VPWR A2 0.018072f
C24 A1 Y 2.43e-19
C25 VPWR VGND 0.114927f
C26 A1 VPWR 0.06146f
C27 VGND A2 0.026246f
C28 A1 A2 0.035119f
C29 A1 VGND 0.032589f
C30 VGND VNB 0.665395f
C31 VPWR VNB 0.590596f
C32 Y VNB 0.023974f
C33 A1 VNB 0.229592f
C34 A2 VNB 0.189182f
C35 A3 VNB 0.235143f
C36 B1 VNB 0.171173f
C37 B2 VNB 0.208909f
C38 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32ai_4 VNB VPB VGND VPWR B2 Y B1 A3 A2 A1
X0 a_1224_297# A1.t0 VPWR.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1825 ps=1.365 w=1 l=0.15
X2 a_27_297.t7 B1.t0 VPWR.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47.t9 A1.t1 VGND.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t1 B2.t0 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t6 B1.t1 a_27_297.t6 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_806_297.t3 A3.t0 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t9 A2.t0 a_27_47.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.20475 ps=1.28 w=0.65 l=0.15
X8 VGND.t10 A2.t1 a_27_47.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47.t3 A3.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.28 as=0.13975 ps=1.08 w=0.65 l=0.15
X10 Y.t3 B2.t1 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_806_297.t2 A3.t2 Y.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y.t10 A3.t3 a_806_297.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47.t18 B1.t2 Y.t15 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_27_297.t2 B2.t2 Y.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47.t6 B2.t3 Y.t8 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47.t12 B2.t4 Y.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_27_47.t17 B1.t3 Y.t14 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t11 A3.t4 a_806_297.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47.t4 A2.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_27_47.t5 A2.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_27_297.t5 B1.t4 VPWR.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 Y.t13 B1.t5 a_27_47.t16 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X23 a_806_297.t6 A2.t4 a_1224_297# VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 Y.t6 B2.t5 a_27_47.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 Y.t12 B1.t6 a_27_47.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t0 B1.t7 a_27_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X27 VGND.t0 A3.t5 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VGND.t1 A3.t6 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_1224_297# A2.t5 a_806_297.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_1224_297# A1.t2 VPWR.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X31 a_806_297.t4 A2.t6 a_1224_297# VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR.t3 A1.t3 a_1224_297# VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 Y.t1 B2.t6 a_27_297.t3 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_27_47.t2 A3.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 VGND.t7 A1.t4 a_27_47.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X36 a_1224_297# A2.t7 a_806_297.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 Y.t5 B2.t7 a_27_47.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 VGND.t6 A1.t5 a_27_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A1.n11 A1.n0 218.507
R1 A1.n2 A1.t2 218.507
R2 A1.n6 A1.t3 218.507
R3 A1.n4 A1.t0 218.507
R4 A1.n12 A1.n11 171.114
R5 A1.n10 A1.n9 152
R6 A1.n8 A1.n7 152
R7 A1.n5 A1.n3 152
R8 A1.n11 A1.n1 146.208
R9 A1.n2 A1.t5 146.208
R10 A1.n6 A1.t1 146.208
R11 A1.n4 A1.t4 146.208
R12 A1.n11 A1.n10 50.6936
R13 A1.n10 A1.n2 34.904
R14 A1.n7 A1.n2 34.904
R15 A1.n7 A1.n6 34.904
R16 A1.n6 A1.n5 34.904
R17 A1.n5 A1.n4 34.904
R18 A1.n8 A1.n3 26.8805
R19 A1.n9 A1 24.6405
R20 A1.n12 A1 22.0805
R21 A1 A1.n12 7.3605
R22 A1.n9 A1 4.8005
R23 A1 A1.n8 2.2405
R24 A1.n3 A1 0.3205
R25 VPWR.n28 VPWR.n1 599.74
R26 VPWR.n26 VPWR.n2 599.74
R27 VPWR.n8 VPWR.t5 342.841
R28 VPWR.n10 VPWR.n9 330.957
R29 VPWR.n13 VPWR.n7 34.6358
R30 VPWR.n14 VPWR.n13 34.6358
R31 VPWR.n15 VPWR.n14 34.6358
R32 VPWR.n15 VPWR.n5 34.6358
R33 VPWR.n19 VPWR.n5 34.6358
R34 VPWR.n20 VPWR.n19 34.6358
R35 VPWR.n21 VPWR.n20 34.6358
R36 VPWR.n21 VPWR.n3 34.6358
R37 VPWR.n25 VPWR.n3 34.6358
R38 VPWR.n28 VPWR.n27 33.8829
R39 VPWR.n1 VPWR.t2 26.5955
R40 VPWR.n1 VPWR.t0 26.5955
R41 VPWR.n2 VPWR.t1 26.5955
R42 VPWR.n2 VPWR.t6 26.5955
R43 VPWR.n9 VPWR.t4 26.5955
R44 VPWR.n9 VPWR.t3 26.5955
R45 VPWR.n8 VPWR.n7 21.0829
R46 VPWR.n11 VPWR.n7 9.3005
R47 VPWR.n13 VPWR.n12 9.3005
R48 VPWR.n14 VPWR.n6 9.3005
R49 VPWR.n16 VPWR.n15 9.3005
R50 VPWR.n17 VPWR.n5 9.3005
R51 VPWR.n19 VPWR.n18 9.3005
R52 VPWR.n20 VPWR.n4 9.3005
R53 VPWR.n22 VPWR.n21 9.3005
R54 VPWR.n23 VPWR.n3 9.3005
R55 VPWR.n25 VPWR.n24 9.3005
R56 VPWR.n27 VPWR.n0 9.3005
R57 VPWR.n10 VPWR.n8 6.87683
R58 VPWR.n29 VPWR.n28 6.11656
R59 VPWR.n26 VPWR.n25 5.27109
R60 VPWR.n27 VPWR.n26 4.51815
R61 VPWR.n11 VPWR.n10 0.681391
R62 VPWR VPWR.n29 0.573095
R63 VPWR.n29 VPWR.n0 0.170228
R64 VPWR.n12 VPWR.n11 0.120292
R65 VPWR.n12 VPWR.n6 0.120292
R66 VPWR.n16 VPWR.n6 0.120292
R67 VPWR.n17 VPWR.n16 0.120292
R68 VPWR.n18 VPWR.n17 0.120292
R69 VPWR.n18 VPWR.n4 0.120292
R70 VPWR.n22 VPWR.n4 0.120292
R71 VPWR.n23 VPWR.n22 0.120292
R72 VPWR.n24 VPWR.n23 0.120292
R73 VPWR.n24 VPWR.n0 0.120292
R74 VPB.t7 VPB.t13 556.386
R75 VPB.t6 VPB.t16 556.386
R76 VPB.t4 VPB.t5 257.478
R77 VPB.t11 VPB.t12 248.599
R78 VPB.t13 VPB.t11 248.599
R79 VPB.t8 VPB.t7 248.599
R80 VPB.t2 VPB.t8 248.599
R81 VPB.t3 VPB.t2 248.599
R82 VPB.t1 VPB.t3 248.599
R83 VPB.t15 VPB.t1 248.599
R84 VPB.t14 VPB.t15 248.599
R85 VPB.t16 VPB.t14 248.599
R86 VPB.t17 VPB.t6 248.599
R87 VPB.t10 VPB.t17 248.599
R88 VPB.t5 VPB.t10 248.599
R89 VPB.t0 VPB.t4 248.599
R90 VPB.t9 VPB.t0 248.599
R91 VPB.t18 VPB.t9 248.599
R92 VPB VPB.t18 189.409
R93 B1.n0 B1.t0 218.507
R94 B1.n6 B1.t1 218.507
R95 B1.n1 B1.t4 218.507
R96 B1.n2 B1.t7 218.507
R97 B1 B1.n3 157.12
R98 B1.n8 B1.n7 152
R99 B1.n5 B1.n4 152
R100 B1.n0 B1.t3 146.208
R101 B1.n6 B1.t6 146.208
R102 B1.n1 B1.t2 146.208
R103 B1.n2 B1.t5 146.208
R104 B1.n6 B1.n5 35.735
R105 B1.n3 B1.n1 35.735
R106 B1.n7 B1.n0 34.904
R107 B1.n7 B1.n6 34.904
R108 B1.n5 B1.n1 34.0729
R109 B1.n3 B1.n2 34.0729
R110 B1.n4 B1 21.7605
R111 B1.n8 B1 19.5205
R112 B1 B1.n8 9.9205
R113 B1.n4 B1 7.6805
R114 a_27_297.n3 a_27_297.n2 585
R115 a_27_297.n4 a_27_297.t7 380.231
R116 a_27_297.n1 a_27_297.n0 297.224
R117 a_27_297.n5 a_27_297.n4 297.224
R118 a_27_297.n1 a_27_297.t3 277.849
R119 a_27_297.n4 a_27_297.n3 75.6711
R120 a_27_297.n3 a_27_297.n1 58.5148
R121 a_27_297.n2 a_27_297.t1 29.5505
R122 a_27_297.n2 a_27_297.t4 26.5955
R123 a_27_297.n0 a_27_297.t0 26.5955
R124 a_27_297.n0 a_27_297.t2 26.5955
R125 a_27_297.t6 a_27_297.n5 26.5955
R126 a_27_297.n5 a_27_297.t5 26.5955
R127 VGND.n8 VGND.t6 242.583
R128 VGND.n10 VGND.n9 207.213
R129 VGND.n16 VGND.n6 207.213
R130 VGND.n18 VGND.n5 207.213
R131 VGND.n1 VGND.n0 207.213
R132 VGND.n25 VGND.n24 199.739
R133 VGND.n24 VGND.t3 39.6928
R134 VGND.n24 VGND.t1 39.6928
R135 VGND.n11 VGND.n7 34.6358
R136 VGND.n15 VGND.n7 34.6358
R137 VGND.n19 VGND.n3 34.6358
R138 VGND.n23 VGND.n3 34.6358
R139 VGND.n26 VGND.n25 33.1299
R140 VGND.n17 VGND.n16 32.0005
R141 VGND.n18 VGND.n17 31.2476
R142 VGND.n11 VGND.n10 30.4946
R143 VGND.n9 VGND.t8 24.9236
R144 VGND.n9 VGND.t7 24.9236
R145 VGND.n6 VGND.t5 24.9236
R146 VGND.n6 VGND.t10 24.9236
R147 VGND.n5 VGND.t4 24.9236
R148 VGND.n5 VGND.t9 24.9236
R149 VGND.n0 VGND.t2 24.9236
R150 VGND.n0 VGND.t0 24.9236
R151 VGND.n26 VGND.n1 23.7181
R152 VGND.n28 VGND.n1 18.5188
R153 VGND.n10 VGND.n8 11.3474
R154 VGND.n25 VGND.n23 11.2946
R155 VGND.n27 VGND.n26 9.3005
R156 VGND.n25 VGND.n2 9.3005
R157 VGND.n12 VGND.n11 9.3005
R158 VGND.n13 VGND.n7 9.3005
R159 VGND.n15 VGND.n14 9.3005
R160 VGND.n17 VGND.n4 9.3005
R161 VGND.n20 VGND.n19 9.3005
R162 VGND.n21 VGND.n3 9.3005
R163 VGND.n23 VGND.n22 9.3005
R164 VGND.n19 VGND.n18 3.38874
R165 VGND.n16 VGND.n15 2.63579
R166 VGND VGND.n28 0.957626
R167 VGND.n12 VGND.n8 0.51599
R168 VGND.n28 VGND.n27 0.147187
R169 VGND.n13 VGND.n12 0.120292
R170 VGND.n14 VGND.n13 0.120292
R171 VGND.n14 VGND.n4 0.120292
R172 VGND.n20 VGND.n4 0.120292
R173 VGND.n21 VGND.n20 0.120292
R174 VGND.n22 VGND.n21 0.120292
R175 VGND.n22 VGND.n2 0.120292
R176 VGND.n27 VGND.n2 0.120292
R177 a_27_47.n5 a_27_47.n4 185
R178 a_27_47.n3 a_27_47.n2 185
R179 a_27_47.n1 a_27_47.n0 185
R180 a_27_47.n1 a_27_47.t14 182.994
R181 a_27_47.n20 a_27_47.n19 152.665
R182 a_27_47.n9 a_27_47.n8 98.9685
R183 a_27_47.n15 a_27_47.n14 98.9685
R184 a_27_47.n11 a_27_47.n10 92.5005
R185 a_27_47.n13 a_27_47.n12 92.5005
R186 a_27_47.n17 a_27_47.n16 92.5005
R187 a_27_47.n19 a_27_47.n18 92.5005
R188 a_27_47.n7 a_27_47.n6 88.1117
R189 a_27_47.n18 a_27_47.n17 66.462
R190 a_27_47.n12 a_27_47.n11 62.7697
R191 a_27_47.n7 a_27_47.n5 55.8227
R192 a_27_47.n18 a_27_47.t8 54.462
R193 a_27_47.n10 a_27_47.n9 53.6968
R194 a_27_47.n5 a_27_47.n3 52.1148
R195 a_27_47.n9 a_27_47.n7 51.2757
R196 a_27_47.n3 a_27_47.n1 51.2005
R197 a_27_47.n15 a_27_47.n13 43.1556
R198 a_27_47.n16 a_27_47.n15 41.6497
R199 a_27_47.n12 a_27_47.t10 28.6159
R200 a_27_47.n2 a_27_47.t16 27.6928
R201 a_27_47.n17 a_27_47.t5 24.9236
R202 a_27_47.n11 a_27_47.t3 24.9236
R203 a_27_47.n6 a_27_47.t0 24.9236
R204 a_27_47.n6 a_27_47.t17 24.9236
R205 a_27_47.n0 a_27_47.t13 24.9236
R206 a_27_47.n0 a_27_47.t6 24.9236
R207 a_27_47.n2 a_27_47.t12 24.9236
R208 a_27_47.n4 a_27_47.t15 24.9236
R209 a_27_47.n4 a_27_47.t18 24.9236
R210 a_27_47.n8 a_27_47.t1 24.9236
R211 a_27_47.n8 a_27_47.t2 24.9236
R212 a_27_47.n14 a_27_47.t11 24.9236
R213 a_27_47.n14 a_27_47.t4 24.9236
R214 a_27_47.n20 a_27_47.t7 24.9236
R215 a_27_47.t9 a_27_47.n20 24.9236
R216 a_27_47.n19 a_27_47.n16 7.08973
R217 a_27_47.n13 a_27_47.n10 6.69588
R218 VNB.t5 VNB.t8 2677.02
R219 VNB.t3 VNB.t10 2221.36
R220 VNB.t1 VNB.t3 1651.78
R221 VNB.t12 VNB.t16 1238.83
R222 VNB.t9 VNB.t7 1196.12
R223 VNB.t8 VNB.t9 1196.12
R224 VNB.t11 VNB.t5 1196.12
R225 VNB.t4 VNB.t11 1196.12
R226 VNB.t10 VNB.t4 1196.12
R227 VNB.t2 VNB.t1 1196.12
R228 VNB.t0 VNB.t2 1196.12
R229 VNB.t17 VNB.t0 1196.12
R230 VNB.t15 VNB.t17 1196.12
R231 VNB.t18 VNB.t15 1196.12
R232 VNB.t16 VNB.t18 1196.12
R233 VNB.t13 VNB.t12 1196.12
R234 VNB.t6 VNB.t13 1196.12
R235 VNB.t14 VNB.t6 1196.12
R236 VNB VNB.t14 911.327
R237 B2.n1 B2.t0 218.507
R238 B2.n3 B2.t1 218.507
R239 B2.n0 B2.t2 218.507
R240 B2.n8 B2.t6 218.507
R241 B2.n9 B2.n8 184.411
R242 B2.n5 B2.n2 178.881
R243 B2.n5 B2.n4 152
R244 B2.n7 B2.n6 152
R245 B2.n1 B2.t4 146.208
R246 B2.n3 B2.t5 146.208
R247 B2.n0 B2.t3 146.208
R248 B2.n8 B2.t7 146.208
R249 B2.n2 B2.n1 34.904
R250 B2.n3 B2.n2 34.904
R251 B2.n4 B2.n3 34.904
R252 B2.n4 B2.n0 34.904
R253 B2.n7 B2.n0 34.904
R254 B2.n8 B2.n7 34.904
R255 B2.n6 B2 24.9605
R256 B2.n9 B2 21.4405
R257 B2 B2.n9 8.0005
R258 B2.n6 B2 4.4805
R259 B2 B2.n5 1.9205
R260 Y.n12 Y.n0 337.264
R261 Y.n3 Y.n1 337.264
R262 Y.n3 Y.n2 298.863
R263 Y.n14 Y.n13 293.327
R264 Y.n6 Y.n4 228.008
R265 Y.n9 Y.n7 228.008
R266 Y.n6 Y.n5 185
R267 Y.n9 Y.n8 185
R268 Y.n11 Y.n3 178.825
R269 Y.n11 Y.n10 48.0005
R270 Y.n13 Y.t4 26.5955
R271 Y.n13 Y.t3 26.5955
R272 Y.n1 Y.t0 26.5955
R273 Y.n1 Y.t10 26.5955
R274 Y.n2 Y.t9 26.5955
R275 Y.n2 Y.t11 26.5955
R276 Y.n0 Y.t2 26.5955
R277 Y.n0 Y.t1 26.5955
R278 Y.n7 Y.t8 24.9236
R279 Y.n7 Y.t5 24.9236
R280 Y.n8 Y.t7 24.9236
R281 Y.n8 Y.t6 24.9236
R282 Y.n5 Y.t15 24.9236
R283 Y.n5 Y.t13 24.9236
R284 Y.n4 Y.t14 24.9236
R285 Y.n4 Y.t12 24.9236
R286 Y.n10 Y.n6 22.0165
R287 Y.n10 Y.n9 21.7605
R288 Y.n12 Y.n11 11.6711
R289 Y.n14 Y.n12 5.26322
R290 Y Y.n14 2.32639
R291 A3.n2 A3.t0 278.341
R292 A3.n3 A3.t3 218.507
R293 A3.n5 A3.t2 218.507
R294 A3.n0 A3.t4 218.507
R295 A3.n12 A3.t5 161.166
R296 A3.n4 A3.n1 152
R297 A3.n8 A3.n7 152
R298 A3.n10 A3.n9 152
R299 A3.n13 A3.n12 152
R300 A3.n11 A3.t7 146.208
R301 A3.n6 A3.t6 146.208
R302 A3.n2 A3.t1 146.208
R303 A3.n5 A3.n4 68.1453
R304 A3.n12 A3.n11 54.8488
R305 A3.n6 A3.n0 53.1867
R306 A3.n8 A3.n1 26.8805
R307 A3.n9 A3 25.2805
R308 A3.n13 A3 22.7205
R309 A3.n7 A3.n6 14.9591
R310 A3.n11 A3.n10 14.9591
R311 A3.n3 A3.n2 9.97291
R312 A3 A3.n13 6.7205
R313 A3.n9 A3 4.1605
R314 A3.n4 A3.n3 1.66257
R315 A3.n7 A3.n5 1.66257
R316 A3.n10 A3.n0 1.66257
R317 A3 A3.n8 1.6005
R318 A3.n1 A3 0.9605
R319 a_806_297.n1 a_806_297.t6 370.428
R320 a_806_297.n3 a_806_297.t0 370.426
R321 a_806_297.n5 a_806_297.n4 297.224
R322 a_806_297.n3 a_806_297.n2 297.224
R323 a_806_297.n1 a_806_297.n0 297.224
R324 a_806_297.n4 a_806_297.n1 51.2005
R325 a_806_297.n4 a_806_297.n3 51.2005
R326 a_806_297.n2 a_806_297.t1 26.5955
R327 a_806_297.n2 a_806_297.t2 26.5955
R328 a_806_297.n0 a_806_297.t7 26.5955
R329 a_806_297.n0 a_806_297.t4 26.5955
R330 a_806_297.n5 a_806_297.t5 26.5955
R331 a_806_297.t3 a_806_297.n5 26.5955
R332 A2.n1 A2.t4 218.507
R333 A2.n0 A2.t5 218.507
R334 A2.n5 A2.t6 218.507
R335 A2.n6 A2.t7 218.507
R336 A2 A2.n2 154.881
R337 A2.n4 A2.n3 152
R338 A2.n8 A2.n7 152
R339 A2.n1 A2.t3 146.208
R340 A2.n0 A2.t1 146.208
R341 A2.n5 A2.t2 146.208
R342 A2.n6 A2.t0 146.208
R343 A2.n2 A2.n1 34.904
R344 A2.n2 A2.n0 34.904
R345 A2.n4 A2.n0 34.904
R346 A2.n5 A2.n4 34.904
R347 A2.n7 A2.n5 34.904
R348 A2.n7 A2.n6 34.904
R349 A2.n3 A2 24.0005
R350 A2.n8 A2 21.4405
R351 A2 A2.n8 8.0005
R352 A2.n3 A2 5.4405
C0 a_1224_297# A2 0.137822f
C1 VPWR a_1224_297# 0.414789f
C2 VPB B2 0.134547f
C3 VGND a_1224_297# 0.010377f
C4 VPB B1 0.122346f
C5 A1 a_1224_297# 0.154463f
C6 B2 B1 0.048281f
C7 VPB A3 0.146712f
C8 Y VPB 0.026461f
C9 VPB A2 0.121951f
C10 Y B2 0.297633f
C11 VPWR VPB 0.205545f
C12 B1 A3 0.052852f
C13 Y B1 0.286943f
C14 VGND VPB 0.017656f
C15 VPWR B2 0.033781f
C16 A1 VPB 0.144732f
C17 Y A3 0.173028f
C18 VPWR B1 0.054201f
C19 VGND B2 0.035355f
C20 A3 A2 0.050706f
C21 VPWR A3 0.032326f
C22 Y A2 0.001732f
C23 VGND B1 0.030602f
C24 Y VPWR 0.057536f
C25 a_1224_297# VPB 0.017023f
C26 VGND A3 0.059304f
C27 VPWR A2 0.034089f
C28 Y VGND 0.0433f
C29 A1 Y 1.23e-19
C30 VGND A2 0.060244f
C31 VPWR VGND 0.192992f
C32 A1 A2 0.022466f
C33 A1 VPWR 0.109425f
C34 a_1224_297# A3 0.001479f
C35 Y a_1224_297# 0.013348f
C36 A1 VGND 0.065627f
C37 VGND VNB 1.07379f
C38 VPWR VNB 0.933389f
C39 Y VNB 0.028851f
C40 A1 VNB 0.432994f
C41 A2 VNB 0.368272f
C42 A3 VNB 0.41177f
C43 B1 VNB 0.353011f
C44 B2 VNB 0.415827f
C45 VPB VNB 2.0223f
C46 a_1224_297# VNB 0.006668f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_1 VPB VNB VGND VPWR X B1 A4 A3 A2 A1
X0 VGND.t0 A4.t0 a_321_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47.t4 A3.t0 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21.t2 B1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t0 a_103_21.t3 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND.t1 a_103_21.t4 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND.t2 A2.t0 a_321_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47.t3 A1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297.t1 A3.t1 a_393_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297.t1 A2.t1 a_511_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47.t1 B1.t1 a_103_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297.t0 A4.t1 a_103_21.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR.t2 A1.t1 a_619_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
R0 A4.n0 A4.t1 233.01
R1 A4 A4.n0 163.055
R2 A4.n0 A4.t0 162.919
R3 a_321_47.n2 a_321_47.n1 259.918
R4 a_321_47.n1 a_321_47.t3 186.724
R5 a_321_47.n1 a_321_47.n0 98.788
R6 a_321_47.n0 a_321_47.t2 36.9236
R7 a_321_47.n0 a_321_47.t4 35.0774
R8 a_321_47.t0 a_321_47.n2 24.9236
R9 a_321_47.n2 a_321_47.t1 24.9236
R10 VGND.n0 VGND.t1 290.289
R11 VGND.n3 VGND.n2 205.167
R12 VGND.n5 VGND.n4 199.739
R13 VGND.n2 VGND.t3 36.0005
R14 VGND.n2 VGND.t2 36.0005
R15 VGND.n4 VGND.t4 35.0774
R16 VGND.n4 VGND.t0 35.0774
R17 VGND.n7 VGND.n6 34.6358
R18 VGND.n6 VGND.n5 33.1299
R19 VGND.n7 VGND.n0 26.3534
R20 VGND.n9 VGND.n0 15.9414
R21 VGND.n8 VGND.n7 9.3005
R22 VGND.n6 VGND.n1 9.3005
R23 VGND.n5 VGND.n3 6.03512
R24 VGND.n3 VGND.n1 0.329556
R25 VGND.n9 VGND.n8 0.141672
R26 VGND VGND.n9 0.121778
R27 VGND.n8 VGND.n1 0.120292
R28 VNB.t2 VNB.t1 2677.02
R29 VNB.t3 VNB.t4 1537.86
R30 VNB.t5 VNB.t3 1537.86
R31 VNB.t0 VNB.t5 1509.39
R32 VNB VNB.t2 1267.31
R33 VNB.t1 VNB.t0 1196.12
R34 A3.n0 A3.t1 236.18
R35 A3.n0 A3.t0 163.881
R36 A3 A3.n0 163.055
R37 B1.n0 B1.t0 262.575
R38 B1.n0 B1.t1 157.308
R39 B1 B1.n0 157.181
R40 VPWR.n1 VPWR.n0 315.889
R41 VPWR.n1 VPWR.t2 250.446
R42 VPWR.n0 VPWR.t1 26.5955
R43 VPWR.n0 VPWR.t0 26.5955
R44 VPWR VPWR.n1 0.243566
R45 a_103_21.n2 a_103_21.n1 235.744
R46 a_103_21.n0 a_103_21.t3 234.173
R47 a_103_21.n0 a_103_21.t4 162.7
R48 a_103_21.n1 a_103_21.n0 154.744
R49 a_103_21.n1 a_103_21.t1 154.456
R50 a_103_21.t0 a_103_21.n2 60.0855
R51 a_103_21.n2 a_103_21.t2 42.3555
R52 VPB.t3 VPB.t1 396.574
R53 VPB VPB.t2 387.695
R54 VPB.t1 VPB.t5 349.221
R55 VPB.t0 VPB.t4 319.627
R56 VPB.t5 VPB.t0 319.627
R57 VPB.t2 VPB.t3 248.599
R58 X.n1 X 589.51
R59 X.n1 X.n0 585
R60 X.n2 X.n1 585
R61 X.n5 X 186.695
R62 X.n6 X.n5 185
R63 X.n1 X.t1 55.1605
R64 X.n5 X.t0 47.0774
R65 X.n6 X 11.1064
R66 X.n4 X 10.4301
R67 X.n4 X 5.68939
R68 X X.n4 4.51815
R69 X.n0 X 4.51098
R70 X.n3 X.n2 4.26717
R71 X.n0 X 3.77955
R72 X.n2 X 3.77955
R73 X X.n6 1.69462
R74 X X.n3 0.474574
R75 X.n3 X 0.24431
R76 A2.n0 A2.t1 236.18
R77 A2.n0 A2.t0 163.881
R78 A2 A2.n0 161.859
R79 A1.n0 A1.t1 236.18
R80 A1.n0 A1.t0 163.881
R81 A1 A1.n0 160.96
R82 a_393_297.t0 a_393_297.t1 86.6805
R83 a_511_297.t0 a_511_297.t1 76.8305
R84 a_619_297.t0 a_619_297.t1 76.8305
C0 X VPWR 0.115292f
C1 X VGND 0.073169f
C2 B1 VPB 0.038249f
C3 A4 VPB 0.039801f
C4 A3 VPB 0.034632f
C5 B1 A4 0.066022f
C6 VPWR VPB 0.095809f
C7 A2 VPB 0.036241f
C8 VGND VPB 0.007783f
C9 A1 VPB 0.036759f
C10 VPWR B1 0.019751f
C11 A4 A3 0.142408f
C12 VPWR A4 0.047227f
C13 VGND B1 0.017222f
C14 X VPB 0.019388f
C15 VPWR A3 0.042939f
C16 VGND A4 0.018823f
C17 A3 A2 0.156111f
C18 X B1 6.86e-19
C19 VGND A3 0.015847f
C20 VPWR A2 0.09531f
C21 VPWR VGND 0.081228f
C22 VPWR A1 0.054343f
C23 VGND A2 0.016385f
C24 A2 A1 0.072316f
C25 VGND A1 0.017159f
C26 VGND VNB 0.493571f
C27 VPWR VNB 0.444338f
C28 X VNB 0.094186f
C29 A1 VNB 0.134954f
C30 A2 VNB 0.101364f
C31 A3 VNB 0.096317f
C32 A4 VNB 0.099398f
C33 B1 VNB 0.112101f
C34 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_2 VNB VPB VGND VPWR A1 A2 A3 A4 B1 X
X0 VGND.t4 A2.t0 a_393_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11375 ps=1 w=0.65 l=0.15
X1 a_496_297.t1 A4.t0 a_79_21.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.3025 ps=1.605 w=1 l=0.15
X2 a_393_47.t2 A3.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.115375 ps=1.005 w=0.65 l=0.15
X3 VPWR.t1 A1.t0 a_697_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=2.82 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR.t2 a_79_21.t3 X.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t2 a_79_21.t4 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_79_21.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3025 pd=1.605 as=0.305 ps=1.61 w=1 l=0.15
X7 VGND.t0 A4.t1 a_393_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.118625 ps=1.015 w=0.65 l=0.15
X8 a_697_297.t0 A2.t1 a_597_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 a_393_47.t4 A1.t1 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.2665 pd=2.12 as=0.11375 ps=1 w=0.65 l=0.15
X10 X.t2 a_79_21.t5 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_393_47.t1 B1.t1 a_79_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.208 ps=1.94 w=0.65 l=0.15
X12 a_597_297.t0 A3.t1 a_496_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.1775 ps=1.355 w=1 l=0.15
X13 X.t0 a_79_21.t6 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t1 239.505
R1 A2.n0 A2.t0 167.204
R2 A2.n1 A2.n0 152
R3 A2.n1 A2 11.055
R4 A2 A2.n1 2.13383
R5 a_393_47.n1 a_393_47.t4 196.954
R6 a_393_47.n2 a_393_47.n1 142.291
R7 a_393_47.n1 a_393_47.n0 99.1759
R8 a_393_47.n0 a_393_47.t3 39.6928
R9 a_393_47.n2 a_393_47.t1 34.1543
R10 a_393_47.t0 a_393_47.n2 33.2313
R11 a_393_47.n0 a_393_47.t2 24.9236
R12 VGND.n3 VGND.n2 210.029
R13 VGND.n5 VGND.n4 203.356
R14 VGND.n10 VGND.t2 155.993
R15 VGND.n12 VGND.t3 154.599
R16 VGND.n4 VGND.t1 40.6159
R17 VGND.n2 VGND.t5 36.0005
R18 VGND.n6 VGND.n1 34.6358
R19 VGND.n6 VGND.n5 31.2476
R20 VGND.n2 VGND.t4 28.6159
R21 VGND.n10 VGND.n1 26.3534
R22 VGND.n12 VGND.n11 25.977
R23 VGND.n4 VGND.t0 24.9236
R24 VGND.n11 VGND.n10 24.4711
R25 VGND.n13 VGND.n12 9.3005
R26 VGND.n7 VGND.n6 9.3005
R27 VGND.n8 VGND.n1 9.3005
R28 VGND.n10 VGND.n9 9.3005
R29 VGND.n11 VGND.n0 9.3005
R30 VGND.n5 VGND.n3 6.53872
R31 VGND.n7 VGND.n3 0.417714
R32 VGND.n8 VGND.n7 0.120292
R33 VGND.n9 VGND.n8 0.120292
R34 VGND.n9 VGND.n0 0.120292
R35 VGND.n13 VGND.n0 0.120292
R36 VGND VGND.n13 0.0213333
R37 VNB.t3 VNB.t1 2847.9
R38 VNB.t1 VNB.t0 1466.67
R39 VNB.t0 VNB.t2 1438.19
R40 VNB.t5 VNB.t6 1423.95
R41 VNB.t2 VNB.t5 1423.95
R42 VNB.t4 VNB.t3 1196.12
R43 VNB VNB.t4 911.327
R44 A4.n0 A4.t0 239.04
R45 A4.n0 A4.t1 166.739
R46 A4.n1 A4.n0 152
R47 A4.n1 A4 11.055
R48 A4 A4.n1 2.13383
R49 a_79_21.n3 a_79_21.n2 223.044
R50 a_79_21.n2 a_79_21.n1 208.891
R51 a_79_21.n1 a_79_21.t3 205.654
R52 a_79_21.n0 a_79_21.t5 205.654
R53 a_79_21.n2 a_79_21.t1 155.144
R54 a_79_21.n1 a_79_21.t4 133.353
R55 a_79_21.n0 a_79_21.t6 133.353
R56 a_79_21.n3 a_79_21.t2 92.5905
R57 a_79_21.n1 a_79_21.n0 54.714
R58 a_79_21.t0 a_79_21.n3 26.5955
R59 a_496_297.t0 a_496_297.t1 69.9355
R60 VPB.t6 VPB.t0 449.844
R61 VPB.t0 VPB.t4 446.885
R62 VPB.t4 VPB.t3 298.911
R63 VPB.t2 VPB.t1 295.95
R64 VPB.t3 VPB.t2 295.95
R65 VPB.t5 VPB.t6 248.599
R66 VPB VPB.t5 189.409
R67 A3.n0 A3.t1 239.505
R68 A3.n0 A3.t0 167.204
R69 A3.n1 A3.n0 152
R70 A3.n1 A3 11.055
R71 A3 A3.n1 2.13383
R72 A1.n0 A1.t0 239.505
R73 A1.n0 A1.t1 167.204
R74 A1 A1.n0 167.105
R75 a_697_297.t0 a_697_297.t1 68.9505
R76 VPWR.n1 VPWR.t1 272.159
R77 VPWR.n5 VPWR.t3 249.362
R78 VPWR.n3 VPWR.n2 126.624
R79 VPWR.n2 VPWR.t0 66.3149
R80 VPWR.n2 VPWR.t2 52.4308
R81 VPWR.n5 VPWR.n4 25.977
R82 VPWR.n4 VPWR.n3 24.4711
R83 VPWR.n4 VPWR.n0 9.3005
R84 VPWR.n6 VPWR.n5 9.3005
R85 VPWR.n3 VPWR.n1 5.5539
R86 VPWR.n1 VPWR.n0 0.179192
R87 VPWR.n6 VPWR.n0 0.120292
R88 VPWR VPWR.n6 0.0213333
R89 X X.n0 593.34
R90 X.n6 X.n0 585
R91 X.n5 X.n0 585
R92 X.n1 X 186.745
R93 X.n2 X.n1 185
R94 X.n0 X.t3 26.5955
R95 X.n0 X.t2 26.5955
R96 X.n1 X.t1 24.9236
R97 X.n1 X.t0 24.9236
R98 X.n2 X 11.4429
R99 X X.n3 10.4732
R100 X.n6 X 8.33989
R101 X.n5 X.n4 6.4005
R102 X.n3 X 5.35323
R103 X X.n6 4.84898
R104 X X.n5 4.84898
R105 X.n3 X 4.46111
R106 X.n4 X 2.32777
R107 X.n4 X 1.93989
R108 X X.n2 1.74595
R109 B1.n0 B1.t0 264.565
R110 B1 B1.n0 162.78
R111 B1.n0 B1.t1 149.421
R112 a_597_297.t0 a_597_297.t1 68.9505
C0 VPWR VPB 0.112815f
C1 A4 B1 0.061147f
C2 VPWR B1 0.012947f
C3 X VGND 0.151826f
C4 A3 A2 0.154008f
C5 VPB X 0.005245f
C6 A3 A1 1.55e-20
C7 VPB VGND 0.008849f
C8 A4 A3 0.154057f
C9 A2 A1 0.078498f
C10 A3 VPWR 0.039499f
C11 B1 VGND 0.021653f
C12 VPB B1 0.046228f
C13 A2 VPWR 0.079841f
C14 A1 VPWR 0.05588f
C15 A4 VPWR 0.040421f
C16 A3 VGND 0.015214f
C17 A3 VPB 0.031018f
C18 A2 VGND 0.015659f
C19 A2 VPB 0.032933f
C20 A1 VGND 0.017271f
C21 VPWR X 0.209267f
C22 A4 VGND 0.017864f
C23 A1 VPB 0.036922f
C24 VPWR VGND 0.106546f
C25 A4 VPB 0.035566f
C26 VGND VNB 0.569697f
C27 X VNB 0.024476f
C28 VPWR VNB 0.519348f
C29 A1 VNB 0.133247f
C30 A2 VNB 0.095692f
C31 A3 VNB 0.091907f
C32 A4 VNB 0.093185f
C33 B1 VNB 0.121943f
C34 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 VPWR VPB VGND VPWRIN A X
X0 a_1028_32.t0 a_620_911.t5 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VGND.t15 A.t0 a_714_58.t3 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND.t17 a_505_297.t2 a_620_911.t3 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X3 X.t0 a_1028_32.t2 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND.t13 A.t1 a_714_58.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_620_911.t4 a_505_297.t3 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_714_58.t0 A.t2 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_714_58.t1 A.t3 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X8 a_1028_32.t1 a_620_911.t6 VGND.t21 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X9 VGND.t3 a_505_297.t4 a_620_911.t0 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 a_505_297.t1 A.t4 VPWRIN.t1 VPWRIN.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X11 VPWR.t0 a_714_58.t5 a_620_911.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1185 pd=1.09 as=0.21725 ps=2.13 w=0.79 l=0.15
X12 X.t1 a_1028_32.t3 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.21725 pd=2.13 as=0.1185 ps=1.09 w=0.79 l=0.15
X13 VPWR.t2 a_620_911.t7 a_714_58.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X14 a_505_297.t0 A.t5 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X15 a_620_911.t1 a_505_297.t5 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t2 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t3 25.8467
R14 a_620_911.n1 a_620_911.t1 25.8467
R15 a_620_911.n0 a_620_911.t0 25.8467
R16 a_620_911.n0 a_620_911.t4 25.8467
R17 VPWR.n2 VPWR.n1 326.825
R18 VPWR.n2 VPWR.n0 325.817
R19 VPWR.n0 VPWR.t3 38.6524
R20 VPWR.n0 VPWR.t2 37.4056
R21 VPWR.n1 VPWR.t1 37.4056
R22 VPWR.n1 VPWR.t0 37.4056
R23 VPWR VPWR.n2 21.8082
R24 a_1028_32.n1 a_1028_32.n0 780.957
R25 a_1028_32.t0 a_1028_32.n1 376.678
R26 a_1028_32.n0 a_1028_32.t2 195.912
R27 a_1028_32.n1 a_1028_32.t1 144.809
R28 a_1028_32.n0 a_1028_32.t3 59.9423
R29 VPB VPB.t2 463.961
R30 VPB.t0 VPB.t1 151.06
R31 VPB.t2 VPB.t0 1.67895
R32 A.n0 A.t0 284.38
R33 A.n3 A.t4 268.313
R34 A.n3 A.t5 165.989
R35 A.n4 A.n3 156.262
R36 A A.n4 154.452
R37 A.n1 A.t1 146.208
R38 A.n0 A.t2 146.208
R39 A.n2 A.t3 146.208
R40 A.n1 A.n0 138.173
R41 A.n2 A.n1 136.774
R42 A.n4 A.n2 87.8489
R43 a_714_58.t4 a_714_58.n3 481.457
R44 a_714_58.n3 a_714_58.t5 446.346
R45 a_714_58.n2 a_714_58.n0 120.412
R46 a_714_58.n2 a_714_58.n1 116.829
R47 a_714_58.n3 a_714_58.n2 95.4968
R48 a_714_58.n1 a_714_58.t2 25.8467
R49 a_714_58.n1 a_714_58.t1 25.8467
R50 a_714_58.n0 a_714_58.t3 25.8467
R51 a_714_58.n0 a_714_58.t0 25.8467
R52 VGND.n54 VGND.n2 9804.72
R53 VGND.n53 VGND.n52 9804.72
R54 VGND.t18 VGND.n2 4955.34
R55 VGND.n55 VGND.n54 4202.78
R56 VGND.n33 VGND.n2 4202.78
R57 VGND.t20 VGND.n51 3839.97
R58 VGND.t0 VGND.n26 3469.08
R59 VGND.n54 VGND.t6 3346.28
R60 VGND.t6 VGND.t10 2947.57
R61 VGND.t16 VGND.t20 2192.88
R62 VGND.t14 VGND.t0 1224.6
R63 VGND.t8 VGND.t14 1224.6
R64 VGND.t12 VGND.t8 1224.6
R65 VGND.t4 VGND.t16 1224.6
R66 VGND.t2 VGND.t18 1224.6
R67 VGND.n53 VGND.t12 882.848
R68 VGND.n52 VGND.t4 768.933
R69 VGND.n52 VGND.t2 455.663
R70 VGND.t10 VGND.n53 341.748
R71 VGND.n14 VGND.t7 249.048
R72 VGND.n22 VGND.n21 203.424
R73 VGND.n42 VGND.t19 154.561
R74 VGND.n8 VGND.t11 139.954
R75 VGND.n29 VGND.n28 122.484
R76 VGND.n4 VGND.n3 114.109
R77 VGND.n50 VGND.n49 59.678
R78 VGND.n49 VGND.t21 57.2313
R79 VGND.n49 VGND.t17 57.2313
R80 VGND.n41 VGND.n31 34.6358
R81 VGND.n37 VGND.n31 34.6358
R82 VGND.n37 VGND.n36 34.6358
R83 VGND.n36 VGND.n35 34.6358
R84 VGND.n44 VGND.n43 34.6358
R85 VGND.n48 VGND.n47 34.6358
R86 VGND.n10 VGND.n9 34.6358
R87 VGND.n10 VGND.n1 34.6358
R88 VGND.n16 VGND.n15 34.6358
R89 VGND.n20 VGND.n6 34.6358
R90 VGND.n24 VGND.n23 34.6358
R91 VGND.n14 VGND.n9 30.8711
R92 VGND.n28 VGND.t5 25.8467
R93 VGND.n28 VGND.t3 25.8467
R94 VGND.n21 VGND.t9 25.8467
R95 VGND.n21 VGND.t13 25.8467
R96 VGND.n3 VGND.t1 25.8467
R97 VGND.n3 VGND.t15 25.8467
R98 VGND.n35 VGND.n33 23.7181
R99 VGND.n55 VGND.n1 23.7181
R100 VGND.n26 VGND.n4 16.2466
R101 VGND.n15 VGND.n14 13.5534
R102 VGND.n47 VGND.n29 10.9181
R103 VGND.n44 VGND.n29 9.41227
R104 VGND.n16 VGND.n8 9.41227
R105 VGND VGND.n55 9.34738
R106 VGND VGND.n33 9.32654
R107 VGND.n12 VGND.n9 9.3005
R108 VGND.n11 VGND.n10 9.3005
R109 VGND.n1 VGND.n0 9.3005
R110 VGND.n14 VGND.n13 9.3005
R111 VGND.n17 VGND.n16 9.3005
R112 VGND.n15 VGND.n7 9.3005
R113 VGND.n20 VGND.n19 9.3005
R114 VGND.n18 VGND.n6 9.3005
R115 VGND.n25 VGND.n24 9.3005
R116 VGND.n23 VGND.n5 9.3005
R117 VGND.n48 VGND.n27 9.3005
R118 VGND.n47 VGND.n46 9.3005
R119 VGND.n45 VGND.n44 9.3005
R120 VGND.n43 VGND.n30 9.3005
R121 VGND.n41 VGND.n40 9.3005
R122 VGND.n39 VGND.n31 9.3005
R123 VGND.n38 VGND.n37 9.3005
R124 VGND.n36 VGND.n32 9.3005
R125 VGND.n35 VGND.n34 9.3005
R126 VGND.n42 VGND.n41 8.65932
R127 VGND.n51 VGND.n50 7.05995
R128 VGND.n43 VGND.n42 6.4005
R129 VGND.n50 VGND.n48 5.64756
R130 VGND.n22 VGND.n20 4.89462
R131 VGND.n23 VGND.n22 4.89462
R132 VGND.n26 VGND.n25 0.878118
R133 VGND.n8 VGND.n6 0.376971
R134 VGND.n24 VGND.n4 0.376971
R135 VGND.n51 VGND.n27 0.314038
R136 VGND.n25 VGND.n5 0.120292
R137 VGND.n19 VGND.n5 0.120292
R138 VGND.n19 VGND.n18 0.120292
R139 VGND.n18 VGND.n17 0.120292
R140 VGND.n17 VGND.n7 0.120292
R141 VGND.n13 VGND.n7 0.120292
R142 VGND.n13 VGND.n12 0.120292
R143 VGND.n12 VGND.n11 0.120292
R144 VGND.n11 VGND.n0 0.120292
R145 VGND.n46 VGND.n27 0.120292
R146 VGND.n46 VGND.n45 0.120292
R147 VGND.n45 VGND.n30 0.120292
R148 VGND.n40 VGND.n30 0.120292
R149 VGND.n40 VGND.n39 0.120292
R150 VGND.n39 VGND.n38 0.120292
R151 VGND.n38 VGND.n32 0.120292
R152 VGND.n34 VGND.n32 0.120292
R153 VGND.n34 VGND 0.09425
R154 VGND VGND.n0 0.0734167
R155 a_505_297.t1 a_505_297.n5 742.867
R156 a_505_297.t1 a_505_297.n6 724.692
R157 a_505_297.n5 a_505_297.n4 311.748
R158 a_505_297.n6 a_505_297.t0 287.401
R159 a_505_297.n0 a_505_297.t2 266.707
R160 a_505_297.n3 a_505_297.t3 137.474
R161 a_505_297.n1 a_505_297.n0 133.353
R162 a_505_297.n0 a_505_297.t5 128.534
R163 a_505_297.n2 a_505_297.t4 117.287
R164 a_505_297.n3 a_505_297.n2 60.56
R165 a_505_297.n4 a_505_297.n1 19.2805
R166 a_505_297.n6 a_505_297.n5 18.1338
R167 a_505_297.n2 a_505_297.n1 14.0588
R168 a_505_297.n4 a_505_297.n3 4.94459
R169 X X.t1 391.517
R170 X X.t0 128.451
R171 X.n0 X 16.7569
R172 X X.n0 0.465955
R173 X.n0 X 0.427167
R174 VPWRIN.n0 VPWRIN.t0 1565.73
R175 VPWRIN.n0 VPWRIN.t1 370.75
R176 VPWRIN VPWRIN.n0 7.13856
C0 VPB VPWRIN 0.106224f
C1 VPB VPWR 0.528032f
C2 VPB X 0.021096f
C3 VPWRIN VPWR 0.771396f
C4 VPWRIN X 0.026094f
C5 VPWR X 0.073906f
C6 VPB A 0.019913f
C7 VPWRIN A 0.089133f
C8 VPWR A 0.004863f
C9 A X 0.002926f
C10 X VGND 0.179867f
C11 A VGND 0.636418f
C12 VPWR VGND 0.267901f
C13 VPWRIN VGND 0.691791f
C14 VPB VGND 1.44754f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 VPWR VPB VGND VPWRIN A X
X0 a_1032_911.t1 a_620_911.t5 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VGND.t15 A.t0 a_714_47.t4 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND.t21 a_505_297.t2 a_620_911.t3 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X3 X.t3 a_1032_911.t2 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.154625 ps=1.325 w=1 l=0.15
X4 VGND.t13 A.t1 a_714_47.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_620_911.t4 a_505_297.t3 VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_714_47.t2 A.t2 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 X.t1 a_1032_911.t3 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_714_47.t1 A.t3 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X9 VPWR.t2 a_1032_911.t4 X.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.185 ps=1.37 w=1 l=0.15
X10 VGND.t1 a_1032_911.t5 X.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.12025 ps=1.02 w=0.65 l=0.15
X11 a_1032_911.t0 a_620_911.t6 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X12 VGND.t17 a_505_297.t4 a_620_911.t1 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_505_297.t0 A.t4 VPWRIN.t1 VPWRIN.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X14 VPWR.t0 a_714_47.t5 a_620_911.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.154625 pd=1.325 as=0.21725 ps=2.13 w=0.79 l=0.15
X15 VPWR.t4 a_620_911.t7 a_714_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X16 a_505_297.t1 A.t5 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X17 a_620_911.t2 a_505_297.t5 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t0 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t3 25.8467
R14 a_620_911.n1 a_620_911.t2 25.8467
R15 a_620_911.n0 a_620_911.t1 25.8467
R16 a_620_911.n0 a_620_911.t4 25.8467
R17 VPWR.n3 VPWR.t2 416.57
R18 VPWR.n2 VPWR.n1 326.825
R19 VPWR.n2 VPWR.n0 325.817
R20 VPWR.n0 VPWR.t3 38.6524
R21 VPWR.n1 VPWR.t1 38.4132
R22 VPWR.n0 VPWR.t4 37.4056
R23 VPWR.n1 VPWR.t0 37.4056
R24 VPWR.n3 VPWR.n2 19.5934
R25 VPWR VPWR.n3 2.21634
R26 a_1032_911.n2 a_1032_911.t4 843.981
R27 a_1032_911.t1 a_1032_911.n2 376.678
R28 a_1032_911.n0 a_1032_911.t2 184.768
R29 a_1032_911.t4 a_1032_911.n1 184.768
R30 a_1032_911.n1 a_1032_911.t5 168.701
R31 a_1032_911.n0 a_1032_911.t3 168.701
R32 a_1032_911.n2 a_1032_911.t0 144.809
R33 a_1032_911.n1 a_1032_911.n0 77.1205
R34 VPB.n0 VPB.t0 550.726
R35 VPB VPB.n0 206.38
R36 VPB.n0 VPB.t2 39.4319
R37 VPB.t0 VPB.t1 11.9753
R38 A.n0 A.t0 302.053
R39 A.n3 A.t4 268.313
R40 A.n3 A.t5 165.989
R41 A.n1 A.t1 163.881
R42 A.n0 A.t2 163.881
R43 A.n2 A.t3 163.881
R44 A.n4 A.n3 156.262
R45 A A.n4 154.452
R46 A.n1 A.n0 138.173
R47 A.n2 A.n1 136.774
R48 A.n4 A.n2 87.8489
R49 a_714_47.t0 a_714_47.n3 481.457
R50 a_714_47.n3 a_714_47.t5 446.346
R51 a_714_47.n2 a_714_47.n0 121.251
R52 a_714_47.n2 a_714_47.n1 117.666
R53 a_714_47.n3 a_714_47.n2 95.4968
R54 a_714_47.n1 a_714_47.t3 25.8467
R55 a_714_47.n1 a_714_47.t1 25.8467
R56 a_714_47.n0 a_714_47.t4 25.8467
R57 a_714_47.n0 a_714_47.t2 25.8467
R58 VGND.n54 VGND.n26 9804.72
R59 VGND.n53 VGND.n52 9804.72
R60 VGND.t22 VGND.n26 4955.34
R61 VGND.t4 VGND.n51 4409.49
R62 VGND.n55 VGND.n54 4202.78
R63 VGND.n33 VGND.n26 4202.78
R64 VGND.n54 VGND.t6 3346.28
R65 VGND.t6 VGND.t8 2947.57
R66 VGND.t20 VGND.t4 2192.88
R67 VGND.t2 VGND.t0 1480.91
R68 VGND.t14 VGND.t2 1338.51
R69 VGND.t10 VGND.t14 1224.6
R70 VGND.t12 VGND.t10 1224.6
R71 VGND.t18 VGND.t20 1224.6
R72 VGND.t16 VGND.t22 1224.6
R73 VGND.n53 VGND.t12 882.848
R74 VGND.n52 VGND.t18 768.933
R75 VGND.n52 VGND.t16 455.663
R76 VGND.t8 VGND.n53 341.748
R77 VGND.n20 VGND.t7 249.048
R78 VGND.n13 VGND.n5 201.292
R79 VGND.n42 VGND.t23 154.561
R80 VGND.n9 VGND.t1 143.803
R81 VGND.n3 VGND.t9 137.821
R82 VGND.n29 VGND.n28 122.484
R83 VGND.n8 VGND.n7 111.975
R84 VGND.n50 VGND.n49 59.678
R85 VGND.n49 VGND.t5 57.2313
R86 VGND.n49 VGND.t21 57.2313
R87 VGND.n41 VGND.n31 34.6358
R88 VGND.n37 VGND.n31 34.6358
R89 VGND.n37 VGND.n36 34.6358
R90 VGND.n36 VGND.n35 34.6358
R91 VGND.n44 VGND.n43 34.6358
R92 VGND.n48 VGND.n47 34.6358
R93 VGND.n24 VGND.n1 34.6358
R94 VGND.n25 VGND.n24 34.6358
R95 VGND.n19 VGND.n18 34.6358
R96 VGND.n15 VGND.n14 34.6358
R97 VGND.n12 VGND.n6 34.6358
R98 VGND.n7 VGND.t3 33.2313
R99 VGND.n20 VGND.n1 30.8711
R100 VGND.n28 VGND.t19 25.8467
R101 VGND.n28 VGND.t17 25.8467
R102 VGND.n5 VGND.t11 25.8467
R103 VGND.n5 VGND.t13 25.8467
R104 VGND.n7 VGND.t15 25.8467
R105 VGND.n35 VGND.n33 23.7181
R106 VGND.n55 VGND.n25 23.7181
R107 VGND.n9 VGND.n8 16.1542
R108 VGND.n20 VGND.n19 13.5534
R109 VGND.n47 VGND.n29 10.9181
R110 VGND.n44 VGND.n29 9.41227
R111 VGND.n18 VGND.n3 9.41227
R112 VGND VGND.n55 9.34738
R113 VGND VGND.n33 9.32654
R114 VGND.n10 VGND.n6 9.3005
R115 VGND.n12 VGND.n11 9.3005
R116 VGND.n14 VGND.n4 9.3005
R117 VGND.n16 VGND.n15 9.3005
R118 VGND.n18 VGND.n17 9.3005
R119 VGND.n19 VGND.n2 9.3005
R120 VGND.n21 VGND.n20 9.3005
R121 VGND.n22 VGND.n1 9.3005
R122 VGND.n24 VGND.n23 9.3005
R123 VGND.n25 VGND.n0 9.3005
R124 VGND.n48 VGND.n27 9.3005
R125 VGND.n47 VGND.n46 9.3005
R126 VGND.n45 VGND.n44 9.3005
R127 VGND.n43 VGND.n30 9.3005
R128 VGND.n41 VGND.n40 9.3005
R129 VGND.n39 VGND.n31 9.3005
R130 VGND.n38 VGND.n37 9.3005
R131 VGND.n36 VGND.n32 9.3005
R132 VGND.n35 VGND.n34 9.3005
R133 VGND.n42 VGND.n41 8.65932
R134 VGND.n51 VGND.n50 7.14073
R135 VGND.n43 VGND.n42 6.4005
R136 VGND.n50 VGND.n48 5.64756
R137 VGND.n14 VGND.n13 4.89462
R138 VGND.n13 VGND.n12 4.89462
R139 VGND.n10 VGND.n9 0.960602
R140 VGND.n15 VGND.n3 0.376971
R141 VGND.n8 VGND.n6 0.376971
R142 VGND.n51 VGND.n27 0.234391
R143 VGND.n11 VGND.n10 0.120292
R144 VGND.n11 VGND.n4 0.120292
R145 VGND.n16 VGND.n4 0.120292
R146 VGND.n17 VGND.n16 0.120292
R147 VGND.n17 VGND.n2 0.120292
R148 VGND.n21 VGND.n2 0.120292
R149 VGND.n22 VGND.n21 0.120292
R150 VGND.n23 VGND.n22 0.120292
R151 VGND.n23 VGND.n0 0.120292
R152 VGND.n46 VGND.n27 0.120292
R153 VGND.n46 VGND.n45 0.120292
R154 VGND.n45 VGND.n30 0.120292
R155 VGND.n40 VGND.n30 0.120292
R156 VGND.n40 VGND.n39 0.120292
R157 VGND.n39 VGND.n38 0.120292
R158 VGND.n38 VGND.n32 0.120292
R159 VGND.n34 VGND.n32 0.120292
R160 VGND.n34 VGND 0.09425
R161 VGND VGND.n0 0.0734167
R162 a_505_297.t0 a_505_297.n5 742.867
R163 a_505_297.t0 a_505_297.n6 724.692
R164 a_505_297.n5 a_505_297.n4 311.748
R165 a_505_297.n6 a_505_297.t1 287.401
R166 a_505_297.n0 a_505_297.t2 266.707
R167 a_505_297.n3 a_505_297.t3 137.474
R168 a_505_297.n1 a_505_297.n0 133.353
R169 a_505_297.n0 a_505_297.t5 128.534
R170 a_505_297.n2 a_505_297.t4 117.287
R171 a_505_297.n3 a_505_297.n2 60.56
R172 a_505_297.n4 a_505_297.n1 19.2805
R173 a_505_297.n6 a_505_297.n5 18.1338
R174 a_505_297.n2 a_505_297.n1 14.0588
R175 a_505_297.n4 a_505_297.n3 4.94459
R176 X X.n1 318.197
R177 X X.n0 104.951
R178 X.n1 X.t2 45.3105
R179 X.n0 X.t0 42.462
R180 X.n1 X.t3 27.5805
R181 X.n0 X.t1 25.8467
R182 X.n2 X 16.7569
R183 X X.n2 0.465955
R184 X.n2 X 0.427167
R185 VPWRIN.n0 VPWRIN.t0 1565.73
R186 VPWRIN.n0 VPWRIN.t1 370.75
R187 VPWRIN VPWRIN.n0 7.13856
C0 A VPB 0.019925f
C1 A X 0.00292f
C2 A VPWRIN 0.089133f
C3 X VPB 0.008022f
C4 VPB VPWRIN 0.103298f
C5 X VPWRIN 0.026823f
C6 A VPWR 0.004863f
C7 VPB VPWR 0.534275f
C8 X VPWR 0.129496f
C9 VPWRIN VPWR 0.805258f
C10 X VGND 0.178135f
C11 A VGND 0.654458f
C12 VPWR VGND 0.29254f
C13 VPWRIN VGND 0.696853f
C14 VPB VGND 1.45906f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 VPWR VPB VGND VPWRIN A X
X0 a_1032_911.t1 a_620_911.t5 VPWR.t6 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VPWR.t0 a_1032_911.t2 X.t7 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2 VGND.t9 A.t0 a_714_47.t3 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VGND.t15 a_505_297.t2 a_620_911.t2 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X4 X.t6 a_1032_911.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.154625 ps=1.325 w=1 l=0.15
X5 VGND.t7 A.t1 a_714_47.t2 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_620_911.t0 a_505_297.t3 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_714_47.t1 A.t2 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 X.t1 a_1032_911.t4 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.104 ps=0.97 w=0.65 l=0.15
X9 VGND.t25 a_1032_911.t5 X.t0 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X10 a_714_47.t0 A.t3 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X11 VPWR.t2 a_1032_911.t6 X.t5 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12 VGND.t23 a_1032_911.t7 X.t3 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12025 ps=1.02 w=0.65 l=0.15
X13 a_1032_911.t0 a_620_911.t6 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X14 VGND.t13 a_505_297.t4 a_620_911.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_505_297.t1 A.t4 VPWRIN.t1 VPWRIN.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X16 VPWR.t4 a_714_47.t5 a_620_911.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.154625 pd=1.325 as=0.21725 ps=2.13 w=0.79 l=0.15
X17 X.t2 a_1032_911.t8 VGND.t21 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VPWR.t5 a_620_911.t7 a_714_47.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X19 X.t4 a_1032_911.t9 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_505_297.t0 A.t5 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X21 a_620_911.t4 a_505_297.t5 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t3 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t2 25.8467
R14 a_620_911.n1 a_620_911.t4 25.8467
R15 a_620_911.n0 a_620_911.t1 25.8467
R16 a_620_911.n0 a_620_911.t0 25.8467
R17 VPWR.n2 VPWR.t0 416.128
R18 VPWR.n3 VPWR.n1 332.486
R19 VPWR.n7 VPWR.n6 326.825
R20 VPWR.n7 VPWR.n5 325.817
R21 VPWR.n5 VPWR.t6 38.6524
R22 VPWR.n6 VPWR.t1 38.4132
R23 VPWR.n5 VPWR.t5 37.4056
R24 VPWR.n6 VPWR.t4 37.4056
R25 VPWR.n8 VPWR.n4 34.6358
R26 VPWR.n1 VPWR.t3 27.5805
R27 VPWR.n1 VPWR.t2 27.5805
R28 VPWR.n3 VPWR.n2 23.1308
R29 VPWR.n4 VPWR.n3 18.0711
R30 VPWR.n8 VPWR.n7 12.8005
R31 VPWR.n4 VPWR.n0 9.3005
R32 VPWR.n9 VPWR.n8 9.3005
R33 VPWR VPWR.n9 1.38004
R34 VPWR.n2 VPWR.n0 1.16591
R35 VPWR.n9 VPWR.n0 0.120292
R36 a_1032_911.n6 a_1032_911.n5 472.841
R37 a_1032_911.n4 a_1032_911.t2 461.113
R38 a_1032_911.t1 a_1032_911.n6 376.678
R39 a_1032_911.n4 a_1032_911.t9 322.94
R40 a_1032_911.n5 a_1032_911.t6 322.94
R41 a_1032_911.n2 a_1032_911.t9 184.768
R42 a_1032_911.n1 a_1032_911.t6 184.768
R43 a_1032_911.n0 a_1032_911.t3 184.768
R44 a_1032_911.t2 a_1032_911.n3 184.768
R45 a_1032_911.n3 a_1032_911.t5 168.701
R46 a_1032_911.n2 a_1032_911.t8 168.701
R47 a_1032_911.n1 a_1032_911.t7 168.701
R48 a_1032_911.n0 a_1032_911.t4 168.701
R49 a_1032_911.n6 a_1032_911.t0 144.809
R50 a_1032_911.n5 a_1032_911.n4 138.173
R51 a_1032_911.n1 a_1032_911.n0 77.1205
R52 a_1032_911.n3 a_1032_911.n2 63.7728
R53 a_1032_911.n2 a_1032_911.n1 63.7728
R54 VPB.n0 VPB.t2 416.839
R55 VPB VPB.n0 206.714
R56 VPB.n0 VPB.t1 29.6401
R57 VPB.t2 VPB.t0 9.03378
R58 X.n6 X.n0 314.94
R59 X.n5 X.n3 314.938
R60 X.n5 X.n4 117.287
R61 X X.n1 104.951
R62 X.n0 X.t5 45.3105
R63 X.n1 X.t3 42.462
R64 X.n6 X.n5 36.2343
R65 X.n3 X.t7 27.5805
R66 X.n3 X.t4 27.5805
R67 X.n0 X.t6 27.5805
R68 X.n1 X.t1 25.8467
R69 X.n4 X.t0 25.8467
R70 X.n4 X.t2 25.8467
R71 X.n6 X.n2 4.88777
R72 X X.n6 3.25868
R73 X.n6 X 2.36358
R74 X.n2 X 0.465955
R75 X.n2 X 0.427167
R76 A.n0 A.t0 302.053
R77 A.n3 A.t4 268.313
R78 A.n3 A.t5 165.989
R79 A.n1 A.t1 163.881
R80 A.n0 A.t2 163.881
R81 A.n2 A.t3 163.881
R82 A.n4 A.n3 156.262
R83 A A.n4 154.452
R84 A.n1 A.n0 138.173
R85 A.n2 A.n1 136.774
R86 A.n4 A.n2 87.8489
R87 a_714_47.t4 a_714_47.n3 481.457
R88 a_714_47.n3 a_714_47.t5 446.346
R89 a_714_47.n2 a_714_47.n0 121.251
R90 a_714_47.n2 a_714_47.n1 117.666
R91 a_714_47.n3 a_714_47.n2 95.4968
R92 a_714_47.n1 a_714_47.t2 25.8467
R93 a_714_47.n1 a_714_47.t0 25.8467
R94 a_714_47.n0 a_714_47.t3 25.8467
R95 a_714_47.n0 a_714_47.t1 25.8467
R96 VGND.n60 VGND.n32 9804.72
R97 VGND.n59 VGND.n58 9804.72
R98 VGND.t16 VGND.n57 7029.87
R99 VGND.t10 VGND.n32 4955.34
R100 VGND.n61 VGND.n60 4202.78
R101 VGND.n39 VGND.n32 4202.78
R102 VGND.n60 VGND.t0 3346.28
R103 VGND.t0 VGND.t2 2947.57
R104 VGND.t14 VGND.t16 2192.88
R105 VGND.t26 VGND.t22 1480.91
R106 VGND.t8 VGND.t26 1338.51
R107 VGND.t20 VGND.t24 1224.6
R108 VGND.t22 VGND.t20 1224.6
R109 VGND.t4 VGND.t8 1224.6
R110 VGND.t6 VGND.t4 1224.6
R111 VGND.t18 VGND.t14 1224.6
R112 VGND.t12 VGND.t10 1224.6
R113 VGND.n59 VGND.t6 882.848
R114 VGND.n58 VGND.t18 768.933
R115 VGND.n58 VGND.t12 455.663
R116 VGND.t2 VGND.n59 341.748
R117 VGND.n26 VGND.t1 249.048
R118 VGND.n19 VGND.n5 201.292
R119 VGND.n48 VGND.t11 154.561
R120 VGND.n9 VGND.t25 151.21
R121 VGND.n3 VGND.t3 137.821
R122 VGND.n35 VGND.n34 122.484
R123 VGND.n13 VGND.n12 111.975
R124 VGND.n10 VGND.n8 111.975
R125 VGND.n56 VGND.n55 59.678
R126 VGND.n55 VGND.t17 57.2313
R127 VGND.n55 VGND.t15 57.2313
R128 VGND.n47 VGND.n37 34.6358
R129 VGND.n43 VGND.n37 34.6358
R130 VGND.n43 VGND.n42 34.6358
R131 VGND.n42 VGND.n41 34.6358
R132 VGND.n50 VGND.n49 34.6358
R133 VGND.n54 VGND.n53 34.6358
R134 VGND.n30 VGND.n1 34.6358
R135 VGND.n31 VGND.n30 34.6358
R136 VGND.n25 VGND.n24 34.6358
R137 VGND.n21 VGND.n20 34.6358
R138 VGND.n18 VGND.n6 34.6358
R139 VGND.n14 VGND.n11 34.6358
R140 VGND.n12 VGND.t27 33.2313
R141 VGND.n26 VGND.n1 30.8711
R142 VGND.n34 VGND.t19 25.8467
R143 VGND.n34 VGND.t13 25.8467
R144 VGND.n5 VGND.t5 25.8467
R145 VGND.n5 VGND.t7 25.8467
R146 VGND.n12 VGND.t9 25.8467
R147 VGND.n8 VGND.t21 25.8467
R148 VGND.n8 VGND.t23 25.8467
R149 VGND.n41 VGND.n39 23.7181
R150 VGND.n61 VGND.n31 23.7181
R151 VGND.n26 VGND.n25 13.5534
R152 VGND.n53 VGND.n35 10.9181
R153 VGND.n10 VGND.n9 10.7918
R154 VGND.n50 VGND.n35 9.41227
R155 VGND.n24 VGND.n3 9.41227
R156 VGND.n14 VGND.n13 9.41227
R157 VGND VGND.n61 9.34738
R158 VGND VGND.n39 9.32654
R159 VGND.n11 VGND.n7 9.3005
R160 VGND.n15 VGND.n14 9.3005
R161 VGND.n16 VGND.n6 9.3005
R162 VGND.n18 VGND.n17 9.3005
R163 VGND.n20 VGND.n4 9.3005
R164 VGND.n22 VGND.n21 9.3005
R165 VGND.n24 VGND.n23 9.3005
R166 VGND.n25 VGND.n2 9.3005
R167 VGND.n27 VGND.n26 9.3005
R168 VGND.n28 VGND.n1 9.3005
R169 VGND.n30 VGND.n29 9.3005
R170 VGND.n31 VGND.n0 9.3005
R171 VGND.n54 VGND.n33 9.3005
R172 VGND.n53 VGND.n52 9.3005
R173 VGND.n51 VGND.n50 9.3005
R174 VGND.n49 VGND.n36 9.3005
R175 VGND.n47 VGND.n46 9.3005
R176 VGND.n45 VGND.n37 9.3005
R177 VGND.n44 VGND.n43 9.3005
R178 VGND.n42 VGND.n38 9.3005
R179 VGND.n41 VGND.n40 9.3005
R180 VGND.n48 VGND.n47 8.65932
R181 VGND.n57 VGND.n56 7.22
R182 VGND.n49 VGND.n48 6.4005
R183 VGND.n56 VGND.n54 5.64756
R184 VGND.n11 VGND.n10 5.64756
R185 VGND.n20 VGND.n19 4.89462
R186 VGND.n19 VGND.n18 4.89462
R187 VGND.n9 VGND.n7 1.07033
R188 VGND.n21 VGND.n3 0.376971
R189 VGND.n13 VGND.n6 0.376971
R190 VGND.n57 VGND.n33 0.155698
R191 VGND.n15 VGND.n7 0.120292
R192 VGND.n16 VGND.n15 0.120292
R193 VGND.n17 VGND.n16 0.120292
R194 VGND.n17 VGND.n4 0.120292
R195 VGND.n22 VGND.n4 0.120292
R196 VGND.n23 VGND.n22 0.120292
R197 VGND.n23 VGND.n2 0.120292
R198 VGND.n27 VGND.n2 0.120292
R199 VGND.n28 VGND.n27 0.120292
R200 VGND.n29 VGND.n28 0.120292
R201 VGND.n29 VGND.n0 0.120292
R202 VGND.n52 VGND.n33 0.120292
R203 VGND.n52 VGND.n51 0.120292
R204 VGND.n51 VGND.n36 0.120292
R205 VGND.n46 VGND.n36 0.120292
R206 VGND.n46 VGND.n45 0.120292
R207 VGND.n45 VGND.n44 0.120292
R208 VGND.n44 VGND.n38 0.120292
R209 VGND.n40 VGND.n38 0.120292
R210 VGND.n40 VGND 0.09425
R211 VGND VGND.n0 0.0734167
R212 a_505_297.t1 a_505_297.n5 742.867
R213 a_505_297.t1 a_505_297.n6 724.692
R214 a_505_297.n5 a_505_297.n4 311.748
R215 a_505_297.n6 a_505_297.t0 287.401
R216 a_505_297.n0 a_505_297.t2 266.707
R217 a_505_297.n3 a_505_297.t3 137.474
R218 a_505_297.n1 a_505_297.n0 133.353
R219 a_505_297.n0 a_505_297.t5 128.534
R220 a_505_297.n2 a_505_297.t4 117.287
R221 a_505_297.n3 a_505_297.n2 60.56
R222 a_505_297.n4 a_505_297.n1 19.2805
R223 a_505_297.n6 a_505_297.n5 18.1338
R224 a_505_297.n2 a_505_297.n1 14.0588
R225 a_505_297.n4 a_505_297.n3 4.94459
R226 VPWRIN.n0 VPWRIN.t0 1565.73
R227 VPWRIN.n0 VPWRIN.t1 370.75
R228 VPWRIN VPWRIN.n0 7.13856
C0 VPWRIN VPWR 0.911213f
C1 A X 0.002945f
C2 VPB A 0.019925f
C3 VPWRIN A 0.089133f
C4 VPB X 0.010944f
C5 VPWRIN X 0.055055f
C6 VPWR A 0.004863f
C7 VPWR X 0.296526f
C8 VPB VPWRIN 0.104184f
C9 VPB VPWR 0.614628f
C10 X VGND 0.348782f
C11 A VGND 0.654476f
C12 VPWR VGND 0.320315f
C13 VPWRIN VGND 0.718335f
C14 VPB VGND 1.76838f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 VPWR VGND LOWLVPWR A X VPB VNB
X0 a_1032_911.t0 a_620_911.t5 VPWR.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VPWR.t0 a_1032_911.t2 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2 VGND A.t0 a_714_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VGND.t0 a_505_297.t2 a_620_911.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X4 X.t2 a_1032_911.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.154625 ps=1.325 w=1 l=0.15
X5 VGND A.t1 a_714_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_620_911.t1 a_505_297.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_714_47.t1 A.t2 VGND VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 X.t7 a_1032_911.t4 VGND VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.104 ps=0.97 w=0.65 l=0.15
X9 VGND a_1032_911.t5 X.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X10 a_714_47.t0 A.t3 VGND VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X11 VPWR.t2 a_1032_911.t6 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12 VGND a_1032_911.t7 X.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12025 ps=1.02 w=0.65 l=0.15
X13 a_1032_911.t1 a_620_911.t6 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X14 VGND.t12 a_505_297.t4 a_620_911.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_505_297.t0 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X16 VPWR.t6 a_714_47.t5 a_620_911.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.154625 pd=1.325 as=0.21725 ps=2.13 w=0.79 l=0.15
X17 X.t4 a_1032_911.t8 VGND VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VPWR.t5 a_620_911.t7 a_714_47.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X19 X.t0 a_1032_911.t9 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_505_297.t1 A.t5 VGND VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X21 a_620_911.t4 a_505_297.t5 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t2 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t0 25.8467
R14 a_620_911.n1 a_620_911.t4 25.8467
R15 a_620_911.n0 a_620_911.t3 25.8467
R16 a_620_911.n0 a_620_911.t1 25.8467
R17 VPWR.n2 VPWR.t0 416.128
R18 VPWR.n3 VPWR.n1 332.486
R19 VPWR.n7 VPWR.n6 326.825
R20 VPWR.n7 VPWR.n5 325.817
R21 VPWR.n5 VPWR.t4 38.6524
R22 VPWR.n6 VPWR.t1 38.4132
R23 VPWR.n5 VPWR.t5 37.4056
R24 VPWR.n6 VPWR.t6 37.4056
R25 VPWR.n8 VPWR.n4 34.6358
R26 VPWR.n1 VPWR.t3 27.5805
R27 VPWR.n1 VPWR.t2 27.5805
R28 VPWR.n3 VPWR.n2 23.1308
R29 VPWR.n4 VPWR.n3 18.0711
R30 VPWR.n8 VPWR.n7 12.8005
R31 VPWR.n4 VPWR.n0 9.3005
R32 VPWR.n9 VPWR.n8 9.3005
R33 VPWR VPWR.n9 1.38004
R34 VPWR.n2 VPWR.n0 1.16591
R35 VPWR.n9 VPWR.n0 0.120292
R36 a_1032_911.n6 a_1032_911.n5 472.841
R37 a_1032_911.n4 a_1032_911.t2 461.113
R38 a_1032_911.t0 a_1032_911.n6 376.678
R39 a_1032_911.n4 a_1032_911.t9 322.94
R40 a_1032_911.n5 a_1032_911.t6 322.94
R41 a_1032_911.n2 a_1032_911.t9 184.768
R42 a_1032_911.n1 a_1032_911.t6 184.768
R43 a_1032_911.n0 a_1032_911.t3 184.768
R44 a_1032_911.t2 a_1032_911.n3 184.768
R45 a_1032_911.n3 a_1032_911.t5 168.701
R46 a_1032_911.n2 a_1032_911.t8 168.701
R47 a_1032_911.n1 a_1032_911.t7 168.701
R48 a_1032_911.n0 a_1032_911.t4 168.701
R49 a_1032_911.n6 a_1032_911.t1 144.809
R50 a_1032_911.n5 a_1032_911.n4 138.173
R51 a_1032_911.n1 a_1032_911.n0 77.1205
R52 a_1032_911.n3 a_1032_911.n2 63.7728
R53 a_1032_911.n2 a_1032_911.n1 63.7728
R54 VPB VPB.t0 290.572
R55 VPB VPB.t2 161.095
R56 VPB.t2 VPB.t1 9.03378
R57 X.n6 X.n0 314.94
R58 X.n5 X.n3 314.938
R59 X.n5 X.n4 117.287
R60 X X.n1 104.951
R61 X.n0 X.t1 45.3105
R62 X.n1 X.t5 42.462
R63 X.n6 X.n5 36.2343
R64 X.n3 X.t3 27.5805
R65 X.n3 X.t0 27.5805
R66 X.n0 X.t2 27.5805
R67 X.n1 X.t7 25.8467
R68 X.n4 X.t6 25.8467
R69 X.n4 X.t4 25.8467
R70 X.n6 X.n2 4.88777
R71 X X.n6 3.25868
R72 X.n6 X 2.36358
R73 X.n2 X 0.465955
R74 X.n2 X 0.427167
R75 A.n0 A.t0 302.053
R76 A.n3 A.t4 268.313
R77 A.n3 A.t5 165.989
R78 A.n1 A.t1 163.881
R79 A.n0 A.t2 163.881
R80 A.n2 A.t3 163.881
R81 A.n4 A.n3 156.262
R82 A A.n4 154.452
R83 A.n1 A.n0 138.173
R84 A.n2 A.n1 136.774
R85 A.n4 A.n2 87.8489
R86 a_714_47.n0 a_714_47.t4 481.457
R87 a_714_47.n0 a_714_47.t5 446.346
R88 a_714_47.n3 a_714_47.n2 121.251
R89 a_714_47.n2 a_714_47.n1 117.666
R90 a_714_47.n2 a_714_47.n0 95.4968
R91 a_714_47.n1 a_714_47.t2 25.8467
R92 a_714_47.n1 a_714_47.t0 25.8467
R93 a_714_47.t3 a_714_47.n3 25.8467
R94 a_714_47.n3 a_714_47.t1 25.8467
R95 VGND.n8 VGND.t1 154.561
R96 VGND.n2 VGND.n1 122.484
R97 VGND.n4 VGND.n3 63.931
R98 VGND.n3 VGND.t7 57.2313
R99 VGND.n3 VGND.t0 57.2313
R100 VGND.n7 VGND.n6 34.6358
R101 VGND.n1 VGND.t13 25.8467
R102 VGND.n1 VGND.t12 25.8467
R103 VGND.n4 VGND.n2 17.8707
R104 VGND.n9 VGND.n8 16.26
R105 VGND.n6 VGND.n2 9.41227
R106 VGND.n6 VGND.n5 9.3005
R107 VGND.n7 VGND.n0 9.3005
R108 VGND.n8 VGND.n7 6.4005
R109 VGND.n5 VGND.n4 0.720832
R110 VGND VGND.n9 0.54977
R111 VGND.n9 VGND.n0 0.147176
R112 VGND.n5 VGND.n0 0.120292
R113 VNB.n2 VNB.t2 13151
R114 VNB.n1 VNB.n0 9804.72
R115 VNB.n2 VNB.t1 4955.34
R116 VNB VNB.n2 3445.95
R117 VNB.t3 VNB.t2 2947.57
R118 VNB.t0 VNB.t7 2192.88
R119 VNB.t11 VNB.t9 1480.91
R120 VNB.t6 VNB.t11 1338.51
R121 VNB.t8 VNB.t10 1224.6
R122 VNB.t9 VNB.t8 1224.6
R123 VNB.t4 VNB.t6 1224.6
R124 VNB.t5 VNB.t4 1224.6
R125 VNB.t13 VNB.t0 1224.6
R126 VNB.t1 VNB.t12 1224.6
R127 VNB.n0 VNB.t5 882.848
R128 VNB.n1 VNB.t13 768.933
R129 VNB.t12 VNB.n1 455.663
R130 VNB.n0 VNB.t3 341.748
R131 a_505_297.t0 a_505_297.n5 742.867
R132 a_505_297.t0 a_505_297.n6 724.692
R133 a_505_297.n5 a_505_297.n4 311.748
R134 a_505_297.n6 a_505_297.t1 287.401
R135 a_505_297.n0 a_505_297.t2 266.707
R136 a_505_297.n3 a_505_297.t3 137.474
R137 a_505_297.n1 a_505_297.n0 133.353
R138 a_505_297.n0 a_505_297.t5 128.534
R139 a_505_297.n2 a_505_297.t4 117.287
R140 a_505_297.n3 a_505_297.n2 60.56
R141 a_505_297.n4 a_505_297.n1 19.2805
R142 a_505_297.n6 a_505_297.n5 18.1338
R143 a_505_297.n2 a_505_297.n1 14.0588
R144 a_505_297.n4 a_505_297.n3 4.94459
R145 LOWLVPWR.n0 LOWLVPWR.t0 1565.73
R146 LOWLVPWR.n0 LOWLVPWR.t1 370.75
R147 LOWLVPWR LOWLVPWR.n0 7.13856
C0 A X 0.002945f
C1 w_n38_261# A 9.27e-19
C2 LOWLVPWR VPB 0.01111f
C3 A VGND 0.112132f
C4 LOWLVPWR VPWR 0.921436f
C5 VPB VPWR 0.103956f
C6 LOWLVPWR X 0.055055f
C7 w_n38_261# LOWLVPWR 0.023199f
C8 VPB X 0.010944f
C9 LOWLVPWR VGND 0.212277f
C10 VPWR X 0.296526f
C11 VPB VGND 0.034255f
C12 w_n38_261# VPWR 0.040297f
C13 LOWLVPWR A 0.089133f
C14 VPWR VGND 0.217594f
C15 VPB A 0.018862f
C16 VPWR A 0.004863f
C17 X VGND 0.311381f
C18 w_n38_261# VGND 0.018561f
C19 VGND VNB 1.982388f
C20 X VNB 0.037401f
C21 A VNB 0.54227f
C22 VPWR VNB 0.301369f
C23 VPB VNB 1.07144f
C24 LOWLVPWR VNB 0.520657f
C25 w_n38_261# VNB 0.285264f $ **FLOATING
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 VPWR VPB VGND LOWLVPWR A X
X0 a_1028_32.t1 a_620_911.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VGND.t15 A.t0 a_714_58.t3 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND.t1 a_505_297.t2 a_620_911.t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X3 X.t0 a_1028_32.t2 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND.t13 A.t1 a_714_58.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_620_911.t2 a_505_297.t3 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_714_58.t0 A.t2 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_714_58.t1 A.t3 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X8 a_1028_32.t0 a_620_911.t6 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X9 VGND.t5 a_505_297.t4 a_620_911.t3 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 a_505_297.t0 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X11 VPWR.t1 a_714_58.t5 a_620_911.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1185 pd=1.09 as=0.21725 ps=2.13 w=0.79 l=0.15
X12 X.t1 a_1028_32.t3 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.21725 pd=2.13 as=0.1185 ps=1.09 w=0.79 l=0.15
X13 VPWR.t3 a_620_911.t7 a_714_58.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X14 a_505_297.t1 A.t5 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X15 a_620_911.t4 a_505_297.t5 VGND.t21 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t1 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t0 25.8467
R14 a_620_911.n1 a_620_911.t4 25.8467
R15 a_620_911.n0 a_620_911.t3 25.8467
R16 a_620_911.n0 a_620_911.t2 25.8467
R17 VPWR.n2 VPWR.n1 326.825
R18 VPWR.n2 VPWR.n0 325.817
R19 VPWR.n0 VPWR.t2 38.6524
R20 VPWR.n0 VPWR.t3 37.4056
R21 VPWR.n1 VPWR.t0 37.4056
R22 VPWR.n1 VPWR.t1 37.4056
R23 VPWR VPWR.n2 21.8082
R24 a_1028_32.n1 a_1028_32.n0 780.957
R25 a_1028_32.t1 a_1028_32.n1 376.678
R26 a_1028_32.n0 a_1028_32.t2 195.912
R27 a_1028_32.n1 a_1028_32.t0 144.809
R28 a_1028_32.n0 a_1028_32.t3 59.9423
R29 VPB VPB.t2 463.961
R30 VPB.t1 VPB.t0 151.06
R31 VPB.t2 VPB.t1 1.67895
R32 A.n0 A.t0 284.38
R33 A.n3 A.t4 268.313
R34 A.n3 A.t5 165.989
R35 A.n4 A.n3 156.262
R36 A A.n4 154.452
R37 A.n1 A.t1 146.208
R38 A.n0 A.t2 146.208
R39 A.n2 A.t3 146.208
R40 A.n1 A.n0 138.173
R41 A.n2 A.n1 136.774
R42 A.n4 A.n2 87.8489
R43 a_714_58.t4 a_714_58.n3 481.457
R44 a_714_58.n3 a_714_58.t5 446.346
R45 a_714_58.n2 a_714_58.n0 120.412
R46 a_714_58.n2 a_714_58.n1 116.829
R47 a_714_58.n3 a_714_58.n2 95.4968
R48 a_714_58.n1 a_714_58.t2 25.8467
R49 a_714_58.n1 a_714_58.t1 25.8467
R50 a_714_58.n0 a_714_58.t3 25.8467
R51 a_714_58.n0 a_714_58.t0 25.8467
R52 VGND.n54 VGND.n2 9804.72
R53 VGND.n53 VGND.n52 9804.72
R54 VGND.t2 VGND.n2 4955.34
R55 VGND.n55 VGND.n54 4202.78
R56 VGND.n33 VGND.n2 4202.78
R57 VGND.t18 VGND.n51 3839.97
R58 VGND.t16 VGND.n26 3469.08
R59 VGND.n54 VGND.t6 3346.28
R60 VGND.t6 VGND.t10 2947.57
R61 VGND.t0 VGND.t18 2192.88
R62 VGND.t14 VGND.t16 1224.6
R63 VGND.t8 VGND.t14 1224.6
R64 VGND.t12 VGND.t8 1224.6
R65 VGND.t20 VGND.t0 1224.6
R66 VGND.t4 VGND.t2 1224.6
R67 VGND.n53 VGND.t12 882.848
R68 VGND.n52 VGND.t20 768.933
R69 VGND.n52 VGND.t4 455.663
R70 VGND.t10 VGND.n53 341.748
R71 VGND.n14 VGND.t7 249.048
R72 VGND.n22 VGND.n21 203.424
R73 VGND.n42 VGND.t3 154.561
R74 VGND.n8 VGND.t11 139.954
R75 VGND.n29 VGND.n28 122.484
R76 VGND.n4 VGND.n3 114.109
R77 VGND.n50 VGND.n49 59.678
R78 VGND.n49 VGND.t19 57.2313
R79 VGND.n49 VGND.t1 57.2313
R80 VGND.n41 VGND.n31 34.6358
R81 VGND.n37 VGND.n31 34.6358
R82 VGND.n37 VGND.n36 34.6358
R83 VGND.n36 VGND.n35 34.6358
R84 VGND.n44 VGND.n43 34.6358
R85 VGND.n48 VGND.n47 34.6358
R86 VGND.n10 VGND.n9 34.6358
R87 VGND.n10 VGND.n1 34.6358
R88 VGND.n16 VGND.n15 34.6358
R89 VGND.n20 VGND.n6 34.6358
R90 VGND.n24 VGND.n23 34.6358
R91 VGND.n14 VGND.n9 30.8711
R92 VGND.n28 VGND.t21 25.8467
R93 VGND.n28 VGND.t5 25.8467
R94 VGND.n21 VGND.t9 25.8467
R95 VGND.n21 VGND.t13 25.8467
R96 VGND.n3 VGND.t17 25.8467
R97 VGND.n3 VGND.t15 25.8467
R98 VGND.n35 VGND.n33 23.7181
R99 VGND.n55 VGND.n1 23.7181
R100 VGND.n26 VGND.n4 16.2466
R101 VGND.n15 VGND.n14 13.5534
R102 VGND.n47 VGND.n29 10.9181
R103 VGND.n44 VGND.n29 9.41227
R104 VGND.n16 VGND.n8 9.41227
R105 VGND VGND.n55 9.34738
R106 VGND VGND.n33 9.32654
R107 VGND.n12 VGND.n9 9.3005
R108 VGND.n11 VGND.n10 9.3005
R109 VGND.n1 VGND.n0 9.3005
R110 VGND.n14 VGND.n13 9.3005
R111 VGND.n17 VGND.n16 9.3005
R112 VGND.n15 VGND.n7 9.3005
R113 VGND.n20 VGND.n19 9.3005
R114 VGND.n18 VGND.n6 9.3005
R115 VGND.n25 VGND.n24 9.3005
R116 VGND.n23 VGND.n5 9.3005
R117 VGND.n48 VGND.n27 9.3005
R118 VGND.n47 VGND.n46 9.3005
R119 VGND.n45 VGND.n44 9.3005
R120 VGND.n43 VGND.n30 9.3005
R121 VGND.n41 VGND.n40 9.3005
R122 VGND.n39 VGND.n31 9.3005
R123 VGND.n38 VGND.n37 9.3005
R124 VGND.n36 VGND.n32 9.3005
R125 VGND.n35 VGND.n34 9.3005
R126 VGND.n42 VGND.n41 8.65932
R127 VGND.n51 VGND.n50 7.05995
R128 VGND.n43 VGND.n42 6.4005
R129 VGND.n50 VGND.n48 5.64756
R130 VGND.n22 VGND.n20 4.89462
R131 VGND.n23 VGND.n22 4.89462
R132 VGND.n26 VGND.n25 0.878118
R133 VGND.n8 VGND.n6 0.376971
R134 VGND.n24 VGND.n4 0.376971
R135 VGND.n51 VGND.n27 0.314038
R136 VGND.n25 VGND.n5 0.120292
R137 VGND.n19 VGND.n5 0.120292
R138 VGND.n19 VGND.n18 0.120292
R139 VGND.n18 VGND.n17 0.120292
R140 VGND.n17 VGND.n7 0.120292
R141 VGND.n13 VGND.n7 0.120292
R142 VGND.n13 VGND.n12 0.120292
R143 VGND.n12 VGND.n11 0.120292
R144 VGND.n11 VGND.n0 0.120292
R145 VGND.n46 VGND.n27 0.120292
R146 VGND.n46 VGND.n45 0.120292
R147 VGND.n45 VGND.n30 0.120292
R148 VGND.n40 VGND.n30 0.120292
R149 VGND.n40 VGND.n39 0.120292
R150 VGND.n39 VGND.n38 0.120292
R151 VGND.n38 VGND.n32 0.120292
R152 VGND.n34 VGND.n32 0.120292
R153 VGND.n34 VGND 0.09425
R154 VGND VGND.n0 0.0734167
R155 a_505_297.t0 a_505_297.n5 742.867
R156 a_505_297.t0 a_505_297.n6 724.692
R157 a_505_297.n5 a_505_297.n4 311.748
R158 a_505_297.n6 a_505_297.t1 287.401
R159 a_505_297.n0 a_505_297.t2 266.707
R160 a_505_297.n3 a_505_297.t3 137.474
R161 a_505_297.n1 a_505_297.n0 133.353
R162 a_505_297.n0 a_505_297.t5 128.534
R163 a_505_297.n2 a_505_297.t4 117.287
R164 a_505_297.n3 a_505_297.n2 60.56
R165 a_505_297.n4 a_505_297.n1 19.2805
R166 a_505_297.n6 a_505_297.n5 18.1338
R167 a_505_297.n2 a_505_297.n1 14.0588
R168 a_505_297.n4 a_505_297.n3 4.94459
R169 X X.t1 391.517
R170 X X.t0 128.451
R171 X.n0 X 16.7569
R172 X X.n0 0.465955
R173 X.n0 X 0.427167
R174 LOWLVPWR.n0 LOWLVPWR.t0 1565.73
R175 LOWLVPWR.n0 LOWLVPWR.t1 370.75
R176 LOWLVPWR LOWLVPWR.n0 7.13856
C0 X VPWR 0.073906f
C1 X A 0.002926f
C2 VPB LOWLVPWR 0.106224f
C3 VPB VPWR 0.528032f
C4 VPB A 0.019913f
C5 LOWLVPWR VPWR 0.771396f
C6 LOWLVPWR A 0.089133f
C7 X VPB 0.021096f
C8 VPWR A 0.004863f
C9 X LOWLVPWR 0.026094f
C10 X VGND 0.179867f
C11 A VGND 0.636418f
C12 VPWR VGND 0.267901f
C13 LOWLVPWR VGND 0.691791f
C14 VPB VGND 1.44754f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 VPWR VPB VGND LOWLVPWR A X
X0 a_1032_911.t1 a_620_911.t5 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VGND.t23 A.t0 a_714_47.t4 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND.t7 a_505_297.t2 a_620_911.t4 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X3 X.t3 a_1032_911.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.154625 ps=1.325 w=1 l=0.15
X4 VGND.t21 A.t1 a_714_47.t3 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_620_911.t1 a_505_297.t3 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_714_47.t2 A.t2 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 X.t1 a_1032_911.t3 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_714_47.t1 A.t3 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X9 VPWR.t2 a_1032_911.t4 X.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.185 ps=1.37 w=1 l=0.15
X10 VGND.t9 a_1032_911.t5 X.t0 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.12025 ps=1.02 w=0.65 l=0.15
X11 a_1032_911.t0 a_620_911.t6 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X12 VGND.t3 a_505_297.t4 a_620_911.t2 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_505_297.t1 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X14 VPWR.t0 a_714_47.t5 a_620_911.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.154625 pd=1.325 as=0.21725 ps=2.13 w=0.79 l=0.15
X15 VPWR.t4 a_620_911.t7 a_714_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X16 a_505_297.t0 A.t5 VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X17 a_620_911.t3 a_505_297.t5 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t0 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t4 25.8467
R14 a_620_911.n1 a_620_911.t3 25.8467
R15 a_620_911.n0 a_620_911.t2 25.8467
R16 a_620_911.n0 a_620_911.t1 25.8467
R17 VPWR.n3 VPWR.t2 416.57
R18 VPWR.n2 VPWR.n1 326.825
R19 VPWR.n2 VPWR.n0 325.817
R20 VPWR.n0 VPWR.t3 38.6524
R21 VPWR.n1 VPWR.t1 38.4132
R22 VPWR.n0 VPWR.t4 37.4056
R23 VPWR.n1 VPWR.t0 37.4056
R24 VPWR.n3 VPWR.n2 19.5934
R25 VPWR VPWR.n3 2.21634
R26 a_1032_911.n2 a_1032_911.t4 843.981
R27 a_1032_911.t1 a_1032_911.n2 376.678
R28 a_1032_911.n0 a_1032_911.t2 184.768
R29 a_1032_911.t4 a_1032_911.n1 184.768
R30 a_1032_911.n1 a_1032_911.t5 168.701
R31 a_1032_911.n0 a_1032_911.t3 168.701
R32 a_1032_911.n2 a_1032_911.t0 144.809
R33 a_1032_911.n1 a_1032_911.n0 77.1205
R34 VPB.n0 VPB.t1 550.726
R35 VPB VPB.n0 206.38
R36 VPB.n0 VPB.t2 39.4319
R37 VPB.t1 VPB.t0 11.9753
R38 A.n0 A.t0 302.053
R39 A.n3 A.t4 268.313
R40 A.n3 A.t5 165.989
R41 A.n1 A.t1 163.881
R42 A.n0 A.t2 163.881
R43 A.n2 A.t3 163.881
R44 A.n4 A.n3 156.262
R45 A A.n4 154.452
R46 A.n1 A.n0 138.173
R47 A.n2 A.n1 136.774
R48 A.n4 A.n2 87.8489
R49 a_714_47.t0 a_714_47.n3 481.457
R50 a_714_47.n3 a_714_47.t5 446.346
R51 a_714_47.n2 a_714_47.n0 121.251
R52 a_714_47.n2 a_714_47.n1 117.666
R53 a_714_47.n3 a_714_47.n2 95.4968
R54 a_714_47.n1 a_714_47.t3 25.8467
R55 a_714_47.n1 a_714_47.t1 25.8467
R56 a_714_47.n0 a_714_47.t4 25.8467
R57 a_714_47.n0 a_714_47.t2 25.8467
R58 VGND.n54 VGND.n26 9804.72
R59 VGND.n53 VGND.n52 9804.72
R60 VGND.t0 VGND.n26 4955.34
R61 VGND.t12 VGND.n51 4409.49
R62 VGND.n55 VGND.n54 4202.78
R63 VGND.n33 VGND.n26 4202.78
R64 VGND.n54 VGND.t14 3346.28
R65 VGND.t14 VGND.t16 2947.57
R66 VGND.t6 VGND.t12 2192.88
R67 VGND.t10 VGND.t8 1480.91
R68 VGND.t22 VGND.t10 1338.51
R69 VGND.t18 VGND.t22 1224.6
R70 VGND.t20 VGND.t18 1224.6
R71 VGND.t4 VGND.t6 1224.6
R72 VGND.t2 VGND.t0 1224.6
R73 VGND.n53 VGND.t20 882.848
R74 VGND.n52 VGND.t4 768.933
R75 VGND.n52 VGND.t2 455.663
R76 VGND.t16 VGND.n53 341.748
R77 VGND.n20 VGND.t15 249.048
R78 VGND.n13 VGND.n5 201.292
R79 VGND.n42 VGND.t1 154.561
R80 VGND.n9 VGND.t9 143.803
R81 VGND.n3 VGND.t17 137.821
R82 VGND.n29 VGND.n28 122.484
R83 VGND.n8 VGND.n7 111.975
R84 VGND.n50 VGND.n49 59.678
R85 VGND.n49 VGND.t13 57.2313
R86 VGND.n49 VGND.t7 57.2313
R87 VGND.n41 VGND.n31 34.6358
R88 VGND.n37 VGND.n31 34.6358
R89 VGND.n37 VGND.n36 34.6358
R90 VGND.n36 VGND.n35 34.6358
R91 VGND.n44 VGND.n43 34.6358
R92 VGND.n48 VGND.n47 34.6358
R93 VGND.n24 VGND.n1 34.6358
R94 VGND.n25 VGND.n24 34.6358
R95 VGND.n19 VGND.n18 34.6358
R96 VGND.n15 VGND.n14 34.6358
R97 VGND.n12 VGND.n6 34.6358
R98 VGND.n7 VGND.t11 33.2313
R99 VGND.n20 VGND.n1 30.8711
R100 VGND.n28 VGND.t5 25.8467
R101 VGND.n28 VGND.t3 25.8467
R102 VGND.n5 VGND.t19 25.8467
R103 VGND.n5 VGND.t21 25.8467
R104 VGND.n7 VGND.t23 25.8467
R105 VGND.n35 VGND.n33 23.7181
R106 VGND.n55 VGND.n25 23.7181
R107 VGND.n9 VGND.n8 16.1542
R108 VGND.n20 VGND.n19 13.5534
R109 VGND.n47 VGND.n29 10.9181
R110 VGND.n44 VGND.n29 9.41227
R111 VGND.n18 VGND.n3 9.41227
R112 VGND VGND.n55 9.34738
R113 VGND VGND.n33 9.32654
R114 VGND.n10 VGND.n6 9.3005
R115 VGND.n12 VGND.n11 9.3005
R116 VGND.n14 VGND.n4 9.3005
R117 VGND.n16 VGND.n15 9.3005
R118 VGND.n18 VGND.n17 9.3005
R119 VGND.n19 VGND.n2 9.3005
R120 VGND.n21 VGND.n20 9.3005
R121 VGND.n22 VGND.n1 9.3005
R122 VGND.n24 VGND.n23 9.3005
R123 VGND.n25 VGND.n0 9.3005
R124 VGND.n48 VGND.n27 9.3005
R125 VGND.n47 VGND.n46 9.3005
R126 VGND.n45 VGND.n44 9.3005
R127 VGND.n43 VGND.n30 9.3005
R128 VGND.n41 VGND.n40 9.3005
R129 VGND.n39 VGND.n31 9.3005
R130 VGND.n38 VGND.n37 9.3005
R131 VGND.n36 VGND.n32 9.3005
R132 VGND.n35 VGND.n34 9.3005
R133 VGND.n42 VGND.n41 8.65932
R134 VGND.n51 VGND.n50 7.14073
R135 VGND.n43 VGND.n42 6.4005
R136 VGND.n50 VGND.n48 5.64756
R137 VGND.n14 VGND.n13 4.89462
R138 VGND.n13 VGND.n12 4.89462
R139 VGND.n10 VGND.n9 0.960602
R140 VGND.n15 VGND.n3 0.376971
R141 VGND.n8 VGND.n6 0.376971
R142 VGND.n51 VGND.n27 0.234391
R143 VGND.n11 VGND.n10 0.120292
R144 VGND.n11 VGND.n4 0.120292
R145 VGND.n16 VGND.n4 0.120292
R146 VGND.n17 VGND.n16 0.120292
R147 VGND.n17 VGND.n2 0.120292
R148 VGND.n21 VGND.n2 0.120292
R149 VGND.n22 VGND.n21 0.120292
R150 VGND.n23 VGND.n22 0.120292
R151 VGND.n23 VGND.n0 0.120292
R152 VGND.n46 VGND.n27 0.120292
R153 VGND.n46 VGND.n45 0.120292
R154 VGND.n45 VGND.n30 0.120292
R155 VGND.n40 VGND.n30 0.120292
R156 VGND.n40 VGND.n39 0.120292
R157 VGND.n39 VGND.n38 0.120292
R158 VGND.n38 VGND.n32 0.120292
R159 VGND.n34 VGND.n32 0.120292
R160 VGND.n34 VGND 0.09425
R161 VGND VGND.n0 0.0734167
R162 a_505_297.t1 a_505_297.n5 742.867
R163 a_505_297.t1 a_505_297.n6 724.692
R164 a_505_297.n5 a_505_297.n4 311.748
R165 a_505_297.n6 a_505_297.t0 287.401
R166 a_505_297.n0 a_505_297.t2 266.707
R167 a_505_297.n3 a_505_297.t3 137.474
R168 a_505_297.n1 a_505_297.n0 133.353
R169 a_505_297.n0 a_505_297.t5 128.534
R170 a_505_297.n2 a_505_297.t4 117.287
R171 a_505_297.n3 a_505_297.n2 60.56
R172 a_505_297.n4 a_505_297.n1 19.2805
R173 a_505_297.n6 a_505_297.n5 18.1338
R174 a_505_297.n2 a_505_297.n1 14.0588
R175 a_505_297.n4 a_505_297.n3 4.94459
R176 X X.n1 318.197
R177 X X.n0 104.951
R178 X.n1 X.t2 45.3105
R179 X.n0 X.t0 42.462
R180 X.n1 X.t3 27.5805
R181 X.n0 X.t1 25.8467
R182 X.n2 X 16.7569
R183 X X.n2 0.465955
R184 X.n2 X 0.427167
R185 LOWLVPWR.n0 LOWLVPWR.t0 1565.73
R186 LOWLVPWR.n0 LOWLVPWR.t1 370.75
R187 LOWLVPWR LOWLVPWR.n0 7.13856
C0 VPB X 0.008022f
C1 VPB LOWLVPWR 0.103298f
C2 LOWLVPWR X 0.026823f
C3 VPB VPWR 0.534275f
C4 VPWR X 0.129496f
C5 LOWLVPWR VPWR 0.805258f
C6 VPB A 0.019925f
C7 A X 0.00292f
C8 LOWLVPWR A 0.089133f
C9 VPWR A 0.004863f
C10 X VGND 0.178135f
C11 A VGND 0.654458f
C12 VPWR VGND 0.29254f
C13 LOWLVPWR VGND 0.696853f
C14 VPB VGND 1.45906f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 VPWR VPB VGND LOWLVPWR A X
X0 a_1032_911.t0 a_620_911.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2133 pd=2.12 as=0.120475 ps=1.095 w=0.79 l=0.15
X1 VPWR.t3 a_1032_911.t2 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2 VGND.t17 A.t0 a_714_47.t3 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VGND.t7 a_505_297.t2 a_620_911.t3 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X4 X.t2 a_1032_911.t3 VPWR.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.154625 ps=1.325 w=1 l=0.15
X5 VGND.t15 A.t1 a_714_47.t2 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_620_911.t1 a_505_297.t3 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_714_47.t1 A.t2 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 X.t7 a_1032_911.t4 VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.104 ps=0.97 w=0.65 l=0.15
X9 VGND.t23 a_1032_911.t5 X.t6 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X10 a_714_47.t4 A.t3 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X11 VPWR.t5 a_1032_911.t6 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12 VGND.t21 a_1032_911.t7 X.t5 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12025 ps=1.02 w=0.65 l=0.15
X13 a_1032_911.t1 a_620_911.t6 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.2015 ps=1.27 w=0.65 l=0.15
X14 VGND.t5 a_505_297.t4 a_620_911.t2 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_505_297.t1 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.275 ps=2.55 w=1 l=0.15
X16 VPWR.t0 a_714_47.t5 a_620_911.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.154625 pd=1.325 as=0.21725 ps=2.13 w=0.79 l=0.15
X17 X.t4 a_1032_911.t8 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VPWR.t2 a_620_911.t7 a_714_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.120475 pd=1.095 as=0.21725 ps=2.13 w=0.79 l=0.15
X19 X.t0 a_1032_911.t9 VPWR.t6 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_505_297.t0 A.t5 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X21 a_620_911.t4 a_505_297.t5 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_620_911.t0 a_620_911.n7 617.596
R1 a_620_911.n6 a_620_911.t5 297.233
R2 a_620_911.n5 a_620_911.t6 244.214
R3 a_620_911.t5 a_620_911.n5 204.048
R4 a_620_911.n7 a_620_911.n6 192.363
R5 a_620_911.n4 a_620_911.n3 174.105
R6 a_620_911.n3 a_620_911.n2 169.738
R7 a_620_911.n2 a_620_911.n0 160.78
R8 a_620_911.n4 a_620_911.t7 155.847
R9 a_620_911.n6 a_620_911.t7 151.028
R10 a_620_911.n7 a_620_911.n3 122.692
R11 a_620_911.n2 a_620_911.n1 120.874
R12 a_620_911.n5 a_620_911.n4 98.0072
R13 a_620_911.n1 a_620_911.t3 25.8467
R14 a_620_911.n1 a_620_911.t4 25.8467
R15 a_620_911.n0 a_620_911.t2 25.8467
R16 a_620_911.n0 a_620_911.t1 25.8467
R17 VPWR.n2 VPWR.t3 416.128
R18 VPWR.n3 VPWR.n1 332.486
R19 VPWR.n7 VPWR.n6 326.825
R20 VPWR.n7 VPWR.n5 325.817
R21 VPWR.n5 VPWR.t1 38.6524
R22 VPWR.n6 VPWR.t4 38.4132
R23 VPWR.n5 VPWR.t2 37.4056
R24 VPWR.n6 VPWR.t0 37.4056
R25 VPWR.n8 VPWR.n4 34.6358
R26 VPWR.n1 VPWR.t6 27.5805
R27 VPWR.n1 VPWR.t5 27.5805
R28 VPWR.n3 VPWR.n2 23.1308
R29 VPWR.n4 VPWR.n3 18.0711
R30 VPWR.n8 VPWR.n7 12.8005
R31 VPWR.n4 VPWR.n0 9.3005
R32 VPWR.n9 VPWR.n8 9.3005
R33 VPWR VPWR.n9 1.38004
R34 VPWR.n2 VPWR.n0 1.16591
R35 VPWR.n9 VPWR.n0 0.120292
R36 a_1032_911.n6 a_1032_911.n5 472.841
R37 a_1032_911.n4 a_1032_911.t2 461.113
R38 a_1032_911.t0 a_1032_911.n6 376.678
R39 a_1032_911.n4 a_1032_911.t9 322.94
R40 a_1032_911.n5 a_1032_911.t6 322.94
R41 a_1032_911.n2 a_1032_911.t9 184.768
R42 a_1032_911.n1 a_1032_911.t6 184.768
R43 a_1032_911.n0 a_1032_911.t3 184.768
R44 a_1032_911.t2 a_1032_911.n3 184.768
R45 a_1032_911.n3 a_1032_911.t5 168.701
R46 a_1032_911.n2 a_1032_911.t8 168.701
R47 a_1032_911.n1 a_1032_911.t7 168.701
R48 a_1032_911.n0 a_1032_911.t4 168.701
R49 a_1032_911.n6 a_1032_911.t1 144.809
R50 a_1032_911.n5 a_1032_911.n4 138.173
R51 a_1032_911.n1 a_1032_911.n0 77.1205
R52 a_1032_911.n3 a_1032_911.n2 63.7728
R53 a_1032_911.n2 a_1032_911.n1 63.7728
R54 VPB.n0 VPB.t2 416.839
R55 VPB VPB.n0 206.714
R56 VPB.n0 VPB.t1 29.6401
R57 VPB.t2 VPB.t0 9.03378
R58 X.n6 X.n0 314.94
R59 X.n5 X.n3 314.938
R60 X.n5 X.n4 117.287
R61 X X.n1 104.951
R62 X.n0 X.t1 45.3105
R63 X.n1 X.t5 42.462
R64 X.n6 X.n5 36.2343
R65 X.n3 X.t3 27.5805
R66 X.n3 X.t0 27.5805
R67 X.n0 X.t2 27.5805
R68 X.n1 X.t7 25.8467
R69 X.n4 X.t6 25.8467
R70 X.n4 X.t4 25.8467
R71 X.n6 X.n2 4.88777
R72 X X.n6 3.25868
R73 X.n6 X 2.36358
R74 X.n2 X 0.465955
R75 X.n2 X 0.427167
R76 A.n0 A.t0 302.053
R77 A.n3 A.t4 268.313
R78 A.n3 A.t5 165.989
R79 A.n1 A.t1 163.881
R80 A.n0 A.t2 163.881
R81 A.n2 A.t3 163.881
R82 A.n4 A.n3 156.262
R83 A A.n4 154.452
R84 A.n1 A.n0 138.173
R85 A.n2 A.n1 136.774
R86 A.n4 A.n2 87.8489
R87 a_714_47.t0 a_714_47.n3 481.457
R88 a_714_47.n3 a_714_47.t5 446.346
R89 a_714_47.n2 a_714_47.n0 121.251
R90 a_714_47.n2 a_714_47.n1 117.666
R91 a_714_47.n3 a_714_47.n2 95.4968
R92 a_714_47.n1 a_714_47.t2 25.8467
R93 a_714_47.n1 a_714_47.t4 25.8467
R94 a_714_47.n0 a_714_47.t3 25.8467
R95 a_714_47.n0 a_714_47.t1 25.8467
R96 VGND.n60 VGND.n32 9804.72
R97 VGND.n59 VGND.n58 9804.72
R98 VGND.t0 VGND.n57 7029.87
R99 VGND.t2 VGND.n32 4955.34
R100 VGND.n61 VGND.n60 4202.78
R101 VGND.n39 VGND.n32 4202.78
R102 VGND.n60 VGND.t8 3346.28
R103 VGND.t8 VGND.t10 2947.57
R104 VGND.t6 VGND.t0 2192.88
R105 VGND.t24 VGND.t20 1480.91
R106 VGND.t16 VGND.t24 1338.51
R107 VGND.t18 VGND.t22 1224.6
R108 VGND.t20 VGND.t18 1224.6
R109 VGND.t12 VGND.t16 1224.6
R110 VGND.t14 VGND.t12 1224.6
R111 VGND.t26 VGND.t6 1224.6
R112 VGND.t4 VGND.t2 1224.6
R113 VGND.n59 VGND.t14 882.848
R114 VGND.n58 VGND.t26 768.933
R115 VGND.n58 VGND.t4 455.663
R116 VGND.t10 VGND.n59 341.748
R117 VGND.n26 VGND.t9 249.048
R118 VGND.n19 VGND.n5 201.292
R119 VGND.n48 VGND.t3 154.561
R120 VGND.n9 VGND.t23 151.21
R121 VGND.n3 VGND.t11 137.821
R122 VGND.n35 VGND.n34 122.484
R123 VGND.n13 VGND.n12 111.975
R124 VGND.n10 VGND.n8 111.975
R125 VGND.n56 VGND.n55 59.678
R126 VGND.n55 VGND.t1 57.2313
R127 VGND.n55 VGND.t7 57.2313
R128 VGND.n47 VGND.n37 34.6358
R129 VGND.n43 VGND.n37 34.6358
R130 VGND.n43 VGND.n42 34.6358
R131 VGND.n42 VGND.n41 34.6358
R132 VGND.n50 VGND.n49 34.6358
R133 VGND.n54 VGND.n53 34.6358
R134 VGND.n30 VGND.n1 34.6358
R135 VGND.n31 VGND.n30 34.6358
R136 VGND.n25 VGND.n24 34.6358
R137 VGND.n21 VGND.n20 34.6358
R138 VGND.n18 VGND.n6 34.6358
R139 VGND.n14 VGND.n11 34.6358
R140 VGND.n12 VGND.t25 33.2313
R141 VGND.n26 VGND.n1 30.8711
R142 VGND.n34 VGND.t27 25.8467
R143 VGND.n34 VGND.t5 25.8467
R144 VGND.n5 VGND.t13 25.8467
R145 VGND.n5 VGND.t15 25.8467
R146 VGND.n12 VGND.t17 25.8467
R147 VGND.n8 VGND.t19 25.8467
R148 VGND.n8 VGND.t21 25.8467
R149 VGND.n41 VGND.n39 23.7181
R150 VGND.n61 VGND.n31 23.7181
R151 VGND.n26 VGND.n25 13.5534
R152 VGND.n53 VGND.n35 10.9181
R153 VGND.n10 VGND.n9 10.7918
R154 VGND.n50 VGND.n35 9.41227
R155 VGND.n24 VGND.n3 9.41227
R156 VGND.n14 VGND.n13 9.41227
R157 VGND VGND.n61 9.34738
R158 VGND VGND.n39 9.32654
R159 VGND.n11 VGND.n7 9.3005
R160 VGND.n15 VGND.n14 9.3005
R161 VGND.n16 VGND.n6 9.3005
R162 VGND.n18 VGND.n17 9.3005
R163 VGND.n20 VGND.n4 9.3005
R164 VGND.n22 VGND.n21 9.3005
R165 VGND.n24 VGND.n23 9.3005
R166 VGND.n25 VGND.n2 9.3005
R167 VGND.n27 VGND.n26 9.3005
R168 VGND.n28 VGND.n1 9.3005
R169 VGND.n30 VGND.n29 9.3005
R170 VGND.n31 VGND.n0 9.3005
R171 VGND.n54 VGND.n33 9.3005
R172 VGND.n53 VGND.n52 9.3005
R173 VGND.n51 VGND.n50 9.3005
R174 VGND.n49 VGND.n36 9.3005
R175 VGND.n47 VGND.n46 9.3005
R176 VGND.n45 VGND.n37 9.3005
R177 VGND.n44 VGND.n43 9.3005
R178 VGND.n42 VGND.n38 9.3005
R179 VGND.n41 VGND.n40 9.3005
R180 VGND.n48 VGND.n47 8.65932
R181 VGND.n57 VGND.n56 7.22
R182 VGND.n49 VGND.n48 6.4005
R183 VGND.n56 VGND.n54 5.64756
R184 VGND.n11 VGND.n10 5.64756
R185 VGND.n20 VGND.n19 4.89462
R186 VGND.n19 VGND.n18 4.89462
R187 VGND.n9 VGND.n7 1.07033
R188 VGND.n21 VGND.n3 0.376971
R189 VGND.n13 VGND.n6 0.376971
R190 VGND.n57 VGND.n33 0.155698
R191 VGND.n15 VGND.n7 0.120292
R192 VGND.n16 VGND.n15 0.120292
R193 VGND.n17 VGND.n16 0.120292
R194 VGND.n17 VGND.n4 0.120292
R195 VGND.n22 VGND.n4 0.120292
R196 VGND.n23 VGND.n22 0.120292
R197 VGND.n23 VGND.n2 0.120292
R198 VGND.n27 VGND.n2 0.120292
R199 VGND.n28 VGND.n27 0.120292
R200 VGND.n29 VGND.n28 0.120292
R201 VGND.n29 VGND.n0 0.120292
R202 VGND.n52 VGND.n33 0.120292
R203 VGND.n52 VGND.n51 0.120292
R204 VGND.n51 VGND.n36 0.120292
R205 VGND.n46 VGND.n36 0.120292
R206 VGND.n46 VGND.n45 0.120292
R207 VGND.n45 VGND.n44 0.120292
R208 VGND.n44 VGND.n38 0.120292
R209 VGND.n40 VGND.n38 0.120292
R210 VGND.n40 VGND 0.09425
R211 VGND VGND.n0 0.0734167
R212 a_505_297.t1 a_505_297.n5 742.867
R213 a_505_297.t1 a_505_297.n6 724.692
R214 a_505_297.n5 a_505_297.n4 311.748
R215 a_505_297.n6 a_505_297.t0 287.401
R216 a_505_297.n0 a_505_297.t2 266.707
R217 a_505_297.n3 a_505_297.t3 137.474
R218 a_505_297.n1 a_505_297.n0 133.353
R219 a_505_297.n0 a_505_297.t5 128.534
R220 a_505_297.n2 a_505_297.t4 117.287
R221 a_505_297.n3 a_505_297.n2 60.56
R222 a_505_297.n4 a_505_297.n1 19.2805
R223 a_505_297.n6 a_505_297.n5 18.1338
R224 a_505_297.n2 a_505_297.n1 14.0588
R225 a_505_297.n4 a_505_297.n3 4.94459
R226 LOWLVPWR.n0 LOWLVPWR.t0 1565.73
R227 LOWLVPWR.n0 LOWLVPWR.t1 370.75
R228 LOWLVPWR LOWLVPWR.n0 7.13856
C0 VPB LOWLVPWR 0.104184f
C1 VPB VPWR 0.614628f
C2 VPB A 0.019925f
C3 LOWLVPWR VPWR 0.911213f
C4 VPB X 0.010944f
C5 LOWLVPWR A 0.089133f
C6 VPWR A 0.004863f
C7 LOWLVPWR X 0.055055f
C8 VPWR X 0.296526f
C9 A X 0.002945f
C10 X VGND 0.348782f
C11 A VGND 0.654476f
C12 VPWR VGND 0.320315f
C13 LOWLVPWR VGND 0.718335f
C14 VPB VGND 1.76838f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y.t3 B.t0 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t1 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t0 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 A.t1 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t5 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND.t0 B.t2 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t3 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297.t1 B.t3 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t0 212.081
R2 B B.n2 182.081
R3 B.n0 B.t2 139.78
R4 B.n1 B.t1 139.78
R5 B.n2 B.n0 30.6732
R6 B.n2 B.n1 30.6732
R7 a_27_297.n0 a_27_297.t1 404.502
R8 a_27_297.n0 a_27_297.t3 301.301
R9 a_27_297.n1 a_27_297.n0 184.905
R10 a_27_297.n1 a_27_297.t2 26.5955
R11 a_27_297.t0 a_27_297.n1 26.5955
R12 Y Y.n0 591.788
R13 Y.n4 Y.n0 585
R14 Y.n3 Y.n1 135.249
R15 Y.n3 Y.n2 98.982
R16 Y.n4 Y.n3 74.7314
R17 Y.n0 Y.t2 26.5955
R18 Y.n0 Y.t3 26.5955
R19 Y.n2 Y.t0 24.9236
R20 Y.n2 Y.t1 24.9236
R21 Y.n1 Y.t4 24.9236
R22 Y.n1 Y.t5 24.9236
R23 Y Y.n4 6.4005
R24 VPB.t2 VPB.t1 248.599
R25 VPB.t0 VPB.t2 248.599
R26 VPB.t3 VPB.t0 248.599
R27 VPB VPB.t3 201.246
R28 VGND.n2 VGND.t0 287.377
R29 VGND.n3 VGND.n1 207.965
R30 VGND.n5 VGND.t3 150.922
R31 VGND.n4 VGND.n3 32.377
R32 VGND.n1 VGND.t1 24.9236
R33 VGND.n1 VGND.t2 24.9236
R34 VGND.n5 VGND.n4 24.4711
R35 VGND.n3 VGND.n2 9.43392
R36 VGND.n6 VGND.n5 9.3005
R37 VGND.n4 VGND.n0 9.3005
R38 VGND.n2 VGND.n0 0.554787
R39 VGND.n6 VGND.n0 0.120292
R40 VGND VGND.n6 0.0213333
R41 VNB.t1 VNB.t0 1196.12
R42 VNB.t2 VNB.t1 1196.12
R43 VNB.t3 VNB.t2 1196.12
R44 VNB VNB.t3 968.285
R45 A.n0 A.t0 212.081
R46 A.n1 A.t3 212.081
R47 A A.n2 183.68
R48 A.n0 A.t1 139.78
R49 A.n1 A.t2 139.78
R50 A.n2 A.n0 38.7066
R51 A.n2 A.n1 22.6399
R52 VPWR VPWR.n0 316.39
R53 VPWR.n0 VPWR.t1 26.5955
R54 VPWR.n0 VPWR.t0 26.5955
C0 VPB A 0.056273f
C1 VPB B 0.056648f
C2 Y VPB 0.009606f
C3 A B 0.071165f
C4 VPB VPWR 0.049962f
C5 VGND VPB 0.006128f
C6 Y A 0.052333f
C7 A VPWR 0.041833f
C8 VGND A 0.059727f
C9 Y B 0.179365f
C10 B VPWR 0.017427f
C11 Y VPWR 0.012692f
C12 VGND B 0.029406f
C13 Y VGND 0.289148f
C14 VGND VPWR 0.046681f
C15 VGND VNB 0.342832f
C16 Y VNB 0.064071f
C17 VPWR VNB 0.248551f
C18 B VNB 0.197736f
C19 A VNB 0.206739f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR.t3 A.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t4 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 B.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47.t1 B.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47.t3 A.t2 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t2 A.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t0 B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t1 B.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n1 A.t1 212.081
R2 A A.n2 152.94
R3 A.n0 A.t2 139.78
R4 A.n1 A.t3 139.78
R5 A.n2 A.n0 30.6732
R6 A.n2 A.n1 30.6732
R7 Y.n3 Y.n1 243.68
R8 Y.n4 Y.n0 206.249
R9 Y.n3 Y.n2 205.28
R10 Y.n1 Y.t1 26.5955
R11 Y.n1 Y.t0 26.5955
R12 Y.n2 Y.t3 26.5955
R13 Y.n2 Y.t4 26.5955
R14 Y Y.n3 24.9955
R15 Y.n0 Y.t5 24.9236
R16 Y.n0 Y.t2 24.9236
R17 Y.n4 Y 14.8576
R18 Y Y.n4 0.686214
R19 VPWR.n2 VPWR.t3 348.959
R20 VPWR.n3 VPWR.n1 320.976
R21 VPWR.n5 VPWR.t0 249.362
R22 VPWR.n4 VPWR.n3 30.8711
R23 VPWR.n1 VPWR.t2 26.5955
R24 VPWR.n1 VPWR.t1 26.5955
R25 VPWR.n5 VPWR.n4 25.977
R26 VPWR.n3 VPWR.n2 10.9193
R27 VPWR.n4 VPWR.n0 9.3005
R28 VPWR.n6 VPWR.n5 9.3005
R29 VPWR.n2 VPWR.n0 0.572285
R30 VPWR.n6 VPWR.n0 0.120292
R31 VPWR VPWR.n6 0.0213333
R32 VPB.t2 VPB.t3 248.599
R33 VPB.t1 VPB.t2 248.599
R34 VPB.t0 VPB.t1 248.599
R35 VPB VPB.t0 189.409
R36 B.n0 B.t0 212.081
R37 B.n1 B.t2 212.081
R38 B B.n2 155.584
R39 B.n0 B.t1 139.78
R40 B.n1 B.t3 139.78
R41 B.n2 B.n0 30.6732
R42 B.n2 B.n1 30.6732
R43 VGND VGND.n0 214.335
R44 VGND.n0 VGND.t0 24.9236
R45 VGND.n0 VGND.t1 24.9236
R46 a_27_47.n0 a_27_47.t3 322.56
R47 a_27_47.n0 a_27_47.t0 188.529
R48 a_27_47.n1 a_27_47.n0 88.3446
R49 a_27_47.n1 a_27_47.t2 24.9236
R50 a_27_47.t1 a_27_47.n1 24.9236
R51 VNB.t2 VNB.t3 1196.12
R52 VNB.t1 VNB.t2 1196.12
R53 VNB.t0 VNB.t1 1196.12
R54 VNB VNB.t0 911.327
C0 Y VGND 0.020763f
C1 VPB VPWR 0.066372f
C2 VPB Y 0.015949f
C3 B VPWR 0.059991f
C4 B Y 0.062045f
C5 A VPWR 0.031531f
C6 VPB VGND 0.005765f
C7 A Y 0.177649f
C8 B VGND 0.02902f
C9 A VGND 0.017966f
C10 VPB B 0.056795f
C11 VPB A 0.057111f
C12 VPWR Y 0.398191f
C13 B A 0.074816f
C14 VPWR VGND 0.047614f
C15 VGND VNB 0.295829f
C16 Y VNB 0.062962f
C17 VPWR VNB 0.309019f
C18 A VNB 0.197653f
C19 B VNB 0.209169f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__conb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
X0 VPWR.t0 HI.t0 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO.t0 VGND.t0 sky130_fd_pr__res_generic_po w=0.48 l=0.045
R0 VPWR VPWR.t0 188.507
R1 HI HI.t0 144.478
R2 LO LO.t0 178.194
R3 VGND VGND.t0 156.286
C0 LO VGND 0.060475f
C1 VPB VGND 0.004789f
C2 HI LO 0.068275f
C3 HI VPB 0.004729f
C4 VGND VPWR 0.031746f
C5 HI VPWR 0.072643f
C6 HI VGND 0.206798f
C7 LO VPB 0.133883f
C8 LO VPWR 0.240897f
C9 VPB VPWR 0.157853f
C10 VGND VNB 0.405957f
C11 LO VNB 0.165803f
C12 HI VNB 0.249567f
C13 VPWR VNB 0.297091f
C14 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__macro_sparecell.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B a_27_47#
X0 VPWR.t1 A.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t2 B.t0 Y.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47.t3 B.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47.t1 A.t2 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t2 A.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t5 B.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t0 B.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n1 A.t1 212.081
R2 A A.n2 152.94
R3 A.n0 A.t2 139.78
R4 A.n1 A.t3 139.78
R5 A.n2 A.n0 30.6732
R6 A.n2 A.n1 30.6732
R7 Y.n3 Y.n1 243.68
R8 Y.n4 Y.n0 206.249
R9 Y.n3 Y.n2 205.28
R10 Y.n1 Y.t4 26.5955
R11 Y.n1 Y.t5 26.5955
R12 Y.n2 Y.t1 26.5955
R13 Y.n2 Y.t0 26.5955
R14 Y Y.n3 24.9955
R15 Y.n0 Y.t3 24.9236
R16 Y.n0 Y.t2 24.9236
R17 Y.n4 Y 14.8576
R18 Y Y.n4 0.686214
R19 VPWR.n2 VPWR.t1 348.959
R20 VPWR.n3 VPWR.n1 320.976
R21 VPWR.n5 VPWR.t3 249.362
R22 VPWR.n4 VPWR.n3 30.8711
R23 VPWR.n1 VPWR.t0 26.5955
R24 VPWR.n1 VPWR.t2 26.5955
R25 VPWR.n5 VPWR.n4 25.977
R26 VPWR.n3 VPWR.n2 10.9193
R27 VPWR.n4 VPWR.n0 9.3005
R28 VPWR.n6 VPWR.n5 9.3005
R29 VPWR.n2 VPWR.n0 0.572285
R30 VPWR.n6 VPWR.n0 0.120292
R31 VPWR VPWR.n6 0.0213333
R32 VPB.t0 VPB.t1 248.599
R33 VPB.t2 VPB.t0 248.599
R34 VPB.t3 VPB.t2 248.599
R35 VPB VPB.t3 189.409
R36 B.n0 B.t0 212.081
R37 B.n1 B.t2 212.081
R38 B B.n2 155.584
R39 B.n0 B.t1 139.78
R40 B.n1 B.t3 139.78
R41 B.n2 B.n0 30.6732
R42 B.n2 B.n1 30.6732
R43 VGND VGND.n0 214.335
R44 VGND.n0 VGND.t1 24.9236
R45 VGND.n0 VGND.t0 24.9236
R46 a_27_47.t1 a_27_47.n1 322.56
R47 a_27_47.n1 a_27_47.t2 188.529
R48 a_27_47.n1 a_27_47.n0 88.3446
R49 a_27_47.n0 a_27_47.t0 24.9236
R50 a_27_47.n0 a_27_47.t3 24.9236
R51 VNB.t0 VNB.t1 1196.12
R52 VNB.t3 VNB.t0 1196.12
R53 VNB.t2 VNB.t3 1196.12
R54 VNB VNB.t2 911.327
C0 VPB B 0.056795f
C1 B Y 0.062045f
C2 A VPWR 0.031531f
C3 VPB A 0.057111f
C4 B VGND 0.02902f
C5 A Y 0.177649f
C6 VPB VPWR 0.066372f
C7 VPWR Y 0.398191f
C8 A VGND 0.017966f
C9 VPB Y 0.015949f
C10 VPWR VGND 0.047614f
C11 VPB VGND 0.005765f
C12 Y VGND 0.020763f
C13 B A 0.074816f
C14 B VPWR 0.059991f
C15 VGND VNB 0.295829f
C16 Y VNB 0.062962f
C17 VPWR VNB 0.309019f
C18 A VNB 0.197653f
C19 B VNB 0.209169f
C20 VPB VNB 0.516168f
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y.t2 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t0 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t0 A.t3 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n0 A.t3 212.081
R1 A.n1 A.t0 212.081
R2 A A.n1 189.073
R3 A.n0 A.t1 139.78
R4 A.n1 A.t2 139.78
R5 A.n1 A.n0 61.346
R6 VPWR.n0 VPWR.t0 262.851
R7 VPWR.n0 VPWR.t1 259.721
R8 VPWR VPWR.n0 0.491471
R9 Y.n2 Y.n1 208.965
R10 Y Y.n0 96.8352
R11 Y.n1 Y.t1 26.5955
R12 Y.n1 Y.t2 26.5955
R13 Y.n0 Y.t3 24.9236
R14 Y.n0 Y.t0 24.9236
R15 Y.n3 Y 11.2645
R16 Y Y.n3 6.1445
R17 Y.n3 Y 4.65505
R18 Y Y.n2 2.0485
R19 Y.n2 Y 1.55202
R20 VPB.t1 VPB.t0 248.599
R21 VPB VPB.t1 198.287
R22 VGND.n0 VGND.t1 169.418
R23 VGND.n0 VGND.t0 166.787
R24 VGND VGND.n0 0.491471
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 954.045
C0 Y VPB 0.006097f
C1 Y VPWR 0.209105f
C2 Y VGND 0.154601f
C3 VPB VPWR 0.052063f
C4 VPB VGND 0.006491f
C5 A Y 0.089386f
C6 VPWR VGND 0.042274f
C7 A VPB 0.074183f
C8 A VPWR 0.06305f
C9 A VGND 0.063754f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A a_27_297#
X0 Y.t4 B.t0 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t2 B.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t3 A.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t0 A.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t1 A.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND.t2 B.t2 Y.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t3 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297.t1 B.t3 Y.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t0 212.081
R2 B B.n2 182.081
R3 B.n0 B.t2 139.78
R4 B.n1 B.t1 139.78
R5 B.n2 B.n0 30.6732
R6 B.n2 B.n1 30.6732
R7 a_27_297.n1 a_27_297.t1 404.502
R8 a_27_297.t0 a_27_297.n1 301.301
R9 a_27_297.n1 a_27_297.n0 184.905
R10 a_27_297.n0 a_27_297.t2 26.5955
R11 a_27_297.n0 a_27_297.t3 26.5955
R12 Y Y.n0 591.788
R13 Y.n4 Y.n0 585
R14 Y.n3 Y.n1 135.249
R15 Y.n3 Y.n2 98.982
R16 Y.n4 Y.n3 74.7314
R17 Y.n0 Y.t3 26.5955
R18 Y.n0 Y.t4 26.5955
R19 Y.n2 Y.t5 24.9236
R20 Y.n2 Y.t2 24.9236
R21 Y.n1 Y.t0 24.9236
R22 Y.n1 Y.t1 24.9236
R23 Y Y.n4 6.4005
R24 VPB.t2 VPB.t1 248.599
R25 VPB.t3 VPB.t2 248.599
R26 VPB.t0 VPB.t3 248.599
R27 VPB VPB.t0 201.246
R28 VGND.n2 VGND.t2 287.377
R29 VGND.n3 VGND.n1 207.965
R30 VGND.n5 VGND.t1 150.922
R31 VGND.n4 VGND.n3 32.377
R32 VGND.n1 VGND.t3 24.9236
R33 VGND.n1 VGND.t0 24.9236
R34 VGND.n5 VGND.n4 24.4711
R35 VGND.n3 VGND.n2 9.43392
R36 VGND.n6 VGND.n5 9.3005
R37 VGND.n4 VGND.n0 9.3005
R38 VGND.n2 VGND.n0 0.554787
R39 VGND.n6 VGND.n0 0.120292
R40 VGND VGND.n6 0.0213333
R41 VNB.t3 VNB.t2 1196.12
R42 VNB.t0 VNB.t3 1196.12
R43 VNB.t1 VNB.t0 1196.12
R44 VNB VNB.t1 968.285
R45 A.n0 A.t0 212.081
R46 A.n1 A.t3 212.081
R47 A A.n2 183.68
R48 A.n0 A.t1 139.78
R49 A.n1 A.t2 139.78
R50 A.n2 A.n0 38.7066
R51 A.n2 A.n1 22.6399
R52 VPWR VPWR.n0 316.39
R53 VPWR.n0 VPWR.t1 26.5955
R54 VPWR.n0 VPWR.t0 26.5955
C0 Y VGND 0.289148f
C1 Y VPB 0.009606f
C2 VPWR A 0.041833f
C3 VGND VPB 0.006128f
C4 Y A 0.052333f
C5 VGND A 0.059727f
C6 VPB A 0.056273f
C7 B VPWR 0.017427f
C8 B Y 0.179365f
C9 B VGND 0.029406f
C10 B VPB 0.056648f
C11 VPWR Y 0.012692f
C12 B A 0.071165f
C13 VPWR VGND 0.046681f
C14 VPWR VPB 0.049962f
C15 VGND VNB 0.342832f
C16 Y VNB 0.064071f
C17 VPWR VNB 0.248551f
C18 B VNB 0.197736f
C19 A VNB 0.206739f
C20 VPB VNB 0.516168f
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
X0 VPWR.t0 HI.t0 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO.t0 VGND.t0 sky130_fd_pr__res_generic_po w=0.48 l=0.045
R0 VPWR VPWR.t0 188.507
R1 HI HI.t0 144.478
R2 LO LO.t0 178.194
R3 VGND VGND.t0 156.286
C0 VGND LO 0.060475f
C1 VPB LO 0.133883f
C2 VPWR VGND 0.031746f
C3 VPWR VPB 0.157853f
C4 VPB VGND 0.004789f
C5 HI LO 0.068275f
C6 VPWR HI 0.072643f
C7 HI VGND 0.206798f
C8 VPB HI 0.004729f
C9 VPWR LO 0.240897f
C10 VGND VNB 0.405957f
C11 LO VNB 0.165803f
C12 HI VNB 0.249567f
C13 VPWR VNB 0.297091f
C14 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__macro_sparecell VGND VPWR LO VNB VPB
Xsky130_fd_sc_hd__nand2_2_1 VPB VNB VGND VPWR sky130_fd_sc_hd__nor2_2_1/B LO LO sky130_fd_sc_hd__nand2_2_1/a_27_47#
+ sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nand2_2_0 VPB VNB VGND VPWR sky130_fd_sc_hd__nor2_2_0/B LO LO sky130_fd_sc_hd__nand2_2_0/a_27_47#
+ sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_0 VPB VNB VPWR VGND sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_2_0/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 VPB VNB VPWR VGND sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_2_0 VPB VNB VGND VPWR sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__inv_2_0/A
+ sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor2_2_0/a_27_297# sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_1 VPB VNB VGND VPWR sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__inv_2_1/A
+ sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__nor2_2_1/a_27_297# sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__conb_1_0 LO sky130_fd_sc_hd__conb_1_0/HI VPB VNB VGND VPWR sky130_fd_sc_hd__conb_1
X0 VPWR LO.t8 sky130_fd_sc_hd__nor2_2_0/B VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
X1 sky130_fd_sc_hd__nor2_2_1/B LO.t6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
X2 sky130_fd_sc_hd__nor2_2_0/B LO.t9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
X3 VPWR LO.t10 sky130_fd_sc_hd__nor2_2_0/B VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
X4 sky130_fd_sc_hd__nor2_2_0/B LO.t14 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
X5 VPWR.t0 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
X6 VPWR LO.t2 sky130_fd_sc_hd__nor2_2_1/B VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
X7 sky130_fd_sc_hd__inv_2_1/Y.t2 sky130_fd_sc_hd__inv_2_1/A VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0 l=0
X8 sky130_fd_sc_hd__nor2_2_1/B LO.t1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
X9 VGND.t0 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0 l=0
X10 VPWR LO.t0 sky130_fd_sc_hd__nor2_2_1/B VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
X11 sky130_fd_sc_hd__inv_2_1/Y.t1 sky130_fd_sc_hd__inv_2_1/A VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
R0 LO.n4 LO.t6 212.081
R1 LO.n5 LO.t2 212.081
R2 LO.n0 LO.t1 212.081
R3 LO.n1 LO.t0 212.081
R4 LO.n10 LO.t10 212.081
R5 LO.n11 LO.t14 212.081
R6 LO.n14 LO.t8 212.081
R7 LO.n15 LO.t9 212.081
R8 LO LO.n12 155.584
R9 LO.n7 LO.n6 152
R10 LO.n3 LO.n2 152
R11 LO.n17 LO.n16 152
R12 LO.n4 LO.t7 139.78
R13 LO.n5 LO.t3 139.78
R14 LO.n0 LO.t5 139.78
R15 LO.n1 LO.t4 139.78
R16 LO.n10 LO.t11 139.78
R17 LO.n11 LO.t15 139.78
R18 LO.n14 LO.t12 139.78
R19 LO.n15 LO.t13 139.78
R20 LO.n8 LO.n7 34.3885
R21 LO.n6 LO.n4 30.6732
R22 LO.n6 LO.n5 30.6732
R23 LO.n2 LO.n0 30.6732
R24 LO.n2 LO.n1 30.6732
R25 LO.n12 LO.n10 30.6732
R26 LO.n12 LO.n11 30.6732
R27 LO.n16 LO.n14 30.6732
R28 LO.n16 LO.n15 30.6732
R29 LO.n8 LO.n3 30.5095
R30 LO.n17 LO.n13 25.839
R31 LO.n13 LO 22.6125
R32 LO.n9 LO 15.5774
R33 LO.n3 LO 9.2165
R34 LO.n7 LO 5.1205
R35 LO LO.n8 0.799413
R36 LO.n13 LO.n9 0.667037
R37 LO LO.n17 0.5125
R38 LO.n9 LO 0.0466957
R39 VPWR.n43 VPWR.t0 253.934
R40 VPWR.n41 VPWR.n3 226.355
R41 VPWR.n13 VPWR.n12 38.6948
R42 VPWR.n36 VPWR.n4 34.6358
R43 VPWR.n40 VPWR.n4 34.6358
R44 VPWR.n29 VPWR.n28 34.6358
R45 VPWR.n30 VPWR.n29 34.6358
R46 VPWR.n23 VPWR.n22 34.6358
R47 VPWR.n17 VPWR.n16 34.6358
R48 VPWR.n18 VPWR.n17 34.6358
R49 VPWR.n34 VPWR.n6 31.624
R50 VPWR.n41 VPWR.n40 26.7299
R51 VPWR.n28 VPWR.n8 25.977
R52 VPWR.n18 VPWR.n10 25.977
R53 VPWR.n42 VPWR.n41 25.224
R54 VPWR.n43 VPWR.n42 25.224
R55 VPWR.n3 VPWR.n2 24.6255
R56 VPWR.n3 VPWR.t1 24.6255
R57 VPWR.n24 VPWR.n8 23.7181
R58 VPWR.n22 VPWR.n10 23.7181
R59 VPWR.n35 VPWR.n34 22.9652
R60 VPWR.n36 VPWR.n35 21.4593
R61 VPWR.n30 VPWR.n6 18.4476
R62 VPWR.n16 VPWR.n12 18.4476
R63 VPWR.n24 VPWR.n23 9.78874
R64 VPWR.n14 VPWR.n12 9.3005
R65 VPWR.n16 VPWR.n15 9.3005
R66 VPWR.n17 VPWR.n11 9.3005
R67 VPWR.n19 VPWR.n18 9.3005
R68 VPWR.n20 VPWR.n10 9.3005
R69 VPWR.n22 VPWR.n21 9.3005
R70 VPWR.n23 VPWR.n9 9.3005
R71 VPWR.n25 VPWR.n24 9.3005
R72 VPWR.n26 VPWR.n8 9.3005
R73 VPWR.n28 VPWR.n27 9.3005
R74 VPWR.n29 VPWR.n7 9.3005
R75 VPWR.n31 VPWR.n30 9.3005
R76 VPWR.n32 VPWR.n6 9.3005
R77 VPWR.n34 VPWR.n33 9.3005
R78 VPWR.n35 VPWR.n5 9.3005
R79 VPWR.n37 VPWR.n36 9.3005
R80 VPWR.n38 VPWR.n4 9.3005
R81 VPWR.n40 VPWR.n39 9.3005
R82 VPWR.n41 VPWR.n1 9.3005
R83 VPWR.n42 VPWR.n0 9.3005
R84 VPWR VPWR.n43 9.3005
R85 VPWR.n13 VPWR 0.542919
R86 VPWR.n15 VPWR.n14 0.120292
R87 VPWR.n15 VPWR.n11 0.120292
R88 VPWR.n19 VPWR.n11 0.120292
R89 VPWR.n20 VPWR.n19 0.120292
R90 VPWR.n21 VPWR.n9 0.120292
R91 VPWR.n25 VPWR.n9 0.120292
R92 VPWR.n27 VPWR.n7 0.120292
R93 VPWR.n31 VPWR.n7 0.120292
R94 VPWR.n32 VPWR.n31 0.120292
R95 VPWR.n33 VPWR.n32 0.120292
R96 VPWR.n37 VPWR.n5 0.120292
R97 VPWR.n38 VPWR.n37 0.120292
R98 VPWR.n39 VPWR.n38 0.120292
R99 VPWR.n39 VPWR.n1 0.120292
R100 VPWR VPWR.n0 0.120292
R101 VPWR.n14 VPWR 0.0994583
R102 VPWR.n21 VPWR 0.0994583
R103 VPWR.n26 VPWR 0.0981562
R104 VPWR VPWR.n0 0.0981562
R105 VPWR.n27 VPWR 0.0968542
R106 VPWR VPWR.n5 0.0968542
R107 VPWR VPWR.n13 0.0585447
R108 VPWR VPWR.n26 0.0239375
R109 VPWR.n33 VPWR 0.0239375
R110 VPWR VPWR.n25 0.0226354
R111 VPWR.n1 VPWR 0.0226354
R112 VPWR VPWR.n20 0.0213333
R113 VPB VPB 1361.37
R114 VPB VPB 1361.37
R115 VPB VPB 1358.41
R116 VPB.n0 VPB 958.879
R117 VPB VPB 819.783
R118 VPB VPB 275.235
R119 VPB.n1 VPB.n0 248.599
R120 VPB.t1 VPB.t0 248.599
R121 VPB.t0 VPB 198.287
R122 VPB VPB.n1 150.935
R123 VPB VPB.t1 97.6641
R124 VGND.n2 VGND.n1 460.262
R125 VGND.n42 VGND.t0 164.136
R126 VGND.n40 VGND.t1 161.679
R127 VGND.n13 VGND.n12 34.6358
R128 VGND.n14 VGND.n13 34.6358
R129 VGND.n14 VGND.n8 34.6358
R130 VGND.n18 VGND.n8 34.6358
R131 VGND.n19 VGND.n18 34.6358
R132 VGND.n23 VGND.n7 34.6358
R133 VGND.n24 VGND.n23 34.6358
R134 VGND.n24 VGND.n6 34.6358
R135 VGND.n28 VGND.n6 34.6358
R136 VGND.n29 VGND.n28 34.6358
R137 VGND.n30 VGND.n29 34.6358
R138 VGND.n35 VGND.n34 34.6358
R139 VGND.n36 VGND.n35 34.6358
R140 VGND.n12 VGND.n10 31.2789
R141 VGND.n41 VGND.n40 25.224
R142 VGND.n42 VGND.n41 25.224
R143 VGND.n34 VGND.n4 24.4711
R144 VGND.n30 VGND.n4 24.0946
R145 VGND.n36 VGND.n2 19.9534
R146 VGND.n40 VGND.n2 19.577
R147 VGND VGND.n42 9.3005
R148 VGND.n12 VGND.n11 9.3005
R149 VGND.n13 VGND.n9 9.3005
R150 VGND.n15 VGND.n14 9.3005
R151 VGND.n16 VGND.n8 9.3005
R152 VGND.n18 VGND.n17 9.3005
R153 VGND.n20 VGND.n19 9.3005
R154 VGND.n21 VGND.n7 9.3005
R155 VGND.n23 VGND.n22 9.3005
R156 VGND.n25 VGND.n24 9.3005
R157 VGND.n26 VGND.n6 9.3005
R158 VGND.n28 VGND.n27 9.3005
R159 VGND.n29 VGND.n5 9.3005
R160 VGND.n31 VGND.n30 9.3005
R161 VGND.n32 VGND.n4 9.3005
R162 VGND.n34 VGND.n33 9.3005
R163 VGND.n35 VGND.n3 9.3005
R164 VGND.n37 VGND.n36 9.3005
R165 VGND.n38 VGND.n2 9.3005
R166 VGND.n40 VGND.n39 9.3005
R167 VGND.n41 VGND.n0 9.3005
R168 VGND.n19 VGND.n7 9.03579
R169 VGND.n10 VGND 0.546583
R170 VGND.n11 VGND.n9 0.120292
R171 VGND.n15 VGND.n9 0.120292
R172 VGND.n16 VGND.n15 0.120292
R173 VGND.n17 VGND.n16 0.120292
R174 VGND.n21 VGND.n20 0.120292
R175 VGND.n22 VGND.n21 0.120292
R176 VGND.n27 VGND.n26 0.120292
R177 VGND.n27 VGND.n5 0.120292
R178 VGND.n31 VGND.n5 0.120292
R179 VGND.n32 VGND.n31 0.120292
R180 VGND.n33 VGND.n3 0.120292
R181 VGND.n37 VGND.n3 0.120292
R182 VGND.n38 VGND.n37 0.120292
R183 VGND.n39 VGND.n38 0.120292
R184 VGND VGND.n0 0.120292
R185 VGND.n11 VGND 0.0994583
R186 VGND.n20 VGND 0.0994583
R187 VGND.n25 VGND 0.0981562
R188 VGND VGND.n0 0.0981562
R189 VGND.n26 VGND 0.0968542
R190 VGND.n33 VGND 0.0968542
R191 VGND VGND.n10 0.0547892
R192 VGND VGND.n25 0.0239375
R193 VGND VGND.n32 0.0239375
R194 VGND.n22 VGND 0.0226354
R195 VGND.n39 VGND 0.0226354
R196 VGND.n17 VGND 0.0213333
R197 VNB VNB 6550.16
R198 VNB VNB 6550.16
R199 VNB VNB 6535.92
R200 VNB VNB.n1 4613.59
R201 VNB VNB 3944.34
R202 VNB VNB 1324.27
R203 VNB.n1 VNB.n0 1196.12
R204 VNB.t0 VNB.t1 1196.12
R205 VNB.t1 VNB 954.045
R206 VNB.n0 VNB 726.215
R207 VNB VNB.t0 469.904
R208 sky130_fd_sc_hd__inv_2_1/Y.n3 sky130_fd_sc_hd__inv_2_1/Y.n2 208.965
R209 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/Y.n0 96.8352
R210 sky130_fd_sc_hd__inv_2_1/Y.n2 sky130_fd_sc_hd__inv_2_1/Y.t1 26.5955
R211 sky130_fd_sc_hd__inv_2_1/Y.n2 sky130_fd_sc_hd__inv_2_1/Y.t0 26.5955
R212 sky130_fd_sc_hd__inv_2_1/Y.n0 sky130_fd_sc_hd__inv_2_1/Y.t2 24.9236
R213 sky130_fd_sc_hd__inv_2_1/Y.n0 sky130_fd_sc_hd__inv_2_1/Y.t3 24.9236
R214 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/Y.n1 11.2645
R215 sky130_fd_sc_hd__inv_2_1/Y.n1 sky130_fd_sc_hd__inv_2_1/Y 6.1445
R216 sky130_fd_sc_hd__inv_2_1/Y.n1 sky130_fd_sc_hd__inv_2_1/Y 4.65505
R217 sky130_fd_sc_hd__inv_2_1/Y.n3 sky130_fd_sc_hd__inv_2_1/Y 2.0485
R218 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/Y.n3 1.55202
C0 VPWR sky130_fd_sc_hd__nor2_2_0/B 0.065017f
C1 VGND LO 0.172883f
C2 VPB VPWR 0.011669f
C3 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__conb_1_0/HI 0.004862f
C4 VGND sky130_fd_sc_hd__inv_2_0/A 0.052251f
C5 VPWR sky130_fd_sc_hd__inv_2_0/Y 0.009521f
C6 sky130_fd_sc_hd__nor2_2_1/B LO 0.047282f
C7 sky130_fd_sc_hd__inv_2_1/A VPWR 0.0422f
C8 VPB sky130_fd_sc_hd__inv_2_1/Y 4.5e-20
C9 VGND sky130_fd_sc_hd__nor2_2_0/B 0.100307f
C10 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y 0.041884f
C11 VPB VGND -0.021231f
C12 VGND sky130_fd_sc_hd__inv_2_0/Y 0.011725f
C13 sky130_fd_sc_hd__inv_2_1/A VGND 0.051792f
C14 LO sky130_fd_sc_hd__conb_1_0/HI 0.092406f
C15 VPB sky130_fd_sc_hd__nor2_2_1/B 0.009162f
C16 VPWR sky130_fd_sc_hd__inv_2_1/Y 0.009774f
C17 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__nor2_2_1/B 0.077645f
C18 LO sky130_fd_sc_hd__inv_2_0/A 1.48e-19
C19 VPWR VGND -0.206828f
C20 sky130_fd_sc_hd__conb_1_0/HI sky130_fd_sc_hd__nor2_2_0/B 3.14e-19
C21 LO sky130_fd_sc_hd__nor2_2_0/B 0.057418f
C22 VPB sky130_fd_sc_hd__conb_1_0/HI 0.001622f
C23 sky130_fd_sc_hd__inv_2_1/Y VGND 0.011876f
C24 VPB LO 0.047615f
C25 VPWR sky130_fd_sc_hd__nor2_2_1/B 0.069576f
C26 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__inv_2_0/A 0.07692f
C27 LO sky130_fd_sc_hd__inv_2_0/Y 9.36e-20
C28 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__conb_1_0/HI 3.74e-19
C29 VPB sky130_fd_sc_hd__inv_2_0/A 0.006695f
C30 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_2_0/Y 0.041494f
C31 VPB sky130_fd_sc_hd__nor2_2_0/B 0.009178f
C32 VGND sky130_fd_sc_hd__nor2_2_1/B 0.099905f
C33 VPWR sky130_fd_sc_hd__conb_1_0/HI 0.017264f
C34 VPWR LO 0.252659f
C35 VPB sky130_fd_sc_hd__inv_2_0/Y 4.5e-20
C36 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__conb_1_0/HI 6.02e-20
C37 VPB sky130_fd_sc_hd__inv_2_1/A 0.006695f
C38 VPWR sky130_fd_sc_hd__inv_2_0/A 0.042174f
C39 VGND sky130_fd_sc_hd__conb_1_0/HI -9.95e-19
C40 sky130_fd_sc_hd__conb_1_0/HI VNB 0.249567f
C41 sky130_fd_sc_hd__nor2_2_1/B VNB 0.384454f
C42 sky130_fd_sc_hd__nor2_2_0/B VNB 0.384527f
C43 VGND VNB 1.697799f
C44 sky130_fd_sc_hd__inv_2_1/Y VNB 0.027809f
C45 VPWR VNB 1.287016f
C46 sky130_fd_sc_hd__inv_2_1/A VNB 0.25725f
C47 VPB VNB 2.642472f
C48 sky130_fd_sc_hd__inv_2_0/Y VNB 0.027809f
C49 sky130_fd_sc_hd__inv_2_0/A VNB 0.257245f
C50 LO VNB 0.777712f
.ends

* NGSPICE file created from sky130_fd_sc_hd__conb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
X0 VPWR.t0 HI.t0 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO.t0 VGND.t0 sky130_fd_pr__res_generic_po w=0.48 l=0.045
R0 VPWR VPWR.t0 188.507
R1 HI HI.t0 144.478
R2 LO LO.t0 178.194
R3 VGND VGND.t0 156.286
C0 LO VGND 0.060475f
C1 VPB VGND 0.004789f
C2 HI LO 0.068275f
C3 HI VPB 0.004729f
C4 VGND VPWR 0.031746f
C5 HI VPWR 0.072643f
C6 HI VGND 0.206798f
C7 LO VPB 0.133883f
C8 LO VPWR 0.240897f
C9 VPB VPWR 0.157853f
C10 VGND VNB 0.405957f
C11 LO VNB 0.165803f
C12 HI VNB 0.249567f
C13 VPWR VNB 0.297091f
C14 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR.t3 A.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t4 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 B.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47.t1 B.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47.t3 A.t2 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t2 A.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t0 B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t1 B.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n1 A.t1 212.081
R2 A A.n2 152.94
R3 A.n0 A.t2 139.78
R4 A.n1 A.t3 139.78
R5 A.n2 A.n0 30.6732
R6 A.n2 A.n1 30.6732
R7 Y.n3 Y.n1 243.68
R8 Y.n4 Y.n0 206.249
R9 Y.n3 Y.n2 205.28
R10 Y.n1 Y.t1 26.5955
R11 Y.n1 Y.t0 26.5955
R12 Y.n2 Y.t3 26.5955
R13 Y.n2 Y.t4 26.5955
R14 Y Y.n3 24.9955
R15 Y.n0 Y.t5 24.9236
R16 Y.n0 Y.t2 24.9236
R17 Y.n4 Y 14.8576
R18 Y Y.n4 0.686214
R19 VPWR.n2 VPWR.t3 348.959
R20 VPWR.n3 VPWR.n1 320.976
R21 VPWR.n5 VPWR.t0 249.362
R22 VPWR.n4 VPWR.n3 30.8711
R23 VPWR.n1 VPWR.t2 26.5955
R24 VPWR.n1 VPWR.t1 26.5955
R25 VPWR.n5 VPWR.n4 25.977
R26 VPWR.n3 VPWR.n2 10.9193
R27 VPWR.n4 VPWR.n0 9.3005
R28 VPWR.n6 VPWR.n5 9.3005
R29 VPWR.n2 VPWR.n0 0.572285
R30 VPWR.n6 VPWR.n0 0.120292
R31 VPWR VPWR.n6 0.0213333
R32 VPB.t2 VPB.t3 248.599
R33 VPB.t1 VPB.t2 248.599
R34 VPB.t0 VPB.t1 248.599
R35 VPB VPB.t0 189.409
R36 B.n0 B.t0 212.081
R37 B.n1 B.t2 212.081
R38 B B.n2 155.584
R39 B.n0 B.t1 139.78
R40 B.n1 B.t3 139.78
R41 B.n2 B.n0 30.6732
R42 B.n2 B.n1 30.6732
R43 VGND VGND.n0 214.335
R44 VGND.n0 VGND.t0 24.9236
R45 VGND.n0 VGND.t1 24.9236
R46 a_27_47.n0 a_27_47.t3 322.56
R47 a_27_47.n0 a_27_47.t0 188.529
R48 a_27_47.n1 a_27_47.n0 88.3446
R49 a_27_47.n1 a_27_47.t2 24.9236
R50 a_27_47.t1 a_27_47.n1 24.9236
R51 VNB.t2 VNB.t3 1196.12
R52 VNB.t1 VNB.t2 1196.12
R53 VNB.t0 VNB.t1 1196.12
R54 VNB VNB.t0 911.327
C0 Y VGND 0.020763f
C1 VPB VPWR 0.066372f
C2 VPB Y 0.015949f
C3 B VPWR 0.059991f
C4 B Y 0.062045f
C5 A VPWR 0.031531f
C6 VPB VGND 0.005765f
C7 A Y 0.177649f
C8 B VGND 0.02902f
C9 A VGND 0.017966f
C10 VPB B 0.056795f
C11 VPB A 0.057111f
C12 VPWR Y 0.398191f
C13 B A 0.074816f
C14 VPWR VGND 0.047614f
C15 VGND VNB 0.295829f
C16 Y VNB 0.062962f
C17 VPWR VNB 0.309019f
C18 A VNB 0.197653f
C19 B VNB 0.209169f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR.t3 A.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t4 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 B.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47.t1 B.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47.t3 A.t2 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t2 A.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t0 B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t1 B.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n1 A.t1 212.081
R2 A A.n2 152.94
R3 A.n0 A.t2 139.78
R4 A.n1 A.t3 139.78
R5 A.n2 A.n0 30.6732
R6 A.n2 A.n1 30.6732
R7 Y.n3 Y.n1 243.68
R8 Y.n4 Y.n0 206.249
R9 Y.n3 Y.n2 205.28
R10 Y.n1 Y.t1 26.5955
R11 Y.n1 Y.t0 26.5955
R12 Y.n2 Y.t3 26.5955
R13 Y.n2 Y.t4 26.5955
R14 Y Y.n3 24.9955
R15 Y.n0 Y.t5 24.9236
R16 Y.n0 Y.t2 24.9236
R17 Y.n4 Y 14.8576
R18 Y Y.n4 0.686214
R19 VPWR.n2 VPWR.t3 348.959
R20 VPWR.n3 VPWR.n1 320.976
R21 VPWR.n5 VPWR.t0 249.362
R22 VPWR.n4 VPWR.n3 30.8711
R23 VPWR.n1 VPWR.t2 26.5955
R24 VPWR.n1 VPWR.t1 26.5955
R25 VPWR.n5 VPWR.n4 25.977
R26 VPWR.n3 VPWR.n2 10.9193
R27 VPWR.n4 VPWR.n0 9.3005
R28 VPWR.n6 VPWR.n5 9.3005
R29 VPWR.n2 VPWR.n0 0.572285
R30 VPWR.n6 VPWR.n0 0.120292
R31 VPWR VPWR.n6 0.0213333
R32 VPB.t2 VPB.t3 248.599
R33 VPB.t1 VPB.t2 248.599
R34 VPB.t0 VPB.t1 248.599
R35 VPB VPB.t0 189.409
R36 B.n0 B.t0 212.081
R37 B.n1 B.t2 212.081
R38 B B.n2 155.584
R39 B.n0 B.t1 139.78
R40 B.n1 B.t3 139.78
R41 B.n2 B.n0 30.6732
R42 B.n2 B.n1 30.6732
R43 VGND VGND.n0 214.335
R44 VGND.n0 VGND.t0 24.9236
R45 VGND.n0 VGND.t1 24.9236
R46 a_27_47.n0 a_27_47.t3 322.56
R47 a_27_47.n0 a_27_47.t0 188.529
R48 a_27_47.n1 a_27_47.n0 88.3446
R49 a_27_47.n1 a_27_47.t2 24.9236
R50 a_27_47.t1 a_27_47.n1 24.9236
R51 VNB.t2 VNB.t3 1196.12
R52 VNB.t1 VNB.t2 1196.12
R53 VNB.t0 VNB.t1 1196.12
R54 VNB VNB.t0 911.327
C0 Y VGND 0.020763f
C1 VPB VPWR 0.066372f
C2 VPB Y 0.015949f
C3 B VPWR 0.059991f
C4 B Y 0.062045f
C5 A VPWR 0.031531f
C6 VPB VGND 0.005765f
C7 A Y 0.177649f
C8 B VGND 0.02902f
C9 A VGND 0.017966f
C10 VPB B 0.056795f
C11 VPB A 0.057111f
C12 VPWR Y 0.398191f
C13 B A 0.074816f
C14 VPWR VGND 0.047614f
C15 VGND VNB 0.295829f
C16 Y VNB 0.062962f
C17 VPWR VNB 0.309019f
C18 A VNB 0.197653f
C19 B VNB 0.209169f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y.t3 B.t0 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t1 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t0 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 A.t1 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t5 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND.t0 B.t2 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t3 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297.t1 B.t3 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t0 212.081
R2 B B.n2 182.081
R3 B.n0 B.t2 139.78
R4 B.n1 B.t1 139.78
R5 B.n2 B.n0 30.6732
R6 B.n2 B.n1 30.6732
R7 a_27_297.n0 a_27_297.t1 404.502
R8 a_27_297.n0 a_27_297.t3 301.301
R9 a_27_297.n1 a_27_297.n0 184.905
R10 a_27_297.n1 a_27_297.t2 26.5955
R11 a_27_297.t0 a_27_297.n1 26.5955
R12 Y Y.n0 591.788
R13 Y.n4 Y.n0 585
R14 Y.n3 Y.n1 135.249
R15 Y.n3 Y.n2 98.982
R16 Y.n4 Y.n3 74.7314
R17 Y.n0 Y.t2 26.5955
R18 Y.n0 Y.t3 26.5955
R19 Y.n2 Y.t0 24.9236
R20 Y.n2 Y.t1 24.9236
R21 Y.n1 Y.t4 24.9236
R22 Y.n1 Y.t5 24.9236
R23 Y Y.n4 6.4005
R24 VPB.t2 VPB.t1 248.599
R25 VPB.t0 VPB.t2 248.599
R26 VPB.t3 VPB.t0 248.599
R27 VPB VPB.t3 201.246
R28 VGND.n2 VGND.t0 287.377
R29 VGND.n3 VGND.n1 207.965
R30 VGND.n5 VGND.t3 150.922
R31 VGND.n4 VGND.n3 32.377
R32 VGND.n1 VGND.t1 24.9236
R33 VGND.n1 VGND.t2 24.9236
R34 VGND.n5 VGND.n4 24.4711
R35 VGND.n3 VGND.n2 9.43392
R36 VGND.n6 VGND.n5 9.3005
R37 VGND.n4 VGND.n0 9.3005
R38 VGND.n2 VGND.n0 0.554787
R39 VGND.n6 VGND.n0 0.120292
R40 VGND VGND.n6 0.0213333
R41 VNB.t1 VNB.t0 1196.12
R42 VNB.t2 VNB.t1 1196.12
R43 VNB.t3 VNB.t2 1196.12
R44 VNB VNB.t3 968.285
R45 A.n0 A.t0 212.081
R46 A.n1 A.t3 212.081
R47 A A.n2 183.68
R48 A.n0 A.t1 139.78
R49 A.n1 A.t2 139.78
R50 A.n2 A.n0 38.7066
R51 A.n2 A.n1 22.6399
R52 VPWR VPWR.n0 316.39
R53 VPWR.n0 VPWR.t1 26.5955
R54 VPWR.n0 VPWR.t0 26.5955
C0 VPB A 0.056273f
C1 VPB B 0.056648f
C2 Y VPB 0.009606f
C3 A B 0.071165f
C4 VPB VPWR 0.049962f
C5 VGND VPB 0.006128f
C6 Y A 0.052333f
C7 A VPWR 0.041833f
C8 VGND A 0.059727f
C9 Y B 0.179365f
C10 B VPWR 0.017427f
C11 Y VPWR 0.012692f
C12 VGND B 0.029406f
C13 Y VGND 0.289148f
C14 VGND VPWR 0.046681f
C15 VGND VNB 0.342832f
C16 Y VNB 0.064071f
C17 VPWR VNB 0.248551f
C18 B VNB 0.197736f
C19 A VNB 0.206739f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y.t3 B.t0 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t1 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t0 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 A.t1 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t5 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND.t0 B.t2 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t3 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297.t1 B.t3 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 B.n0 B.t3 212.081
R1 B.n1 B.t0 212.081
R2 B B.n2 182.081
R3 B.n0 B.t2 139.78
R4 B.n1 B.t1 139.78
R5 B.n2 B.n0 30.6732
R6 B.n2 B.n1 30.6732
R7 a_27_297.n0 a_27_297.t1 404.502
R8 a_27_297.n0 a_27_297.t3 301.301
R9 a_27_297.n1 a_27_297.n0 184.905
R10 a_27_297.n1 a_27_297.t2 26.5955
R11 a_27_297.t0 a_27_297.n1 26.5955
R12 Y Y.n0 591.788
R13 Y.n4 Y.n0 585
R14 Y.n3 Y.n1 135.249
R15 Y.n3 Y.n2 98.982
R16 Y.n4 Y.n3 74.7314
R17 Y.n0 Y.t2 26.5955
R18 Y.n0 Y.t3 26.5955
R19 Y.n2 Y.t0 24.9236
R20 Y.n2 Y.t1 24.9236
R21 Y.n1 Y.t4 24.9236
R22 Y.n1 Y.t5 24.9236
R23 Y Y.n4 6.4005
R24 VPB.t2 VPB.t1 248.599
R25 VPB.t0 VPB.t2 248.599
R26 VPB.t3 VPB.t0 248.599
R27 VPB VPB.t3 201.246
R28 VGND.n2 VGND.t0 287.377
R29 VGND.n3 VGND.n1 207.965
R30 VGND.n5 VGND.t3 150.922
R31 VGND.n4 VGND.n3 32.377
R32 VGND.n1 VGND.t1 24.9236
R33 VGND.n1 VGND.t2 24.9236
R34 VGND.n5 VGND.n4 24.4711
R35 VGND.n3 VGND.n2 9.43392
R36 VGND.n6 VGND.n5 9.3005
R37 VGND.n4 VGND.n0 9.3005
R38 VGND.n2 VGND.n0 0.554787
R39 VGND.n6 VGND.n0 0.120292
R40 VGND VGND.n6 0.0213333
R41 VNB.t1 VNB.t0 1196.12
R42 VNB.t2 VNB.t1 1196.12
R43 VNB.t3 VNB.t2 1196.12
R44 VNB VNB.t3 968.285
R45 A.n0 A.t0 212.081
R46 A.n1 A.t3 212.081
R47 A A.n2 183.68
R48 A.n0 A.t1 139.78
R49 A.n1 A.t2 139.78
R50 A.n2 A.n0 38.7066
R51 A.n2 A.n1 22.6399
R52 VPWR VPWR.n0 316.39
R53 VPWR.n0 VPWR.t1 26.5955
R54 VPWR.n0 VPWR.t0 26.5955
C0 VPB A 0.056273f
C1 VPB B 0.056648f
C2 Y VPB 0.009606f
C3 A B 0.071165f
C4 VPB VPWR 0.049962f
C5 VGND VPB 0.006128f
C6 Y A 0.052333f
C7 A VPWR 0.041833f
C8 VGND A 0.059727f
C9 Y B 0.179365f
C10 B VPWR 0.017427f
C11 Y VPWR 0.012692f
C12 VGND B 0.029406f
C13 Y VGND 0.289148f
C14 VGND VPWR 0.046681f
C15 VGND VNB 0.342832f
C16 Y VNB 0.064071f
C17 VPWR VNB 0.248551f
C18 B VNB 0.197736f
C19 A VNB 0.206739f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t0 A.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n0 A.t3 212.081
R1 A.n1 A.t0 212.081
R2 A A.n1 189.073
R3 A.n0 A.t1 139.78
R4 A.n1 A.t2 139.78
R5 A.n1 A.n0 61.346
R6 VPWR.n0 VPWR.t0 262.851
R7 VPWR.n0 VPWR.t1 259.721
R8 VPWR VPWR.n0 0.491471
R9 Y.n2 Y.n1 208.965
R10 Y Y.n0 96.8352
R11 Y.n1 Y.t0 26.5955
R12 Y.n1 Y.t1 26.5955
R13 Y.n0 Y.t3 24.9236
R14 Y.n0 Y.t2 24.9236
R15 Y.n3 Y 11.2645
R16 Y Y.n3 6.1445
R17 Y.n3 Y 4.65505
R18 Y Y.n2 2.0485
R19 Y.n2 Y 1.55202
R20 VPB.t1 VPB.t0 248.599
R21 VPB VPB.t1 198.287
R22 VGND.n0 VGND.t1 169.418
R23 VGND.n0 VGND.t0 166.787
R24 VGND VGND.n0 0.491471
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 954.045
C0 Y VGND 0.154601f
C1 VPB A 0.074183f
C2 VPB VPWR 0.052063f
C3 A VPWR 0.06305f
C4 VGND VPB 0.006491f
C5 VGND A 0.063754f
C6 VGND VPWR 0.042274f
C7 Y VPB 0.006097f
C8 Y A 0.089386f
C9 Y VPWR 0.209105f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t0 A.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n0 A.t3 212.081
R1 A.n1 A.t0 212.081
R2 A A.n1 189.073
R3 A.n0 A.t1 139.78
R4 A.n1 A.t2 139.78
R5 A.n1 A.n0 61.346
R6 VPWR.n0 VPWR.t0 262.851
R7 VPWR.n0 VPWR.t1 259.721
R8 VPWR VPWR.n0 0.491471
R9 Y.n2 Y.n1 208.965
R10 Y Y.n0 96.8352
R11 Y.n1 Y.t0 26.5955
R12 Y.n1 Y.t1 26.5955
R13 Y.n0 Y.t3 24.9236
R14 Y.n0 Y.t2 24.9236
R15 Y.n3 Y 11.2645
R16 Y Y.n3 6.1445
R17 Y.n3 Y 4.65505
R18 Y Y.n2 2.0485
R19 Y.n2 Y 1.55202
R20 VPB.t1 VPB.t0 248.599
R21 VPB VPB.t1 198.287
R22 VGND.n0 VGND.t1 169.418
R23 VGND.n0 VGND.t0 166.787
R24 VGND VGND.n0 0.491471
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 954.045
C0 Y VGND 0.154601f
C1 VPB A 0.074183f
C2 VPB VPWR 0.052063f
C3 A VPWR 0.06305f
C4 VGND VPB 0.006491f
C5 VGND A 0.063754f
C6 VGND VPWR 0.042274f
C7 Y VPB 0.006097f
C8 Y A 0.089386f
C9 Y VPWR 0.209105f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends


* NGSPICE file created from sky130_fd_sc_hd__maj3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_1 VPB VNB VGND VPWR X C A B
X0 X.t0 a_27_47.t6 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.23725 pd=2.03 as=0.1474 ps=1.215 w=0.65 l=0.15
X1 X.t1 a_27_47.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=2.73 as=0.2492 ps=1.565 w=1 l=0.15
X2 a_109_341.t0 C.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_27_47.t4 B.t0 a_265_341.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VGND.t2 A.t0 a_109_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_265_341.t0 A.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR.t3 A.t2 a_109_341.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_421_47.t1 B.t1 a_27_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_265_47.t1 A.t3 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND.t1 C.t1 a_421_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1474 pd=1.215 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_27_47.t1 B.t2 a_265_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR.t1 C.t2 a_421_341.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2492 pd=1.565 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 a_421_341.t1 B.t3 a_27_47.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_109_47.t0 C.t3 a_27_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t0 a_27_47.n5 706.168
R1 a_27_47.n2 a_27_47.n0 612.717
R2 a_27_47.n5 a_27_47.t3 238.095
R3 a_27_47.n2 a_27_47.n1 236.481
R4 a_27_47.n1 a_27_47.t7 236.18
R5 a_27_47.n4 a_27_47.n3 185
R6 a_27_47.n1 a_27_47.t6 163.881
R7 a_27_47.n5 a_27_47.n4 98.5764
R8 a_27_47.n4 a_27_47.n2 66.2609
R9 a_27_47.n0 a_27_47.t2 63.3219
R10 a_27_47.n0 a_27_47.t4 63.3219
R11 a_27_47.n3 a_27_47.t5 38.5719
R12 a_27_47.n3 a_27_47.t1 38.5719
R13 VGND.n2 VGND.n0 205.996
R14 VGND.n2 VGND.n1 205.696
R15 VGND.n1 VGND.t0 78.7917
R16 VGND.n1 VGND.t1 70.0005
R17 VGND.n0 VGND.t3 38.5719
R18 VGND.n0 VGND.t2 38.5719
R19 VGND VGND.n2 0.274268
R20 X.n3 X.n2 585
R21 X.n2 X 304.101
R22 X.n0 X 186.695
R23 X.n1 X.n0 185
R24 X.n2 X.t1 47.2805
R25 X.n0 X.t0 44.3082
R26 X.n5 X 15.9294
R27 X.n1 X 11.1064
R28 X.n4 X.n3 6.4005
R29 X.n3 X 4.84898
R30 X X.n5 3.41383
R31 X X.n4 2.84494
R32 X.n5 X 2.25932
R33 X.n4 X 1.93989
R34 X X.n1 1.69462
R35 VNB.t1 VNB.t0 2036.25
R36 VNB.t2 VNB.t5 1196.12
R37 VNB.t3 VNB.t6 1196.12
R38 VNB.t5 VNB.t1 1025.24
R39 VNB.t6 VNB.t2 1025.24
R40 VNB.t4 VNB.t3 1025.24
R41 VNB VNB.t4 911.327
R42 VPWR.n2 VPWR.n0 632.029
R43 VPWR.n2 VPWR.n1 322.767
R44 VPWR.n1 VPWR.t1 106.186
R45 VPWR.n0 VPWR.t2 63.3219
R46 VPWR.n0 VPWR.t3 63.3219
R47 VPWR.n1 VPWR.t0 57.2545
R48 VPWR VPWR.n2 0.282199
R49 VPB.t2 VPB.t0 423.209
R50 VPB.t5 VPB.t3 248.599
R51 VPB.t6 VPB.t4 248.599
R52 VPB.t3 VPB.t2 213.084
R53 VPB.t4 VPB.t5 213.084
R54 VPB.t1 VPB.t6 213.084
R55 VPB VPB.t1 189.409
R56 C.t2 C.t0 970.428
R57 C.t0 C.t3 472.361
R58 C.n0 C.t2 208.3
R59 C.n0 C.t1 195.446
R60 C C.n0 154.857
R61 a_109_341.t0 a_109_341.t1 98.5005
R62 B.n0 B.t3 189.588
R63 B.n1 B.t0 189.588
R64 B.n0 B.t1 176.733
R65 B.n1 B.t2 176.733
R66 B B.n2 157.988
R67 B.n2 B.n0 30.6732
R68 B.n2 B.n1 30.6732
R69 a_265_341.t0 a_265_341.t1 98.5005
R70 A.n0 A.t1 189.588
R71 A.n1 A.t2 189.588
R72 A.n0 A.t3 176.733
R73 A.n1 A.t0 176.733
R74 A A.n2 168.679
R75 A.n2 A.n0 30.6732
R76 A.n2 A.n1 30.6732
R77 a_109_47.t0 a_109_47.t1 60.0005
R78 a_421_47.t0 a_421_47.t1 60.0005
R79 a_265_47.t0 a_265_47.t1 60.0005
R80 a_421_341.t0 a_421_341.t1 98.5005
C0 B VGND 0.019483f
C1 VPWR X 0.087666f
C2 A VPB 0.082062f
C3 VPWR VGND 0.07394f
C4 A C 0.148433f
C5 X VGND 0.065924f
C6 B VPB 0.073834f
C7 VPWR VPB 0.097459f
C8 B C 0.127365f
C9 VPWR C 0.090262f
C10 X VPB 0.011741f
C11 X C 0.011556f
C12 VGND VPB 0.011198f
C13 A B 0.132046f
C14 VGND C 0.054519f
C15 A VPWR 0.121153f
C16 A VGND 0.032104f
C17 B VPWR 0.016556f
C18 VPB C 0.266419f
C19 B X 2.05e-19
C20 VGND VNB 0.442359f
C21 X VNB 0.09315f
C22 VPWR VNB 0.370922f
C23 B VNB 0.174586f
C24 A VNB 0.185641f
C25 C VNB 0.341798f
C26 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__maj3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_2 VNB VPB VGND VPWR X A B C
X0 VGND.t4 C.t0 a_441_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.162225 pd=1.25 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_285_369.t0 A.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 a_47_47.t2 B.t0 a_285_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR.t2 A.t1 a_129_369.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X4 a_129_47.t1 C.t1 a_47_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR.t4 C.t2 a_441_369.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.237 pd=1.6 as=0.0672 ps=0.85 w=0.64 l=0.15
X6 VPWR.t3 a_47_47.t6 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t3 a_47_47.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.162225 ps=1.25 w=0.65 l=0.15
X8 a_129_369.t1 C.t3 a_47_47.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 X.t0 a_47_47.t8 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.237 ps=1.6 w=1 l=0.15
X10 VGND.t0 A.t2 a_129_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 a_441_369.t0 B.t1 a_47_47.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 a_47_47.t1 B.t2 a_285_369.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X13 a_441_47.t0 B.t3 a_47_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VGND.t3 a_47_47.t9 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_285_47.t1 A.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 C.n1 C.t0 321.772
R1 C.n0 C.t3 299.377
R2 C C.n0 292.378
R3 C.n0 C.t1 206.19
R4 C.n1 C.t2 183.599
R5 C.n2 C.n1 152
R6 C C.n2 16.3845
R7 C.n2 C 6.9125
R8 a_441_47.t0 a_441_47.t1 60.0005
R9 VGND.n3 VGND.n2 199.739
R10 VGND.n10 VGND.n9 198.964
R11 VGND.n4 VGND.t3 160.034
R12 VGND.n2 VGND.t2 88.1104
R13 VGND.n2 VGND.t4 67.1434
R14 VGND.n9 VGND.t1 38.5719
R15 VGND.n9 VGND.t0 38.5719
R16 VGND.n7 VGND.n1 34.6358
R17 VGND.n8 VGND.n7 34.6358
R18 VGND.n10 VGND.n8 22.9652
R19 VGND.n8 VGND.n0 9.3005
R20 VGND.n7 VGND.n6 9.3005
R21 VGND.n5 VGND.n1 9.3005
R22 VGND.n4 VGND.n3 9.11771
R23 VGND.n3 VGND.n1 7.90638
R24 VGND.n11 VGND.n10 7.02387
R25 VGND.n5 VGND.n4 0.503351
R26 VGND VGND.n11 0.228883
R27 VGND.n11 VGND.n0 0.154841
R28 VGND.n6 VGND.n5 0.120292
R29 VGND.n6 VGND.n0 0.120292
R30 VNB.t7 VNB.t2 2135.92
R31 VNB VNB.t6 1210.36
R32 VNB.t2 VNB.t3 1196.12
R33 VNB.t5 VNB.t4 1196.12
R34 VNB.t0 VNB.t1 1196.12
R35 VNB.t4 VNB.t7 1025.24
R36 VNB.t1 VNB.t5 1025.24
R37 VNB.t6 VNB.t0 1025.24
R38 A.n0 A.t0 269.921
R39 A.n1 A.t1 269.921
R40 A.n0 A.t3 176.733
R41 A.n1 A.t2 176.733
R42 A.n3 A.n2 152
R43 A.n2 A.n0 30.6732
R44 A.n2 A.n1 30.6732
R45 A.n3 A 14.9338
R46 A A.n3 2.90959
R47 VPWR.n1 VPWR.n0 599.74
R48 VPWR.n4 VPWR.n3 310.777
R49 VPWR.n5 VPWR.t3 255.394
R50 VPWR.n3 VPWR.t0 133.184
R51 VPWR.n0 VPWR.t1 41.5552
R52 VPWR.n0 VPWR.t2 41.5552
R53 VPWR.n3 VPWR.t4 41.5552
R54 VPWR.n8 VPWR.n7 34.6358
R55 VPWR.n9 VPWR.n8 34.6358
R56 VPWR.n9 VPWR.n1 22.9652
R57 VPWR.n5 VPWR.n4 17.0236
R58 VPWR.n7 VPWR.n6 9.3005
R59 VPWR.n8 VPWR.n2 9.3005
R60 VPWR.n10 VPWR.n9 9.3005
R61 VPWR.n11 VPWR.n1 7.02387
R62 VPWR.n6 VPWR.n5 0.503351
R63 VPWR.n7 VPWR.n4 0.376971
R64 VPWR VPWR.n11 0.228883
R65 VPWR.n11 VPWR.n10 0.154841
R66 VPWR.n6 VPWR.n2 0.120292
R67 VPWR.n10 VPWR.n2 0.120292
R68 a_285_369.t0 a_285_369.t1 64.6411
R69 VPB.t5 VPB.t0 443.925
R70 VPB VPB.t4 251.559
R71 VPB.t0 VPB.t3 248.599
R72 VPB.t7 VPB.t6 248.599
R73 VPB.t1 VPB.t2 248.599
R74 VPB.t6 VPB.t5 213.084
R75 VPB.t2 VPB.t7 213.084
R76 VPB.t4 VPB.t1 213.084
R77 B.n0 B.t1 269.921
R78 B.n1 B.t2 269.921
R79 B.n0 B.t3 176.733
R80 B.n1 B.t0 176.733
R81 B B.n2 154.429
R82 B.n2 B.n1 35.055
R83 B.n2 B.n0 26.2914
R84 a_285_47.t0 a_285_47.t1 60.0005
R85 a_47_47.n6 a_47_47.n5 384.7
R86 a_47_47.n5 a_47_47.t4 360.846
R87 a_47_47.n3 a_47_47.n1 268.699
R88 a_47_47.n4 a_47_47.t5 232.154
R89 a_47_47.n0 a_47_47.t6 221.72
R90 a_47_47.n1 a_47_47.t8 221.72
R91 a_47_47.n3 a_47_47.n2 199.739
R92 a_47_47.n0 a_47_47.t9 149.421
R93 a_47_47.n1 a_47_47.t7 149.421
R94 a_47_47.n4 a_47_47.n3 92.6123
R95 a_47_47.n5 a_47_47.n4 80.5731
R96 a_47_47.n1 a_47_47.n0 74.9783
R97 a_47_47.n6 a_47_47.t3 41.5552
R98 a_47_47.t1 a_47_47.n6 41.5552
R99 a_47_47.n2 a_47_47.t0 38.5719
R100 a_47_47.n2 a_47_47.t2 38.5719
R101 a_129_369.t0 a_129_369.t1 64.6411
R102 a_129_47.t0 a_129_47.t1 60.0005
R103 a_441_369.t0 a_441_369.t1 64.6411
R104 X.n1 X.n0 259.401
R105 X X.n2 185.97
R106 X.n2 X.n1 185
R107 X.n0 X.t1 26.5955
R108 X.n0 X.t0 26.5955
R109 X.n2 X.t2 24.9236
R110 X.n2 X.t3 24.9236
R111 X X.n1 12.2187
C0 VPB A 0.085303f
C1 C A 0.216633f
C2 VPB B 0.084464f
C3 C B 0.161534f
C4 VPB VPWR 0.09607f
C5 C VPWR 0.085287f
C6 A B 0.146077f
C7 VPB X 0.009436f
C8 C X 0.020273f
C9 A VPWR 0.031744f
C10 VPB VGND 0.010399f
C11 B VPWR 0.023811f
C12 C VGND 0.029213f
C13 A X 2.74e-19
C14 B X 0.00232f
C15 A VGND 0.032512f
C16 VPWR X 0.162928f
C17 B VGND 0.021529f
C18 VPWR VGND 0.095199f
C19 X VGND 0.116907f
C20 VPB C 0.142127f
C21 VGND VNB 0.51576f
C22 X VNB 0.023995f
C23 VPWR VNB 0.443473f
C24 B VNB 0.189444f
C25 A VNB 0.189624f
C26 C VNB 0.262485f
C27 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__maj3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_4 VPB VNB VGND VPWR A X B C
X0 X.t3 a_47_297.t6 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.157625 ps=1.135 w=0.65 l=0.15
X1 a_151_297.t0 C.t0 a_47_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1225 pd=1.245 as=0.37 ps=2.74 w=1 l=0.15
X2 VPWR.t1 A.t0 a_151_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1225 ps=1.245 w=1 l=0.15
X3 VGND.t0 A.t1 a_151_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.079625 ps=0.895 w=0.65 l=0.15
X4 VGND.t5 a_47_297.t7 X.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t4 a_47_297.t8 X.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 C.t1 a_482_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.105 ps=1.21 w=1 l=0.15
X7 a_314_47.t0 A.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_482_47.t1 B.t0 a_47_297.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X.t0 a_47_297.t9 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR.t6 a_47_297.t10 X.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_482_297.t1 B.t1 a_47_297.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t2 C.t2 a_482_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.157625 pd=1.135 as=0.06825 ps=0.86 w=0.65 l=0.15
X13 X.t6 a_47_297.t11 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_47_297.t0 B.t2 a_314_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t4 a_47_297.t12 X.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_47_297.t4 B.t3 a_314_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_314_297.t0 A.t3 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_151_47.t0 C.t3 a_47_297.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.079625 pd=0.895 as=0.182 ps=1.86 w=0.65 l=0.15
X19 X.t4 a_47_297.t13 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2425 ps=1.485 w=1 l=0.15
R0 a_47_297.n13 a_47_297.n12 361.783
R1 a_47_297.n11 a_47_297.t2 296.728
R2 a_47_297.n1 a_47_297.t10 212.081
R3 a_47_297.n3 a_47_297.t11 212.081
R4 a_47_297.n5 a_47_297.t12 212.081
R5 a_47_297.n6 a_47_297.t13 212.081
R6 a_47_297.n2 a_47_297.n0 177.601
R7 a_47_297.n8 a_47_297.n7 152
R8 a_47_297.n4 a_47_297.n0 152
R9 a_47_297.n1 a_47_297.t8 139.78
R10 a_47_297.n3 a_47_297.t9 139.78
R11 a_47_297.n5 a_47_297.t7 139.78
R12 a_47_297.n6 a_47_297.t6 139.78
R13 a_47_297.n11 a_47_297.t3 131.942
R14 a_47_297.n10 a_47_297.n8 104.712
R15 a_47_297.n10 a_47_297.n9 97.6244
R16 a_47_297.n12 a_47_297.n11 60.8716
R17 a_47_297.n2 a_47_297.n1 30.6732
R18 a_47_297.n3 a_47_297.n2 30.6732
R19 a_47_297.n4 a_47_297.n3 30.6732
R20 a_47_297.n5 a_47_297.n4 30.6732
R21 a_47_297.n7 a_47_297.n5 30.6732
R22 a_47_297.n7 a_47_297.n6 30.6732
R23 a_47_297.n13 a_47_297.t5 26.5955
R24 a_47_297.t0 a_47_297.n13 26.5955
R25 a_47_297.n8 a_47_297.n0 25.6005
R26 a_47_297.n9 a_47_297.t1 24.9236
R27 a_47_297.n9 a_47_297.t4 24.9236
R28 a_47_297.n12 a_47_297.n10 14.5072
R29 VGND.n5 VGND.t4 297.377
R30 VGND.n4 VGND.n3 207.213
R31 VGND.n17 VGND.n16 199.739
R32 VGND.n10 VGND.n9 199.1
R33 VGND.n9 VGND.t2 47.0774
R34 VGND.n9 VGND.t6 42.462
R35 VGND.n5 VGND.n4 36.5149
R36 VGND.n8 VGND.n7 34.6358
R37 VGND.n14 VGND.n1 34.6358
R38 VGND.n15 VGND.n14 34.6358
R39 VGND.n3 VGND.t3 24.9236
R40 VGND.n3 VGND.t5 24.9236
R41 VGND.n16 VGND.t1 24.9236
R42 VGND.n16 VGND.t0 24.9236
R43 VGND.n10 VGND.n1 24.8476
R44 VGND.n10 VGND.n8 18.4476
R45 VGND.n17 VGND.n15 12.0476
R46 VGND.n7 VGND.n6 9.3005
R47 VGND.n8 VGND.n2 9.3005
R48 VGND.n11 VGND.n10 9.3005
R49 VGND.n12 VGND.n1 9.3005
R50 VGND.n14 VGND.n13 9.3005
R51 VGND.n15 VGND.n0 9.3005
R52 VGND.n18 VGND.n17 7.52635
R53 VGND.n7 VGND.n4 3.76521
R54 VGND.n6 VGND.n5 2.15642
R55 VGND VGND.n18 0.237813
R56 VGND.n18 VGND.n0 0.147328
R57 VGND.n6 VGND.n2 0.120292
R58 VGND.n11 VGND.n2 0.120292
R59 VGND.n12 VGND.n11 0.120292
R60 VGND.n13 VGND.n12 0.120292
R61 VGND.n13 VGND.n0 0.120292
R62 X.n5 X.n3 243.843
R63 X.n5 X.n4 205.442
R64 X.n2 X.n0 134.6
R65 X.n2 X.n1 98.4002
R66 X.n3 X.t5 26.5955
R67 X.n3 X.t4 26.5955
R68 X.n4 X.t7 26.5955
R69 X.n4 X.t6 26.5955
R70 X.n0 X.t2 24.9236
R71 X.n0 X.t3 24.9236
R72 X.n1 X.t1 24.9236
R73 X.n1 X.t0 24.9236
R74 X X.n5 17.4774
R75 X.n6 X 14.5236
R76 X.n6 X.n2 11.4531
R77 X X.n6 2.21588
R78 VNB.t3 VNB.t9 1808.41
R79 VNB VNB.t4 1537.86
R80 VNB.t6 VNB.t7 1196.12
R81 VNB.t8 VNB.t6 1196.12
R82 VNB.t9 VNB.t8 1196.12
R83 VNB.t5 VNB.t0 1196.12
R84 VNB.t2 VNB.t5 1196.12
R85 VNB.t1 VNB.t2 1196.12
R86 VNB.t4 VNB.t1 1124.92
R87 VNB.t0 VNB.t3 1025.24
R88 C C.n0 444.661
R89 C.n0 C.t1 236.552
R90 C.n1 C.t0 236.18
R91 C.n0 C.t2 164.251
R92 C.n1 C.t3 163.881
R93 C C.n1 152.915
R94 a_151_297.t0 a_151_297.t1 48.2655
R95 VPB.t1 VPB.t6 375.858
R96 VPB VPB.t2 319.627
R97 VPB.t8 VPB.t9 248.599
R98 VPB.t7 VPB.t8 248.599
R99 VPB.t6 VPB.t7 248.599
R100 VPB.t0 VPB.t4 248.599
R101 VPB.t5 VPB.t0 248.599
R102 VPB.t3 VPB.t5 248.599
R103 VPB.t2 VPB.t3 233.802
R104 VPB.t4 VPB.t1 213.084
R105 A.n0 A.t3 212.081
R106 A.n1 A.t0 212.081
R107 A.n3 A.n2 152
R108 A.n0 A.t2 139.78
R109 A.n1 A.t1 139.78
R110 A.n2 A.n0 30.6732
R111 A.n2 A.n1 30.6732
R112 A.n3 A 9.35435
R113 A A.n3 1.80563
R114 VPWR.n1 VPWR.n0 599.74
R115 VPWR.n7 VPWR.t6 353.411
R116 VPWR.n8 VPWR.n6 321.695
R117 VPWR.n4 VPWR.n3 217.581
R118 VPWR.n3 VPWR.t3 48.2655
R119 VPWR.n3 VPWR.t0 47.2805
R120 VPWR.n8 VPWR.n7 36.2765
R121 VPWR.n15 VPWR.n14 34.6358
R122 VPWR.n16 VPWR.n15 34.6358
R123 VPWR.n10 VPWR.n9 34.6358
R124 VPWR.n0 VPWR.t2 26.5955
R125 VPWR.n0 VPWR.t1 26.5955
R126 VPWR.n6 VPWR.t5 26.5955
R127 VPWR.n6 VPWR.t4 26.5955
R128 VPWR.n14 VPWR.n4 23.7181
R129 VPWR.n10 VPWR.n4 20.7064
R130 VPWR.n16 VPWR.n1 12.0476
R131 VPWR.n9 VPWR.n5 9.3005
R132 VPWR.n11 VPWR.n10 9.3005
R133 VPWR.n12 VPWR.n4 9.3005
R134 VPWR.n14 VPWR.n13 9.3005
R135 VPWR.n15 VPWR.n2 9.3005
R136 VPWR.n17 VPWR.n16 9.3005
R137 VPWR.n18 VPWR.n1 7.52635
R138 VPWR.n9 VPWR.n8 3.76521
R139 VPWR.n7 VPWR.n5 2.08078
R140 VPWR VPWR.n18 0.237813
R141 VPWR.n18 VPWR.n17 0.147328
R142 VPWR.n11 VPWR.n5 0.120292
R143 VPWR.n12 VPWR.n11 0.120292
R144 VPWR.n13 VPWR.n12 0.120292
R145 VPWR.n13 VPWR.n2 0.120292
R146 VPWR.n17 VPWR.n2 0.120292
R147 a_151_47.t0 a_151_47.t1 45.2313
R148 a_482_297.t0 a_482_297.t1 41.3705
R149 a_314_47.t0 a_314_47.t1 49.8467
R150 B.n0 B.t1 212.081
R151 B.n1 B.t2 212.081
R152 B B.n2 159.424
R153 B.n0 B.t0 139.78
R154 B.n1 B.t3 139.78
R155 B.n2 B.n0 30.6732
R156 B.n2 B.n1 30.6732
R157 a_482_47.t0 a_482_47.t1 38.7697
R158 a_314_297.t0 a_314_297.t1 53.1905
C0 X VPWR 0.399413f
C1 X VGND 0.256905f
C2 VPB C 0.073395f
C3 VPB A 0.052198f
C4 VPB B 0.050258f
C5 C A 0.156669f
C6 C B 0.119365f
C7 VPB VPWR 0.104504f
C8 VGND VPB 0.006661f
C9 C VPWR 0.295422f
C10 A B 0.050963f
C11 VGND C 0.032063f
C12 X VPB 0.01284f
C13 A VPWR 0.03279f
C14 VGND A 0.029635f
C15 X C 0.002415f
C16 B VPWR 0.020256f
C17 VGND B 0.025551f
C18 VGND VPWR 0.101493f
C19 X B 1.54e-19
C20 VGND VNB 0.583547f
C21 X VNB 0.058681f
C22 VPWR VNB 0.502341f
C23 B VNB 0.165877f
C24 A VNB 0.167306f
C25 C VNB 0.224552f
C26 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR.t3 a_505_21.t2 a_535_374.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21.t1 S.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374.t0 S.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND.t2 a_505_21.t3 a_439_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199.t2 A0.t0 a_218_374.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21.t0 S.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47.t1 A0.t1 a_76_199.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374.t1 A1.t0 a_76_199.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199.t1 A1.t1 a_218_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47.t0 S.t3 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR.t2 a_76_199.t4 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND.t3 a_76_199.t5 X.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_505_21.n1 a_505_21.t1 703.471
R1 a_505_21.n0 a_505_21.t2 329.805
R2 a_505_21.t0 a_505_21.n1 246.56
R3 a_505_21.n0 a_505_21.t3 209.597
R4 a_505_21.n1 a_505_21.n0 202.071
R5 a_535_374.t0 a_535_374.t1 98.5005
R6 VPWR.n2 VPWR.n0 642.889
R7 VPWR.n2 VPWR.n1 242.226
R8 VPWR.n1 VPWR.t0 123.507
R9 VPWR.n0 VPWR.t3 86.7743
R10 VPWR.n0 VPWR.t1 68.0124
R11 VPWR.n1 VPWR.t2 28.752
R12 VPWR VPWR.n2 0.145102
R13 VPB.t5 VPB.t4 633.333
R14 VPB.t2 VPB.t0 322.587
R15 VPB.t0 VPB.t5 304.829
R16 VPB.t3 VPB.t1 284.113
R17 VPB.t4 VPB.t3 213.084
R18 VPB VPB.t2 59.1905
R19 S S.n1 428.005
R20 S.n0 S.t2 329.902
R21 S.n1 S.t1 272.062
R22 S.n1 S.t3 206.19
R23 S S.n0 152.674
R24 S.n0 S.t0 148.35
R25 a_218_374.t0 a_218_374.t1 171.202
R26 a_439_47.t0 a_439_47.t1 94.2862
R27 VGND.n13 VGND.n12 199.739
R28 VGND.n3 VGND.n2 187.565
R29 VGND.n5 VGND.n4 185
R30 VGND.n4 VGND.n3 97.1434
R31 VGND.n12 VGND.t1 74.2862
R32 VGND.n4 VGND.t2 61.4291
R33 VGND.n3 VGND.t0 38.5719
R34 VGND.n6 VGND.n1 34.6358
R35 VGND.n10 VGND.n1 34.6358
R36 VGND.n11 VGND.n10 34.6358
R37 VGND.n12 VGND.t3 25.4291
R38 VGND.n13 VGND.n11 22.9652
R39 VGND.n6 VGND.n5 22.2496
R40 VGND.n11 VGND.n0 9.3005
R41 VGND.n10 VGND.n9 9.3005
R42 VGND.n8 VGND.n1 9.3005
R43 VGND.n7 VGND.n6 9.3005
R44 VGND.n14 VGND.n13 7.12063
R45 VGND.n7 VGND.n2 5.59093
R46 VGND.n5 VGND.n2 3.03853
R47 VGND.n14 VGND.n0 0.148519
R48 VGND.n8 VGND.n7 0.120292
R49 VGND.n9 VGND.n8 0.120292
R50 VGND.n9 VGND.n0 0.120292
R51 VGND VGND.n14 0.11354
R52 VNB.t2 VNB.t1 2392.23
R53 VNB.t5 VNB.t4 1779.94
R54 VNB.t3 VNB.t0 1552.1
R55 VNB.t4 VNB.t2 1366.99
R56 VNB.t0 VNB.t5 1366.99
R57 VNB VNB.t3 142.395
R58 A0.n0 A0.t0 471.289
R59 A0 A0.n0 154.097
R60 A0.n0 A0.t1 148.35
R61 a_76_199.n3 a_76_199.n2 390.017
R62 a_76_199.n0 a_76_199.t4 241.536
R63 a_76_199.n2 a_76_199.n0 223.53
R64 a_76_199.t0 a_76_199.n3 214.52
R65 a_76_199.n2 a_76_199.n1 206.403
R66 a_76_199.n3 a_76_199.t2 194.49
R67 a_76_199.n0 a_76_199.t5 169.237
R68 a_76_199.n1 a_76_199.t3 94.2862
R69 a_76_199.n1 a_76_199.t1 41.4291
R70 A1.n0 A1.t1 414.432
R71 A1.n0 A1.t0 300.349
R72 A1 A1.n0 29.6426
R73 a_218_47.t0 a_218_47.t1 94.2862
R74 X X.n0 593.216
R75 X.n3 X.n0 585
R76 X.n2 X.n0 585
R77 X.n1 X.t0 209.923
R78 X.n2 X.n1 74.3207
R79 X.n0 X.t1 26.5955
R80 X.n3 X 8.21543
R81 X X.n3 4.77662
R82 X X.n2 4.77662
R83 X.n1 X 2.5103
C0 A1 VGND 0.075211f
C1 VPB VGND 0.013448f
C2 VPWR A0 0.007316f
C3 VPB X 0.012046f
C4 S A0 0.034107f
C5 X VGND 0.058643f
C6 VPWR A1 0.011366f
C7 VPB VPWR 0.10994f
C8 S A1 0.087223f
C9 VPWR VGND 0.080355f
C10 VPB S 0.168493f
C11 X VPWR 0.12783f
C12 S VGND 0.032964f
C13 X S 0.00823f
C14 VPWR S 0.392437f
C15 A0 A1 0.266805f
C16 VPB A0 0.106597f
C17 A0 VGND 0.043233f
C18 VPB A1 0.072083f
C19 VGND VNB 0.498664f
C20 A1 VNB 0.140423f
C21 A0 VNB 0.13429f
C22 S VNB 0.268143f
C23 VPWR VNB 0.419248f
C24 X VNB 0.092356f
C25 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR.t1 S.t0 a_591_369.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369.t0 A0.t0 a_79_21.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X2 VPWR.t3 a_79_21.t4 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21.t3 A1.t0 a_306_369.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4 VGND.t4 a_79_21.t5 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t1 S.t1 a_578_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X6 a_306_369.t0 a_257_199.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X7 a_79_21.t1 A0.t1 a_288_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8 a_288_47.t1 a_257_199.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199.t1 S.t2 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47.t1 A1.t1 a_79_21.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11 X.t2 a_79_21.t6 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199.t0 S.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X.t0 a_79_21.t7 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 S.n0 S.t3 269.921
R1 S.n1 S.t0 269.921
R2 S.n0 S.t2 176.733
R3 S.n1 S.t1 176.733
R4 S.n3 S.n2 152
R5 S.n2 S.n1 31.4035
R6 S.n2 S.n0 29.9429
R7 S.n3 S 19.2005
R8 S S.n3 3.70576
R9 a_591_369.t0 a_591_369.t1 64.6411
R10 VPWR.n2 VPWR.n1 613.683
R11 VPWR.n4 VPWR.n3 601.773
R12 VPWR.n6 VPWR.t4 249.901
R13 VPWR.n3 VPWR.t0 70.7974
R14 VPWR.n3 VPWR.t3 46.9964
R15 VPWR.n1 VPWR.t2 41.5552
R16 VPWR.n1 VPWR.t1 41.5552
R17 VPWR.n6 VPWR.n5 25.977
R18 VPWR.n5 VPWR.n4 25.224
R19 VPWR.n5 VPWR.n0 9.3005
R20 VPWR.n7 VPWR.n6 9.3005
R21 VPWR.n4 VPWR.n2 7.06091
R22 VPWR.n2 VPWR.n0 0.157826
R23 VPWR.n7 VPWR.n0 0.120292
R24 VPWR VPWR.n7 0.0213333
R25 VPB.t0 VPB.t6 511.995
R26 VPB.t4 VPB.t0 334.425
R27 VPB.t6 VPB.t1 331.464
R28 VPB.t3 VPB.t2 248.599
R29 VPB.t5 VPB.t4 248.599
R30 VPB.t1 VPB.t3 213.084
R31 VPB VPB.t5 189.409
R32 A0.n1 A0.t0 367.733
R33 A0.n0 A0.t1 284.283
R34 A0.n1 A0 14.0392
R35 A0 A0.n1 4.95534
R36 A0 A0.n0 3.55606
R37 A0.n0 A0 3.35288
R38 a_79_21.n4 a_79_21.n3 765.742
R39 a_79_21.n2 a_79_21.t4 212.081
R40 a_79_21.n1 a_79_21.t6 212.081
R41 a_79_21.n3 a_79_21.n0 181.423
R42 a_79_21.n3 a_79_21.n2 159.304
R43 a_79_21.n2 a_79_21.t5 139.78
R44 a_79_21.n1 a_79_21.t7 139.78
R45 a_79_21.n0 a_79_21.t2 109.231
R46 a_79_21.n0 a_79_21.t1 87.5389
R47 a_79_21.n4 a_79_21.t3 72.3364
R48 a_79_21.n2 a_79_21.n1 61.346
R49 a_79_21.t0 a_79_21.n4 53.8677
R50 X.n0 X 592.226
R51 X.n1 X.n0 585
R52 X X.n2 273.365
R53 X.n0 X.t3 26.5955
R54 X.n0 X.t2 26.5955
R55 X.n2 X.t1 24.9236
R56 X.n2 X.t0 24.9236
R57 X X.n1 7.22631
R58 X.n1 X 6.8134
R59 A1.n0 A1.t0 457.024
R60 A1 A1.n0 157.298
R61 A1.n0 A1.t1 135.399
R62 a_306_369.t0 a_306_369.t1 220.087
R63 VGND.n2 VGND.n1 218.51
R64 VGND.n4 VGND.n3 199.739
R65 VGND.n6 VGND.t3 155.046
R66 VGND.n3 VGND.t0 54.2862
R67 VGND.n1 VGND.t2 38.5719
R68 VGND.n1 VGND.t1 38.5719
R69 VGND.n6 VGND.n5 25.977
R70 VGND.n3 VGND.t4 25.9346
R71 VGND.n5 VGND.n4 18.4476
R72 VGND.n7 VGND.n6 9.3005
R73 VGND.n5 VGND.n0 9.3005
R74 VGND.n4 VGND.n2 7.25702
R75 VGND.n2 VGND.n0 0.154487
R76 VGND.n7 VGND.n0 0.120292
R77 VGND VGND.n7 0.0213333
R78 VNB.t3 VNB.t6 2776.7
R79 VNB.t0 VNB.t3 1352.75
R80 VNB.t5 VNB.t0 1352.75
R81 VNB.t6 VNB.t2 1210.36
R82 VNB.t2 VNB.t1 1196.12
R83 VNB.t4 VNB.t5 1196.12
R84 VNB VNB.t4 911.327
R85 a_578_47.t0 a_578_47.t1 78.5719
R86 a_257_199.n1 a_257_199.n0 362.825
R87 a_257_199.t0 a_257_199.n1 360.752
R88 a_257_199.n0 a_257_199.t2 299.377
R89 a_257_199.n1 a_257_199.t1 284.562
R90 a_257_199.n0 a_257_199.t3 206.19
R91 a_288_47.t0 a_288_47.t1 92.8576
C0 VPB A1 0.058508f
C1 VPB A0 0.072912f
C2 VPB X 0.004573f
C3 A1 A0 0.157881f
C4 VPB S 0.098742f
C5 VPB VGND 0.011037f
C6 VPB VPWR 0.09532f
C7 A1 S 0.066236f
C8 A1 VGND 0.049662f
C9 A1 VPWR 0.009938f
C10 A0 S 0.084169f
C11 A0 VGND 0.018476f
C12 A0 VPWR 0.017749f
C13 X VGND 0.108904f
C14 VPWR X 0.149294f
C15 S VGND 0.056865f
C16 S VPWR 0.032955f
C17 VPWR VGND 0.092236f
C18 VGND VNB 0.515723f
C19 X VNB 0.024395f
C20 VPWR VNB 0.440866f
C21 S VNB 0.243683f
C22 A0 VNB 0.128792f
C23 A1 VNB 0.161724f
C24 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_4 VNB VPB VPWR VGND X S A1 A0
X0 a_204_297.t0 A1.t0 a_396_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR.t5 a_396_47.t4 X.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X.t2 a_396_47.t5 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t1 S.t0 a_314_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297.t1 a_27_47.t2 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_396_47.t3 A0.t0 a_314_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47.t0 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.108875 ps=0.985 w=0.65 l=0.15
X7 X.t7 a_396_47.t6 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X.t6 a_396_47.t7 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t3 a_396_47.t8 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47.t0 A1.t1 a_396_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND.t2 S.t1 a_490_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.274625 ps=1.495 w=0.65 l=0.15
X12 VGND.t4 a_396_47.t9 X.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_396_47.t2 A0.t1 a_206_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND.t3 a_396_47.t10 X.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR.t6 S.t2 a_27_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X16 X.t0 a_396_47.t11 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t1 S.t3 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t0 241.536
R1 A1.n0 A1.t1 169.237
R2 A1 A1.n0 166.352
R3 a_396_47.n13 a_396_47.n12 724.672
R4 a_396_47.n12 a_396_47.n0 331.825
R5 a_396_47.n3 a_396_47.t8 212.081
R6 a_396_47.n2 a_396_47.t11 212.081
R7 a_396_47.n7 a_396_47.t4 212.081
R8 a_396_47.n9 a_396_47.t5 212.081
R9 a_396_47.n5 a_396_47.n4 177.601
R10 a_396_47.n11 a_396_47.n10 152
R11 a_396_47.n8 a_396_47.n1 152
R12 a_396_47.n6 a_396_47.n5 152
R13 a_396_47.n3 a_396_47.t10 139.78
R14 a_396_47.n2 a_396_47.t7 139.78
R15 a_396_47.n7 a_396_47.t9 139.78
R16 a_396_47.n9 a_396_47.t6 139.78
R17 a_396_47.n10 a_396_47.n8 49.6611
R18 a_396_47.n7 a_396_47.n6 46.0096
R19 a_396_47.n4 a_396_47.n2 34.3247
R20 a_396_47.n13 a_396_47.t3 32.5055
R21 a_396_47.t0 a_396_47.n13 30.5355
R22 a_396_47.n0 a_396_47.t1 29.539
R23 a_396_47.n0 a_396_47.t2 29.539
R24 a_396_47.n4 a_396_47.n3 27.0217
R25 a_396_47.n5 a_396_47.n1 25.6005
R26 a_396_47.n11 a_396_47.n1 25.6005
R27 a_396_47.n6 a_396_47.n2 15.3369
R28 a_396_47.n12 a_396_47.n11 14.6829
R29 a_396_47.n10 a_396_47.n9 8.03383
R30 a_396_47.n8 a_396_47.n7 3.65202
R31 a_204_297.t0 a_204_297.t1 1249.63
R32 VPB.t0 VPB.t2 588.942
R33 VPB.t1 VPB.t3 568.225
R34 VPB.t8 VPB.t1 281.154
R35 VPB.t3 VPB.t0 278.193
R36 VPB.t4 VPB.t5 248.599
R37 VPB.t7 VPB.t4 248.599
R38 VPB.t6 VPB.t7 248.599
R39 VPB.t2 VPB.t6 248.599
R40 VPB VPB.t8 189.409
R41 X.n2 X.n1 378.2
R42 X.n2 X.n0 314.952
R43 X.n5 X.n4 264.435
R44 X.n5 X.n3 201.189
R45 X X.n2 39.0716
R46 X X.n5 29.6107
R47 X.n0 X.t1 26.5955
R48 X.n0 X.t0 26.5955
R49 X.n1 X.t3 26.5955
R50 X.n1 X.t2 26.5955
R51 X.n4 X.t5 24.9236
R52 X.n4 X.t7 24.9236
R53 X.n3 X.t4 24.9236
R54 X.n3 X.t6 24.9236
R55 VPWR.n11 VPWR.n5 599.74
R56 VPWR.n8 VPWR.t3 343.545
R57 VPWR.n19 VPWR.n1 311.973
R58 VPWR.n7 VPWR.n6 310.502
R59 VPWR.n1 VPWR.t0 37.4305
R60 VPWR.n13 VPWR.n12 34.6358
R61 VPWR.n13 VPWR.n2 34.6358
R62 VPWR.n17 VPWR.n2 34.6358
R63 VPWR.n18 VPWR.n17 34.6358
R64 VPWR.n12 VPWR.n11 32.0005
R65 VPWR.n1 VPWR.t6 26.5955
R66 VPWR.n5 VPWR.t4 26.5955
R67 VPWR.n5 VPWR.t1 26.5955
R68 VPWR.n6 VPWR.t2 26.5955
R69 VPWR.n6 VPWR.t5 26.5955
R70 VPWR.n10 VPWR.n7 25.977
R71 VPWR.n19 VPWR.n18 24.8476
R72 VPWR.n11 VPWR.n10 12.424
R73 VPWR.n10 VPWR.n9 9.3005
R74 VPWR.n11 VPWR.n4 9.3005
R75 VPWR.n12 VPWR.n3 9.3005
R76 VPWR.n14 VPWR.n13 9.3005
R77 VPWR.n15 VPWR.n2 9.3005
R78 VPWR.n17 VPWR.n16 9.3005
R79 VPWR.n18 VPWR.n0 9.3005
R80 VPWR.n20 VPWR.n19 7.12063
R81 VPWR.n8 VPWR.n7 6.18988
R82 VPWR.n9 VPWR.n8 0.755914
R83 VPWR.n20 VPWR.n0 0.148519
R84 VPWR.n9 VPWR.n4 0.120292
R85 VPWR.n4 VPWR.n3 0.120292
R86 VPWR.n14 VPWR.n3 0.120292
R87 VPWR.n15 VPWR.n14 0.120292
R88 VPWR.n16 VPWR.n15 0.120292
R89 VPWR.n16 VPWR.n0 0.120292
R90 VPWR VPWR.n20 0.11354
R91 S S.n1 351.533
R92 S.n1 S.t2 241.536
R93 S.n0 S.t0 212.081
R94 S.n1 S.t3 169.237
R95 S.n0 S.t1 139.78
R96 S S.n0 102.284
R97 a_314_297.t0 a_314_297.t1 1560.26
R98 a_27_47.t0 a_27_47.n1 342.377
R99 a_27_47.n1 a_27_47.t1 287.978
R100 a_27_47.n0 a_27_47.t2 241.536
R101 a_27_47.n1 a_27_47.n0 226.166
R102 a_27_47.n0 a_27_47.t3 169.237
R103 A0.n0 A0.t0 229.754
R104 A0.n0 A0.t1 157.453
R105 A0.n1 A0.n0 152
R106 A0.n1 A0 13.5116
R107 A0 A0.n1 2.60791
R108 VGND.n7 VGND.t3 289.265
R109 VGND.n6 VGND.n5 199.739
R110 VGND.n10 VGND.n4 199.739
R111 VGND.n19 VGND.n18 199.739
R112 VGND.n18 VGND.t0 36.9236
R113 VGND.n12 VGND.n11 34.6358
R114 VGND.n12 VGND.n1 34.6358
R115 VGND.n16 VGND.n1 34.6358
R116 VGND.n17 VGND.n16 34.6358
R117 VGND.n11 VGND.n10 32.0005
R118 VGND.n6 VGND.n3 25.977
R119 VGND.n5 VGND.t5 24.9236
R120 VGND.n5 VGND.t4 24.9236
R121 VGND.n4 VGND.t6 24.9236
R122 VGND.n4 VGND.t2 24.9236
R123 VGND.n18 VGND.t1 24.9236
R124 VGND.n19 VGND.n17 22.9652
R125 VGND.n10 VGND.n3 12.424
R126 VGND.n8 VGND.n3 9.3005
R127 VGND.n10 VGND.n9 9.3005
R128 VGND.n11 VGND.n2 9.3005
R129 VGND.n13 VGND.n12 9.3005
R130 VGND.n14 VGND.n1 9.3005
R131 VGND.n16 VGND.n15 9.3005
R132 VGND.n17 VGND.n0 9.3005
R133 VGND.n20 VGND.n19 7.12063
R134 VGND.n7 VGND.n6 6.18988
R135 VGND.n8 VGND.n7 0.755914
R136 VGND.n20 VGND.n0 0.148519
R137 VGND.n9 VGND.n8 0.120292
R138 VGND.n9 VGND.n2 0.120292
R139 VGND.n13 VGND.n2 0.120292
R140 VGND.n14 VGND.n13 0.120292
R141 VGND.n15 VGND.n14 0.120292
R142 VGND.n15 VGND.n0 0.120292
R143 VGND VGND.n20 0.11354
R144 a_206_47.t0 a_206_47.t1 147.692
R145 VNB.t1 VNB.t3 2833.66
R146 VNB.t0 VNB.t4 2705.5
R147 VNB.t2 VNB.t0 1381.23
R148 VNB.t4 VNB.t1 1338.51
R149 VNB.t7 VNB.t5 1196.12
R150 VNB.t6 VNB.t7 1196.12
R151 VNB.t8 VNB.t6 1196.12
R152 VNB.t3 VNB.t8 1196.12
R153 VNB VNB.t2 911.327
R154 a_490_47.t0 a_490_47.t1 156
C0 VPB VGND 0.011308f
C1 S X 0.001879f
C2 A0 VPWR 0.011515f
C3 S VGND 0.132851f
C4 A0 X 5.48e-20
C5 A1 VPWR 0.009275f
C6 A1 X 8.93e-20
C7 A0 VGND 0.015119f
C8 VPWR X 0.299151f
C9 A1 VGND 0.010789f
C10 VPWR VGND 0.107914f
C11 X VGND 0.221702f
C12 VPB S 0.08369f
C13 VPB A0 0.047471f
C14 S A0 0.03575f
C15 VPB A1 0.03248f
C16 S A1 0.094243f
C17 VPB VPWR 0.11878f
C18 S VPWR 0.040338f
C19 VPB X 0.011848f
C20 A0 A1 0.081182f
C21 VGND VNB 0.632032f
C22 X VNB 0.075034f
C23 VPWR VNB 0.536034f
C24 A1 VNB 0.098044f
C25 A0 VNB 0.115452f
C26 S VNB 0.264681f
C27 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_8 S A1 VPWR VGND VPB VNB A0 X
X0 VGND.t11 a_79_21.t8 X.t15 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t10 a_79_21.t9 X.t14 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_79_21.t2 A0.t0 a_792_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.5375 ps=2.075 w=1 l=0.15
X3 X.t7 a_79_21.t10 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t11 a_79_21.t11 X.t6 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1259_199.t0 S.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11325 ps=1 w=0.65 l=0.15
X6 X.t5 a_79_21.t12 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1302_47.t1 A0.t1 a_79_21.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.336 pd=1.69 as=0.0864 ps=0.91 w=0.64 l=0.15
X8 VPWR.t9 a_79_21.t13 X.t4 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_792_297.t0 S.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.5375 pd=2.075 as=0.1625 ps=1.325 w=1 l=0.15
X10 a_1259_199.t1 S.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X11 VGND.t9 a_79_21.t14 X.t13 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t8 a_79_21.t15 X.t12 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t12 a_1259_199.t2 a_1302_47.t3 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.11325 pd=1 as=0.336 ps=1.69 w=0.64 l=0.15
X14 a_79_21.t7 A1.t0 a_792_47.t3 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0944 ps=0.935 w=0.64 l=0.15
X15 a_79_21.t5 A0.t2 a_1302_47.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.1552 ps=1.125 w=0.64 l=0.15
X16 VPWR.t8 a_79_21.t16 X.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR.t2 S.t3 a_792_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1675 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X18 X.t11 a_79_21.t17 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_792_297.t2 A0.t3 a_79_21.t6 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 X.t10 a_79_21.t18 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 X.t2 a_79_21.t19 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1302_47.t2 a_1259_199.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1552 pd=1.125 as=0.1072 ps=0.975 w=0.64 l=0.15
X23 VPWR.t3 a_1259_199.t4 a_1302_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X24 X.t9 a_79_21.t20 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_1302_297.t0 a_1259_199.t5 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.6325 pd=2.265 as=0.1675 ps=1.335 w=1 l=0.15
X26 a_792_47.t2 A1.t1 a_79_21.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.336 pd=1.69 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 VPWR.t6 a_79_21.t21 X.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1302_297.t3 A1.t2 a_79_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND.t1 S.t4 a_792_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1072 pd=0.975 as=0.336 ps=1.69 w=0.64 l=0.15
X30 X.t0 a_79_21.t22 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 a_79_21.t4 A1.t3 a_1302_297.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.6325 ps=2.265 w=1 l=0.15
X32 X.t8 a_79_21.t23 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X33 a_792_47.t0 S.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0944 pd=0.935 as=0.10525 ps=0.975 w=0.64 l=0.15
R0 a_79_21.n27 a_79_21.n26 791.307
R1 a_79_21.n26 a_79_21.n25 585
R2 a_79_21.n2 a_79_21.n0 257.908
R3 a_79_21.n4 a_79_21.t16 205.654
R4 a_79_21.n21 a_79_21.t19 205.654
R5 a_79_21.n19 a_79_21.t21 205.654
R6 a_79_21.n7 a_79_21.t10 205.654
R7 a_79_21.n13 a_79_21.t11 205.654
R8 a_79_21.n11 a_79_21.t12 205.654
R9 a_79_21.n9 a_79_21.t13 205.654
R10 a_79_21.n8 a_79_21.t22 205.654
R11 a_79_21.n2 a_79_21.n1 185
R12 a_79_21.n26 a_79_21.n24 178.447
R13 a_79_21.n10 a_79_21.n6 177.601
R14 a_79_21.n12 a_79_21.n6 152
R15 a_79_21.n15 a_79_21.n14 152
R16 a_79_21.n16 a_79_21.n5 152
R17 a_79_21.n18 a_79_21.n17 152
R18 a_79_21.n20 a_79_21.n3 152
R19 a_79_21.n23 a_79_21.n22 152
R20 a_79_21.n4 a_79_21.t9 139.78
R21 a_79_21.n21 a_79_21.t20 139.78
R22 a_79_21.n19 a_79_21.t8 139.78
R23 a_79_21.n7 a_79_21.t18 139.78
R24 a_79_21.n13 a_79_21.t15 139.78
R25 a_79_21.n11 a_79_21.t17 139.78
R26 a_79_21.n9 a_79_21.t14 139.78
R27 a_79_21.n8 a_79_21.t23 139.78
R28 a_79_21.n24 a_79_21.n2 95.624
R29 a_79_21.n9 a_79_21.n8 57.8405
R30 a_79_21.n18 a_79_21.n5 46.8234
R31 a_79_21.n14 a_79_21.n7 44.0691
R32 a_79_21.n20 a_79_21.n19 38.5605
R33 a_79_21.n10 a_79_21.n9 35.8062
R34 a_79_21.n13 a_79_21.n12 33.0519
R35 a_79_21.n22 a_79_21.n4 30.2976
R36 a_79_21.n22 a_79_21.n21 27.5434
R37 a_79_21.n25 a_79_21.t6 26.5955
R38 a_79_21.n25 a_79_21.t2 26.5955
R39 a_79_21.t1 a_79_21.n27 26.5955
R40 a_79_21.n27 a_79_21.t4 26.5955
R41 a_79_21.n24 a_79_21.n23 26.3534
R42 a_79_21.n23 a_79_21.n3 25.6005
R43 a_79_21.n17 a_79_21.n3 25.6005
R44 a_79_21.n17 a_79_21.n16 25.6005
R45 a_79_21.n16 a_79_21.n15 25.6005
R46 a_79_21.n15 a_79_21.n6 25.6005
R47 a_79_21.n1 a_79_21.t0 25.313
R48 a_79_21.n1 a_79_21.t7 25.313
R49 a_79_21.n0 a_79_21.t3 25.313
R50 a_79_21.n0 a_79_21.t5 25.313
R51 a_79_21.n12 a_79_21.n11 24.7891
R52 a_79_21.n11 a_79_21.n10 22.0348
R53 a_79_21.n21 a_79_21.n20 19.2805
R54 a_79_21.n14 a_79_21.n13 13.7719
R55 a_79_21.n19 a_79_21.n18 8.26336
R56 a_79_21.n7 a_79_21.n5 2.75479
R57 X.n3 X.n2 378.199
R58 X.n6 X.n5 319.899
R59 X.n3 X.n1 314.952
R60 X.n4 X.n0 314.952
R61 X.n10 X.n9 261.425
R62 X.n13 X.n12 206.135
R63 X.n10 X.n8 201.189
R64 X.n11 X.n7 198.177
R65 X.n4 X.n3 63.2476
R66 X.n11 X.n10 63.2476
R67 X.n6 X.n4 53.0829
R68 X.n13 X.n11 53.0829
R69 X X.n6 32.2914
R70 X.n2 X.t3 26.5955
R71 X.n2 X.t2 26.5955
R72 X.n1 X.t1 26.5955
R73 X.n1 X.t7 26.5955
R74 X.n0 X.t6 26.5955
R75 X.n0 X.t5 26.5955
R76 X.n5 X.t4 26.5955
R77 X.n5 X.t0 26.5955
R78 X.n7 X.t12 24.9236
R79 X.n7 X.t11 24.9236
R80 X.n8 X.t15 24.9236
R81 X.n8 X.t10 24.9236
R82 X.n9 X.t14 24.9236
R83 X.n9 X.t9 24.9236
R84 X.n12 X.t13 24.9236
R85 X.n12 X.t8 24.9236
R86 X X.n13 22.4005
R87 VGND.n34 VGND.t4 282.596
R88 VGND.n8 VGND.n7 206.168
R89 VGND.n10 VGND.n9 199.739
R90 VGND.n18 VGND.n17 199.739
R91 VGND.n25 VGND.n24 199.739
R92 VGND.n28 VGND.n27 199.739
R93 VGND.n32 VGND.n2 199.739
R94 VGND.n7 VGND.t12 40.313
R95 VGND.n9 VGND.t1 37.5005
R96 VGND.n17 VGND.t2 35.6255
R97 VGND.n11 VGND.n6 34.6358
R98 VGND.n15 VGND.n6 34.6358
R99 VGND.n16 VGND.n15 34.6358
R100 VGND.n19 VGND.n16 34.6358
R101 VGND.n23 VGND.n4 34.6358
R102 VGND.n28 VGND.n26 32.0005
R103 VGND.n32 VGND.n1 25.977
R104 VGND.n9 VGND.t3 25.313
R105 VGND.n24 VGND.t5 24.9236
R106 VGND.n24 VGND.t11 24.9236
R107 VGND.n27 VGND.t6 24.9236
R108 VGND.n27 VGND.t8 24.9236
R109 VGND.n2 VGND.t7 24.9236
R110 VGND.n2 VGND.t9 24.9236
R111 VGND.n11 VGND.n10 23.3417
R112 VGND.n7 VGND.t0 22.1675
R113 VGND.n17 VGND.t10 22.1675
R114 VGND.n34 VGND.n33 19.9534
R115 VGND.n33 VGND.n32 18.4476
R116 VGND.n28 VGND.n1 12.424
R117 VGND.n19 VGND.n18 9.41227
R118 VGND.n35 VGND.n34 9.3005
R119 VGND.n12 VGND.n11 9.3005
R120 VGND.n13 VGND.n6 9.3005
R121 VGND.n15 VGND.n14 9.3005
R122 VGND.n16 VGND.n5 9.3005
R123 VGND.n20 VGND.n19 9.3005
R124 VGND.n21 VGND.n4 9.3005
R125 VGND.n23 VGND.n22 9.3005
R126 VGND.n26 VGND.n3 9.3005
R127 VGND.n29 VGND.n28 9.3005
R128 VGND.n30 VGND.n1 9.3005
R129 VGND.n32 VGND.n31 9.3005
R130 VGND.n33 VGND.n0 9.3005
R131 VGND.n10 VGND.n8 6.99647
R132 VGND.n26 VGND.n25 6.4005
R133 VGND.n25 VGND.n23 3.38874
R134 VGND.n18 VGND.n4 0.376971
R135 VGND.n12 VGND.n8 0.157005
R136 VGND.n13 VGND.n12 0.120292
R137 VGND.n14 VGND.n13 0.120292
R138 VGND.n14 VGND.n5 0.120292
R139 VGND.n20 VGND.n5 0.120292
R140 VGND.n21 VGND.n20 0.120292
R141 VGND.n22 VGND.n21 0.120292
R142 VGND.n22 VGND.n3 0.120292
R143 VGND.n29 VGND.n3 0.120292
R144 VGND.n30 VGND.n29 0.120292
R145 VGND.n31 VGND.n30 0.120292
R146 VGND.n31 VGND.n0 0.120292
R147 VGND.n35 VGND.n0 0.120292
R148 VGND VGND.n35 0.0213333
R149 VNB.t5 VNB.t15 3417.48
R150 VNB.t3 VNB.t1 3417.48
R151 VNB.t4 VNB.t14 1808.41
R152 VNB.t15 VNB.t0 1423.95
R153 VNB.t1 VNB.t4 1381.23
R154 VNB.t12 VNB.t2 1352.75
R155 VNB.t2 VNB.t16 1267.31
R156 VNB.t14 VNB.t5 1196.12
R157 VNB.t16 VNB.t3 1196.12
R158 VNB.t7 VNB.t12 1196.12
R159 VNB.t13 VNB.t7 1196.12
R160 VNB.t8 VNB.t13 1196.12
R161 VNB.t10 VNB.t8 1196.12
R162 VNB.t9 VNB.t10 1196.12
R163 VNB.t11 VNB.t9 1196.12
R164 VNB.t6 VNB.t11 1196.12
R165 VNB VNB.t6 911.327
R166 A0.n2 A0.n0 279.625
R167 A0.n1 A0.t3 215.546
R168 A0.n2 A0.n1 202.825
R169 A0.n1 A0.t0 202.769
R170 A0.n0 A0.t1 180.321
R171 A0.n0 A0.t2 135.423
R172 A0 A0.n2 4.81418
R173 a_792_297.n1 a_792_297.n0 1291.98
R174 a_792_297.n0 a_792_297.t3 180.256
R175 a_792_297.n0 a_792_297.t0 31.5205
R176 a_792_297.n1 a_792_297.t1 26.5955
R177 a_792_297.t2 a_792_297.n1 26.5955
R178 VPB.t7 VPB.t8 837.539
R179 VPB.t0 VPB.t4 725.078
R180 VPB.t6 VPB.t1 295.95
R181 VPB.t2 VPB.t7 287.072
R182 VPB.t12 VPB.t0 281.154
R183 VPB.t5 VPB.t6 248.599
R184 VPB.t8 VPB.t5 248.599
R185 VPB.t3 VPB.t2 248.599
R186 VPB.t4 VPB.t3 248.599
R187 VPB.t11 VPB.t12 248.599
R188 VPB.t10 VPB.t11 248.599
R189 VPB.t16 VPB.t10 248.599
R190 VPB.t15 VPB.t16 248.599
R191 VPB.t14 VPB.t15 248.599
R192 VPB.t13 VPB.t14 248.599
R193 VPB.t9 VPB.t13 248.599
R194 VPB VPB.t9 189.409
R195 VPWR.n14 VPWR.n13 607.212
R196 VPWR.n12 VPWR.n11 606.178
R197 VPWR.n8 VPWR.n7 599.74
R198 VPWR.n34 VPWR.t5 336.827
R199 VPWR.n32 VPWR.n2 310.502
R200 VPWR.n4 VPWR.n3 310.502
R201 VPWR.n26 VPWR.n6 310.502
R202 VPWR.n11 VPWR.t3 42.3555
R203 VPWR.n13 VPWR.t4 39.4005
R204 VPWR.n7 VPWR.t0 37.4305
R205 VPWR.n25 VPWR.n24 34.6358
R206 VPWR.n15 VPWR.n10 34.6358
R207 VPWR.n19 VPWR.n10 34.6358
R208 VPWR.n20 VPWR.n19 34.6358
R209 VPWR.n21 VPWR.n20 34.6358
R210 VPWR.n27 VPWR.n4 32.0005
R211 VPWR.n15 VPWR.n14 30.8711
R212 VPWR.n2 VPWR.t10 26.5955
R213 VPWR.n2 VPWR.t9 26.5955
R214 VPWR.n3 VPWR.t12 26.5955
R215 VPWR.n3 VPWR.t11 26.5955
R216 VPWR.n6 VPWR.t7 26.5955
R217 VPWR.n6 VPWR.t6 26.5955
R218 VPWR.n7 VPWR.t8 26.5955
R219 VPWR.n13 VPWR.t2 26.5955
R220 VPWR.n11 VPWR.t1 26.5955
R221 VPWR.n32 VPWR.n31 25.977
R222 VPWR.n34 VPWR.n33 19.9534
R223 VPWR.n33 VPWR.n32 18.4476
R224 VPWR.n31 VPWR.n4 12.424
R225 VPWR.n14 VPWR.n12 11.3655
R226 VPWR.n21 VPWR.n8 9.41227
R227 VPWR.n16 VPWR.n15 9.3005
R228 VPWR.n17 VPWR.n10 9.3005
R229 VPWR.n19 VPWR.n18 9.3005
R230 VPWR.n20 VPWR.n9 9.3005
R231 VPWR.n22 VPWR.n21 9.3005
R232 VPWR.n24 VPWR.n23 9.3005
R233 VPWR.n25 VPWR.n5 9.3005
R234 VPWR.n28 VPWR.n27 9.3005
R235 VPWR.n29 VPWR.n4 9.3005
R236 VPWR.n31 VPWR.n30 9.3005
R237 VPWR.n32 VPWR.n1 9.3005
R238 VPWR.n33 VPWR.n0 9.3005
R239 VPWR.n35 VPWR.n34 9.3005
R240 VPWR.n27 VPWR.n26 6.4005
R241 VPWR.n26 VPWR.n25 3.38874
R242 VPWR.n24 VPWR.n8 0.376971
R243 VPWR.n16 VPWR.n12 0.147508
R244 VPWR.n17 VPWR.n16 0.120292
R245 VPWR.n18 VPWR.n17 0.120292
R246 VPWR.n18 VPWR.n9 0.120292
R247 VPWR.n22 VPWR.n9 0.120292
R248 VPWR.n23 VPWR.n22 0.120292
R249 VPWR.n23 VPWR.n5 0.120292
R250 VPWR.n28 VPWR.n5 0.120292
R251 VPWR.n29 VPWR.n28 0.120292
R252 VPWR.n30 VPWR.n29 0.120292
R253 VPWR.n30 VPWR.n1 0.120292
R254 VPWR.n1 VPWR.n0 0.120292
R255 VPWR.n35 VPWR.n0 0.120292
R256 VPWR VPWR.n35 0.0213333
R257 S.n3 S.n1 313.753
R258 S.n2 S.t3 241.536
R259 S.n1 S.t1 241
R260 S.n0 S.t2 236.934
R261 S S.n0 177.4
R262 S.n2 S.t4 170.843
R263 S.n1 S.t5 170.308
R264 S.n3 S.n2 164.976
R265 S.n0 S.t0 164.633
R266 S S.n3 12.4298
R267 a_1259_199.t1 a_1259_199.n3 389.348
R268 a_1259_199.n3 a_1259_199.n2 353.413
R269 a_1259_199.n1 a_1259_199.t0 297.264
R270 a_1259_199.n0 a_1259_199.t4 239.505
R271 a_1259_199.n2 a_1259_199.t5 235.821
R272 a_1259_199.n0 a_1259_199.t2 168.811
R273 a_1259_199.n2 a_1259_199.t3 165.127
R274 a_1259_199.n1 a_1259_199.n0 152
R275 a_1259_199.n3 a_1259_199.n1 25.224
R276 a_1302_47.n1 a_1302_47.n0 442.283
R277 a_1302_47.n1 a_1302_47.t3 171.562
R278 a_1302_47.n0 a_1302_47.t0 47.813
R279 a_1302_47.n0 a_1302_47.t2 43.1255
R280 a_1302_47.t1 a_1302_47.n1 25.313
R281 A1.n0 A1.t3 220.772
R282 A1.n0 A1.t2 197.543
R283 A1.n1 A1.t1 177.68
R284 A1 A1.n1 166.506
R285 A1 A1.n0 165.808
R286 A1.n1 A1.t0 138.064
R287 a_792_47.n1 a_792_47.n0 433.248
R288 a_792_47.t1 a_792_47.n1 171.562
R289 a_792_47.n0 a_792_47.t0 30.0005
R290 a_792_47.n0 a_792_47.t3 25.313
R291 a_792_47.n1 a_792_47.t2 25.313
R292 a_1302_297.n1 a_1302_297.n0 1308.16
R293 a_1302_297.n0 a_1302_297.t2 222.611
R294 a_1302_297.n0 a_1302_297.t0 26.5955
R295 a_1302_297.t1 a_1302_297.n1 26.5955
R296 a_1302_297.n1 a_1302_297.t3 26.5955
C0 VGND X 0.389518f
C1 VPB A0 0.088435f
C2 S A0 0.164422f
C3 VPB A1 0.090738f
C4 S A1 0.39222f
C5 VPB VPWR 0.18344f
C6 VPB X 0.014424f
C7 S VPWR 0.213383f
C8 A0 A1 0.118497f
C9 A0 VPWR 0.019456f
C10 S X 0.001709f
C11 A0 X 0.00226f
C12 A1 VPWR 0.058061f
C13 VGND VPB 0.009144f
C14 A1 X 3.67e-19
C15 VGND S 0.086288f
C16 VPWR X 0.590589f
C17 VGND A0 0.122959f
C18 VGND A1 0.061491f
C19 VGND VPWR 0.098398f
C20 VPB S 0.116855f
C21 VGND VNB 1.05453f
C22 X VNB 0.077793f
C23 VPWR VNB 0.880479f
C24 A1 VNB 0.266859f
C25 A0 VNB 0.267924f
C26 S VNB 0.353746f
C27 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2i_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2i_1 VPB VNB VGND VPWR A0 Y A1 S
X0 a_27_297.t1 S.t0 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=1.6 w=1 l=0.15
X1 VGND.t1 S.t1 a_283_205.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_204_297.t1 A1.t0 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.395 as=0.1525 ps=1.305 w=1 l=0.15
X3 a_193_47.t0 A1.t1 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t0 A0.t0 a_27_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.28 ps=2.56 w=1 l=0.15
X5 VPWR.t0 a_283_205.t2 a_204_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=1.6 as=0.1975 ps=1.395 w=1 l=0.15
X6 VPWR.t2 S.t2 a_283_205.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.29 ps=2.58 w=1 l=0.15
X7 VGND.t0 a_283_205.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_193_47.t1 S.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t1 A0.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 S.n1 S.t2 234.573
R1 S.n1 S.n0 225.369
R2 S.n0 S.t0 211.863
R3 S.n0 S.t3 194.407
R4 S.n2 S.t1 191.194
R5 S.n3 S.n2 173.583
R6 S.n2 S.n1 32.1338
R7 S.n3 S 10.8901
R8 S S.n3 2.10199
R9 VPWR.n1 VPWR.t2 346.673
R10 VPWR.n1 VPWR.n0 326.284
R11 VPWR.n0 VPWR.t1 65.9955
R12 VPWR.n0 VPWR.t0 52.2055
R13 VPWR VPWR.n1 0.488797
R14 a_27_297.t0 a_27_297.t1 653.557
R15 VPB.t4 VPB.t3 574.144
R16 VPB.t1 VPB.t4 443.925
R17 VPB.t0 VPB.t1 322.587
R18 VPB.t2 VPB.t0 269.315
R19 VPB VPB.t2 204.207
R20 a_283_205.t1 a_283_205.n1 255.047
R21 a_283_205.n0 a_283_205.t2 237.787
R22 a_283_205.n1 a_283_205.n0 218.452
R23 a_283_205.n0 a_283_205.t3 197.62
R24 a_283_205.n1 a_283_205.t0 155.744
R25 VGND.n1 VGND.t1 297.724
R26 VGND.n1 VGND.n0 214.089
R27 VGND.n0 VGND.t2 24.9236
R28 VGND.n0 VGND.t0 24.9236
R29 VGND VGND.n1 0.5538
R30 VNB.t2 VNB.t0 2733.98
R31 VNB.t3 VNB.t4 2677.02
R32 VNB.t0 VNB.t3 1196.12
R33 VNB.t1 VNB.t2 1196.12
R34 VNB VNB.t1 925.567
R35 A1.n0 A1.t0 234.173
R36 A1 A1.n0 169.483
R37 A1.n0 A1.t1 161.873
R38 Y Y.n0 593.961
R39 Y.n2 Y.n0 585
R40 Y.n2 Y.n1 240.269
R41 Y.n0 Y.t2 33.4905
R42 Y.n0 Y.t0 26.5955
R43 Y.n1 Y.t3 24.9236
R44 Y.n1 Y.t1 24.9236
R45 Y Y.n2 8.4485
R46 a_204_297.t0 a_204_297.t1 77.8155
R47 a_193_47.t0 a_193_47.t1 576.511
R48 A0.n0 A0.t1 1554.35
R49 A0.n0 A0.t0 229.369
R50 A0 A0.n0 158.258
R51 a_27_47.t0 a_27_47.t1 491.416
C0 A0 VPWR 0.010531f
C1 A1 Y 0.103049f
C2 A0 VGND 0.010876f
C3 A1 VPWR 0.013451f
C4 S Y 1.79e-19
C5 A1 VGND 0.011828f
C6 S VPWR 0.072039f
C7 S VGND 0.062246f
C8 Y VPWR 0.008136f
C9 A0 VPB 0.039826f
C10 Y VGND 0.007539f
C11 A1 VPB 0.035899f
C12 VPWR VGND 0.073802f
C13 S VPB 0.113347f
C14 Y VPB 0.003301f
C15 VPWR VPB 0.087399f
C16 A0 A1 0.050532f
C17 VGND VPB 0.007946f
C18 A1 S 6.46e-19
C19 A0 Y 0.036639f
C20 VGND VNB 0.453067f
C21 VPWR VNB 0.388182f
C22 Y VNB 0.016962f
C23 S VNB 0.319014f
C24 A1 VNB 0.104015f
C25 A0 VNB 0.143714f
C26 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2i_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2i_2 VNB VPB VPWR VGND S A0 A1 Y
X0 a_361_47.t3 A0.t0 Y.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y.t5 A0.t1 a_193_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t2 a_27_47.t2 a_361_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_361_297.t2 a_27_47.t3 VPWR.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t4 S.t0 a_193_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t7 A0.t2 a_361_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_193_297.t2 S.t1 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_361_297.t0 A1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.155 ps=1.31 w=1 l=0.15
X8 a_193_47.t3 S.t2 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_361_47.t0 a_27_47.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_193_297.t0 A0.t3 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y.t1 A1.t1 a_361_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.455 pd=2.91 as=0.1375 ps=1.275 w=1 l=0.15
X12 Y.t2 A1.t2 a_193_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.29575 pd=2.21 as=0.089375 ps=0.925 w=0.65 l=0.15
X13 VGND.t4 S.t3 a_193_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t0 a_27_47.t5 a_361_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_193_47.t0 A1.t3 Y.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.10075 ps=0.96 w=0.65 l=0.15
X16 VPWR.t0 S.t4 a_27_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VGND.t3 S.t5 a_27_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A0.n1 A0.t1 212.081
R1 A0.n4 A0.t3 212.081
R2 A0.n3 A0.n2 206.627
R3 A0.n6 A0.n5 152
R4 A0.n3 A0.n0 152
R5 A0.n1 A0.t2 139.78
R6 A0.n4 A0.t0 139.78
R7 A0.n5 A0.n4 32.8641
R8 A0.n5 A0.n1 28.4823
R9 A0.n6 A0.n0 21.7605
R10 A0.n2 A0 18.8805
R11 A0.n4 A0.n3 17.3817
R12 A0.n2 A0 10.5605
R13 A0 A0.n6 4.8005
R14 A0 A0.n0 2.8805
R15 Y.n1 Y.t4 918.735
R16 Y.n2 Y.t1 738.703
R17 Y.n1 Y.n0 585
R18 Y.n4 Y.t6 331.325
R19 Y.n5 Y.t2 245.923
R20 Y.n4 Y.n3 185
R21 Y Y.n5 106.165
R22 Y.n5 Y.n4 81.3181
R23 Y.n2 Y.n1 65.5064
R24 Y.n3 Y.t3 32.3082
R25 Y.n0 Y.t0 30.5355
R26 Y.n0 Y.t5 30.5355
R27 Y.n3 Y.t7 24.9236
R28 Y Y.n2 22.7728
R29 a_361_47.n1 a_361_47.n0 489.13
R30 a_361_47.n0 a_361_47.t1 24.9236
R31 a_361_47.n0 a_361_47.t0 24.9236
R32 a_361_47.t2 a_361_47.n1 24.9236
R33 a_361_47.n1 a_361_47.t3 24.9236
R34 VNB.t3 VNB.t6 2677.02
R35 VNB.t5 VNB.t1 1310.03
R36 VNB.t1 VNB.t0 1210.36
R37 VNB.t6 VNB.t5 1196.12
R38 VNB.t2 VNB.t3 1196.12
R39 VNB.t4 VNB.t2 1196.12
R40 VNB.t7 VNB.t4 1196.12
R41 VNB.t8 VNB.t7 1196.12
R42 VNB VNB.t8 911.327
R43 a_193_297.n1 a_193_297.n0 1345.62
R44 a_193_297.n0 a_193_297.t3 26.5955
R45 a_193_297.n0 a_193_297.t2 26.5955
R46 a_193_297.t1 a_193_297.n1 26.5955
R47 a_193_297.n1 a_193_297.t0 26.5955
R48 VPB.t7 VPB.t3 556.386
R49 VPB.t4 VPB.t0 272.274
R50 VPB.t0 VPB.t1 251.559
R51 VPB.t3 VPB.t4 248.599
R52 VPB.t8 VPB.t7 248.599
R53 VPB.t6 VPB.t8 248.599
R54 VPB.t5 VPB.t6 248.599
R55 VPB.t2 VPB.t5 248.599
R56 VPB VPB.t2 189.409
R57 a_27_47.t0 a_27_47.n3 872.39
R58 a_27_47.n3 a_27_47.t1 288.187
R59 a_27_47.n3 a_27_47.n2 278.284
R60 a_27_47.n0 a_27_47.t2 212.081
R61 a_27_47.n1 a_27_47.t3 212.081
R62 a_27_47.n0 a_27_47.t5 149.421
R63 a_27_47.n1 a_27_47.t4 149.421
R64 a_27_47.n2 a_27_47.n0 53.0205
R65 a_27_47.n2 a_27_47.n1 14.4605
R66 a_361_297.n1 a_361_297.n0 1349.97
R67 a_361_297.t0 a_361_297.n1 27.5805
R68 a_361_297.n0 a_361_297.t3 26.5955
R69 a_361_297.n0 a_361_297.t2 26.5955
R70 a_361_297.n1 a_361_297.t1 26.5955
R71 VPWR.n2 VPWR.t2 879.044
R72 VPWR.n6 VPWR.n1 599.74
R73 VPWR.n4 VPWR.n3 599.74
R74 VPWR.n1 VPWR.t3 26.5955
R75 VPWR.n1 VPWR.t0 26.5955
R76 VPWR.n3 VPWR.t1 26.5955
R77 VPWR.n3 VPWR.t4 26.5955
R78 VPWR.n6 VPWR.n5 22.9652
R79 VPWR.n5 VPWR.n4 15.4358
R80 VPWR.n5 VPWR.n0 9.3005
R81 VPWR.n7 VPWR.n6 7.12063
R82 VPWR.n4 VPWR.n2 6.88313
R83 VPWR.n2 VPWR.n0 0.619932
R84 VPWR.n7 VPWR.n0 0.148519
R85 VPWR VPWR.n7 0.11354
R86 S.n0 S.t0 212.081
R87 S.n1 S.t1 212.081
R88 S.n2 S.t4 212.081
R89 S S.n3 155.685
R90 S.n0 S.t3 139.78
R91 S.n1 S.t2 139.78
R92 S.n2 S.t5 139.78
R93 S.n1 S.n0 61.346
R94 S.n3 S.n1 54.7732
R95 S.n3 S.n2 6.57323
R96 A1.n1 A1.t1 212.081
R97 A1.n0 A1.t0 212.081
R98 A1.n2 A1.n1 174.639
R99 A1.n1 A1.t2 139.78
R100 A1.n0 A1.t3 139.78
R101 A1.n1 A1.n0 62.0763
R102 A1.n2 A1 11.2251
R103 A1 A1.n2 2.16665
R104 VGND.n1 VGND.t0 301.7
R105 VGND.n6 VGND.n5 200.201
R106 VGND.n3 VGND.n2 116.112
R107 VGND.n2 VGND.t1 24.9236
R108 VGND.n2 VGND.t4 24.9236
R109 VGND.n5 VGND.t2 24.9236
R110 VGND.n5 VGND.t3 24.9236
R111 VGND.n6 VGND.n4 23.7181
R112 VGND.n4 VGND.n3 21.4593
R113 VGND.n4 VGND.n0 9.3005
R114 VGND.n7 VGND.n6 7.12063
R115 VGND.n3 VGND.n1 6.65102
R116 VGND.n1 VGND.n0 0.892006
R117 VGND.n7 VGND.n0 0.148519
R118 VGND VGND.n7 0.11354
R119 a_193_47.n1 a_193_47.n0 410.267
R120 a_193_47.t1 a_193_47.n1 25.8467
R121 a_193_47.n0 a_193_47.t2 24.9236
R122 a_193_47.n0 a_193_47.t3 24.9236
R123 a_193_47.n1 a_193_47.t0 24.9236
C0 A0 A1 0.057658f
C1 A0 VPB 0.085382f
C2 A0 VPWR 0.0186f
C3 A0 S 3.64e-19
C4 A1 VPB 0.07355f
C5 A1 VPWR 0.01686f
C6 A0 Y 0.032763f
C7 VPWR VPB 0.101697f
C8 A1 S 7.14e-19
C9 VPB S 0.087264f
C10 A0 VGND 0.013618f
C11 A1 Y 0.120815f
C12 VPWR S 0.051139f
C13 Y VPB 0.014943f
C14 VPWR Y 0.241738f
C15 A1 VGND 0.015967f
C16 VGND VPB 0.004732f
C17 Y S 3.9e-19
C18 VPWR VGND 0.039222f
C19 VGND S 0.082942f
C20 Y VGND 0.236205f
C21 VGND VNB 0.577021f
C22 Y VNB 0.107908f
C23 VPWR VNB 0.479572f
C24 A1 VNB 0.220681f
C25 A0 VNB 0.23234f
C26 S VNB 0.290862f
C27 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR.t0 A.t0 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t0 A.t1 a_113_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47.t1 B.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y.t2 B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R0 A.n0 A.t0 230.155
R1 A.n0 A.t1 157.856
R2 A A.n0 154.102
R3 Y Y.n0 237.577
R4 Y.n1 Y.t0 140.53
R5 Y.n0 Y.t1 26.5955
R6 Y.n0 Y.t2 26.5955
R7 Y.n1 Y 16.5652
R8 Y Y.n1 9.03579
R9 Y.n1 Y 1.72748
R10 VPWR.n0 VPWR.t0 256.344
R11 VPWR.n0 VPWR.t1 254.13
R12 VPWR VPWR.n0 0.493374
R13 VPB.t1 VPB.t0 248.599
R14 VPB VPB.t1 207.166
R15 a_113_47.t0 a_113_47.t1 49.8467
R16 VNB.t1 VNB.t0 1196.12
R17 VNB VNB.t1 996.764
R18 B.n0 B.t1 229.369
R19 B B.n0 157.927
R20 B.n0 B.t0 157.07
R21 VGND VGND.t0 158.046
C0 B Y 0.048071f
C1 VPB VGND 0.004396f
C2 B VGND 0.054404f
C3 A Y 0.085479f
C4 VPWR Y 0.211407f
C5 A VGND 0.009489f
C6 VPWR VGND 0.032185f
C7 Y VGND 0.138901f
C8 VPB B 0.039072f
C9 VPB A 0.037877f
C10 B A 0.050963f
C11 VPB VPWR 0.050862f
C12 B VPWR 0.047843f
C13 A VPWR 0.04444f
C14 VPB Y 0.006185f
C15 VGND VNB 0.23167f
C16 Y VNB 0.055661f
C17 VPWR VNB 0.245114f
C18 A VNB 0.143376f
C19 B VNB 0.145827f
C20 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_4 VPB VNB VGND VPWR B Y A
X0 a_27_47.t6 A.t0 Y.t10 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47.t5 A.t1 Y.t9 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t6 A.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t0 B.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t11 B.t1 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t1 B.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47.t0 B.t3 VGND.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47.t1 B.t4 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t5 A.t3 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t1 B.t5 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t8 A.t4 a_27_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y.t4 A.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y.t7 A.t6 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR.t3 A.t7 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t2 B.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t0 B.t7 a_27_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n1 A.t3 212.081
R1 A.n3 A.t5 212.081
R2 A.n5 A.t7 212.081
R3 A.n4 A.t2 212.081
R4 A A.n6 158.656
R5 A.n2 A.n0 152
R6 A.n1 A.t1 139.78
R7 A.n3 A.t6 139.78
R8 A.n5 A.t0 139.78
R9 A.n4 A.t4 139.78
R10 A.n5 A.n4 61.346
R11 A.n2 A.n1 30.6732
R12 A.n3 A.n2 30.6732
R13 A.n6 A.n3 30.6732
R14 A.n6 A.n5 30.6732
R15 A A.n0 14.8485
R16 A.n0 A 8.7045
R17 Y.n2 Y.n1 256.103
R18 Y.n5 Y.n3 243.68
R19 Y.n9 Y.n7 241.847
R20 Y.n5 Y.n4 205.28
R21 Y.n2 Y.n0 202.095
R22 Y.n9 Y.n8 185
R23 Y.n0 Y.t3 26.5955
R24 Y.n0 Y.t6 26.5955
R25 Y.n3 Y.t1 26.5955
R26 Y.n3 Y.t2 26.5955
R27 Y.n4 Y.t0 26.5955
R28 Y.n4 Y.t11 26.5955
R29 Y.n1 Y.t5 26.5955
R30 Y.n1 Y.t4 26.5955
R31 Y.n8 Y.t10 24.9236
R32 Y.n8 Y.t8 24.9236
R33 Y.n7 Y.t9 24.9236
R34 Y.n7 Y.t7 24.9236
R35 Y Y.n5 22.9652
R36 Y Y.n9 18.8943
R37 Y.n6 Y.n2 13.9299
R38 Y.n6 Y 13.9299
R39 Y Y.n6 1.19676
R40 a_27_47.n5 a_27_47.n4 185
R41 a_27_47.n4 a_27_47.t5 183.096
R42 a_27_47.n1 a_27_47.t7 172.548
R43 a_27_47.n1 a_27_47.n0 99.1759
R44 a_27_47.n3 a_27_47.n2 88.3446
R45 a_27_47.n4 a_27_47.n3 55.3569
R46 a_27_47.n3 a_27_47.n1 47.2798
R47 a_27_47.n2 a_27_47.t4 24.9236
R48 a_27_47.n2 a_27_47.t1 24.9236
R49 a_27_47.n0 a_27_47.t2 24.9236
R50 a_27_47.n0 a_27_47.t0 24.9236
R51 a_27_47.n5 a_27_47.t3 24.9236
R52 a_27_47.t6 a_27_47.n5 24.9236
R53 VNB.t3 VNB.t5 1196.12
R54 VNB.t6 VNB.t3 1196.12
R55 VNB.t4 VNB.t6 1196.12
R56 VNB.t1 VNB.t4 1196.12
R57 VNB.t2 VNB.t1 1196.12
R58 VNB.t0 VNB.t2 1196.12
R59 VNB.t7 VNB.t0 1196.12
R60 VNB VNB.t7 911.327
R61 VPWR.n5 VPWR.t5 350.045
R62 VPWR.n15 VPWR.n1 320.976
R63 VPWR.n9 VPWR.n8 320.976
R64 VPWR.n6 VPWR.n4 320.976
R65 VPWR.n17 VPWR.t2 249.901
R66 VPWR.n10 VPWR.n7 34.6358
R67 VPWR.n14 VPWR.n2 34.6358
R68 VPWR.n16 VPWR.n15 30.8711
R69 VPWR.n1 VPWR.t7 26.5955
R70 VPWR.n1 VPWR.t1 26.5955
R71 VPWR.n8 VPWR.t6 26.5955
R72 VPWR.n8 VPWR.t0 26.5955
R73 VPWR.n4 VPWR.t4 26.5955
R74 VPWR.n4 VPWR.t3 26.5955
R75 VPWR.n17 VPWR.n16 25.977
R76 VPWR.n9 VPWR.n2 24.8476
R77 VPWR.n6 VPWR.n5 22.4624
R78 VPWR.n7 VPWR.n6 18.824
R79 VPWR.n10 VPWR.n9 9.78874
R80 VPWR.n7 VPWR.n3 9.3005
R81 VPWR.n11 VPWR.n10 9.3005
R82 VPWR.n12 VPWR.n2 9.3005
R83 VPWR.n14 VPWR.n13 9.3005
R84 VPWR.n16 VPWR.n0 9.3005
R85 VPWR.n18 VPWR.n17 9.3005
R86 VPWR.n15 VPWR.n14 3.76521
R87 VPWR.n5 VPWR.n3 1.07033
R88 VPWR.n11 VPWR.n3 0.120292
R89 VPWR.n12 VPWR.n11 0.120292
R90 VPWR.n13 VPWR.n12 0.120292
R91 VPWR.n13 VPWR.n0 0.120292
R92 VPWR.n18 VPWR.n0 0.120292
R93 VPWR VPWR.n18 0.0213333
R94 VPB.t4 VPB.t5 248.599
R95 VPB.t3 VPB.t4 248.599
R96 VPB.t6 VPB.t3 248.599
R97 VPB.t0 VPB.t6 248.599
R98 VPB.t7 VPB.t0 248.599
R99 VPB.t1 VPB.t7 248.599
R100 VPB.t2 VPB.t1 248.599
R101 VPB VPB.t2 189.409
R102 B.n2 B.t0 212.081
R103 B.n1 B.t1 212.081
R104 B.n7 B.t2 212.081
R105 B.n9 B.t6 212.081
R106 B.n10 B.n9 180.482
R107 B.n4 B.n3 152
R108 B.n6 B.n5 152
R109 B.n8 B.n0 152
R110 B.n2 B.t4 139.78
R111 B.n1 B.t5 139.78
R112 B.n7 B.t3 139.78
R113 B.n9 B.t7 139.78
R114 B.n3 B.n2 30.6732
R115 B.n3 B.n1 30.6732
R116 B.n6 B.n1 30.6732
R117 B.n7 B.n6 30.6732
R118 B.n8 B.n7 30.6732
R119 B.n9 B.n8 30.6732
R120 B.n5 B.n4 21.5045
R121 B B.n0 19.9685
R122 B B.n10 17.1525
R123 B.n10 B 6.4005
R124 B B.n0 3.5845
R125 B.n5 B 1.5365
R126 B.n4 B 0.5125
R127 VGND.n2 VGND.n1 217.232
R128 VGND.n2 VGND.n0 213.804
R129 VGND.n1 VGND.t2 24.9236
R130 VGND.n1 VGND.t1 24.9236
R131 VGND.n0 VGND.t3 24.9236
R132 VGND.n0 VGND.t0 24.9236
R133 VGND VGND.n2 0.53334
C0 Y VGND 0.024648f
C1 VPB A 0.127754f
C2 B A 0.050963f
C3 VPB VPWR 0.105197f
C4 B VPWR 0.094712f
C5 A VPWR 0.07227f
C6 Y VPB 0.019848f
C7 VGND VPB 0.009063f
C8 Y B 0.200103f
C9 VGND B 0.059788f
C10 Y A 0.263237f
C11 Y VPWR 0.730648f
C12 VGND A 0.039395f
C13 VGND VPWR 0.084054f
C14 VPB B 0.13391f
C15 VGND VNB 0.481506f
C16 Y VNB 0.030628f
C17 VPWR VNB 0.468596f
C18 A VNB 0.396805f
C19 B VNB 0.41776f
C20 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_8 VNB VPB VGND VPWR A Y B
X0 a_27_47.t9 B.t0 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y.t15 A.t0 VPWR.t14 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47.t8 B.t1 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_47.t11 A.t1 Y.t23 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47.t12 A.t2 Y.t22 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t7 B.t2 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t6 B.t3 Y.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t21 A.t3 a_27_47.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t20 A.t4 a_27_47.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t19 A.t5 a_27_47.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t5 B.t4 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR.t13 A.t6 Y.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y.t13 A.t7 VPWR.t12 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR.t4 B.t5 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t11 A.t8 Y.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47.t7 B.t6 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47.t6 B.t7 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_27_47.t0 A.t9 Y.t18 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t11 A.t10 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t3 B.t8 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t3 B.t9 a_27_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t2 B.t10 a_27_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t2 B.t11 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t9 A.t11 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND.t1 B.t12 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 Y.t17 A.t12 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t1 B.t13 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t9 A.t13 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y.t0 B.t14 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 VPWR.t15 A.t14 Y.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND.t0 B.t15 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_27_47.t10 A.t15 Y.t16 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B.n3 B.t8 221.72
R1 B.n5 B.t11 221.72
R2 B.n2 B.t13 221.72
R3 B.n10 B.t2 221.72
R4 B.n12 B.t3 221.72
R5 B.n18 B.t4 221.72
R6 B.n16 B.t5 221.72
R7 B.n13 B.t14 221.72
R8 B.n4 B 168.874
R9 B.n7 B.n6 152
R10 B.n9 B.n8 152
R11 B.n11 B.n0 152
R12 B.n20 B.n19 152
R13 B.n17 B.n1 152
R14 B.n15 B.n14 152
R15 B.n3 B.t1 149.421
R16 B.n5 B.t12 149.421
R17 B.n2 B.t0 149.421
R18 B.n10 B.t10 149.421
R19 B.n12 B.t7 149.421
R20 B.n18 B.t9 149.421
R21 B.n16 B.t6 149.421
R22 B.n13 B.t15 149.421
R23 B.n16 B.n15 38.382
R24 B.n4 B.n3 37.4894
R25 B.n5 B.n4 37.4894
R26 B.n6 B.n5 37.4894
R27 B.n6 B.n2 37.4894
R28 B.n9 B.n2 37.4894
R29 B.n10 B.n9 37.4894
R30 B.n11 B.n10 37.4894
R31 B.n12 B.n11 37.4894
R32 B.n19 B.n12 37.4894
R33 B.n19 B.n18 37.4894
R34 B.n18 B.n17 37.4894
R35 B.n17 B.n16 37.4894
R36 B.n15 B.n13 36.5968
R37 B.n20 B.n1 24.4369
R38 B B.n0 23.855
R39 B.n14 B 22.9823
R40 B.n8 B 21.5278
R41 B B.n7 19.2005
R42 B.n7 B 7.56414
R43 B.n8 B 5.23686
R44 B.n14 B 3.78232
R45 B B.n0 2.90959
R46 B B.n1 1.74595
R47 B B.n20 0.582318
R48 VGND.n7 VGND.n6 220.403
R49 VGND.n8 VGND.n5 208.719
R50 VGND.n3 VGND.n2 208.719
R51 VGND.n15 VGND.n1 208.719
R52 VGND.n16 VGND.n15 43.1829
R53 VGND.n10 VGND.n9 34.6358
R54 VGND.n14 VGND.n13 34.6358
R55 VGND.n13 VGND.n3 27.8593
R56 VGND.n6 VGND.t6 24.9236
R57 VGND.n6 VGND.t1 24.9236
R58 VGND.n5 VGND.t7 24.9236
R59 VGND.n5 VGND.t2 24.9236
R60 VGND.n2 VGND.t4 24.9236
R61 VGND.n2 VGND.t3 24.9236
R62 VGND.n1 VGND.t5 24.9236
R63 VGND.n1 VGND.t0 24.9236
R64 VGND.n9 VGND.n8 21.8358
R65 VGND.n8 VGND.n7 19.5455
R66 VGND.n9 VGND.n4 9.3005
R67 VGND.n11 VGND.n10 9.3005
R68 VGND.n13 VGND.n12 9.3005
R69 VGND.n14 VGND.n0 9.3005
R70 VGND.n10 VGND.n3 6.77697
R71 VGND.n7 VGND.n4 1.00279
R72 VGND.n15 VGND.n14 0.753441
R73 VGND.n11 VGND.n4 0.120292
R74 VGND.n12 VGND.n11 0.120292
R75 VGND.n12 VGND.n0 0.120292
R76 VGND.n16 VGND.n0 0.120292
R77 VGND VGND.n16 0.0213333
R78 a_27_47.n5 a_27_47.n4 185
R79 a_27_47.n7 a_27_47.n6 185
R80 a_27_47.n9 a_27_47.n8 185
R81 a_27_47.n5 a_27_47.t0 181.739
R82 a_27_47.n1 a_27_47.t2 176.43
R83 a_27_47.n1 a_27_47.n0 98.788
R84 a_27_47.n3 a_27_47.n2 98.788
R85 a_27_47.n13 a_27_47.n12 98.788
R86 a_27_47.n11 a_27_47.n10 88.3446
R87 a_27_47.n11 a_27_47.n9 51.8673
R88 a_27_47.n12 a_27_47.n11 50.8099
R89 a_27_47.n7 a_27_47.n5 46.7483
R90 a_27_47.n9 a_27_47.n7 46.7483
R91 a_27_47.n3 a_27_47.n1 38.4005
R92 a_27_47.n12 a_27_47.n3 38.4005
R93 a_27_47.n10 a_27_47.t1 24.9236
R94 a_27_47.n10 a_27_47.t8 24.9236
R95 a_27_47.n8 a_27_47.t15 24.9236
R96 a_27_47.n8 a_27_47.t12 24.9236
R97 a_27_47.n6 a_27_47.t13 24.9236
R98 a_27_47.n6 a_27_47.t10 24.9236
R99 a_27_47.n4 a_27_47.t14 24.9236
R100 a_27_47.n4 a_27_47.t11 24.9236
R101 a_27_47.n0 a_27_47.t5 24.9236
R102 a_27_47.n0 a_27_47.t7 24.9236
R103 a_27_47.n2 a_27_47.t4 24.9236
R104 a_27_47.n2 a_27_47.t6 24.9236
R105 a_27_47.n13 a_27_47.t3 24.9236
R106 a_27_47.t9 a_27_47.n13 24.9236
R107 VNB.t14 VNB.t0 1196.12
R108 VNB.t11 VNB.t14 1196.12
R109 VNB.t13 VNB.t11 1196.12
R110 VNB.t10 VNB.t13 1196.12
R111 VNB.t15 VNB.t10 1196.12
R112 VNB.t12 VNB.t15 1196.12
R113 VNB.t1 VNB.t12 1196.12
R114 VNB.t8 VNB.t1 1196.12
R115 VNB.t3 VNB.t8 1196.12
R116 VNB.t9 VNB.t3 1196.12
R117 VNB.t4 VNB.t9 1196.12
R118 VNB.t6 VNB.t4 1196.12
R119 VNB.t5 VNB.t6 1196.12
R120 VNB.t7 VNB.t5 1196.12
R121 VNB.t2 VNB.t7 1196.12
R122 VNB VNB.t2 911.327
R123 A.n1 A.t11 221.72
R124 A.n2 A.t13 221.72
R125 A.n4 A.t14 221.72
R126 A.n6 A.t0 221.72
R127 A.n14 A.t6 221.72
R128 A.n7 A.t7 221.72
R129 A.n9 A.t8 221.72
R130 A.n8 A.t10 221.72
R131 A.n3 A 152.641
R132 A.n5 A.n0 152
R133 A.n16 A.n15 152
R134 A.n13 A.n12 152
R135 A.n11 A.n10 152
R136 A.n1 A.t9 149.421
R137 A.n2 A.t4 149.421
R138 A.n4 A.t1 149.421
R139 A.n6 A.t3 149.421
R140 A.n14 A.t15 149.421
R141 A.n7 A.t5 149.421
R142 A.n9 A.t2 149.421
R143 A.n8 A.t12 149.421
R144 A.n2 A.n1 74.9783
R145 A.n9 A.n8 74.9783
R146 A.n3 A.n2 37.4894
R147 A.n4 A.n3 37.4894
R148 A.n5 A.n4 37.4894
R149 A.n6 A.n5 37.4894
R150 A.n15 A.n6 37.4894
R151 A.n15 A.n14 37.4894
R152 A.n14 A.n13 37.4894
R153 A.n13 A.n7 37.4894
R154 A.n10 A.n7 37.4894
R155 A.n10 A.n9 37.4894
R156 A A.n0 26.2405
R157 A A.n16 23.6805
R158 A.n12 A 21.1205
R159 A A.n11 18.5605
R160 A.n11 A 10.8805
R161 A.n12 A 8.3205
R162 A.n16 A 5.7605
R163 A A.n0 3.2005
R164 VPWR.n37 VPWR.n1 320.976
R165 VPWR.n31 VPWR.n30 320.976
R166 VPWR.n28 VPWR.n4 320.976
R167 VPWR.n22 VPWR.n21 320.976
R168 VPWR.n19 VPWR.n7 320.976
R169 VPWR.n13 VPWR.n12 320.976
R170 VPWR.n11 VPWR.n10 320.976
R171 VPWR.n9 VPWR.t9 268.26
R172 VPWR.n39 VPWR.t0 249.901
R173 VPWR.n18 VPWR.n8 34.6358
R174 VPWR.n23 VPWR.n20 34.6358
R175 VPWR.n27 VPWR.n5 34.6358
R176 VPWR.n32 VPWR.n29 34.6358
R177 VPWR.n36 VPWR.n2 34.6358
R178 VPWR.n14 VPWR.n13 33.8829
R179 VPWR.n38 VPWR.n37 30.8711
R180 VPWR.n14 VPWR.n11 29.3652
R181 VPWR.n19 VPWR.n18 27.8593
R182 VPWR.n1 VPWR.t5 26.5955
R183 VPWR.n1 VPWR.t4 26.5955
R184 VPWR.n30 VPWR.t7 26.5955
R185 VPWR.n30 VPWR.t6 26.5955
R186 VPWR.n4 VPWR.t2 26.5955
R187 VPWR.n4 VPWR.t1 26.5955
R188 VPWR.n21 VPWR.t10 26.5955
R189 VPWR.n21 VPWR.t3 26.5955
R190 VPWR.n7 VPWR.t12 26.5955
R191 VPWR.n7 VPWR.t11 26.5955
R192 VPWR.n12 VPWR.t14 26.5955
R193 VPWR.n12 VPWR.t13 26.5955
R194 VPWR.n10 VPWR.t8 26.5955
R195 VPWR.n10 VPWR.t15 26.5955
R196 VPWR.n39 VPWR.n38 25.977
R197 VPWR.n31 VPWR.n2 24.8476
R198 VPWR.n23 VPWR.n22 21.8358
R199 VPWR.n29 VPWR.n28 18.824
R200 VPWR.n28 VPWR.n27 15.8123
R201 VPWR.n22 VPWR.n5 12.8005
R202 VPWR.n11 VPWR.n9 12.4252
R203 VPWR.n32 VPWR.n31 9.78874
R204 VPWR.n15 VPWR.n14 9.3005
R205 VPWR.n16 VPWR.n8 9.3005
R206 VPWR.n18 VPWR.n17 9.3005
R207 VPWR.n20 VPWR.n6 9.3005
R208 VPWR.n24 VPWR.n23 9.3005
R209 VPWR.n25 VPWR.n5 9.3005
R210 VPWR.n27 VPWR.n26 9.3005
R211 VPWR.n29 VPWR.n3 9.3005
R212 VPWR.n33 VPWR.n32 9.3005
R213 VPWR.n34 VPWR.n2 9.3005
R214 VPWR.n36 VPWR.n35 9.3005
R215 VPWR.n38 VPWR.n0 9.3005
R216 VPWR.n40 VPWR.n39 9.3005
R217 VPWR.n20 VPWR.n19 6.77697
R218 VPWR.n37 VPWR.n36 3.76521
R219 VPWR.n13 VPWR.n8 0.753441
R220 VPWR.n15 VPWR.n9 0.572285
R221 VPWR.n16 VPWR.n15 0.120292
R222 VPWR.n17 VPWR.n16 0.120292
R223 VPWR.n17 VPWR.n6 0.120292
R224 VPWR.n24 VPWR.n6 0.120292
R225 VPWR.n25 VPWR.n24 0.120292
R226 VPWR.n26 VPWR.n25 0.120292
R227 VPWR.n26 VPWR.n3 0.120292
R228 VPWR.n33 VPWR.n3 0.120292
R229 VPWR.n34 VPWR.n33 0.120292
R230 VPWR.n35 VPWR.n34 0.120292
R231 VPWR.n35 VPWR.n0 0.120292
R232 VPWR.n40 VPWR.n0 0.120292
R233 VPWR VPWR.n40 0.0213333
R234 Y.n2 Y.n0 238.502
R235 Y.n2 Y.n1 205.863
R236 Y.n4 Y.n3 205.863
R237 Y.n6 Y.n5 205.863
R238 Y.n11 Y.n10 205.863
R239 Y.n13 Y.n12 205.863
R240 Y.n15 Y.n14 205.863
R241 Y.n9 Y.n8 202.095
R242 Y.n17 Y.n16 185
R243 Y.n19 Y.n18 185
R244 Y.n21 Y.n20 185
R245 Y.n23 Y.n22 185
R246 Y.n11 Y.n9 43.2005
R247 Y.n19 Y.n17 43.0085
R248 Y.n21 Y.n19 43.0085
R249 Y.n23 Y.n21 43.0085
R250 Y.n17 Y.n15 34.5993
R251 Y.n4 Y.n2 32.6405
R252 Y.n6 Y.n4 32.6405
R253 Y.n13 Y.n11 32.6405
R254 Y.n15 Y.n13 32.6405
R255 Y Y.n6 29.7605
R256 Y.n14 Y.t10 26.5955
R257 Y.n14 Y.t9 26.5955
R258 Y.n8 Y.t12 26.5955
R259 Y.n8 Y.t11 26.5955
R260 Y.n0 Y.t4 26.5955
R261 Y.n0 Y.t0 26.5955
R262 Y.n1 Y.t6 26.5955
R263 Y.n1 Y.t5 26.5955
R264 Y.n3 Y.t1 26.5955
R265 Y.n3 Y.t7 26.5955
R266 Y.n5 Y.t3 26.5955
R267 Y.n5 Y.t2 26.5955
R268 Y.n10 Y.t14 26.5955
R269 Y.n10 Y.t13 26.5955
R270 Y.n12 Y.t8 26.5955
R271 Y.n12 Y.t15 26.5955
R272 Y.n22 Y.t22 24.9236
R273 Y.n22 Y.t17 24.9236
R274 Y.n20 Y.t16 24.9236
R275 Y.n20 Y.t19 24.9236
R276 Y.n18 Y.t23 24.9236
R277 Y.n18 Y.t21 24.9236
R278 Y.n16 Y.t18 24.9236
R279 Y.n16 Y.t20 24.9236
R280 Y Y.n23 11.9861
R281 Y.n9 Y.n7 10.2405
R282 Y.n7 Y 3.2005
R283 Y Y.n7 0.533833
R284 VPB.t9 VPB.t10 248.599
R285 VPB.t8 VPB.t9 248.599
R286 VPB.t15 VPB.t8 248.599
R287 VPB.t14 VPB.t15 248.599
R288 VPB.t13 VPB.t14 248.599
R289 VPB.t12 VPB.t13 248.599
R290 VPB.t11 VPB.t12 248.599
R291 VPB.t3 VPB.t11 248.599
R292 VPB.t2 VPB.t3 248.599
R293 VPB.t1 VPB.t2 248.599
R294 VPB.t7 VPB.t1 248.599
R295 VPB.t6 VPB.t7 248.599
R296 VPB.t5 VPB.t6 248.599
R297 VPB.t4 VPB.t5 248.599
R298 VPB.t0 VPB.t4 248.599
R299 VPB VPB.t0 189.409
C0 VPB B 0.247918f
C1 VPB A 0.247231f
C2 B A 0.050963f
C3 VPB VPWR 0.156716f
C4 VPB Y 0.036586f
C5 B VPWR 0.117991f
C6 VPB VGND 0.010109f
C7 B Y 0.413143f
C8 A VPWR 0.128592f
C9 A Y 0.643618f
C10 B VGND 0.107679f
C11 A VGND 0.064532f
C12 VPWR Y 1.48567f
C13 VPWR VGND 0.14858f
C14 Y VGND 0.055934f
C15 VGND VNB 0.796973f
C16 Y VNB 0.044568f
C17 VPWR VNB 0.753023f
C18 A VNB 0.746105f
C19 B VNB 0.757847f
C20 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_1 VPB VNB VGND VPWR A_N B Y
X0 VGND.t0 A_N.t0 a_27_93.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y.t1 a_27_93.t2 a_206_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47.t1 B.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR.t0 a_27_93.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t2 B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR.t2 A_N.t1 a_27_93.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A_N A_N.n0 158.667
R1 A_N.n0 A_N.t1 137.177
R2 A_N.n0 A_N.t0 121.109
R3 a_27_93.t0 a_27_93.n1 744.056
R4 a_27_93.n1 a_27_93.t1 319.224
R5 a_27_93.n0 a_27_93.t3 236.18
R6 a_27_93.n0 a_27_93.t2 163.881
R7 a_27_93.n1 a_27_93.n0 152
R8 VGND VGND.n0 208.192
R9 VGND.n0 VGND.t0 58.5719
R10 VGND.n0 VGND.t1 24.0005
R11 VNB.t1 VNB.t2 1381.23
R12 VNB.t2 VNB.t0 1196.12
R13 VNB VNB.t1 911.327
R14 a_206_47.t0 a_206_47.t1 49.8467
R15 Y Y.n0 338.923
R16 Y Y.t1 278.432
R17 Y.n0 Y.t0 26.5955
R18 Y.n0 Y.t2 26.5955
R19 B.n0 B.t1 236.18
R20 B B.n0 168.534
R21 B.n0 B.t0 163.881
R22 VPWR.n1 VPWR.t0 877.471
R23 VPWR.n1 VPWR.n0 323.575
R24 VPWR.n0 VPWR.t2 96.1553
R25 VPWR.n0 VPWR.t1 25.6105
R26 VPWR VPWR.n1 0.450714
R27 VPB.t2 VPB.t1 287.072
R28 VPB.t1 VPB.t0 248.599
R29 VPB VPB.t2 189.409
C0 VPB VGND 0.009422f
C1 B Y 0.009537f
C2 VPWR A_N 0.008355f
C3 VPWR Y 0.183529f
C4 B VGND 0.018122f
C5 VPWR VGND 0.046752f
C6 A_N Y 0.001943f
C7 A_N VGND 0.011824f
C8 Y VGND 0.109422f
C9 VPB B 0.03218f
C10 VPB VPWR 0.07884f
C11 B VPWR 0.017592f
C12 VPB A_N 0.044474f
C13 B A_N 0.060249f
C14 VPB Y 0.026386f
C15 VGND VNB 0.312047f
C16 Y VNB 0.094349f
C17 A_N VNB 0.145084f
C18 VPWR VNB 0.278655f
C19 B VNB 0.101877f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2i_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2i_4 VNB VPB VGND VPWR Y A0 A1 S
X0 Y.t5 A1.t0 a_445_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y.t4 A1.t1 a_445_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t8 a_1191_21.t2 a_445_297.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.1625 ps=1.325 w=1 l=0.15
X3 a_445_297.t3 A1.t2 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t14 A0.t0 a_109_297.t3 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_445_297.t4 a_1191_21.t3 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6 a_1191_21.t1 S.t0 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X7 VPWR.t6 a_1191_21.t4 a_445_297.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_445_47.t4 S.t1 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_297.t2 A0.t1 Y.t15 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_445_297.t6 a_1191_21.t5 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_445_47.t5 S.t2 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_109_47.t7 a_1191_21.t6 VGND.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t11 A0.t2 a_109_297.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t12 A0.t3 a_109_47.t3 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y.t13 A0.t4 a_109_47.t2 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_1191_21.t0 S.t3 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X17 VGND.t5 S.t4 a_445_47.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t6 A1.t3 a_445_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t4 S.t5 a_445_47.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND.t2 a_1191_21.t7 a_109_47.t6 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_109_47.t1 A0.t5 Y.t8 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_445_47.t1 A1.t4 Y.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_445_297.t1 A1.t5 Y.t7 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t4 S.t6 a_109_297.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_445_47.t0 A1.t6 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VGND.t1 a_1191_21.t8 a_109_47.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.105625 ps=0.975 w=0.65 l=0.15
X27 Y.t0 A1.t7 a_445_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_109_297.t4 S.t7 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR.t1 S.t8 a_109_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_109_47.t4 a_1191_21.t9 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_109_297.t0 A0.t6 Y.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_109_297.t6 S.t9 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_109_47.t0 A0.t7 Y.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n1 A1.t3 212.081
R1 A1.n9 A1.t5 212.081
R2 A1.n2 A1.t7 212.081
R3 A1.n3 A1.t2 212.081
R4 A1.n11 A1.n10 152
R5 A1.n8 A1.n0 152
R6 A1.n7 A1.n6 152
R7 A1.n5 A1.n4 152
R8 A1.n1 A1.t1 139.78
R9 A1.n9 A1.t6 139.78
R10 A1.n2 A1.t0 139.78
R11 A1.n3 A1.t4 139.78
R12 A1.n8 A1.n7 49.6611
R13 A1.n4 A1.n2 48.2005
R14 A1.n10 A1.n9 39.4369
R15 A1.n10 A1.n1 21.9096
R16 A1.n11 A1.n0 13.1884
R17 A1.n4 A1.n3 13.146
R18 A1.n6 A1 12.8005
R19 A1.n9 A1.n8 10.2247
R20 A1.n5 A1 9.69747
R21 A1 A1.n5 8.14595
R22 A1.n6 A1 5.04292
R23 A1 A1.n11 4.26717
R24 A1.n7 A1.n2 1.46111
R25 A1 A1.n0 0.388379
R26 a_445_47.n2 a_445_47.n1 265.942
R27 a_445_47.n4 a_445_47.n3 248.248
R28 a_445_47.n2 a_445_47.n0 202.695
R29 a_445_47.n5 a_445_47.n4 185
R30 a_445_47.n4 a_445_47.n2 102.4
R31 a_445_47.n3 a_445_47.t3 24.9236
R32 a_445_47.n3 a_445_47.t1 24.9236
R33 a_445_47.n0 a_445_47.t7 24.9236
R34 a_445_47.n0 a_445_47.t5 24.9236
R35 a_445_47.n1 a_445_47.t6 24.9236
R36 a_445_47.n1 a_445_47.t4 24.9236
R37 a_445_47.n5 a_445_47.t2 24.9236
R38 a_445_47.t0 a_445_47.n5 24.9236
R39 Y.n1 Y.t6 917.229
R40 Y.n6 Y.t9 853.981
R41 Y.n1 Y.n0 585
R42 Y.n3 Y.n2 585
R43 Y.n5 Y.n4 585
R44 Y.n8 Y.t4 322.094
R45 Y.n13 Y.t10 258.846
R46 Y.n8 Y.n7 185
R47 Y.n10 Y.n9 185
R48 Y.n12 Y.n11 185
R49 Y.n3 Y.n1 63.2476
R50 Y.n5 Y.n3 63.2476
R51 Y.n10 Y.n8 63.2476
R52 Y.n12 Y.n10 63.2476
R53 Y.n6 Y.n5 58.7299
R54 Y.n13 Y.n12 58.7299
R55 Y.n4 Y.t15 26.5955
R56 Y.n4 Y.t11 26.5955
R57 Y.n2 Y.t1 26.5955
R58 Y.n2 Y.t14 26.5955
R59 Y.n0 Y.t7 26.5955
R60 Y.n0 Y.t0 26.5955
R61 Y.n11 Y.t8 24.9236
R62 Y.n11 Y.t12 24.9236
R63 Y.n9 Y.t3 24.9236
R64 Y.n9 Y.t13 24.9236
R65 Y.n7 Y.t2 24.9236
R66 Y.n7 Y.t5 24.9236
R67 Y Y.n13 20.7649
R68 Y Y.n6 12.2316
R69 VNB.t6 VNB.t9 2677.02
R70 VNB.t3 VNB.t2 1352.75
R71 VNB.t2 VNB.t12 1324.27
R72 VNB.t1 VNB.t3 1196.12
R73 VNB.t0 VNB.t1 1196.12
R74 VNB.t10 VNB.t0 1196.12
R75 VNB.t8 VNB.t10 1196.12
R76 VNB.t11 VNB.t8 1196.12
R77 VNB.t9 VNB.t11 1196.12
R78 VNB.t4 VNB.t6 1196.12
R79 VNB.t7 VNB.t4 1196.12
R80 VNB.t5 VNB.t7 1196.12
R81 VNB.t16 VNB.t5 1196.12
R82 VNB.t13 VNB.t16 1196.12
R83 VNB.t15 VNB.t13 1196.12
R84 VNB.t14 VNB.t15 1196.12
R85 VNB VNB.t14 911.327
R86 a_1191_21.t0 a_1191_21.n5 406.478
R87 a_1191_21.n5 a_1191_21.t1 265.37
R88 a_1191_21.n0 a_1191_21.t2 212.081
R89 a_1191_21.n3 a_1191_21.t3 212.081
R90 a_1191_21.n2 a_1191_21.t4 212.081
R91 a_1191_21.n1 a_1191_21.t5 212.081
R92 a_1191_21.n5 a_1191_21.n4 140.978
R93 a_1191_21.n0 a_1191_21.t8 139.78
R94 a_1191_21.n3 a_1191_21.t9 139.78
R95 a_1191_21.n2 a_1191_21.t7 139.78
R96 a_1191_21.n1 a_1191_21.t6 139.78
R97 a_1191_21.n3 a_1191_21.n2 61.346
R98 a_1191_21.n2 a_1191_21.n1 61.346
R99 a_1191_21.n4 a_1191_21.n0 33.977
R100 a_1191_21.n4 a_1191_21.n3 28.1978
R101 a_445_297.n5 a_445_297.n4 648.247
R102 a_445_297.n4 a_445_297.n3 585
R103 a_445_297.n2 a_445_297.n1 359.74
R104 a_445_297.n2 a_445_297.n0 296.493
R105 a_445_297.n4 a_445_297.n2 228.894
R106 a_445_297.n1 a_445_297.t5 37.4305
R107 a_445_297.n3 a_445_297.t2 26.5955
R108 a_445_297.n3 a_445_297.t1 26.5955
R109 a_445_297.n0 a_445_297.t7 26.5955
R110 a_445_297.n0 a_445_297.t6 26.5955
R111 a_445_297.n1 a_445_297.t4 26.5955
R112 a_445_297.n5 a_445_297.t0 26.5955
R113 a_445_297.t3 a_445_297.n5 26.5955
R114 VPWR.n0 VPWR.t2 868.721
R115 VPWR.n6 VPWR.n5 605.277
R116 VPWR.n14 VPWR.n2 599.74
R117 VPWR.n4 VPWR.n3 599.74
R118 VPWR.n8 VPWR.n7 599.74
R119 VPWR.n5 VPWR.t8 35.4605
R120 VPWR.n15 VPWR.n14 33.5064
R121 VPWR.n13 VPWR.n4 27.4829
R122 VPWR.n2 VPWR.t0 26.5955
R123 VPWR.n2 VPWR.t1 26.5955
R124 VPWR.n3 VPWR.t5 26.5955
R125 VPWR.n3 VPWR.t4 26.5955
R126 VPWR.n7 VPWR.t7 26.5955
R127 VPWR.n7 VPWR.t6 26.5955
R128 VPWR.n5 VPWR.t3 26.5955
R129 VPWR.n9 VPWR.n8 21.4593
R130 VPWR.n9 VPWR.n4 16.9417
R131 VPWR.n17 VPWR.n0 12.4952
R132 VPWR.n14 VPWR.n13 10.9181
R133 VPWR.n10 VPWR.n9 9.3005
R134 VPWR.n11 VPWR.n4 9.3005
R135 VPWR.n13 VPWR.n12 9.3005
R136 VPWR.n14 VPWR.n1 9.3005
R137 VPWR.n16 VPWR.n15 9.3005
R138 VPWR.n8 VPWR.n6 6.68038
R139 VPWR.n15 VPWR.n0 4.89462
R140 VPWR VPWR.n17 0.957626
R141 VPWR.n10 VPWR.n6 0.551658
R142 VPWR.n17 VPWR.n16 0.147187
R143 VPWR.n11 VPWR.n10 0.120292
R144 VPWR.n12 VPWR.n11 0.120292
R145 VPWR.n12 VPWR.n1 0.120292
R146 VPWR.n16 VPWR.n1 0.120292
R147 VPB.t2 VPB.t6 556.386
R148 VPB.t11 VPB.t12 281.154
R149 VPB.t12 VPB.t7 275.235
R150 VPB.t10 VPB.t11 248.599
R151 VPB.t9 VPB.t10 248.599
R152 VPB.t8 VPB.t9 248.599
R153 VPB.t4 VPB.t8 248.599
R154 VPB.t5 VPB.t4 248.599
R155 VPB.t6 VPB.t5 248.599
R156 VPB.t1 VPB.t2 248.599
R157 VPB.t0 VPB.t1 248.599
R158 VPB.t3 VPB.t0 248.599
R159 VPB.t15 VPB.t3 248.599
R160 VPB.t16 VPB.t15 248.599
R161 VPB.t14 VPB.t16 248.599
R162 VPB.t13 VPB.t14 248.599
R163 VPB VPB.t13 189.409
R164 A0.n1 A0.t0 212.081
R165 A0.n2 A0.t1 212.081
R166 A0.n4 A0.t2 212.081
R167 A0.n5 A0.t6 212.081
R168 A0.n3 A0.n0 152
R169 A0.n7 A0.n6 152
R170 A0.n1 A0.t4 139.78
R171 A0.n2 A0.t5 139.78
R172 A0.n4 A0.t3 139.78
R173 A0.n5 A0.t7 139.78
R174 A0.n2 A0.n1 61.346
R175 A0.n3 A0.n2 47.4702
R176 A0.n6 A0.n4 35.7853
R177 A0.n6 A0.n5 25.5611
R178 A0.n4 A0.n3 13.8763
R179 A0.n7 A0.n0 13.1884
R180 A0.n0 A0 11.5798
R181 A0 A0.n7 1.35808
R182 a_109_297.n2 a_109_297.n0 648.247
R183 a_109_297.n4 a_109_297.n3 648.247
R184 a_109_297.n2 a_109_297.n1 585
R185 a_109_297.n5 a_109_297.n4 585
R186 a_109_297.n4 a_109_297.n2 228.894
R187 a_109_297.n3 a_109_297.t1 26.5955
R188 a_109_297.n3 a_109_297.t0 26.5955
R189 a_109_297.n1 a_109_297.t5 26.5955
R190 a_109_297.n1 a_109_297.t6 26.5955
R191 a_109_297.n0 a_109_297.t7 26.5955
R192 a_109_297.n0 a_109_297.t4 26.5955
R193 a_109_297.t3 a_109_297.n5 26.5955
R194 a_109_297.n5 a_109_297.t2 26.5955
R195 S S.n0 335.911
R196 S.n0 S.t3 241.536
R197 S.n1 S.t6 212.081
R198 S.n11 S.t7 212.081
R199 S.n3 S.t8 212.081
R200 S.n5 S.t9 212.081
R201 S.n5 S.n4 179.752
R202 S.n0 S.t0 169.237
R203 S.n13 S.n12 152
R204 S.n10 S.n9 152
R205 S.n8 S.n2 152
R206 S.n7 S.n6 152
R207 S.n1 S.t4 139.78
R208 S.n11 S.t1 139.78
R209 S.n3 S.t5 139.78
R210 S.n5 S.t2 139.78
R211 S.n10 S.n2 49.6611
R212 S.n12 S.n11 48.2005
R213 S.n6 S.n3 39.4369
R214 S.n6 S.n5 21.9096
R215 S.n9 S.n8 20.2424
R216 S.n4 S 18.4563
R217 S.n13 S 17.2656
R218 S S.n7 16.0749
R219 S.n12 S.n1 13.146
R220 S.n7 S 11.3121
R221 S.n3 S.n2 10.2247
R222 S S.n13 10.1214
R223 S.n4 S 8.93073
R224 S.n8 S 4.16794
R225 S.n9 S 2.97724
R226 S.n11 S.n10 1.46111
R227 VGND.n0 VGND.t6 282.817
R228 VGND.n5 VGND.n4 205.304
R229 VGND.n7 VGND.n6 204.457
R230 VGND.n3 VGND.n2 201.738
R231 VGND.n14 VGND.n13 199.739
R232 VGND.n15 VGND.n14 33.5064
R233 VGND.n4 VGND.t1 33.2313
R234 VGND.n12 VGND.n3 27.4829
R235 VGND.n8 VGND.n7 25.224
R236 VGND.n4 VGND.t8 24.9236
R237 VGND.n6 VGND.t0 24.9236
R238 VGND.n6 VGND.t2 24.9236
R239 VGND.n2 VGND.t3 24.9236
R240 VGND.n2 VGND.t5 24.9236
R241 VGND.n13 VGND.t7 24.9236
R242 VGND.n13 VGND.t4 24.9236
R243 VGND.n8 VGND.n3 17.3181
R244 VGND.n17 VGND.n0 12.4952
R245 VGND.n14 VGND.n12 10.9181
R246 VGND.n16 VGND.n15 9.3005
R247 VGND.n14 VGND.n1 9.3005
R248 VGND.n12 VGND.n11 9.3005
R249 VGND.n10 VGND.n3 9.3005
R250 VGND.n9 VGND.n8 9.3005
R251 VGND.n7 VGND.n5 6.82214
R252 VGND.n15 VGND.n0 4.89462
R253 VGND VGND.n17 0.957626
R254 VGND.n9 VGND.n5 0.52835
R255 VGND.n17 VGND.n16 0.147187
R256 VGND.n10 VGND.n9 0.120292
R257 VGND.n11 VGND.n10 0.120292
R258 VGND.n11 VGND.n1 0.120292
R259 VGND.n16 VGND.n1 0.120292
R260 a_109_47.n5 a_109_47.n4 243.367
R261 a_109_47.n2 a_109_47.n1 242.964
R262 a_109_47.n2 a_109_47.n0 206.577
R263 a_109_47.n4 a_109_47.n3 185
R264 a_109_47.n1 a_109_47.t5 35.0774
R265 a_109_47.n4 a_109_47.n2 26.967
R266 a_109_47.n3 a_109_47.t2 24.9236
R267 a_109_47.n3 a_109_47.t1 24.9236
R268 a_109_47.n0 a_109_47.t6 24.9236
R269 a_109_47.n0 a_109_47.t7 24.9236
R270 a_109_47.n1 a_109_47.t4 24.9236
R271 a_109_47.t3 a_109_47.n5 24.9236
R272 a_109_47.n5 a_109_47.t0 24.9236
C0 A0 VPWR 0.034775f
C1 VPB VGND 0.005597f
C2 A1 Y 0.066272f
C3 S Y 0.001828f
C4 A1 VPWR 0.028431f
C5 A0 VGND 0.03469f
C6 A1 VGND 0.020527f
C7 S VPWR 0.119081f
C8 Y VPWR 0.37433f
C9 S VGND 0.091216f
C10 Y VGND 0.353044f
C11 VPWR VGND 0.06614f
C12 VPB A0 0.118755f
C13 VPB A1 0.12186f
C14 VPB S 0.180058f
C15 A0 A1 0.068801f
C16 A0 S 1.23e-19
C17 VPB Y 0.01933f
C18 VPB VPWR 0.152099f
C19 A1 S 0.037819f
C20 A0 Y 0.116232f
C21 VGND VNB 0.882559f
C22 VPWR VNB 0.743574f
C23 Y VNB 0.1105f
C24 S VNB 0.515601f
C25 A1 VNB 0.363133f
C26 A0 VNB 0.37923f
C27 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux4_1 VNB VPB VGND VPWR A1 A0 S0 A3 A2 S1 X
X0 a_277_47.t1 a_247_21.t2 a_27_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND.t6 S0.t0 a_247_21.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_834_97.t0 a_247_21.t3 a_750_97.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND.t1 A3.t0 a_668_97.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X4 a_1290_413.t0 S1.t0 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_834_97.t1 A2.t0 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97.t4 S0.t1 a_757_363.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7 a_27_47.t1 S0.t2 a_277_47.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X8 X.t1 a_1478_413.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR.t3 A1.t0 a_27_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR.t6 S0.t3 a_247_21.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X11 X.t0 a_1478_413.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47.t1 A0.t0 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1478_413.t1 S1.t1 a_277_47.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_1290_413.t1 S1.t2 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_277_47.t0 a_247_21.t4 a_193_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_750_97.t3 S0.t4 a_668_97.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 a_923_363.t0 a_247_21.t5 a_750_97.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_757_363.t0 A2.t1 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR.t2 A3.t1 a_923_363.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X20 a_277_47.t5 a_1290_413.t2 a_1478_413.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X21 a_193_413.t0 A0.t1 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_193_413.t1 S0.t5 a_277_47.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 VGND.t0 A1.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_1478_413.t0 S1.t3 a_750_97.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_247_21.n0 a_247_21.t1 694.98
R1 a_247_21.n1 a_247_21.t4 404.88
R2 a_247_21.n2 a_247_21.t5 296.717
R3 a_247_21.n0 a_247_21.n1 262.856
R4 a_247_21.t0 a_247_21.n0 244.727
R5 a_247_21.n1 a_247_21.t2 221.72
R6 a_247_21.n0 a_247_21.n2 182.435
R7 a_247_21.n2 a_247_21.t3 137.428
R8 a_27_413.t0 a_27_413.t1 1424.27
R9 a_277_47.n1 a_277_47.t4 762.566
R10 a_277_47.n2 a_277_47.n0 691.061
R11 a_277_47.n1 a_277_47.t5 248.65
R12 a_277_47.n3 a_277_47.n2 196.034
R13 a_277_47.t0 a_277_47.n3 74.1148
R14 a_277_47.n0 a_277_47.t3 63.3219
R15 a_277_47.n0 a_277_47.t1 63.3219
R16 a_277_47.n3 a_277_47.t2 37.1434
R17 a_277_47.n2 a_277_47.n1 14.1278
R18 VPB.t6 VPB.t0 1109.81
R19 VPB.t5 VPB.t6 556.386
R20 VPB.t9 VPB.t5 556.386
R21 VPB.t4 VPB.t11 556.386
R22 VPB.t8 VPB.t2 556.386
R23 VPB.t11 VPB.t3 550.467
R24 VPB.t1 VPB.t10 281.154
R25 VPB.t10 VPB.t9 248.599
R26 VPB.t3 VPB.t1 248.599
R27 VPB.t2 VPB.t4 248.599
R28 VPB.t7 VPB.t8 248.599
R29 VPB VPB.t7 192.369
R30 S0.t0 S0.t2 547.874
R31 S0.n0 S0.t1 377.241
R32 S0.n1 S0.t5 223.327
R33 S0.n0 S0.t3 173.996
R34 S0 S0.n3 163.308
R35 S0.n3 S0.t4 130.27
R36 S0.n2 S0.t0 123.43
R37 S0.n2 S0.n1 41.3757
R38 S0.n3 S0.n2 24.7519
R39 S0.n1 S0.n0 1.78419
R40 VGND.n8 VGND.t4 297.955
R41 VGND.n19 VGND.t6 251.821
R42 VGND.n7 VGND.t2 238.311
R43 VGND.n12 VGND.n5 207.213
R44 VGND.n27 VGND.n26 199.739
R45 VGND.n5 VGND.t5 38.5719
R46 VGND.n5 VGND.t1 38.5719
R47 VGND.n26 VGND.t3 38.5719
R48 VGND.n26 VGND.t0 38.5719
R49 VGND.n11 VGND.n6 34.6358
R50 VGND.n14 VGND.n13 34.6358
R51 VGND.n14 VGND.n3 34.6358
R52 VGND.n18 VGND.n3 34.6358
R53 VGND.n20 VGND.n1 34.6358
R54 VGND.n24 VGND.n1 34.6358
R55 VGND.n25 VGND.n24 34.6358
R56 VGND.n13 VGND.n12 30.4946
R57 VGND.n19 VGND.n18 27.1064
R58 VGND.n27 VGND.n25 22.9652
R59 VGND.n20 VGND.n19 20.3299
R60 VGND.n7 VGND.n6 19.577
R61 VGND.n25 VGND.n0 9.3005
R62 VGND.n24 VGND.n23 9.3005
R63 VGND.n22 VGND.n1 9.3005
R64 VGND.n21 VGND.n20 9.3005
R65 VGND.n19 VGND.n2 9.3005
R66 VGND.n9 VGND.n6 9.3005
R67 VGND.n11 VGND.n10 9.3005
R68 VGND.n13 VGND.n4 9.3005
R69 VGND.n15 VGND.n14 9.3005
R70 VGND.n16 VGND.n3 9.3005
R71 VGND.n18 VGND.n17 9.3005
R72 VGND.n8 VGND.n7 7.20364
R73 VGND.n28 VGND.n27 7.12063
R74 VGND.n12 VGND.n11 4.14168
R75 VGND.n9 VGND.n8 0.153669
R76 VGND.n28 VGND.n0 0.148519
R77 VGND.n10 VGND.n9 0.120292
R78 VGND.n10 VGND.n4 0.120292
R79 VGND.n15 VGND.n4 0.120292
R80 VGND.n16 VGND.n15 0.120292
R81 VGND.n17 VGND.n16 0.120292
R82 VGND.n17 VGND.n2 0.120292
R83 VGND.n21 VGND.n2 0.120292
R84 VGND.n22 VGND.n21 0.120292
R85 VGND.n23 VGND.n22 0.120292
R86 VGND.n23 VGND.n0 0.120292
R87 VGND VGND.n28 0.114842
R88 VNB.t8 VNB.t6 3132.69
R89 VNB.t4 VNB.t9 2677.02
R90 VNB.t7 VNB.t4 2677.02
R91 VNB.t12 VNB.t10 2677.02
R92 VNB.t11 VNB.t12 2677.02
R93 VNB.t2 VNB.t3 2648.54
R94 VNB.t9 VNB.t8 2178.64
R95 VNB.t1 VNB.t11 1381.23
R96 VNB.t3 VNB.t7 1196.12
R97 VNB.t10 VNB.t2 1196.12
R98 VNB.t5 VNB.t1 1196.12
R99 VNB.t0 VNB.t5 1196.12
R100 VNB VNB.t0 925.567
R101 a_750_97.n2 a_750_97.n1 591.595
R102 a_750_97.n1 a_750_97.t2 369.337
R103 a_750_97.n1 a_750_97.n0 270.195
R104 a_750_97.t0 a_750_97.n2 63.3219
R105 a_750_97.n2 a_750_97.t4 63.3219
R106 a_750_97.n0 a_750_97.t1 38.5719
R107 a_750_97.n0 a_750_97.t3 38.5719
R108 a_834_97.n0 a_834_97.t1 518.242
R109 a_834_97.n0 a_834_97.t0 27.6928
R110 A3.n0 A3.t1 310.457
R111 A3.n0 A3.t0 220.484
R112 A3 A3.n0 155.304
R113 a_668_97.n0 a_668_97.t1 522.929
R114 a_668_97.n0 a_668_97.t0 30.0005
R115 S1.n1 S1.t0 322.747
R116 S1.n0 S1.t1 305.267
R117 S1.n1 S1.t2 194.213
R118 S1.n0 S1.t3 179.823
R119 S1 S1.n1 154.429
R120 S1.n1 S1.n0 126.803
R121 VPWR.n9 VPWR.t0 875.153
R122 VPWR.n18 VPWR.t6 665.163
R123 VPWR.n8 VPWR.t1 662.22
R124 VPWR.n26 VPWR.n1 599.74
R125 VPWR.n12 VPWR.n7 599.74
R126 VPWR.n1 VPWR.t4 63.3219
R127 VPWR.n1 VPWR.t3 63.3219
R128 VPWR.n7 VPWR.t5 63.3219
R129 VPWR.n7 VPWR.t2 63.3219
R130 VPWR.n20 VPWR.n19 34.6358
R131 VPWR.n20 VPWR.n2 34.6358
R132 VPWR.n24 VPWR.n2 34.6358
R133 VPWR.n25 VPWR.n24 34.6358
R134 VPWR.n13 VPWR.n5 34.6358
R135 VPWR.n17 VPWR.n5 34.6358
R136 VPWR.n12 VPWR.n11 27.1064
R137 VPWR.n18 VPWR.n17 25.977
R138 VPWR.n26 VPWR.n25 22.9652
R139 VPWR.n19 VPWR.n18 18.4476
R140 VPWR.n13 VPWR.n12 17.3181
R141 VPWR.n11 VPWR.n8 17.3181
R142 VPWR.n11 VPWR.n10 9.3005
R143 VPWR.n12 VPWR.n6 9.3005
R144 VPWR.n14 VPWR.n13 9.3005
R145 VPWR.n15 VPWR.n5 9.3005
R146 VPWR.n17 VPWR.n16 9.3005
R147 VPWR.n18 VPWR.n4 9.3005
R148 VPWR.n19 VPWR.n3 9.3005
R149 VPWR.n21 VPWR.n20 9.3005
R150 VPWR.n22 VPWR.n2 9.3005
R151 VPWR.n24 VPWR.n23 9.3005
R152 VPWR.n25 VPWR.n0 9.3005
R153 VPWR.n9 VPWR.n8 7.24059
R154 VPWR.n27 VPWR.n26 7.12063
R155 VPWR.n10 VPWR.n9 0.153169
R156 VPWR.n27 VPWR.n0 0.148519
R157 VPWR.n10 VPWR.n6 0.120292
R158 VPWR.n14 VPWR.n6 0.120292
R159 VPWR.n15 VPWR.n14 0.120292
R160 VPWR.n16 VPWR.n15 0.120292
R161 VPWR.n16 VPWR.n4 0.120292
R162 VPWR.n4 VPWR.n3 0.120292
R163 VPWR.n21 VPWR.n3 0.120292
R164 VPWR.n22 VPWR.n21 0.120292
R165 VPWR.n23 VPWR.n22 0.120292
R166 VPWR.n23 VPWR.n0 0.120292
R167 VPWR VPWR.n27 0.114842
R168 a_1290_413.t0 a_1290_413.n2 728.242
R169 a_1290_413.n1 a_1290_413.n0 312.229
R170 a_1290_413.n2 a_1290_413.t1 273.274
R171 a_1290_413.n2 a_1290_413.n1 234.885
R172 a_1290_413.n1 a_1290_413.t2 115.68
R173 A2.n0 A2.t1 315.442
R174 A2.n0 A2.t0 225.47
R175 A2 A2.n0 156.335
R176 a_757_363.t0 a_757_363.t1 1486.6
R177 a_27_47.t0 a_27_47.t1 619.567
R178 a_1478_413.n1 a_1478_413.t1 834.532
R179 a_1478_413.n2 a_1478_413.n1 319.776
R180 a_1478_413.n0 a_1478_413.t4 233.576
R181 a_1478_413.n0 a_1478_413.t3 161.275
R182 a_1478_413.n1 a_1478_413.n0 152
R183 a_1478_413.n2 a_1478_413.t2 121.85
R184 a_1478_413.t0 a_1478_413.n2 118.572
R185 X X.t0 849.028
R186 X X.t1 266.601
R187 A1.n0 A1.t0 334.723
R188 A1.n0 A1.t1 206.19
R189 A1.n1 A1.n0 152
R190 A1.n1 A1 10.5744
R191 A1 A1.n1 2.04108
R192 A0.n0 A0.t1 334.723
R193 A0.n0 A0.t0 206.19
R194 A0.n1 A0.n0 152
R195 A0.n1 A0 8.38671
R196 A0 A0.n1 1.61889
R197 a_193_47.t0 a_193_47.t1 77.1434
R198 a_923_363.t0 a_923_363.t1 204.174
R199 a_193_413.t0 a_193_413.t1 1426.37
C0 VPB A1 0.074097f
C1 VGND VPWR 0.058958f
C2 S1 A3 1.18e-19
C3 VPB A0 0.080186f
C4 VGND S0 0.066755f
C5 S1 A2 0.068534f
C6 A1 A0 0.141225f
C7 VPB VPWR 0.226889f
C8 VGND A3 0.011612f
C9 A1 VPWR 0.017122f
C10 VPB S0 0.310736f
C11 VGND A2 0.012202f
C12 VPB A3 0.072523f
C13 A0 VPWR 0.01747f
C14 S1 X 2.3e-19
C15 A0 S0 0.00186f
C16 VPB A2 0.078716f
C17 S1 VGND 0.04087f
C18 VPWR S0 0.068699f
C19 X VGND 0.059393f
C20 S1 VPB 0.215337f
C21 VPWR A3 0.012005f
C22 X VPB 0.011812f
C23 VPWR A2 0.012899f
C24 S0 A3 0.003168f
C25 VGND VPB 0.013874f
C26 S1 VPWR 0.040895f
C27 VGND A1 0.017046f
C28 A3 A2 0.154918f
C29 VGND A0 0.017092f
C30 X VPWR 0.059373f
C31 VGND VNB 1.07507f
C32 X VNB 0.092356f
C33 S1 VNB 0.320621f
C34 A2 VNB 0.11249f
C35 A3 VNB 0.119256f
C36 S0 VNB 0.464858f
C37 VPWR VNB 0.868874f
C38 A0 VNB 0.102565f
C39 A1 VNB 0.175855f
C40 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux4_2 VNB VPB VGND VPWR S0 A2 A3 S1 A1 A0 X
X0 a_600_345.t1 S1.t0 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_788_316.t2 S1.t1 a_288_47.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t7 A3.t0 a_372_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1645 ps=1.33 w=0.64 l=0.15
X3 a_872_316.t1 a_600_345.t2 a_788_316.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X4 VPWR.t4 S0.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VGND.t2 a_788_316.t4 X.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_1060_369.t0 A1.t0 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.13775 pd=1.165 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_193_47.t0 A2.t0 VGND.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_1064_47.t0 A1.t1 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_1281_47.t0 a_27_47.t2 a_872_316.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X10 a_872_316.t2 S1.t2 a_788_316.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1404 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X11 X.t0 a_788_316.t5 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X12 a_788_316.t0 a_600_345.t3 a_288_47.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.1404 ps=1.6 w=0.54 l=0.15
X13 a_372_413.t0 a_27_47.t3 a_288_47.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1645 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VGND.t7 A3.t1 a_397_47.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.06705 ps=0.75 w=0.42 l=0.15
X15 a_600_345.t0 S1.t3 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X16 a_193_369.t0 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X17 VPWR.t2 a_788_316.t6 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.135 ps=1.27 w=1 l=0.15
X18 a_288_47.t2 S0.t1 a_193_369.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X19 VGND.t0 A0.t0 a_1281_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.066 ps=0.745 w=0.42 l=0.15
X20 a_397_47.t0 S0.t2 a_288_47.t0 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X21 X.t2 a_788_316.t7 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X22 a_288_47.t1 a_27_47.t4 a_193_47.t1 VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X23 VGND.t5 S0.t3 a_27_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VPWR.t1 A0.t1 a_1279_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.10535 ps=0.995 w=0.64 l=0.15
R0 S1.t0 S1.t2 769.593
R1 S1.n0 S1.t1 367.928
R2 S1.n1 S1.t0 350.712
R3 S1.n2 S1.n1 152
R4 S1.n0 S1.t3 112.237
R5 S1.n1 S1.n0 34.4291
R6 S1.n2 S1 7.72464
R7 S1 S1.n2 7.28326
R8 VPWR.n18 VPWR.t6 644.364
R9 VPWR.n25 VPWR.n4 612.827
R10 VPWR.n32 VPWR.n1 599.74
R11 VPWR.n11 VPWR.n9 320.976
R12 VPWR.n10 VPWR.t2 273.318
R13 VPWR.n9 VPWR.t1 61.563
R14 VPWR.n1 VPWR.t0 41.5552
R15 VPWR.n1 VPWR.t4 41.5552
R16 VPWR.n4 VPWR.t5 41.5552
R17 VPWR.n4 VPWR.t7 41.5552
R18 VPWR.n26 VPWR.n2 34.6358
R19 VPWR.n30 VPWR.n2 34.6358
R20 VPWR.n31 VPWR.n30 34.6358
R21 VPWR.n19 VPWR.n5 34.6358
R22 VPWR.n23 VPWR.n5 34.6358
R23 VPWR.n24 VPWR.n23 34.6358
R24 VPWR.n13 VPWR.n12 34.6358
R25 VPWR.n13 VPWR.n7 34.6358
R26 VPWR.n17 VPWR.n7 34.6358
R27 VPWR.n12 VPWR.n11 32.377
R28 VPWR.n9 VPWR.t3 30.5947
R29 VPWR.n19 VPWR.n18 28.9887
R30 VPWR.n32 VPWR.n31 22.9652
R31 VPWR.n18 VPWR.n17 14.3064
R32 VPWR.n25 VPWR.n24 12.424
R33 VPWR.n11 VPWR.n10 9.50159
R34 VPWR.n12 VPWR.n8 9.3005
R35 VPWR.n14 VPWR.n13 9.3005
R36 VPWR.n15 VPWR.n7 9.3005
R37 VPWR.n17 VPWR.n16 9.3005
R38 VPWR.n18 VPWR.n6 9.3005
R39 VPWR.n20 VPWR.n19 9.3005
R40 VPWR.n21 VPWR.n5 9.3005
R41 VPWR.n23 VPWR.n22 9.3005
R42 VPWR.n24 VPWR.n3 9.3005
R43 VPWR.n27 VPWR.n26 9.3005
R44 VPWR.n28 VPWR.n2 9.3005
R45 VPWR.n30 VPWR.n29 9.3005
R46 VPWR.n31 VPWR.n0 9.3005
R47 VPWR.n33 VPWR.n32 7.12063
R48 VPWR.n26 VPWR.n25 4.89462
R49 VPWR.n10 VPWR.n8 0.497031
R50 VPWR.n33 VPWR.n0 0.148519
R51 VPWR.n14 VPWR.n8 0.120292
R52 VPWR.n15 VPWR.n14 0.120292
R53 VPWR.n16 VPWR.n15 0.120292
R54 VPWR.n16 VPWR.n6 0.120292
R55 VPWR.n20 VPWR.n6 0.120292
R56 VPWR.n21 VPWR.n20 0.120292
R57 VPWR.n22 VPWR.n21 0.120292
R58 VPWR.n22 VPWR.n3 0.120292
R59 VPWR.n27 VPWR.n3 0.120292
R60 VPWR.n28 VPWR.n27 0.120292
R61 VPWR.n29 VPWR.n28 0.120292
R62 VPWR.n29 VPWR.n0 0.120292
R63 VPWR VPWR.n33 0.114842
R64 a_600_345.t1 a_600_345.n1 758.737
R65 a_600_345.n0 a_600_345.t2 337.937
R66 a_600_345.n1 a_600_345.t0 293.769
R67 a_600_345.n1 a_600_345.n0 235.905
R68 a_600_345.n0 a_600_345.t3 157.453
R69 VPB.t10 VPB.t1 947.042
R70 VPB.t8 VPB.t10 556.386
R71 VPB.t9 VPB.t6 556.386
R72 VPB.t7 VPB.t11 426.168
R73 VPB.t1 VPB.t3 287.072
R74 VPB.t0 VPB.t5 281.154
R75 VPB.t3 VPB.t2 248.599
R76 VPB.t6 VPB.t8 248.599
R77 VPB.t11 VPB.t9 248.599
R78 VPB.t5 VPB.t7 248.599
R79 VPB.t4 VPB.t0 248.599
R80 VPB VPB.t4 192.369
R81 a_288_47.t3 a_288_47.n3 634.25
R82 a_288_47.n2 a_288_47.n1 622.271
R83 a_288_47.n2 a_288_47.n0 337.471
R84 a_288_47.n3 a_288_47.t5 326.3
R85 a_288_47.n0 a_288_47.t0 66.6672
R86 a_288_47.n0 a_288_47.t1 65.0005
R87 a_288_47.n1 a_288_47.t4 63.3219
R88 a_288_47.n1 a_288_47.t2 63.3219
R89 a_288_47.n3 a_288_47.n2 40.1862
R90 a_788_316.n5 a_788_316.n4 585
R91 a_788_316.n4 a_788_316.n2 313.687
R92 a_788_316.n4 a_788_316.n3 266.853
R93 a_788_316.n0 a_788_316.t6 212.081
R94 a_788_316.n1 a_788_316.t7 212.081
R95 a_788_316.n0 a_788_316.t4 139.78
R96 a_788_316.n1 a_788_316.t5 139.78
R97 a_788_316.n2 a_788_316.n0 56.9641
R98 a_788_316.n5 a_788_316.t3 49.2505
R99 a_788_316.t0 a_788_316.n5 49.2505
R100 a_788_316.n3 a_788_316.t2 40.0005
R101 a_788_316.n3 a_788_316.t1 38.5719
R102 a_788_316.n2 a_788_316.n1 4.38232
R103 VNB.t8 VNB.t0 3089.97
R104 VNB.t10 VNB.t11 2705.5
R105 VNB.t4 VNB.t8 2677.02
R106 VNB.t3 VNB.t1 1552.1
R107 VNB.t12 VNB.t10 1537.86
R108 VNB.t5 VNB.t6 1438.19
R109 VNB.t1 VNB.t12 1366.99
R110 VNB.t0 VNB.t5 1352.75
R111 VNB.t9 VNB.t3 1352.75
R112 VNB.t11 VNB.t4 1210.36
R113 VNB.t6 VNB.t7 1196.12
R114 VNB.t2 VNB.t9 1196.12
R115 VNB VNB.t2 925.567
R116 A3.n0 A3.t0 313.805
R117 A3.n1 A3.n0 152
R118 A3.n0 A3.t1 132.282
R119 A3 A3.n1 8.52135
R120 A3.n1 A3 5.6325
R121 a_372_413.t1 a_372_413.t0 245.006
R122 a_372_413.n0 a_372_413.t1 101.897
R123 a_872_316.t2 a_872_316.n0 639.64
R124 a_872_316.n0 a_872_316.t0 445.173
R125 a_872_316.n0 a_872_316.t1 313.389
R126 S0.n3 S0.t2 459.507
R127 S0.n2 S0.n1 432.193
R128 S0.n5 S0.t0 287.995
R129 S0.n3 S0.t1 265.101
R130 S0.n2 S0.n0 254.389
R131 S0.n5 S0.t3 194.809
R132 S0.n4 S0.n3 172.971
R133 S0.n4 S0.n2 171.157
R134 S0.n6 S0.n5 152
R135 S0 S0.n6 20.2672
R136 S0 S0.n4 16.0651
R137 S0.n6 S0 3.91161
R138 a_27_47.t1 a_27_47.n4 663.449
R139 a_27_47.n4 a_27_47.t0 336.815
R140 a_27_47.n2 a_27_47.t4 322.296
R141 a_27_47.n1 a_27_47.t2 314.822
R142 a_27_47.n2 a_27_47.t3 300.252
R143 a_27_47.n1 a_27_47.n0 300.252
R144 a_27_47.n4 a_27_47.n3 67.3887
R145 a_27_47.n3 a_27_47.n1 27.9335
R146 a_27_47.n3 a_27_47.n2 4.89462
R147 a_1279_413.n0 a_1279_413.t0 111.359
R148 X.n0 X 590.152
R149 X.n1 X.n0 585
R150 X.n4 X.n3 185
R151 X.n4 X 81.3936
R152 X.n0 X.t3 26.5955
R153 X.n0 X.t2 26.5955
R154 X.n3 X.t1 24.9236
R155 X.n3 X.t0 24.9236
R156 X.n1 X 6.4005
R157 X.n2 X.n1 2.65416
R158 X X.n2 2.06502
R159 X.n2 X 1.56148
R160 X X.n4 0.194439
R161 VGND.n16 VGND.t3 238.311
R162 VGND.n9 VGND.n8 211.601
R163 VGND.n24 VGND.n23 199.739
R164 VGND.n31 VGND.n30 199.739
R165 VGND.n7 VGND.t2 162.327
R166 VGND.n8 VGND.t0 62.3526
R167 VGND.n23 VGND.t6 57.1434
R168 VGND.n23 VGND.t7 54.2862
R169 VGND.n30 VGND.t4 38.5719
R170 VGND.n30 VGND.t5 38.5719
R171 VGND.n11 VGND.n10 34.6358
R172 VGND.n11 VGND.n5 34.6358
R173 VGND.n15 VGND.n5 34.6358
R174 VGND.n17 VGND.n3 34.6358
R175 VGND.n21 VGND.n3 34.6358
R176 VGND.n22 VGND.n21 34.6358
R177 VGND.n28 VGND.n1 34.6358
R178 VGND.n29 VGND.n28 34.6358
R179 VGND.n17 VGND.n16 32.0005
R180 VGND.n24 VGND.n1 28.6123
R181 VGND.n10 VGND.n9 25.977
R182 VGND.n8 VGND.t1 24.9241
R183 VGND.n31 VGND.n29 22.9652
R184 VGND.n24 VGND.n22 15.8123
R185 VGND.n16 VGND.n15 12.424
R186 VGND.n29 VGND.n0 9.3005
R187 VGND.n28 VGND.n27 9.3005
R188 VGND.n26 VGND.n1 9.3005
R189 VGND.n25 VGND.n24 9.3005
R190 VGND.n22 VGND.n2 9.3005
R191 VGND.n21 VGND.n20 9.3005
R192 VGND.n19 VGND.n3 9.3005
R193 VGND.n18 VGND.n17 9.3005
R194 VGND.n16 VGND.n4 9.3005
R195 VGND.n15 VGND.n14 9.3005
R196 VGND.n13 VGND.n5 9.3005
R197 VGND.n12 VGND.n11 9.3005
R198 VGND.n10 VGND.n6 9.3005
R199 VGND.n32 VGND.n31 7.12063
R200 VGND.n9 VGND.n7 6.73566
R201 VGND.n7 VGND.n6 0.589728
R202 VGND.n32 VGND.n0 0.148519
R203 VGND.n12 VGND.n6 0.120292
R204 VGND.n13 VGND.n12 0.120292
R205 VGND.n14 VGND.n13 0.120292
R206 VGND.n14 VGND.n4 0.120292
R207 VGND.n18 VGND.n4 0.120292
R208 VGND.n19 VGND.n18 0.120292
R209 VGND.n20 VGND.n19 0.120292
R210 VGND.n20 VGND.n2 0.120292
R211 VGND.n25 VGND.n2 0.120292
R212 VGND.n26 VGND.n25 0.120292
R213 VGND.n27 VGND.n26 0.120292
R214 VGND.n27 VGND.n0 0.120292
R215 VGND VGND.n32 0.114842
R216 A1.n0 A1.t0 266.14
R217 A1.n0 A1.t1 217.94
R218 A1 A1.n0 156.325
R219 a_1060_369.n0 a_1060_369.t0 41.2767
R220 A2.n0 A2.t1 372.868
R221 A2 A2.n0 157.625
R222 A2.n0 A2.t0 132.282
R223 a_193_47.n0 a_193_47.t1 66.6672
R224 a_193_47.n0 a_193_47.t0 26.3935
R225 a_193_47.n1 a_193_47.n0 14.4005
R226 a_1064_47.n0 a_1064_47.t0 38.9529
R227 a_1281_47.t1 a_1281_47.t0 93.0601
R228 a_397_47.t1 a_397_47.t0 93.5174
R229 a_193_369.t0 a_193_369.t1 132.286
R230 A0.n0 A0.t1 299.377
R231 A0.n0 A0.t0 206.19
R232 A0 A0.n0 181.006
C0 VGND A3 0.041113f
C1 X VPWR 0.191335f
C2 S0 A0 0.053348f
C3 VPWR S1 0.055891f
C4 VGND X 0.143747f
C5 VGND S1 0.035291f
C6 A3 S1 0.132409f
C7 VPWR A1 0.012097f
C8 VGND A1 0.049336f
C9 X S1 1.11e-19
C10 VPWR A0 0.012367f
C11 VGND A0 0.084706f
C12 S1 A1 0.006345f
C13 VPB S0 0.274332f
C14 X A0 0.007586f
C15 VPB A2 0.042858f
C16 S0 A2 0.169993f
C17 VPB VPWR 0.18178f
C18 VGND VPB 0.013573f
C19 VPB A3 0.061927f
C20 S0 VPWR 0.098721f
C21 VGND S0 0.235037f
C22 X VPB 0.005146f
C23 S0 A3 0.063625f
C24 A2 VPWR 0.013413f
C25 VPB S1 0.20632f
C26 X S0 0.001187f
C27 VGND A2 0.049946f
C28 VPB A1 0.078954f
C29 S0 S1 0.020079f
C30 VGND VPWR 0.053361f
C31 VPWR A3 0.018882f
C32 S0 A1 0.060803f
C33 VPB A0 0.057378f
C34 X VNB 0.025732f
C35 VGND VNB 0.969275f
C36 A0 VNB 0.129327f
C37 A1 VNB 0.140821f
C38 S1 VNB 0.29851f
C39 A3 VNB 0.118003f
C40 VPWR VNB 0.799468f
C41 A2 VNB 0.113101f
C42 S0 VNB 0.489648f
C43 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux4_4 VNB VPB VGND VPWR S0 A2 A3 S1 A1 A0 X
X0 X.t3 a_789_316.t4 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X1 X.t7 a_789_316.t5 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X2 VPWR.t7 A0.t0 a_1280_413.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.10535 ps=0.995 w=0.64 l=0.15
X3 a_873_316.t2 a_601_345.t2 a_789_316.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X4 a_601_345.t0 S1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VPWR.t9 S0.t0 a_27_47.t0 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 VGND.t4 a_789_316.t6 X.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.21775 pd=1.97 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t3 a_789_316.t7 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t2 A3.t0 a_373_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1645 ps=1.33 w=0.64 l=0.15
X9 a_1280_413.t1 S0.t1 a_873_316.t4 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.10535 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_1065_47.t0 A1.t0 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_1282_47.t1 a_27_47.t2 a_873_316.t1 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X12 a_193_47.t0 A2.t0 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_873_316.t5 S0.t2 a_1065_47.t1 VNB.t13 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0786 ps=0.805 w=0.36 l=0.15
X14 X.t0 a_789_316.t8 VGND.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X15 a_1061_369.t0 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.13775 pd=1.165 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 a_873_316.t0 a_27_47.t3 a_1061_369.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.13775 ps=1.165 w=0.42 l=0.15
X17 VPWR.t5 a_789_316.t9 X.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.135 ps=1.27 w=1 l=0.15
X18 X.t5 a_789_316.t10 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X19 VGND.t2 A3.t1 a_398_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.06705 ps=0.75 w=0.42 l=0.15
X20 a_601_345.t1 S1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 a_873_316.t3 S1.t2 a_789_316.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1404 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X22 a_193_369.t0 A2.t1 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.09735 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_789_316.t2 a_601_345.t3 a_288_47.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.1404 ps=1.6 w=0.54 l=0.15
X24 a_398_47.t0 S0.t3 a_288_47.t1 VNB.t14 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X25 VGND.t0 A0.t1 a_1282_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.066 ps=0.745 w=0.42 l=0.15
X26 a_373_413.t1 a_27_47.t4 a_288_47.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1645 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X27 a_288_47.t2 a_27_47.t5 a_193_47.t1 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X28 VPWR.t3 a_789_316.t11 X.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X29 a_288_47.t0 S0.t4 a_193_369.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09735 ps=0.97 w=0.42 l=0.15
X30 VGND.t9 S0.t5 a_27_47.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_789_316.t0 S1.t3 a_288_47.t5 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_789_316.n7 a_789_316.n6 585
R1 a_789_316.n6 a_789_316.n4 313.687
R2 a_789_316.n6 a_789_316.n5 266.853
R3 a_789_316.n0 a_789_316.t9 212.081
R4 a_789_316.n1 a_789_316.t10 212.081
R5 a_789_316.n2 a_789_316.t11 212.081
R6 a_789_316.n3 a_789_316.t5 212.081
R7 a_789_316.n0 a_789_316.t6 139.78
R8 a_789_316.n1 a_789_316.t4 139.78
R9 a_789_316.n2 a_789_316.t7 139.78
R10 a_789_316.n3 a_789_316.t8 139.78
R11 a_789_316.n2 a_789_316.n1 73.0308
R12 a_789_316.n1 a_789_316.n0 61.346
R13 a_789_316.n4 a_789_316.n2 56.9641
R14 a_789_316.n7 a_789_316.t3 49.2505
R15 a_789_316.t2 a_789_316.n7 49.2505
R16 a_789_316.n5 a_789_316.t0 40.0005
R17 a_789_316.n5 a_789_316.t1 38.5719
R18 a_789_316.n4 a_789_316.n3 4.38232
R19 VGND.n21 VGND.t8 238.311
R20 VGND.n14 VGND.n8 211.601
R21 VGND.n29 VGND.n28 199.739
R22 VGND.n36 VGND.n35 199.739
R23 VGND.n11 VGND.t4 161.858
R24 VGND.n10 VGND.n9 116.112
R25 VGND.n8 VGND.t0 62.3526
R26 VGND.n28 VGND.t1 57.1434
R27 VGND.n28 VGND.t2 54.2862
R28 VGND.n9 VGND.t3 39.6928
R29 VGND.n35 VGND.t7 38.5719
R30 VGND.n35 VGND.t9 38.5719
R31 VGND.n16 VGND.n15 34.6358
R32 VGND.n16 VGND.n5 34.6358
R33 VGND.n20 VGND.n5 34.6358
R34 VGND.n22 VGND.n3 34.6358
R35 VGND.n26 VGND.n3 34.6358
R36 VGND.n27 VGND.n26 34.6358
R37 VGND.n33 VGND.n1 34.6358
R38 VGND.n34 VGND.n33 34.6358
R39 VGND.n22 VGND.n21 32.377
R40 VGND.n29 VGND.n1 28.9887
R41 VGND.n10 VGND.n7 26.3534
R42 VGND.n15 VGND.n14 26.3534
R43 VGND.n8 VGND.t6 24.9241
R44 VGND.n9 VGND.t5 24.9236
R45 VGND.n14 VGND.n7 24.0946
R46 VGND.n36 VGND.n34 22.9652
R47 VGND.n29 VGND.n27 15.4358
R48 VGND.n21 VGND.n20 12.0476
R49 VGND.n34 VGND.n0 9.3005
R50 VGND.n33 VGND.n32 9.3005
R51 VGND.n31 VGND.n1 9.3005
R52 VGND.n30 VGND.n29 9.3005
R53 VGND.n27 VGND.n2 9.3005
R54 VGND.n26 VGND.n25 9.3005
R55 VGND.n24 VGND.n3 9.3005
R56 VGND.n23 VGND.n22 9.3005
R57 VGND.n21 VGND.n4 9.3005
R58 VGND.n20 VGND.n19 9.3005
R59 VGND.n18 VGND.n5 9.3005
R60 VGND.n17 VGND.n16 9.3005
R61 VGND.n15 VGND.n6 9.3005
R62 VGND.n14 VGND.n13 9.3005
R63 VGND.n12 VGND.n7 9.3005
R64 VGND.n37 VGND.n36 7.12063
R65 VGND.n11 VGND.n10 6.71203
R66 VGND.n12 VGND.n11 0.594047
R67 VGND.n37 VGND.n0 0.148519
R68 VGND.n13 VGND.n12 0.120292
R69 VGND.n13 VGND.n6 0.120292
R70 VGND.n17 VGND.n6 0.120292
R71 VGND.n18 VGND.n17 0.120292
R72 VGND.n19 VGND.n18 0.120292
R73 VGND.n19 VGND.n4 0.120292
R74 VGND.n23 VGND.n4 0.120292
R75 VGND.n24 VGND.n23 0.120292
R76 VGND.n25 VGND.n24 0.120292
R77 VGND.n25 VGND.n2 0.120292
R78 VGND.n30 VGND.n2 0.120292
R79 VGND.n31 VGND.n30 0.120292
R80 VGND.n32 VGND.n31 0.120292
R81 VGND.n32 VGND.n0 0.120292
R82 VGND VGND.n37 0.11354
R83 X.n6 X 591.499
R84 X.n7 X.n6 585
R85 X.n2 X.n0 326.36
R86 X.n2 X.n1 217
R87 X.n4 X.n3 185
R88 X.n5 X.n2 36.0005
R89 X.n6 X.t6 26.5955
R90 X.n6 X.t5 26.5955
R91 X.n0 X.t4 26.5955
R92 X.n0 X.t7 26.5955
R93 X.n3 X.t2 24.9236
R94 X.n3 X.t3 24.9236
R95 X.n1 X.t1 24.9236
R96 X.n1 X.t0 24.9236
R97 X X.n5 10.2405
R98 X.n7 X 8.46819
R99 X X.n4 8.07435
R100 X.n4 X 5.31742
R101 X X.n7 4.92358
R102 X.n5 X 3.15127
R103 VNB.t2 VNB.t0 2705.5
R104 VNB.t9 VNB.t12 2677.02
R105 VNB.t13 VNB.t11 1566.34
R106 VNB.t8 VNB.t14 1566.34
R107 VNB.t3 VNB.t2 1537.86
R108 VNB.t12 VNB.t13 1523.62
R109 VNB.t1 VNB.t4 1438.19
R110 VNB.t5 VNB.t7 1423.95
R111 VNB.t14 VNB.t3 1366.99
R112 VNB.t11 VNB.t1 1352.75
R113 VNB.t10 VNB.t8 1352.75
R114 VNB.t0 VNB.t9 1210.36
R115 VNB.t7 VNB.t6 1196.12
R116 VNB.t4 VNB.t5 1196.12
R117 VNB.t15 VNB.t10 1196.12
R118 VNB VNB.t15 911.327
R119 VPWR.n24 VPWR.t1 646.962
R120 VPWR.n31 VPWR.n4 612.827
R121 VPWR.n38 VPWR.n1 599.74
R122 VPWR.n17 VPWR.n9 320.976
R123 VPWR.n13 VPWR.t5 272.214
R124 VPWR.n12 VPWR.n11 223.869
R125 VPWR.n9 VPWR.t7 61.563
R126 VPWR.n11 VPWR.t3 42.3555
R127 VPWR.n1 VPWR.t8 41.5552
R128 VPWR.n1 VPWR.t9 41.5552
R129 VPWR.n4 VPWR.t0 41.5552
R130 VPWR.n4 VPWR.t2 41.5552
R131 VPWR.n32 VPWR.n2 34.6358
R132 VPWR.n36 VPWR.n2 34.6358
R133 VPWR.n37 VPWR.n36 34.6358
R134 VPWR.n25 VPWR.n5 34.6358
R135 VPWR.n29 VPWR.n5 34.6358
R136 VPWR.n30 VPWR.n29 34.6358
R137 VPWR.n16 VPWR.n10 34.6358
R138 VPWR.n19 VPWR.n18 34.6358
R139 VPWR.n19 VPWR.n7 34.6358
R140 VPWR.n23 VPWR.n7 34.6358
R141 VPWR.n18 VPWR.n17 32.7534
R142 VPWR.n9 VPWR.t6 30.5947
R143 VPWR.n25 VPWR.n24 29.3652
R144 VPWR.n11 VPWR.t4 26.5955
R145 VPWR.n12 VPWR.n10 26.3534
R146 VPWR.n38 VPWR.n37 22.9652
R147 VPWR.n24 VPWR.n23 13.9299
R148 VPWR.n31 VPWR.n30 12.0476
R149 VPWR.n14 VPWR.n10 9.3005
R150 VPWR.n16 VPWR.n15 9.3005
R151 VPWR.n18 VPWR.n8 9.3005
R152 VPWR.n20 VPWR.n19 9.3005
R153 VPWR.n21 VPWR.n7 9.3005
R154 VPWR.n23 VPWR.n22 9.3005
R155 VPWR.n24 VPWR.n6 9.3005
R156 VPWR.n26 VPWR.n25 9.3005
R157 VPWR.n27 VPWR.n5 9.3005
R158 VPWR.n29 VPWR.n28 9.3005
R159 VPWR.n30 VPWR.n3 9.3005
R160 VPWR.n33 VPWR.n32 9.3005
R161 VPWR.n34 VPWR.n2 9.3005
R162 VPWR.n36 VPWR.n35 9.3005
R163 VPWR.n37 VPWR.n0 9.3005
R164 VPWR.n39 VPWR.n38 7.12063
R165 VPWR.n13 VPWR.n12 6.71203
R166 VPWR.n32 VPWR.n31 5.27109
R167 VPWR.n17 VPWR.n16 1.88285
R168 VPWR.n14 VPWR.n13 0.594047
R169 VPWR.n39 VPWR.n0 0.148519
R170 VPWR.n15 VPWR.n14 0.120292
R171 VPWR.n15 VPWR.n8 0.120292
R172 VPWR.n20 VPWR.n8 0.120292
R173 VPWR.n21 VPWR.n20 0.120292
R174 VPWR.n22 VPWR.n21 0.120292
R175 VPWR.n22 VPWR.n6 0.120292
R176 VPWR.n26 VPWR.n6 0.120292
R177 VPWR.n27 VPWR.n26 0.120292
R178 VPWR.n28 VPWR.n27 0.120292
R179 VPWR.n28 VPWR.n3 0.120292
R180 VPWR.n33 VPWR.n3 0.120292
R181 VPWR.n34 VPWR.n33 0.120292
R182 VPWR.n35 VPWR.n34 0.120292
R183 VPWR.n35 VPWR.n0 0.120292
R184 VPWR VPWR.n39 0.11354
R185 VPB.t12 VPB.t1 556.386
R186 VPB.t0 VPB.t9 556.386
R187 VPB.t8 VPB.t2 426.168
R188 VPB.t1 VPB.t7 399.534
R189 VPB.t14 VPB.t10 298.911
R190 VPB.t3 VPB.t4 295.95
R191 VPB.t10 VPB.t6 287.072
R192 VPB.t11 VPB.t15 284.113
R193 VPB.t4 VPB.t5 248.599
R194 VPB.t6 VPB.t3 248.599
R195 VPB.t7 VPB.t14 248.599
R196 VPB.t9 VPB.t12 248.599
R197 VPB.t2 VPB.t0 248.599
R198 VPB.t15 VPB.t8 248.599
R199 VPB.t13 VPB.t11 248.599
R200 VPB VPB.t13 189.409
R201 A0.n0 A0.t0 299.377
R202 A0.n0 A0.t1 206.19
R203 A0 A0.n0 181.006
R204 a_1280_413.n0 a_1280_413.t1 100.846
R205 a_1280_413.n1 a_1280_413.n0 77.3934
R206 a_1280_413.n0 a_1280_413.t0 33.966
R207 a_601_345.t0 a_601_345.n1 758.737
R208 a_601_345.n0 a_601_345.t2 337.937
R209 a_601_345.n1 a_601_345.t1 293.769
R210 a_601_345.n1 a_601_345.n0 235.905
R211 a_601_345.n0 a_601_345.t3 157.453
R212 a_873_316.n2 a_873_316.n0 669.33
R213 a_873_316.t3 a_873_316.n3 639.64
R214 a_873_316.n2 a_873_316.n1 316.389
R215 a_873_316.n3 a_873_316.t2 313.389
R216 a_873_316.n1 a_873_316.t1 66.6672
R217 a_873_316.n1 a_873_316.t5 66.6672
R218 a_873_316.n0 a_873_316.t4 63.3219
R219 a_873_316.n0 a_873_316.t0 63.3219
R220 a_873_316.n3 a_873_316.n2 62.1181
R221 S1.t0 S1.t2 769.593
R222 S1.n0 S1.t3 367.928
R223 S1.n1 S1.t0 350.712
R224 S1.n2 S1.n1 152
R225 S1.n0 S1.t1 112.237
R226 S1.n1 S1.n0 34.4291
R227 S1.n2 S1 7.72464
R228 S1 S1.n2 7.28326
R229 S0.n1 S0.t3 459.507
R230 S0.n0 S0.t2 432.193
R231 S0.n3 S0.t0 287.995
R232 S0.n1 S0.t4 265.101
R233 S0.n0 S0.t1 254.389
R234 S0.n3 S0.t5 194.809
R235 S0.n2 S0.n1 172.971
R236 S0.n2 S0.n0 171.157
R237 S0.n4 S0.n3 152
R238 S0 S0.n4 20.2672
R239 S0 S0.n2 16.0651
R240 S0.n4 S0 3.91161
R241 a_27_47.t0 a_27_47.n3 660.813
R242 a_27_47.n3 a_27_47.t1 334.63
R243 a_27_47.n1 a_27_47.t5 321.947
R244 a_27_47.n0 a_27_47.t2 314.822
R245 a_27_47.n1 a_27_47.t4 300.252
R246 a_27_47.n0 a_27_47.t3 300.252
R247 a_27_47.n3 a_27_47.n2 67.3887
R248 a_27_47.n2 a_27_47.n0 27.9335
R249 a_27_47.n2 a_27_47.n1 4.89462
R250 A3.n0 A3.t0 313.805
R251 A3.n1 A3.n0 152
R252 A3.n0 A3.t1 132.282
R253 A3 A3.n1 8.52135
R254 A3.n1 A3 5.6325
R255 a_373_413.t0 a_373_413.t1 245.006
R256 a_373_413.n0 a_373_413.t0 101.897
R257 A1.n0 A1.t1 282.238
R258 A1.n0 A1.t0 247.428
R259 A1 A1.n0 173.731
R260 a_1065_47.n0 a_1065_47.t1 76.6672
R261 a_1065_47.n0 a_1065_47.t0 27.34
R262 a_1065_47.n1 a_1065_47.n0 11.6134
R263 a_1282_47.t0 a_1282_47.t1 93.0601
R264 A2.n0 A2.t1 373.283
R265 A2 A2.n0 157.625
R266 A2.n0 A2.t0 132.282
R267 a_193_47.n0 a_193_47.t1 66.6672
R268 a_193_47.n0 a_193_47.t0 26.3935
R269 a_193_47.n1 a_193_47.n0 14.4005
R270 a_1061_369.t0 a_1061_369.t1 226.096
R271 a_398_47.t1 a_398_47.t0 93.5174
R272 a_193_369.t0 a_193_369.t1 134.631
R273 a_288_47.t4 a_288_47.n3 634.25
R274 a_288_47.n2 a_288_47.n1 622.271
R275 a_288_47.n2 a_288_47.n0 337.471
R276 a_288_47.n3 a_288_47.t5 326.466
R277 a_288_47.n0 a_288_47.t1 66.6672
R278 a_288_47.n0 a_288_47.t2 66.6672
R279 a_288_47.n1 a_288_47.t3 63.3219
R280 a_288_47.n1 a_288_47.t0 63.3219
R281 a_288_47.n3 a_288_47.n2 40.7986
C0 S0 A2 0.168608f
C1 VPB VPWR 0.198756f
C2 A0 S0 0.053348f
C3 VGND VPB 0.014118f
C4 S0 VPWR 0.098521f
C5 VPB A3 0.061928f
C6 VGND S0 0.234501f
C7 X VPB 0.010946f
C8 VPB S1 0.206585f
C9 A2 VPWR 0.013392f
C10 S0 A3 0.063625f
C11 VGND A2 0.049706f
C12 A0 VPWR 0.012617f
C13 X S0 0.001624f
C14 A0 VGND 0.084882f
C15 S0 S1 0.020079f
C16 VPB A1 0.07876f
C17 VGND VPWR 0.072981f
C18 A0 X 0.008147f
C19 S0 A1 0.060338f
C20 VPWR A3 0.018691f
C21 X VPWR 0.431355f
C22 VGND A3 0.040974f
C23 VGND X 0.328367f
C24 VPWR S1 0.055682f
C25 VGND S1 0.034993f
C26 A3 S1 0.132409f
C27 VPWR A1 0.011926f
C28 VGND A1 0.049089f
C29 X S1 1.64e-19
C30 S1 A1 0.006345f
C31 VPB S0 0.275045f
C32 VPB A2 0.042784f
C33 A0 VPB 0.058697f
C34 X VNB 0.031735f
C35 VGND VNB 1.06029f
C36 A0 VNB 0.128008f
C37 A1 VNB 0.140821f
C38 S1 VNB 0.298245f
C39 A3 VNB 0.118001f
C40 VPWR VNB 0.873943f
C41 A2 VNB 0.113118f
C42 S0 VNB 0.487986f
C43 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_2 VNB VPB VGND VPWR A_N Y B
X0 Y.t2 B.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND.t2 A_N.t0 a_27_93.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND.t0 B.t1 a_229_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t4 a_27_93.t2 a_229_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47.t2 a_27_93.t3 Y.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t0 a_27_93.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X6 VPWR.t3 a_27_93.t5 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR.t1 B.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47.t0 B.t3 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t4 A_N.t1 a_27_93.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 B.n0 B.t3 869.207
R1 B.n2 B.t0 232.431
R2 B.n1 B.t2 218.507
R3 B.n0 B 164.889
R4 B.n4 B.n3 152
R5 B.n2 B.t1 149.421
R6 B.n3 B.n1 37.0112
R7 B.n1 B.n0 36.1505
R8 B.n4 B 28.1605
R9 B.n3 B.n2 26.7783
R10 B B.n4 1.2805
R11 VPWR.n3 VPWR.n2 585
R12 VPWR.n5 VPWR.n4 585
R13 VPWR.n10 VPWR.n1 317.478
R14 VPWR.n6 VPWR.t1 250.245
R15 VPWR.n1 VPWR.t4 98.5005
R16 VPWR.n4 VPWR.n3 66.9805
R17 VPWR.n4 VPWR.t2 38.4155
R18 VPWR.n9 VPWR.n8 30.5125
R19 VPWR.n3 VPWR.t3 26.5955
R20 VPWR.n1 VPWR.t0 25.6105
R21 VPWR.n10 VPWR.n9 23.7181
R22 VPWR.n8 VPWR.n7 9.3005
R23 VPWR.n9 VPWR.n0 9.3005
R24 VPWR.n6 VPWR.n5 8.71508
R25 VPWR.n11 VPWR.n10 7.35738
R26 VPWR.n5 VPWR.n2 6.90844
R27 VPWR.n8 VPWR.n2 0.813198
R28 VPWR.n7 VPWR.n6 0.565684
R29 VPWR.n11 VPWR.n0 0.145509
R30 VPWR.n7 VPWR.n0 0.120292
R31 VPWR VPWR.n11 0.11659
R32 Y.n2 Y.n0 311.288
R33 Y.n2 Y.n1 234.264
R34 Y Y.n3 187.058
R35 Y.n0 Y.t3 32.5055
R36 Y.n0 Y.t0 32.5055
R37 Y.n1 Y.t1 26.5955
R38 Y.n1 Y.t2 26.5955
R39 Y.n3 Y.t5 24.9236
R40 Y.n3 Y.t4 24.9236
R41 Y Y.n2 6.17193
R42 VPB.t3 VPB.t2 485.358
R43 VPB.t4 VPB.t0 290.031
R44 VPB.t0 VPB.t3 284.113
R45 VPB.t2 VPB.t1 248.599
R46 VPB VPB.t4 189.409
R47 A_N A_N.n0 154.715
R48 A_N.n0 A_N.t1 147.298
R49 A_N.n0 A_N.t0 131.231
R50 a_27_93.t0 a_27_93.n3 648.322
R51 a_27_93.n3 a_27_93.t1 284.156
R52 a_27_93.n2 a_27_93.t4 263.673
R53 a_27_93.n0 a_27_93.t3 224.399
R54 a_27_93.n1 a_27_93.t5 221.72
R55 a_27_93.n3 a_27_93.n2 220.234
R56 a_27_93.n0 a_27_93.t2 149.421
R57 a_27_93.n2 a_27_93.n1 43.7375
R58 a_27_93.n1 a_27_93.n0 7.14124
R59 VGND.n1 VGND.n0 212.631
R60 VGND.n1 VGND.t2 168.487
R61 VGND.n0 VGND.t1 24.9236
R62 VGND.n0 VGND.t0 24.9236
R63 VGND VGND.n1 0.155311
R64 VNB.t4 VNB.t3 2876.38
R65 VNB.t1 VNB.t0 1196.12
R66 VNB.t2 VNB.t1 1196.12
R67 VNB.t3 VNB.t2 1196.12
R68 VNB VNB.t4 911.327
R69 a_229_47.n0 a_229_47.t3 186.775
R70 a_229_47.n0 a_229_47.t0 181.044
R71 a_229_47.n1 a_229_47.n0 88.3446
R72 a_229_47.t1 a_229_47.n1 24.9236
R73 a_229_47.n1 a_229_47.t2 24.9236
C0 B VPB 0.082971f
C1 VPWR VPB 0.092473f
C2 A_N VPB 0.037697f
C3 B VPWR 0.071341f
C4 Y VPB 0.006317f
C5 VGND VPB 0.007778f
C6 B Y 0.136294f
C7 VPWR A_N 0.008542f
C8 B VGND 0.031145f
C9 VPWR Y 0.367782f
C10 A_N Y 0.00387f
C11 VPWR VGND 0.066989f
C12 A_N VGND 0.042341f
C13 Y VGND 0.011854f
C14 VGND VNB 0.411323f
C15 Y VNB 0.009401f
C16 A_N VNB 0.124489f
C17 VPWR VNB 0.375429f
C18 B VNB 0.245378f
C19 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_4 VNB VPB VGND VPWR A_N Y B
X0 VGND.t4 B.t0 a_215_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X1 Y.t9 B.t1 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X2 Y.t1 a_27_47.t2 a_215_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VGND.t3 B.t2 a_215_47.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t10 a_27_47.t3 a_215_47.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_215_47.t7 a_27_47.t4 Y.t11 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_215_47.t3 B.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t7 B.t4 Y.t8 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t0 a_27_47.t5 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t7 B.t5 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t5 B.t6 Y.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y.t2 a_27_47.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR.t3 a_27_47.t7 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_215_47.t2 B.t7 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_215_47.t1 a_27_47.t8 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y.t5 a_27_47.t9 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR.t1 A_N.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X17 VGND.t0 A_N.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n1 B.t4 221.72
R1 B.n5 B.t5 221.72
R2 B.n7 B.t6 221.72
R3 B.n8 B.t1 221.72
R4 B.n2 B.n1 194.845
R5 B B.n9 156.481
R6 B.n4 B.n3 152
R7 B.n6 B.n0 152
R8 B.n1 B.t3 149.421
R9 B.n5 B.t2 149.421
R10 B.n7 B.t7 149.421
R11 B.n8 B.t0 149.421
R12 B.n4 B.n1 38.382
R13 B.n9 B.n8 38.382
R14 B.n6 B.n5 37.4894
R15 B.n7 B.n6 37.4894
R16 B.n5 B.n4 36.5968
R17 B.n9 B.n7 36.5968
R18 B B.n0 22.0805
R19 B.n3 B 19.2005
R20 B B.n2 18.8805
R21 B.n2 B 10.5605
R22 B.n3 B 10.2405
R23 B B.n0 7.3605
R24 a_215_47.n1 a_215_47.t3 186.175
R25 a_215_47.n5 a_215_47.n4 185
R26 a_215_47.t0 a_215_47.n5 183.096
R27 a_215_47.n1 a_215_47.n0 99.1759
R28 a_215_47.n3 a_215_47.n2 88.3446
R29 a_215_47.n5 a_215_47.n3 56.2712
R30 a_215_47.n3 a_215_47.n1 47.2798
R31 a_215_47.n2 a_215_47.t7 27.6928
R32 a_215_47.n4 a_215_47.t6 24.9236
R33 a_215_47.n4 a_215_47.t1 24.9236
R34 a_215_47.n2 a_215_47.t5 24.9236
R35 a_215_47.n0 a_215_47.t4 24.9236
R36 a_215_47.n0 a_215_47.t2 24.9236
R37 VGND.n14 VGND.t0 293.022
R38 VGND.n5 VGND.n4 212.31
R39 VGND.n6 VGND.n3 207.213
R40 VGND.n8 VGND.n7 34.6358
R41 VGND.n8 VGND.n1 34.6358
R42 VGND.n12 VGND.n1 34.6358
R43 VGND.n13 VGND.n12 34.6358
R44 VGND.n14 VGND.n13 27.1064
R45 VGND.n4 VGND.t2 24.9236
R46 VGND.n4 VGND.t3 24.9236
R47 VGND.n3 VGND.t1 24.9236
R48 VGND.n3 VGND.t4 24.9236
R49 VGND.n7 VGND.n6 24.4711
R50 VGND.n6 VGND.n5 17.1176
R51 VGND.n7 VGND.n2 9.3005
R52 VGND.n9 VGND.n8 9.3005
R53 VGND.n10 VGND.n1 9.3005
R54 VGND.n12 VGND.n11 9.3005
R55 VGND.n13 VGND.n0 9.3005
R56 VGND.n15 VGND.n14 7.4049
R57 VGND.n5 VGND.n2 0.765894
R58 VGND.n15 VGND.n0 0.144904
R59 VGND.n9 VGND.n2 0.120292
R60 VGND.n10 VGND.n9 0.120292
R61 VGND.n11 VGND.n10 0.120292
R62 VGND.n11 VGND.n0 0.120292
R63 VGND VGND.n15 0.117202
R64 VNB.t2 VNB.t0 2677.02
R65 VNB.t8 VNB.t6 1238.83
R66 VNB.t5 VNB.t4 1196.12
R67 VNB.t3 VNB.t5 1196.12
R68 VNB.t6 VNB.t3 1196.12
R69 VNB.t7 VNB.t8 1196.12
R70 VNB.t1 VNB.t7 1196.12
R71 VNB.t0 VNB.t1 1196.12
R72 VNB VNB.t2 911.327
R73 VPWR.n16 VPWR.n2 320.976
R74 VPWR.n10 VPWR.n9 320.976
R75 VPWR.n7 VPWR.n5 320.976
R76 VPWR.n1 VPWR.t1 318.582
R77 VPWR.n6 VPWR.t7 271.024
R78 VPWR.n1 VPWR.t4 223.397
R79 VPWR.n11 VPWR.n8 34.6358
R80 VPWR.n15 VPWR.n3 34.6358
R81 VPWR.n17 VPWR.n16 32.377
R82 VPWR.n9 VPWR.t0 29.5505
R83 VPWR.n10 VPWR.n3 27.4829
R84 VPWR.n2 VPWR.t2 26.5955
R85 VPWR.n2 VPWR.t3 26.5955
R86 VPWR.n9 VPWR.t8 26.5955
R87 VPWR.n5 VPWR.t6 26.5955
R88 VPWR.n5 VPWR.t5 26.5955
R89 VPWR.n18 VPWR.n17 24.4711
R90 VPWR.n8 VPWR.n7 21.4593
R91 VPWR.n7 VPWR.n6 20.204
R92 VPWR.n8 VPWR.n4 9.3005
R93 VPWR.n12 VPWR.n11 9.3005
R94 VPWR.n13 VPWR.n3 9.3005
R95 VPWR.n15 VPWR.n14 9.3005
R96 VPWR.n17 VPWR.n0 9.3005
R97 VPWR.n18 VPWR.n1 9.12091
R98 VPWR.n11 VPWR.n10 7.15344
R99 VPWR.n19 VPWR.n18 4.0883
R100 VPWR.n16 VPWR.n15 2.25932
R101 VPWR.n6 VPWR.n4 0.680746
R102 VPWR.n19 VPWR.n0 0.200784
R103 VPWR VPWR.n19 0.18088
R104 VPWR.n12 VPWR.n4 0.120292
R105 VPWR.n13 VPWR.n12 0.120292
R106 VPWR.n14 VPWR.n13 0.120292
R107 VPWR.n14 VPWR.n0 0.120292
R108 Y.n9 Y.n4 235.923
R109 Y.n7 Y.n5 235.923
R110 Y.n2 Y.n0 224.822
R111 Y.n7 Y.n6 206.25
R112 Y.n9 Y.n8 205.768
R113 Y.n2 Y.n1 185
R114 Y.n9 Y.n7 29.6732
R115 Y.n8 Y.t0 26.5955
R116 Y.n8 Y.t2 26.5955
R117 Y.n5 Y.t8 26.5955
R118 Y.n5 Y.t7 26.5955
R119 Y.n6 Y.t6 26.5955
R120 Y.n6 Y.t9 26.5955
R121 Y.n4 Y.t3 26.5955
R122 Y.n4 Y.t5 26.5955
R123 Y.n0 Y.t4 24.9236
R124 Y.n0 Y.t1 24.9236
R125 Y.n1 Y.t11 24.9236
R126 Y.n1 Y.t10 24.9236
R127 Y Y.n3 9.66088
R128 Y.n3 Y 6.76276
R129 Y Y.n9 4.08166
R130 Y.n3 Y 1.65976
R131 Y Y.n2 0.474574
R132 VPB.t1 VPB.t4 556.386
R133 VPB.t0 VPB.t8 257.478
R134 VPB.t6 VPB.t7 248.599
R135 VPB.t5 VPB.t6 248.599
R136 VPB.t8 VPB.t5 248.599
R137 VPB.t2 VPB.t0 248.599
R138 VPB.t3 VPB.t2 248.599
R139 VPB.t4 VPB.t3 248.599
R140 VPB VPB.t1 189.409
R141 a_27_47.t0 a_27_47.n8 261.188
R142 a_27_47.n1 a_27_47.t5 221.72
R143 a_27_47.n2 a_27_47.t6 221.72
R144 a_27_47.n4 a_27_47.t7 221.72
R145 a_27_47.n6 a_27_47.t9 221.72
R146 a_27_47.n7 a_27_47.n6 194.845
R147 a_27_47.n3 a_27_47.n0 178.881
R148 a_27_47.n8 a_27_47.t1 169.179
R149 a_27_47.n5 a_27_47.n0 152
R150 a_27_47.n1 a_27_47.t4 149.421
R151 a_27_47.n2 a_27_47.t3 149.421
R152 a_27_47.n4 a_27_47.t8 149.421
R153 a_27_47.n6 a_27_47.t2 149.421
R154 a_27_47.n2 a_27_47.n1 74.9783
R155 a_27_47.n3 a_27_47.n2 37.4894
R156 a_27_47.n4 a_27_47.n3 37.4894
R157 a_27_47.n5 a_27_47.n4 37.4894
R158 a_27_47.n6 a_27_47.n5 37.4894
R159 a_27_47.n8 a_27_47.n7 30.4005
R160 a_27_47.n7 a_27_47.n0 28.8005
R161 A_N.n0 A_N.t0 234.573
R162 A_N.n0 A_N.t1 162.274
R163 A_N A_N.n0 160
C0 VPB A_N 0.042542f
C1 B VPWR 0.092841f
C2 B Y 0.187688f
C3 B VGND 0.056199f
C4 VPWR Y 0.75829f
C5 VPWR VGND 0.104185f
C6 VPB B 0.139195f
C7 Y VGND 0.026845f
C8 VPB VPWR 0.124282f
C9 VPB Y 0.018025f
C10 A_N VPWR 0.017658f
C11 VPB VGND 0.009599f
C12 A_N VGND 0.014953f
C13 VGND VNB 0.5839f
C14 Y VNB 0.018254f
C15 VPWR VNB 0.516766f
C16 B VNB 0.423282f
C17 A_N VNB 0.147431f
C18 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR.t2 B.t0 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t2 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47.t1 B.t1 a_109_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t1 A.t1 a_193_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y.t0 C.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47.t0 C.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t0 241.536
R1 B.n0 B.t1 169.237
R2 B B.n0 154.744
R3 Y.n1 Y.t2 274.793
R4 Y.n1 Y.n0 205.28
R5 Y Y.t1 169.452
R6 Y Y.n1 67.4857
R7 Y.n0 Y.t3 26.5955
R8 Y.n0 Y.t0 26.5955
R9 VPWR.n1 VPWR.n0 324.12
R10 VPWR.n1 VPWR.t0 256.774
R11 VPWR.n0 VPWR.t1 38.4155
R12 VPWR.n0 VPWR.t2 26.5955
R13 VPWR VPWR.n1 0.418937
R14 VPB.t2 VPB.t1 284.113
R15 VPB.t0 VPB.t2 248.599
R16 VPB VPB.t0 189.409
R17 A.n0 A.t0 232.214
R18 A.n0 A.t1 159.915
R19 A A.n0 154.272
R20 a_109_47.t0 a_109_47.t1 49.8467
R21 a_193_47.t0 a_193_47.t1 60.9236
R22 VNB.t2 VNB.t1 1366.99
R23 VNB.t0 VNB.t2 1196.12
R24 VNB VNB.t0 911.327
R25 C.n0 C.t0 230.363
R26 C.n0 C.t1 158.064
R27 C C.n0 154.097
R28 VGND VGND.t0 282.123
C0 VPB Y 0.016577f
C1 C VPWR 0.041384f
C2 B A 0.082275f
C3 VPB VGND 0.005189f
C4 B VPWR 0.016994f
C5 C Y 0.072383f
C6 A VPWR 0.018588f
C7 B Y 0.149015f
C8 C VGND 0.041475f
C9 A Y 0.090927f
C10 B VGND 0.011586f
C11 VPWR Y 0.316891f
C12 A VGND 0.010023f
C13 VPWR VGND 0.041611f
C14 Y VGND 0.180582f
C15 VPB C 0.037322f
C16 VPB B 0.026782f
C17 VPB A 0.036833f
C18 C B 0.050963f
C19 VPB VPWR 0.050636f
C20 VGND VNB 0.263199f
C21 Y VNB 0.081638f
C22 VPWR VNB 0.246778f
C23 A VNB 0.142578f
C24 B VNB 0.097586f
C25 C VNB 0.157001f
C26 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_2 VNB VPB VGND VPWR C A Y B
X0 VGND.t1 C.t0 a_277_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR.t1 B.t0 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47.t2 C.t1 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y.t0 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t3 A.t0 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47.t3 A.t1 Y.t5 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47.t1 B.t2 a_277_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t5 C.t2 Y.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t7 C.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47.t1 B.t3 a_27_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t2 A.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y.t4 A.t3 a_27_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C.n1 C.t2 237.934
R1 C.n2 C.t3 218.507
R2 C.n1 C.t0 166.51
R3 C.n1 C.n0 152
R4 C.n4 C.n3 152
R5 C.n2 C.t1 146.208
R6 C.n3 C.n1 42.3833
R7 C C.n4 18.5605
R8 C.n0 C 16.0005
R9 C.n3 C.n2 14.9591
R10 C.n0 C 13.1205
R11 C.n4 C 10.8805
R12 a_277_47.n1 a_277_47.n0 434.474
R13 a_277_47.n0 a_277_47.t3 24.9236
R14 a_277_47.n0 a_277_47.t2 24.9236
R15 a_277_47.t0 a_277_47.n1 24.9236
R16 a_277_47.n1 a_277_47.t1 24.9236
R17 VGND.n0 VGND.t0 288.012
R18 VGND.n0 VGND.t1 145.041
R19 VGND VGND.n0 1.00936
R20 VNB.t2 VNB.t4 2677.02
R21 VNB.t4 VNB.t5 1196.12
R22 VNB.t3 VNB.t2 1196.12
R23 VNB.t1 VNB.t3 1196.12
R24 VNB.t0 VNB.t1 1196.12
R25 VNB VNB.t0 911.327
R26 B.n3 B.t0 218.507
R27 B.n0 B.t1 218.507
R28 B.n4 B.n3 166.959
R29 B.n2 B.n1 152
R30 B.n3 B.t2 146.208
R31 B.n0 B.t3 146.208
R32 B.n3 B.n2 64.8212
R33 B.n4 B 18.5605
R34 B.n1 B 17.2805
R35 B.n1 B 12.1605
R36 B B.n4 10.8805
R37 B.n2 B.n0 4.98671
R38 Y.n2 Y.n0 266.178
R39 Y.n4 Y.n3 206.25
R40 Y.n2 Y.n1 206.25
R41 Y Y.n5 186.745
R42 Y.n4 Y.n2 29.6732
R43 Y.n3 Y.t3 26.5955
R44 Y.n3 Y.t2 26.5955
R45 Y.n0 Y.t6 26.5955
R46 Y.n0 Y.t7 26.5955
R47 Y.n1 Y.t1 26.5955
R48 Y.n1 Y.t0 26.5955
R49 Y.n5 Y.t5 24.9236
R50 Y.n5 Y.t4 24.9236
R51 Y Y.n4 4.26717
R52 VPWR.n9 VPWR.n1 320.976
R53 VPWR.n3 VPWR.t4 319.096
R54 VPWR.n3 VPWR.t1 319.096
R55 VPWR.n5 VPWR.t5 253.244
R56 VPWR.n11 VPWR.t2 249.901
R57 VPWR.n8 VPWR.n2 34.6358
R58 VPWR.n10 VPWR.n9 30.8711
R59 VPWR.n1 VPWR.t0 26.5955
R60 VPWR.n1 VPWR.t3 26.5955
R61 VPWR.n11 VPWR.n10 25.977
R62 VPWR.n4 VPWR.n2 18.4476
R63 VPWR.n6 VPWR.n2 9.3005
R64 VPWR.n8 VPWR.n7 9.3005
R65 VPWR.n10 VPWR.n0 9.3005
R66 VPWR.n12 VPWR.n11 9.3005
R67 VPWR.n4 VPWR.n3 8.61052
R68 VPWR.n5 VPWR.n4 3.87951
R69 VPWR.n9 VPWR.n8 3.76521
R70 VPWR.n6 VPWR.n5 0.450477
R71 VPWR.n7 VPWR.n6 0.120292
R72 VPWR.n7 VPWR.n0 0.120292
R73 VPWR.n12 VPWR.n0 0.120292
R74 VPWR VPWR.n12 0.0213333
R75 VPB.t1 VPB.t4 556.386
R76 VPB.t4 VPB.t5 248.599
R77 VPB.t0 VPB.t1 248.599
R78 VPB.t3 VPB.t0 248.599
R79 VPB.t2 VPB.t3 248.599
R80 VPB VPB.t2 189.409
R81 A.n0 A.t0 212.081
R82 A.n1 A.t2 212.081
R83 A A.n1 188.548
R84 A.n0 A.t1 139.78
R85 A.n1 A.t3 139.78
R86 A.n1 A.n0 61.346
R87 a_27_47.t1 a_27_47.n1 331.325
R88 a_27_47.n1 a_27_47.t2 273.296
R89 a_27_47.n1 a_27_47.n0 185
R90 a_27_47.n0 a_27_47.t0 24.9236
R91 a_27_47.n0 a_27_47.t3 24.9236
C0 C VPWR 0.076304f
C1 B Y 0.151516f
C2 A VGND 0.019146f
C3 C Y 0.081859f
C4 B VGND 0.021269f
C5 C VGND 0.075502f
C6 VPWR Y 0.627912f
C7 VPWR VGND 0.077629f
C8 Y VGND 0.016488f
C9 VPB A 0.068652f
C10 VPB B 0.069242f
C11 A B 0.057811f
C12 VPB C 0.071885f
C13 VPB VPWR 0.10162f
C14 B C 0.031389f
C15 VPB Y 0.020026f
C16 A VPWR 0.05789f
C17 VPB VGND 0.00687f
C18 B VPWR 0.033809f
C19 A Y 0.095774f
C20 VGND VNB 0.46594f
C21 Y VNB 0.024821f
C22 VPWR VNB 0.435692f
C23 C VNB 0.236469f
C24 B VNB 0.204852f
C25 A VNB 0.236265f
C26 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_4 VNB VPB VGND VPWR C A Y B
X0 a_27_47.t7 B.t0 a_445_47.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47.t6 B.t1 a_445_47.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t12 B.t2 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t0 C.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t3 A.t0 a_445_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t1 C.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t4 A.t1 a_445_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR.t6 C.t2 Y.t8 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47.t0 C.t3 VGND.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47.t1 C.t4 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_445_47.t6 A.t2 Y.t13 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t9 B.t3 Y.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47.t7 A.t3 Y.t14 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t1 C.t5 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_445_47.t3 B.t4 a_27_47.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y.t10 B.t5 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR.t11 A.t4 Y.t15 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X17 a_445_47.t2 B.t6 a_27_47.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t7 B.t7 Y.t9 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y.t5 A.t5 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t4 A.t6 Y.t6 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 Y.t2 C.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 Y.t7 A.t7 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VGND.t0 C.t7 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n1 B.t3 221.72
R1 B.n0 B.t5 221.72
R2 B.n6 B.t7 221.72
R3 B.n7 B.t2 221.72
R4 B.n3 B.n2 152
R5 B.n5 B.n4 152
R6 B.n9 B.n8 152
R7 B.n1 B.t1 149.421
R8 B.n0 B.t6 149.421
R9 B.n6 B.t0 149.421
R10 B.n7 B.t4 149.421
R11 B.n2 B.n1 37.4894
R12 B.n2 B.n0 37.4894
R13 B.n5 B.n0 37.4894
R14 B.n6 B.n5 37.4894
R15 B.n8 B.n6 37.4894
R16 B.n8 B.n7 37.4894
R17 B B.n9 23.6805
R18 B.n4 B 21.1205
R19 B B.n3 18.5605
R20 B.n3 B 10.8805
R21 B.n4 B 8.3205
R22 B.n9 B 5.7605
R23 a_445_47.n4 a_445_47.t6 302.86
R24 a_445_47.n3 a_445_47.t1 258.846
R25 a_445_47.n2 a_445_47.n0 231.749
R26 a_445_47.n2 a_445_47.n1 185
R27 a_445_47.n5 a_445_47.n4 185
R28 a_445_47.n3 a_445_47.n2 52.3135
R29 a_445_47.n4 a_445_47.n3 46.7483
R30 a_445_47.n0 a_445_47.t5 24.9236
R31 a_445_47.n0 a_445_47.t3 24.9236
R32 a_445_47.n1 a_445_47.t4 24.9236
R33 a_445_47.n1 a_445_47.t2 24.9236
R34 a_445_47.t0 a_445_47.n5 24.9236
R35 a_445_47.n5 a_445_47.t7 24.9236
R36 a_27_47.t6 a_27_47.n5 323.373
R37 a_27_47.n3 a_27_47.n2 185
R38 a_27_47.n5 a_27_47.n4 185
R39 a_27_47.n1 a_27_47.t3 176.43
R40 a_27_47.n1 a_27_47.n0 98.788
R41 a_27_47.n5 a_27_47.n3 55.2965
R42 a_27_47.n3 a_27_47.n1 46.8485
R43 a_27_47.n4 a_27_47.t4 24.9236
R44 a_27_47.n4 a_27_47.t7 24.9236
R45 a_27_47.n2 a_27_47.t5 24.9236
R46 a_27_47.n2 a_27_47.t1 24.9236
R47 a_27_47.n0 a_27_47.t2 24.9236
R48 a_27_47.n0 a_27_47.t0 24.9236
R49 VNB.t8 VNB.t5 2677.02
R50 VNB.t4 VNB.t10 1196.12
R51 VNB.t11 VNB.t4 1196.12
R52 VNB.t5 VNB.t11 1196.12
R53 VNB.t6 VNB.t8 1196.12
R54 VNB.t9 VNB.t6 1196.12
R55 VNB.t7 VNB.t9 1196.12
R56 VNB.t1 VNB.t7 1196.12
R57 VNB.t2 VNB.t1 1196.12
R58 VNB.t0 VNB.t2 1196.12
R59 VNB.t3 VNB.t0 1196.12
R60 VNB VNB.t3 911.327
R61 VPWR.n10 VPWR.t11 346.161
R62 VPWR.n28 VPWR.n1 320.976
R63 VPWR.n22 VPWR.n21 320.976
R64 VPWR.n19 VPWR.n4 320.976
R65 VPWR.n9 VPWR.n8 320.976
R66 VPWR.n7 VPWR.t5 319.096
R67 VPWR.n7 VPWR.t9 319.096
R68 VPWR.n30 VPWR.t2 249.901
R69 VPWR.n18 VPWR.n5 34.6358
R70 VPWR.n23 VPWR.n20 34.6358
R71 VPWR.n27 VPWR.n2 34.6358
R72 VPWR.n13 VPWR.n12 34.6358
R73 VPWR.n29 VPWR.n28 30.8711
R74 VPWR.n10 VPWR.n9 29.6092
R75 VPWR.n1 VPWR.t1 26.5955
R76 VPWR.n1 VPWR.t6 26.5955
R77 VPWR.n21 VPWR.t10 26.5955
R78 VPWR.n21 VPWR.t0 26.5955
R79 VPWR.n4 VPWR.t8 26.5955
R80 VPWR.n4 VPWR.t7 26.5955
R81 VPWR.n8 VPWR.t3 26.5955
R82 VPWR.n8 VPWR.t4 26.5955
R83 VPWR.n30 VPWR.n29 25.977
R84 VPWR.n22 VPWR.n2 24.8476
R85 VPWR.n20 VPWR.n19 18.824
R86 VPWR.n19 VPWR.n18 15.8123
R87 VPWR.n12 VPWR.n9 11.2946
R88 VPWR.n14 VPWR.n13 10.9181
R89 VPWR.n23 VPWR.n22 9.78874
R90 VPWR.n12 VPWR.n11 9.3005
R91 VPWR.n13 VPWR.n6 9.3005
R92 VPWR.n15 VPWR.n14 9.3005
R93 VPWR.n16 VPWR.n5 9.3005
R94 VPWR.n18 VPWR.n17 9.3005
R95 VPWR.n20 VPWR.n3 9.3005
R96 VPWR.n24 VPWR.n23 9.3005
R97 VPWR.n25 VPWR.n2 9.3005
R98 VPWR.n27 VPWR.n26 9.3005
R99 VPWR.n29 VPWR.n0 9.3005
R100 VPWR.n31 VPWR.n30 9.3005
R101 VPWR.n14 VPWR.n7 8.61052
R102 VPWR.n14 VPWR.n5 6.4005
R103 VPWR.n28 VPWR.n27 3.76521
R104 VPWR.n11 VPWR.n10 1.41422
R105 VPWR.n11 VPWR.n6 0.120292
R106 VPWR.n15 VPWR.n6 0.120292
R107 VPWR.n16 VPWR.n15 0.120292
R108 VPWR.n17 VPWR.n16 0.120292
R109 VPWR.n17 VPWR.n3 0.120292
R110 VPWR.n24 VPWR.n3 0.120292
R111 VPWR.n25 VPWR.n24 0.120292
R112 VPWR.n26 VPWR.n25 0.120292
R113 VPWR.n26 VPWR.n0 0.120292
R114 VPWR.n31 VPWR.n0 0.120292
R115 VPWR VPWR.n31 0.0213333
R116 Y.n5 Y.n3 235.923
R117 Y.n2 Y.n0 228.008
R118 Y.n5 Y.n4 206.25
R119 Y.n7 Y.n6 206.25
R120 Y.n9 Y.n8 206.25
R121 Y.n11 Y.n10 206.25
R122 Y.n13 Y.n12 206.25
R123 Y.n2 Y.n1 185
R124 Y.n11 Y.n9 59.9278
R125 Y Y.n13 38.7041
R126 Y Y.n2 37.1205
R127 Y.n7 Y.n5 29.6732
R128 Y.n9 Y.n7 29.6732
R129 Y.n13 Y.n11 29.6732
R130 Y.n3 Y.t8 26.5955
R131 Y.n3 Y.t2 26.5955
R132 Y.n4 Y.t0 26.5955
R133 Y.n4 Y.t1 26.5955
R134 Y.n6 Y.t9 26.5955
R135 Y.n6 Y.t12 26.5955
R136 Y.n8 Y.t11 26.5955
R137 Y.n8 Y.t10 26.5955
R138 Y.n10 Y.t6 26.5955
R139 Y.n10 Y.t7 26.5955
R140 Y.n12 Y.t15 26.5955
R141 Y.n12 Y.t5 26.5955
R142 Y.n0 Y.t14 24.9236
R143 Y.n0 Y.t4 24.9236
R144 Y.n1 Y.t13 24.9236
R145 Y.n1 Y.t3 24.9236
R146 Y.n14 Y 11.1309
R147 Y Y.n14 7.7918
R148 Y.n14 Y 5.8885
R149 VPB.t9 VPB.t5 556.386
R150 VPB.t3 VPB.t11 248.599
R151 VPB.t4 VPB.t3 248.599
R152 VPB.t5 VPB.t4 248.599
R153 VPB.t8 VPB.t9 248.599
R154 VPB.t7 VPB.t8 248.599
R155 VPB.t10 VPB.t7 248.599
R156 VPB.t0 VPB.t10 248.599
R157 VPB.t1 VPB.t0 248.599
R158 VPB.t6 VPB.t1 248.599
R159 VPB.t2 VPB.t6 248.599
R160 VPB VPB.t2 189.409
R161 C.n9 C.t6 234.573
R162 C.n2 C.t0 221.72
R163 C.n4 C.t1 221.72
R164 C.n0 C.t2 221.72
R165 C.n9 C.t7 162.274
R166 C.n3 C.n1 152
R167 C.n6 C.n5 152
R168 C.n8 C.n7 152
R169 C.n10 C.n9 152
R170 C.n2 C.t4 149.421
R171 C.n4 C.t5 149.421
R172 C.n0 C.t3 149.421
R173 C.n3 C.n2 37.4894
R174 C.n4 C.n3 37.4894
R175 C.n5 C.n4 37.4894
R176 C.n5 C.n0 37.4894
R177 C.n8 C.n0 37.4894
R178 C.n6 C.n1 26.8805
R179 C.n7 C 24.9605
R180 C.n9 C.n8 24.1005
R181 C.n10 C 21.4405
R182 C C.n10 8.0005
R183 C.n7 C 4.4805
R184 C C.n6 1.9205
R185 C.n1 C 0.6405
R186 A.n1 A.t4 221.72
R187 A.n3 A.t5 221.72
R188 A.n0 A.t6 221.72
R189 A.n8 A.t7 221.72
R190 A.n9 A.n8 194.845
R191 A.n2 A 162.881
R192 A.n5 A.n4 152
R193 A.n7 A.n6 152
R194 A.n1 A.t2 149.421
R195 A.n3 A.t0 149.421
R196 A.n0 A.t3 149.421
R197 A.n8 A.t1 149.421
R198 A.n7 A.n0 38.382
R199 A.n2 A.n1 37.4894
R200 A.n3 A.n2 37.4894
R201 A.n4 A.n3 37.4894
R202 A.n4 A.n0 37.4894
R203 A.n8 A.n7 36.5968
R204 A A.n9 16.6405
R205 A.n5 A 16.0005
R206 A.n6 A 15.6805
R207 A.n6 A 13.7605
R208 A A.n5 13.4405
R209 A.n9 A 12.8005
R210 VGND.n2 VGND.n1 218.738
R211 VGND.n2 VGND.n0 215.31
R212 VGND.n1 VGND.t2 24.9236
R213 VGND.n1 VGND.t1 24.9236
R214 VGND.n0 VGND.t3 24.9236
R215 VGND.n0 VGND.t0 24.9236
R216 VGND VGND.n2 0.53334
C0 A Y 0.372238f
C1 B VGND 0.033261f
C2 A VGND 0.033556f
C3 VPWR Y 1.1919f
C4 VPWR VGND 0.128935f
C5 VPB C 0.13304f
C6 Y VGND 0.054374f
C7 VPB B 0.121158f
C8 VPB A 0.143027f
C9 VPB VPWR 0.155326f
C10 C B 0.064343f
C11 VPB Y 0.045077f
C12 VPB VGND 0.011581f
C13 C VPWR 0.094929f
C14 B A 0.033231f
C15 C Y 0.176232f
C16 B VPWR 0.050458f
C17 A VPWR 0.059042f
C18 B Y 0.212024f
C19 C VGND 0.060637f
C20 VGND VNB 0.712848f
C21 Y VNB 0.077614f
C22 VPWR VNB 0.661943f
C23 A VNB 0.423631f
C24 B VNB 0.363154f
C25 C VNB 0.416992f
C26 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_1 VPB VNB VGND VPWR Y B C A_N
X0 Y.t2 a_53_93.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47.t1 C.t0 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR.t2 B.t0 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t0 A_N.t0 a_53_93.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND.t0 A_N.t1 a_53_93.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_316_47.t1 B.t1 a_232_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t3 a_53_93.t3 a_316_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X7 Y.t0 C.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
R0 a_53_93.n1 a_53_93.t1 722.242
R1 a_53_93.n1 a_53_93.n0 303.243
R2 a_53_93.n0 a_53_93.t2 236.18
R3 a_53_93.t0 a_53_93.n1 223.571
R4 a_53_93.n0 a_53_93.t3 163.881
R5 VPWR.n2 VPWR.n1 319.389
R6 VPWR.n2 VPWR.n0 230.242
R7 VPWR.n0 VPWR.t0 95.3969
R8 VPWR.n1 VPWR.t2 38.4155
R9 VPWR.n1 VPWR.t3 37.4305
R10 VPWR.n0 VPWR.t1 26.3637
R11 VPWR VPWR.n2 0.493918
R12 Y.n4 Y.n3 585
R13 Y.n5 Y.n4 292.933
R14 Y Y.t3 272.084
R15 Y.n2 Y.n0 252.339
R16 Y.n4 Y.t2 26.5955
R17 Y.n0 Y.t1 26.5955
R18 Y.n0 Y.t0 26.5955
R19 Y.n5 Y 5.95827
R20 Y.n3 Y 2.82084
R21 Y.n1 Y 2.2074
R22 Y.n2 Y.n1 1.84457
R23 Y.n3 Y.n2 1.62762
R24 Y Y.n5 1.41325
R25 Y.n1 Y 1.08525
R26 VPB.t2 VPB.t3 316.668
R27 VPB.t0 VPB.t1 287.072
R28 VPB VPB.t0 269.315
R29 VPB.t1 VPB.t2 248.599
R30 C.n0 C.t1 236.18
R31 C.n0 C.t0 163.881
R32 C C.n0 154.607
R33 VGND VGND.n0 208.304
R34 VGND.n0 VGND.t0 58.5719
R35 VGND.n0 VGND.t1 24.0005
R36 a_232_47.t0 a_232_47.t1 49.8467
R37 VNB.t1 VNB.t2 1523.62
R38 VNB.t0 VNB.t3 1381.23
R39 VNB VNB.t0 1295.79
R40 VNB.t3 VNB.t1 1196.12
R41 B.n0 B.t0 236.18
R42 B.n0 B.t1 163.881
R43 B B.n0 154.522
R44 A_N A_N.n0 155.685
R45 A_N.n0 A_N.t0 142.994
R46 A_N.n0 A_N.t1 126.927
R47 a_316_47.t0 a_316_47.t1 71.0774
C0 VPWR A_N 0.02091f
C1 Y VGND 0.084616f
C2 Y VPB 0.027316f
C3 Y C 0.020663f
C4 VGND VPB 0.007843f
C5 Y B 0.046906f
C6 VGND C 0.014636f
C7 VPB C 0.031831f
C8 Y VPWR 0.357261f
C9 VGND B 0.012548f
C10 VPB B 0.029981f
C11 Y A_N 0.001234f
C12 VGND VPWR 0.055361f
C13 VPB VPWR 0.077773f
C14 C B 0.082225f
C15 VGND A_N 0.010189f
C16 VPB A_N 0.04217f
C17 C VPWR 0.02217f
C18 C A_N 0.065966f
C19 B VPWR 0.017594f
C20 VGND VNB 0.355372f
C21 Y VNB 0.10206f
C22 A_N VNB 0.125463f
C23 VPWR VNB 0.306818f
C24 B VNB 0.095312f
C25 C VNB 0.100588f
C26 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_2 VNB VPB VGND VPWR A_N C B Y
X0 a_408_47.t1 B.t0 a_218_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_408_47.t3 a_27_47.t2 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t2 a_27_47.t3 a_408_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t6 A_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND.t1 C.t0 a_218_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t3 B.t1 Y.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47.t3 C.t1 VGND.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11975 ps=1.045 w=0.65 l=0.15
X7 Y.t4 B.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t5 C.t2 Y.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR.t1 a_27_47.t4 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47.t1 B.t3 a_408_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y.t6 C.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17575 ps=1.395 w=1 l=0.15
X12 Y.t0 a_27_47.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND.t2 A_N.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 B.n3 B.t2 268.135
R1 B.n2 B.t1 221.72
R2 B.n0 B.t0 206.547
R3 B.n4 B.n0 175.041
R4 B.n4 B.n3 152
R5 B.n1 B.t3 149.421
R6 B.n3 B.n2 28.5635
R7 B.n1 B.n0 17.8524
R8 B.n2 B.n1 17.8524
R9 B B.n4 2.5605
R10 a_218_47.n1 a_218_47.n0 353.003
R11 a_218_47.n0 a_218_47.t2 24.9236
R12 a_218_47.n0 a_218_47.t1 24.9236
R13 a_218_47.t0 a_218_47.n1 24.9236
R14 a_218_47.n1 a_218_47.t3 24.9236
R15 a_408_47.n0 a_408_47.t0 319.277
R16 a_408_47.n0 a_408_47.t3 319.277
R17 a_408_47.n1 a_408_47.n0 97.0637
R18 a_408_47.n1 a_408_47.t2 24.9236
R19 a_408_47.t1 a_408_47.n1 24.9236
R20 VNB.t0 VNB.t1 2677.02
R21 VNB.t6 VNB.t5 1552.1
R22 VNB.t3 VNB.t4 1196.12
R23 VNB.t2 VNB.t3 1196.12
R24 VNB.t1 VNB.t2 1196.12
R25 VNB.t5 VNB.t0 1196.12
R26 VNB VNB.t6 911.327
R27 a_27_47.t0 a_27_47.n3 691.605
R28 a_27_47.n3 a_27_47.n2 403.151
R29 a_27_47.n3 a_27_47.t1 292.454
R30 a_27_47.n0 a_27_47.t4 221.72
R31 a_27_47.n1 a_27_47.t5 221.72
R32 a_27_47.n0 a_27_47.t2 149.421
R33 a_27_47.n1 a_27_47.t3 149.421
R34 a_27_47.n2 a_27_47.n1 48.2005
R35 a_27_47.n2 a_27_47.n0 26.7783
R36 Y.n3 Y.n1 329.507
R37 Y.n4 Y.n0 300.116
R38 Y.n3 Y.n2 299.834
R39 Y Y.n5 222.69
R40 Y.n4 Y.n3 79.8031
R41 Y Y.n4 47.3605
R42 Y.n0 Y.t1 26.5955
R43 Y.n0 Y.t0 26.5955
R44 Y.n2 Y.t5 26.5955
R45 Y.n2 Y.t4 26.5955
R46 Y.n1 Y.t7 26.5955
R47 Y.n1 Y.t6 26.5955
R48 Y.n5 Y.t3 24.9236
R49 Y.n5 Y.t2 24.9236
R50 A_N.n0 A_N.t0 329.007
R51 A_N.n0 A_N.t1 200.475
R52 A_N A_N.n0 154.012
R53 VPWR.n5 VPWR.t1 877.606
R54 VPWR.n7 VPWR.t3 873.438
R55 VPWR.n6 VPWR.t0 873.438
R56 VPWR.n3 VPWR.n2 607.212
R57 VPWR.n13 VPWR.n1 310.486
R58 VPWR.n1 VPWR.t6 101.733
R59 VPWR.n1 VPWR.t4 39.7937
R60 VPWR.n12 VPWR.n11 34.6358
R61 VPWR.n8 VPWR.n3 32.0005
R62 VPWR.n2 VPWR.t2 26.5955
R63 VPWR.n2 VPWR.t5 26.5955
R64 VPWR.n8 VPWR.n7 24.8476
R65 VPWR.n13 VPWR.n12 19.577
R66 VPWR.n7 VPWR.n6 14.3064
R67 VPWR.n7 VPWR.n4 9.3005
R68 VPWR.n9 VPWR.n8 9.3005
R69 VPWR.n11 VPWR.n10 9.3005
R70 VPWR.n12 VPWR.n0 9.3005
R71 VPWR.n14 VPWR.n13 7.35738
R72 VPWR.n6 VPWR.n5 6.85691
R73 VPWR.n11 VPWR.n3 2.63579
R74 VPWR.n5 VPWR.n4 0.588885
R75 VPWR.n14 VPWR.n0 0.145509
R76 VPWR.n9 VPWR.n4 0.120292
R77 VPWR.n10 VPWR.n9 0.120292
R78 VPWR.n10 VPWR.n0 0.120292
R79 VPWR VPWR.n14 0.11659
R80 VPB.t3 VPB.t0 556.386
R81 VPB.t6 VPB.t4 322.587
R82 VPB.t0 VPB.t1 248.599
R83 VPB.t2 VPB.t3 248.599
R84 VPB.t5 VPB.t2 248.599
R85 VPB.t4 VPB.t5 248.599
R86 VPB VPB.t6 189.409
R87 C.n0 C.t2 221.72
R88 C.n1 C.t3 221.72
R89 C C.n2 161.921
R90 C.n0 C.t0 149.421
R91 C.n1 C.t1 149.421
R92 C.n2 C.n0 37.4894
R93 C.n2 C.n1 37.4894
R94 VGND.n1 VGND.t1 293.288
R95 VGND.n1 VGND.n0 118.659
R96 VGND.n0 VGND.t2 61.6309
R97 VGND.n0 VGND.t0 34.8099
R98 VGND VGND.n1 0.444038
C0 VPB A_N 0.091314f
C1 VPB C 0.053576f
C2 A_N C 0.060294f
C3 VPB B 0.082027f
C4 VPB VPWR 0.096085f
C5 VPB Y 0.020121f
C6 A_N VPWR 0.023045f
C7 C B 0.058257f
C8 C VPWR 0.03203f
C9 A_N Y 0.003022f
C10 VPB VGND 0.008769f
C11 A_N VGND 0.045949f
C12 C Y 0.023214f
C13 B VPWR 0.030525f
C14 B Y 0.031005f
C15 C VGND 0.034844f
C16 VPWR Y 0.457314f
C17 B VGND 0.022341f
C18 VPWR VGND 0.083448f
C19 Y VGND 0.017637f
C20 VGND VNB 0.48281f
C21 Y VNB 0.068514f
C22 VPWR VNB 0.409991f
C23 B VNB 0.226562f
C24 C VNB 0.176474f
C25 A_N VNB 0.17071f
C26 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_4 VNB VPB VGND VPWR B C A_N Y
X0 VGND.t3 C.t0 a_633_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y.t11 B.t0 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t0 a_27_47.t2 a_215_47.t7 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y.t1 a_27_47.t3 a_215_47.t6 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_633_47.t4 B.t1 a_215_47.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t6 B.t2 Y.t10 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t15 C.t1 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_633_47.t5 B.t3 a_215_47.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t10 C.t2 Y.t14 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_215_47.t5 a_27_47.t4 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t13 C.t3 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_215_47.t1 B.t4 a_633_47.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_215_47.t0 B.t5 a_633_47.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t9 B.t6 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t0 a_27_47.t5 Y.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y.t4 a_27_47.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_633_47.t2 C.t4 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_633_47.t1 C.t5 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t2 a_27_47.t7 Y.t5 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t8 C.t6 Y.t12 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X20 a_215_47.t4 a_27_47.t8 Y.t6 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t7 a_27_47.t9 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 VPWR.t12 A_N.t0 a_27_47.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X23 VGND.t0 C.t7 a_633_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VPWR.t4 B.t7 Y.t8 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND.t4 A_N.t1 a_27_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C.n0 C.t6 221.72
R1 C.n2 C.t1 221.72
R2 C.n7 C.t2 221.72
R3 C.n3 C.t3 221.72
R4 C.n4 C.n3 194.845
R5 C C.n1 162.56
R6 C.n9 C.n8 152
R7 C.n6 C.n5 152
R8 C.n0 C.t0 149.421
R9 C.n2 C.t5 149.421
R10 C.n7 C.t7 149.421
R11 C.n3 C.t4 149.421
R12 C.n1 C.n0 38.382
R13 C.n8 C.n2 37.4894
R14 C.n8 C.n7 37.4894
R15 C.n7 C.n6 37.4894
R16 C.n6 C.n3 37.4894
R17 C.n2 C.n1 36.5968
R18 C.n4 C 16.6405
R19 C C.n9 16.0005
R20 C.n5 C 16.0005
R21 C.n9 C 13.4405
R22 C.n5 C 13.4405
R23 C C.n4 12.8005
R24 a_633_47.n2 a_633_47.n0 224.822
R25 a_633_47.n2 a_633_47.n1 185
R26 a_633_47.n4 a_633_47.n3 133.534
R27 a_633_47.n5 a_633_47.n4 99.1759
R28 a_633_47.n4 a_633_47.n2 68.8286
R29 a_633_47.n3 a_633_47.t3 24.9236
R30 a_633_47.n3 a_633_47.t1 24.9236
R31 a_633_47.n0 a_633_47.t6 24.9236
R32 a_633_47.n0 a_633_47.t4 24.9236
R33 a_633_47.n1 a_633_47.t7 24.9236
R34 a_633_47.n1 a_633_47.t5 24.9236
R35 a_633_47.t0 a_633_47.n5 24.9236
R36 a_633_47.n5 a_633_47.t2 24.9236
R37 VGND.n12 VGND.t2 287.534
R38 VGND.n26 VGND.t4 287.534
R39 VGND.n7 VGND.n6 207.213
R40 VGND.n8 VGND.t3 154.691
R41 VGND.n11 VGND.n5 34.6358
R42 VGND.n14 VGND.n13 34.6358
R43 VGND.n14 VGND.n3 34.6358
R44 VGND.n18 VGND.n3 34.6358
R45 VGND.n19 VGND.n18 34.6358
R46 VGND.n20 VGND.n19 34.6358
R47 VGND.n20 VGND.n1 34.6358
R48 VGND.n24 VGND.n1 34.6358
R49 VGND.n25 VGND.n24 34.6358
R50 VGND.n8 VGND.n7 28.26
R51 VGND.n6 VGND.t1 24.9236
R52 VGND.n6 VGND.t0 24.9236
R53 VGND.n26 VGND.n25 22.9652
R54 VGND.n7 VGND.n5 12.8005
R55 VGND.n12 VGND.n11 9.41227
R56 VGND.n25 VGND.n0 9.3005
R57 VGND.n24 VGND.n23 9.3005
R58 VGND.n22 VGND.n1 9.3005
R59 VGND.n21 VGND.n20 9.3005
R60 VGND.n19 VGND.n2 9.3005
R61 VGND.n18 VGND.n17 9.3005
R62 VGND.n16 VGND.n3 9.3005
R63 VGND.n15 VGND.n14 9.3005
R64 VGND.n13 VGND.n4 9.3005
R65 VGND.n11 VGND.n10 9.3005
R66 VGND.n9 VGND.n5 9.3005
R67 VGND.n27 VGND.n26 7.4049
R68 VGND.n13 VGND.n12 6.4005
R69 VGND.n9 VGND.n8 1.27836
R70 VGND.n27 VGND.n0 0.144904
R71 VGND.n10 VGND.n9 0.120292
R72 VGND.n10 VGND.n4 0.120292
R73 VGND.n15 VGND.n4 0.120292
R74 VGND.n16 VGND.n15 0.120292
R75 VGND.n17 VGND.n16 0.120292
R76 VGND.n17 VGND.n2 0.120292
R77 VGND.n21 VGND.n2 0.120292
R78 VGND.n22 VGND.n21 0.120292
R79 VGND.n23 VGND.n22 0.120292
R80 VGND.n23 VGND.n0 0.120292
R81 VGND VGND.n27 0.117202
R82 VNB.t12 VNB.t6 2677.02
R83 VNB.t10 VNB.t0 2677.02
R84 VNB.t5 VNB.t7 1196.12
R85 VNB.t4 VNB.t5 1196.12
R86 VNB.t6 VNB.t4 1196.12
R87 VNB.t9 VNB.t12 1196.12
R88 VNB.t11 VNB.t9 1196.12
R89 VNB.t8 VNB.t11 1196.12
R90 VNB.t2 VNB.t8 1196.12
R91 VNB.t1 VNB.t2 1196.12
R92 VNB.t3 VNB.t1 1196.12
R93 VNB.t0 VNB.t3 1196.12
R94 VNB VNB.t10 911.327
R95 B.n0 B.t7 221.72
R96 B.n3 B.t0 221.72
R97 B.n4 B.t2 221.72
R98 B.n5 B.t6 221.72
R99 B.n2 B.n1 152
R100 B.n7 B.n6 152
R101 B.n0 B.t5 149.421
R102 B.n3 B.t3 149.421
R103 B.n4 B.t4 149.421
R104 B.n5 B.t1 149.421
R105 B.n4 B.n3 74.9783
R106 B.n6 B.n5 61.5894
R107 B.n2 B.n0 41.9524
R108 B.n3 B.n2 33.0264
R109 B.n7 B 26.5605
R110 B.n1 B 16.9605
R111 B.n6 B.n4 13.3894
R112 B.n1 B 12.4805
R113 B B.n7 2.8805
R114 VPWR.n23 VPWR.n22 607.212
R115 VPWR.n29 VPWR.n2 320.976
R116 VPWR.n20 VPWR.n5 320.976
R117 VPWR.n10 VPWR.n9 320.976
R118 VPWR.n8 VPWR.t9 319.096
R119 VPWR.n8 VPWR.t4 319.096
R120 VPWR.n11 VPWR.t8 263.849
R121 VPWR.n1 VPWR.t12 221.597
R122 VPWR.n1 VPWR.t3 221.596
R123 VPWR.n19 VPWR.n6 34.6358
R124 VPWR.n24 VPWR.n21 34.6358
R125 VPWR.n28 VPWR.n3 34.6358
R126 VPWR.n14 VPWR.n13 34.6358
R127 VPWR.n30 VPWR.n29 32.377
R128 VPWR.n11 VPWR.n10 28.26
R129 VPWR.n2 VPWR.t1 26.5955
R130 VPWR.n2 VPWR.t2 26.5955
R131 VPWR.n22 VPWR.t5 26.5955
R132 VPWR.n22 VPWR.t0 26.5955
R133 VPWR.n5 VPWR.t7 26.5955
R134 VPWR.n5 VPWR.t6 26.5955
R135 VPWR.n9 VPWR.t11 26.5955
R136 VPWR.n9 VPWR.t10 26.5955
R137 VPWR.n23 VPWR.n3 26.3534
R138 VPWR.n31 VPWR.n30 24.4711
R139 VPWR.n21 VPWR.n20 20.3299
R140 VPWR.n20 VPWR.n19 14.3064
R141 VPWR.n13 VPWR.n10 12.8005
R142 VPWR.n31 VPWR.n1 10.4861
R143 VPWR.n15 VPWR.n14 9.41227
R144 VPWR.n13 VPWR.n12 9.3005
R145 VPWR.n14 VPWR.n7 9.3005
R146 VPWR.n16 VPWR.n15 9.3005
R147 VPWR.n17 VPWR.n6 9.3005
R148 VPWR.n19 VPWR.n18 9.3005
R149 VPWR.n21 VPWR.n4 9.3005
R150 VPWR.n25 VPWR.n24 9.3005
R151 VPWR.n26 VPWR.n3 9.3005
R152 VPWR.n28 VPWR.n27 9.3005
R153 VPWR.n30 VPWR.n0 9.3005
R154 VPWR.n15 VPWR.n8 8.61052
R155 VPWR.n24 VPWR.n23 8.28285
R156 VPWR.n15 VPWR.n6 7.90638
R157 VPWR.n32 VPWR.n31 4.0883
R158 VPWR.n29 VPWR.n28 2.25932
R159 VPWR.n12 VPWR.n11 1.27836
R160 VPWR.n32 VPWR.n0 0.200784
R161 VPWR VPWR.n32 0.18088
R162 VPWR.n12 VPWR.n7 0.120292
R163 VPWR.n16 VPWR.n7 0.120292
R164 VPWR.n17 VPWR.n16 0.120292
R165 VPWR.n18 VPWR.n17 0.120292
R166 VPWR.n18 VPWR.n4 0.120292
R167 VPWR.n25 VPWR.n4 0.120292
R168 VPWR.n26 VPWR.n25 0.120292
R169 VPWR.n27 VPWR.n26 0.120292
R170 VPWR.n27 VPWR.n0 0.120292
R171 Y.n9 Y.n8 239.695
R172 Y.n2 Y.n0 235.923
R173 Y.n13 Y.n11 224.822
R174 Y.n2 Y.n1 206.25
R175 Y.n4 Y.n3 206.25
R176 Y.n6 Y.n5 196.423
R177 Y.n9 Y.n7 196.423
R178 Y.n13 Y.n12 185
R179 Y.n4 Y.n2 59.9278
R180 Y Y.n13 33.9706
R181 Y.n6 Y.n4 33.4447
R182 Y.n7 Y.t3 26.5955
R183 Y.n7 Y.t4 26.5955
R184 Y.n5 Y.t10 26.5955
R185 Y.n5 Y.t9 26.5955
R186 Y.n8 Y.t5 26.5955
R187 Y.n8 Y.t7 26.5955
R188 Y.n0 Y.t12 26.5955
R189 Y.n0 Y.t15 26.5955
R190 Y.n1 Y.t14 26.5955
R191 Y.n1 Y.t13 26.5955
R192 Y.n3 Y.t8 26.5955
R193 Y.n3 Y.t11 26.5955
R194 Y.n11 Y.t6 24.9236
R195 Y.n11 Y.t0 24.9236
R196 Y.n12 Y.t2 24.9236
R197 Y.n12 Y.t1 24.9236
R198 Y Y.n10 14.2694
R199 Y Y.n9 10.7434
R200 Y.n10 Y.n6 8.11479
R201 Y.n10 Y 0.343357
R202 VPB.t4 VPB.t9 556.386
R203 VPB.t12 VPB.t3 556.386
R204 VPB.t11 VPB.t8 248.599
R205 VPB.t10 VPB.t11 248.599
R206 VPB.t9 VPB.t10 248.599
R207 VPB.t7 VPB.t4 248.599
R208 VPB.t6 VPB.t7 248.599
R209 VPB.t5 VPB.t6 248.599
R210 VPB.t0 VPB.t5 248.599
R211 VPB.t1 VPB.t0 248.599
R212 VPB.t2 VPB.t1 248.599
R213 VPB.t3 VPB.t2 248.599
R214 VPB VPB.t12 189.409
R215 a_27_47.t0 a_27_47.n10 279.733
R216 a_27_47.n2 a_27_47.t5 221.72
R217 a_27_47.n1 a_27_47.t6 221.72
R218 a_27_47.n6 a_27_47.t7 221.72
R219 a_27_47.n8 a_27_47.t9 221.72
R220 a_27_47.n9 a_27_47.n8 194.845
R221 a_27_47.n4 a_27_47.n3 178.881
R222 a_27_47.n7 a_27_47.n0 152
R223 a_27_47.n5 a_27_47.n4 152
R224 a_27_47.n2 a_27_47.t4 149.421
R225 a_27_47.n1 a_27_47.t3 149.421
R226 a_27_47.n6 a_27_47.t8 149.421
R227 a_27_47.n8 a_27_47.t2 149.421
R228 a_27_47.n10 a_27_47.t1 138.095
R229 a_27_47.n10 a_27_47.n9 55.0742
R230 a_27_47.n3 a_27_47.n2 37.4894
R231 a_27_47.n3 a_27_47.n1 37.4894
R232 a_27_47.n5 a_27_47.n1 37.4894
R233 a_27_47.n6 a_27_47.n5 37.4894
R234 a_27_47.n7 a_27_47.n6 37.4894
R235 a_27_47.n8 a_27_47.n7 37.4894
R236 a_27_47.n4 a_27_47.n0 26.8805
R237 a_27_47.n9 a_27_47.n0 22.1262
R238 a_215_47.n3 a_215_47.t7 319.277
R239 a_215_47.n1 a_215_47.t0 319.277
R240 a_215_47.n1 a_215_47.n0 185
R241 a_215_47.n3 a_215_47.n2 185
R242 a_215_47.n5 a_215_47.n4 185
R243 a_215_47.n4 a_215_47.n1 51.2005
R244 a_215_47.n4 a_215_47.n3 51.2005
R245 a_215_47.n2 a_215_47.t6 24.9236
R246 a_215_47.n2 a_215_47.t4 24.9236
R247 a_215_47.n0 a_215_47.t2 24.9236
R248 a_215_47.n0 a_215_47.t1 24.9236
R249 a_215_47.t3 a_215_47.n5 24.9236
R250 a_215_47.n5 a_215_47.t5 24.9236
R251 A_N.n0 A_N.t0 237.655
R252 A_N.n0 A_N.t1 165.356
R253 A_N A_N.n0 154.012
C0 VPWR VGND 0.16685f
C1 Y VGND 0.038593f
C2 VPB A_N 0.039378f
C3 VPB B 0.120652f
C4 VPB C 0.142934f
C5 VPB VPWR 0.178217f
C6 B C 0.033231f
C7 A_N VPWR 0.041327f
C8 VPB Y 0.031453f
C9 A_N Y 2.4e-19
C10 B VPWR 0.048702f
C11 VPB VGND 0.014069f
C12 B Y 0.221701f
C13 A_N VGND 0.015614f
C14 C VPWR 0.064148f
C15 B VGND 0.031015f
C16 C Y 0.220297f
C17 C VGND 0.059214f
C18 VPWR Y 1.13685f
C19 VGND VNB 0.851911f
C20 Y VNB 0.018998f
C21 VPWR VNB 0.717408f
C22 C VNB 0.42729f
C23 B VNB 0.361267f
C24 A_N VNB 0.130941f
C25 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_1 VPB VNB VPWR VGND A C D Y B
X0 Y.t1 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t2 A.t0 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR.t3 C.t0 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47.t1 C.t1 a_109_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t3 A.t1 a_277_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_277_47.t1 B.t1 a_193_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t0 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47.t1 D.t1 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t0 241.536
R1 B B.n0 184.056
R2 B.n0 B.t1 169.237
R3 VPWR.n2 VPWR.t2 347.216
R4 VPWR.n3 VPWR.n1 320.976
R5 VPWR.n5 VPWR.t0 249.362
R6 VPWR.n4 VPWR.n3 30.8711
R7 VPWR.n1 VPWR.t1 26.5955
R8 VPWR.n1 VPWR.t3 26.5955
R9 VPWR.n5 VPWR.n4 25.977
R10 VPWR.n3 VPWR.n2 10.9762
R11 VPWR.n4 VPWR.n0 9.3005
R12 VPWR.n6 VPWR.n5 9.3005
R13 VPWR.n2 VPWR.n0 0.523738
R14 VPWR.n6 VPWR.n0 0.120292
R15 VPWR VPWR.n6 0.0213333
R16 Y.n2 Y.n1 258.363
R17 Y.n2 Y.n0 202.095
R18 Y.n3 Y.t3 132.982
R19 Y.n3 Y.n2 62.4946
R20 Y.n0 Y.t2 32.5055
R21 Y.n0 Y.t1 32.5055
R22 Y.n1 Y.t4 26.5955
R23 Y.n1 Y.t0 26.5955
R24 Y Y.n3 4.04261
R25 VPB.t1 VPB.t2 284.113
R26 VPB.t3 VPB.t1 248.599
R27 VPB.t0 VPB.t3 248.599
R28 VPB VPB.t0 189.409
R29 A.n0 A.t0 228.649
R30 A.n0 A.t1 156.35
R31 A A.n0 153.434
R32 C.n0 C.t0 241.536
R33 C.n0 C.t1 169.237
R34 C C.n0 162.862
R35 a_109_47.t0 a_109_47.t1 49.8467
R36 a_193_47.t0 a_193_47.t1 49.8467
R37 VNB.t1 VNB.t0 1366.99
R38 VNB.t2 VNB.t1 1196.12
R39 VNB.t3 VNB.t2 1196.12
R40 VNB VNB.t3 911.327
R41 a_277_47.t0 a_277_47.t1 60.9236
R42 D.n0 D.t0 231.017
R43 D.n0 D.t1 158.716
R44 D D.n0 156.268
R45 VGND VGND.t0 156.477
C0 VPB A 0.044229f
C1 C B 0.141978f
C2 VPB VPWR 0.06379f
C3 VPB Y 0.009854f
C4 D VPWR 0.043786f
C5 D Y 0.01167f
C6 B A 0.05084f
C7 C VPWR 0.017084f
C8 VPB VGND 0.005518f
C9 C Y 0.05106f
C10 B VPWR 0.018371f
C11 D VGND 0.05031f
C12 B Y 0.135767f
C13 C VGND 0.087258f
C14 A VPWR 0.044315f
C15 A Y 0.114624f
C16 B VGND 0.05182f
C17 VPWR Y 0.362705f
C18 A VGND 0.009735f
C19 VPB D 0.036864f
C20 VPWR VGND 0.050206f
C21 VPB C 0.02565f
C22 Y VGND 0.096772f
C23 VPB B 0.026752f
C24 D C 0.091581f
C25 VGND VNB 0.318472f
C26 Y VNB 0.046422f
C27 VPWR VNB 0.309872f
C28 A VNB 0.162204f
C29 B VNB 0.091902f
C30 C VNB 0.096347f
C31 D VNB 0.143483f
C32 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_2 VNB VPB VGND VPWR D C Y B A
X0 VPWR.t5 C.t0 Y.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_47.t3 B.t0 a_277_47.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t6 C.t1 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t2 D.t0 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t0 A.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47.t3 D.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47.t1 C.t2 a_277_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t1 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X8 a_277_47.t3 B.t1 a_471_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VPWR.t6 B.t2 Y.t8 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X10 Y.t2 A.t2 a_471_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_277_47.t0 C.t3 a_27_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y.t9 B.t3 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X13 a_471_47.t1 A.t3 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t5 D.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t0 D.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C.n0 C.t0 221.72
R1 C.n1 C.t1 221.72
R2 C.n3 C.n2 152
R3 C.n0 C.t2 149.421
R4 C.n1 C.t3 149.421
R5 C.n2 C.n0 37.4894
R6 C.n2 C.n1 37.4894
R7 C C.n3 28.8005
R8 C.n3 C 0.6405
R9 Y.n3 Y.n1 235.923
R10 Y.n3 Y.n2 206.25
R11 Y.n5 Y.n4 206.25
R12 Y.n6 Y.n0 204.565
R13 Y Y.n7 199.148
R14 Y.n5 Y.n3 38.9823
R15 Y.n6 Y 26.7641
R16 Y.n1 Y.t3 26.5955
R17 Y.n1 Y.t5 26.5955
R18 Y.n2 Y.t7 26.5955
R19 Y.n2 Y.t6 26.5955
R20 Y.n4 Y.t8 26.5955
R21 Y.n4 Y.t9 26.5955
R22 Y.n0 Y.t0 26.5955
R23 Y.n0 Y.t1 26.5955
R24 Y.n7 Y.t4 24.9236
R25 Y.n7 Y.t2 24.9236
R26 Y Y.n5 13.0914
R27 Y.n5 Y 4.26717
R28 Y Y.n6 2.53744
R29 VPWR.n16 VPWR.n1 320.976
R30 VPWR.n11 VPWR.n4 310.502
R31 VPWR.n6 VPWR.n5 310.502
R32 VPWR.n7 VPWR.t0 265.426
R33 VPWR.n18 VPWR.t3 249.901
R34 VPWR.n5 VPWR.t6 69.9355
R35 VPWR.n5 VPWR.t1 62.0555
R36 VPWR.n4 VPWR.t7 42.3555
R37 VPWR.n4 VPWR.t5 42.3555
R38 VPWR.n15 VPWR.n2 34.6358
R39 VPWR.n10 VPWR.n9 34.6358
R40 VPWR.n17 VPWR.n16 30.8711
R41 VPWR.n1 VPWR.t4 26.5955
R42 VPWR.n1 VPWR.t2 26.5955
R43 VPWR.n18 VPWR.n17 25.977
R44 VPWR.n11 VPWR.n10 25.977
R45 VPWR.n11 VPWR.n2 18.4476
R46 VPWR.n7 VPWR.n6 16.4929
R47 VPWR.n9 VPWR.n8 9.3005
R48 VPWR.n10 VPWR.n3 9.3005
R49 VPWR.n12 VPWR.n11 9.3005
R50 VPWR.n13 VPWR.n2 9.3005
R51 VPWR.n15 VPWR.n14 9.3005
R52 VPWR.n17 VPWR.n0 9.3005
R53 VPWR.n19 VPWR.n18 9.3005
R54 VPWR.n16 VPWR.n15 3.76521
R55 VPWR.n8 VPWR.n7 0.634969
R56 VPWR.n9 VPWR.n6 0.376971
R57 VPWR.n8 VPWR.n3 0.120292
R58 VPWR.n12 VPWR.n3 0.120292
R59 VPWR.n13 VPWR.n12 0.120292
R60 VPWR.n14 VPWR.n13 0.120292
R61 VPWR.n14 VPWR.n0 0.120292
R62 VPWR.n19 VPWR.n0 0.120292
R63 VPWR VPWR.n19 0.0213333
R64 VPB.t6 VPB.t1 485.358
R65 VPB.t5 VPB.t7 343.303
R66 VPB.t1 VPB.t0 248.599
R67 VPB.t7 VPB.t6 248.599
R68 VPB.t4 VPB.t5 248.599
R69 VPB.t2 VPB.t4 248.599
R70 VPB.t3 VPB.t2 248.599
R71 VPB VPB.t3 189.409
R72 B.n4 B.t3 237.787
R73 B.n2 B.t2 221.72
R74 B.n1 B.t0 192.264
R75 B B.n4 155.201
R76 B.n1 B.n0 152
R77 B.n3 B.t1 149.421
R78 B.n4 B.n3 55.3412
R79 B.n2 B.n1 28.5635
R80 B B.n0 28.1605
R81 B.n3 B.n2 3.57087
R82 B.n0 B 1.2805
R83 a_277_47.n1 a_277_47.n0 436.37
R84 a_277_47.n0 a_277_47.t2 24.9236
R85 a_277_47.n0 a_277_47.t3 24.9236
R86 a_277_47.n1 a_277_47.t1 24.9236
R87 a_277_47.t0 a_277_47.n1 24.9236
R88 a_471_47.t2 a_471_47.n1 314.562
R89 a_471_47.n1 a_471_47.t1 182.172
R90 a_471_47.n1 a_471_47.n0 97.0637
R91 a_471_47.n0 a_471_47.t0 24.9236
R92 a_471_47.n0 a_471_47.t3 24.9236
R93 VNB.t5 VNB.t6 2790.94
R94 VNB.t0 VNB.t1 1196.12
R95 VNB.t7 VNB.t0 1196.12
R96 VNB.t6 VNB.t7 1196.12
R97 VNB.t4 VNB.t5 1196.12
R98 VNB.t3 VNB.t4 1196.12
R99 VNB.t2 VNB.t3 1196.12
R100 VNB VNB.t2 911.327
R101 D.n2 D.t2 234.573
R102 D.n0 D.t0 221.72
R103 D.n2 D.t3 162.274
R104 D.n1 D 156.481
R105 D.n3 D.n2 152
R106 D.n0 D.t1 149.421
R107 D.n1 D.n0 37.4894
R108 D.n2 D.n1 24.1005
R109 D.n3 D 21.4405
R110 D D.n3 8.0005
R111 A.n0 A.t1 221.72
R112 A.n1 A.t0 218.507
R113 A A.n1 213.969
R114 A.n0 A.t2 149.421
R115 A.n1 A.t3 146.208
R116 A.n1 A.n0 74.0549
R117 VGND VGND.n0 214.335
R118 VGND.n0 VGND.t1 24.9236
R119 VGND.n0 VGND.t0 24.9236
R120 a_27_47.t1 a_27_47.n1 318.719
R121 a_27_47.n1 a_27_47.t2 190.405
R122 a_27_47.n1 a_27_47.n0 88.3446
R123 a_27_47.n0 a_27_47.t0 24.9236
R124 a_27_47.n0 a_27_47.t3 24.9236
C0 VPB D 0.069252f
C1 VPB C 0.054058f
C2 D C 0.067173f
C3 VPB B 0.076937f
C4 VPWR VPB 0.109103f
C5 VPB A 0.08242f
C6 VPWR D 0.058844f
C7 Y VPB 0.021153f
C8 C B 0.03543f
C9 Y D 0.063269f
C10 VPWR C 0.033381f
C11 VGND VPB 0.00787f
C12 VGND D 0.029651f
C13 Y C 0.09522f
C14 VPWR B 0.038579f
C15 B A 0.039642f
C16 VPWR A 0.065928f
C17 Y B 0.133834f
C18 VGND C 0.017465f
C19 VPWR Y 0.787425f
C20 VGND B 0.01908f
C21 Y A 0.08649f
C22 VPWR VGND 0.095336f
C23 VGND A 0.018365f
C24 Y VGND 0.020194f
C25 VGND VNB 0.525212f
C26 Y VNB 0.028202f
C27 VPWR VNB 0.508353f
C28 A VNB 0.246867f
C29 B VNB 0.216473f
C30 C VNB 0.178935f
C31 D VNB 0.232315f
C32 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_4 A D C B Y VPWR VGND VPB VNB
X0 a_27_47.t3 C.t0 a_445_47.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47.t2 C.t1 a_445_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t10 C.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t7 D.t0 Y.t11 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t11 A.t0 Y.t15 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t6 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_47.t0 B.t0 a_803_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t12 D.t1 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_445_47.t7 B.t1 a_803_47.t2 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR.t9 D.t2 Y.t13 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t0 A.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47.t4 D.t3 VGND.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_47.t5 D.t4 VGND.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t1 A.t3 a_803_47.t7 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X14 Y.t2 A.t4 a_803_47.t6 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_803_47.t1 B.t2 a_445_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t5 C.t3 Y.t9 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47.t0 B.t3 a_445_47.t6 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t1 D.t5 a_27_47.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_445_47.t4 C.t4 a_27_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y.t8 C.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_803_47.t5 A.t5 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t12 B.t4 Y.t16 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X23 Y.t4 A.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X24 a_445_47.t3 C.t6 a_27_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_803_47.t4 A.t7 Y.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t3 C.t7 Y.t7 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t17 B.t5 VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VPWR.t14 B.t6 Y.t18 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y.t14 D.t6 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 Y.t19 B.t7 VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND.t0 D.t7 a_27_47.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C.n0 C.t3 221.72
R1 C.n7 C.t5 221.72
R2 C.n1 C.t7 221.72
R3 C.n2 C.t2 221.72
R4 C.n9 C.n8 152
R5 C.n6 C.n5 152
R6 C.n4 C.n3 152
R7 C.n0 C.t1 149.421
R8 C.n7 C.t6 149.421
R9 C.n1 C.t0 149.421
R10 C.n2 C.t4 149.421
R11 C.n3 C.n1 38.382
R12 C.n8 C.n0 37.4894
R13 C.n8 C.n7 37.4894
R14 C.n7 C.n6 37.4894
R15 C.n6 C.n1 37.4894
R16 C.n3 C.n2 36.5968
R17 C.n4 C 23.3605
R18 C.n5 C 21.1205
R19 C.n9 C 18.5605
R20 C C.n9 10.8805
R21 C.n5 C 8.3205
R22 C C.n4 6.0805
R23 a_445_47.n5 a_445_47.n4 228.008
R24 a_445_47.n2 a_445_47.n0 228.008
R25 a_445_47.n4 a_445_47.n3 185
R26 a_445_47.n2 a_445_47.n1 185
R27 a_445_47.n4 a_445_47.n2 69.6325
R28 a_445_47.n0 a_445_47.t2 24.9236
R29 a_445_47.n0 a_445_47.t4 24.9236
R30 a_445_47.n1 a_445_47.t1 24.9236
R31 a_445_47.n1 a_445_47.t3 24.9236
R32 a_445_47.n3 a_445_47.t6 24.9236
R33 a_445_47.n3 a_445_47.t7 24.9236
R34 a_445_47.n5 a_445_47.t5 24.9236
R35 a_445_47.t0 a_445_47.n5 24.9236
R36 a_27_47.n4 a_27_47.t2 305.594
R37 a_27_47.n1 a_27_47.t7 256.36
R38 a_27_47.n1 a_27_47.n0 187.26
R39 a_27_47.n3 a_27_47.n2 185
R40 a_27_47.n5 a_27_47.n4 185
R41 a_27_47.n4 a_27_47.n3 57.2895
R42 a_27_47.n3 a_27_47.n1 45.2673
R43 a_27_47.n2 a_27_47.t1 24.9236
R44 a_27_47.n2 a_27_47.t5 24.9236
R45 a_27_47.n0 a_27_47.t6 24.9236
R46 a_27_47.n0 a_27_47.t4 24.9236
R47 a_27_47.n5 a_27_47.t0 24.9236
R48 a_27_47.t3 a_27_47.n5 24.9236
R49 VNB.t7 VNB.t15 2677.02
R50 VNB.t13 VNB.t0 1366.99
R51 VNB.t1 VNB.t3 1196.12
R52 VNB.t2 VNB.t1 1196.12
R53 VNB.t0 VNB.t2 1196.12
R54 VNB.t4 VNB.t13 1196.12
R55 VNB.t14 VNB.t4 1196.12
R56 VNB.t15 VNB.t14 1196.12
R57 VNB.t5 VNB.t7 1196.12
R58 VNB.t8 VNB.t5 1196.12
R59 VNB.t6 VNB.t8 1196.12
R60 VNB.t10 VNB.t6 1196.12
R61 VNB.t11 VNB.t10 1196.12
R62 VNB.t9 VNB.t11 1196.12
R63 VNB.t12 VNB.t9 1196.12
R64 VNB VNB.t12 911.327
R65 VPWR.n40 VPWR.n1 320.976
R66 VPWR.n34 VPWR.n33 320.976
R67 VPWR.n31 VPWR.n4 320.976
R68 VPWR.n9 VPWR.n8 320.976
R69 VPWR.n19 VPWR.n11 320.976
R70 VPWR.n14 VPWR.n13 320.976
R71 VPWR.n15 VPWR.t11 254.838
R72 VPWR.n42 VPWR.t10 249.901
R73 VPWR.n26 VPWR.n7 133.066
R74 VPWR.n7 VPWR.t5 70.1844
R75 VPWR.n7 VPWR.t15 70.1841
R76 VPWR.n15 VPWR.n14 36.2765
R77 VPWR.n30 VPWR.n5 34.6358
R78 VPWR.n35 VPWR.n32 34.6358
R79 VPWR.n39 VPWR.n2 34.6358
R80 VPWR.n18 VPWR.n12 34.6358
R81 VPWR.n21 VPWR.n20 34.6358
R82 VPWR.n25 VPWR.n24 34.6358
R83 VPWR.n11 VPWR.t12 33.4905
R84 VPWR.n11 VPWR.t1 31.5205
R85 VPWR.n41 VPWR.n40 30.8711
R86 VPWR.n19 VPWR.n18 26.7299
R87 VPWR.n1 VPWR.t8 26.5955
R88 VPWR.n1 VPWR.t9 26.5955
R89 VPWR.n33 VPWR.t6 26.5955
R90 VPWR.n33 VPWR.t7 26.5955
R91 VPWR.n4 VPWR.t4 26.5955
R92 VPWR.n4 VPWR.t3 26.5955
R93 VPWR.n8 VPWR.t13 26.5955
R94 VPWR.n8 VPWR.t14 26.5955
R95 VPWR.n13 VPWR.t2 26.5955
R96 VPWR.n13 VPWR.t0 26.5955
R97 VPWR.n42 VPWR.n41 25.977
R98 VPWR.n34 VPWR.n2 24.8476
R99 VPWR.n21 VPWR.n9 23.3417
R100 VPWR.n32 VPWR.n31 18.824
R101 VPWR.n31 VPWR.n30 15.8123
R102 VPWR.n24 VPWR.n9 11.2946
R103 VPWR.n26 VPWR.n25 10.9181
R104 VPWR.n35 VPWR.n34 9.78874
R105 VPWR.n16 VPWR.n12 9.3005
R106 VPWR.n18 VPWR.n17 9.3005
R107 VPWR.n20 VPWR.n10 9.3005
R108 VPWR.n22 VPWR.n21 9.3005
R109 VPWR.n24 VPWR.n23 9.3005
R110 VPWR.n25 VPWR.n6 9.3005
R111 VPWR.n27 VPWR.n26 9.3005
R112 VPWR.n28 VPWR.n5 9.3005
R113 VPWR.n30 VPWR.n29 9.3005
R114 VPWR.n32 VPWR.n3 9.3005
R115 VPWR.n36 VPWR.n35 9.3005
R116 VPWR.n37 VPWR.n2 9.3005
R117 VPWR.n39 VPWR.n38 9.3005
R118 VPWR.n41 VPWR.n0 9.3005
R119 VPWR.n43 VPWR.n42 9.3005
R120 VPWR.n20 VPWR.n19 7.90638
R121 VPWR.n26 VPWR.n5 6.4005
R122 VPWR.n40 VPWR.n39 3.76521
R123 VPWR.n14 VPWR.n12 3.76521
R124 VPWR.n16 VPWR.n15 2.08078
R125 VPWR.n17 VPWR.n16 0.120292
R126 VPWR.n17 VPWR.n10 0.120292
R127 VPWR.n22 VPWR.n10 0.120292
R128 VPWR.n23 VPWR.n22 0.120292
R129 VPWR.n23 VPWR.n6 0.120292
R130 VPWR.n27 VPWR.n6 0.120292
R131 VPWR.n28 VPWR.n27 0.120292
R132 VPWR.n29 VPWR.n28 0.120292
R133 VPWR.n29 VPWR.n3 0.120292
R134 VPWR.n36 VPWR.n3 0.120292
R135 VPWR.n37 VPWR.n36 0.120292
R136 VPWR.n38 VPWR.n37 0.120292
R137 VPWR.n38 VPWR.n0 0.120292
R138 VPWR.n43 VPWR.n0 0.120292
R139 VPWR VPWR.n43 0.0213333
R140 Y.n2 Y.n1 245.523
R141 Y.n5 Y.n3 235.923
R142 Y.n17 Y.n15 228.008
R143 Y.n5 Y.n4 206.25
R144 Y.n7 Y.n6 206.25
R145 Y.n9 Y.n8 206.25
R146 Y.n11 Y.n10 206.25
R147 Y.n13 Y.n12 206.25
R148 Y.n2 Y.n0 202.095
R149 Y.n17 Y.n16 185
R150 Y.n11 Y.n9 59.9278
R151 Y.n14 Y.n13 36.946
R152 Y.n7 Y.n5 29.6732
R153 Y.n9 Y.n7 29.6732
R154 Y.n13 Y.n11 29.6732
R155 Y.n0 Y.t0 26.5955
R156 Y.n0 Y.t4 26.5955
R157 Y.n3 Y.t13 26.5955
R158 Y.n3 Y.t14 26.5955
R159 Y.n4 Y.t11 26.5955
R160 Y.n4 Y.t12 26.5955
R161 Y.n6 Y.t7 26.5955
R162 Y.n6 Y.t10 26.5955
R163 Y.n8 Y.t9 26.5955
R164 Y.n8 Y.t8 26.5955
R165 Y.n10 Y.t18 26.5955
R166 Y.n10 Y.t19 26.5955
R167 Y.n12 Y.t16 26.5955
R168 Y.n12 Y.t17 26.5955
R169 Y.n1 Y.t15 26.5955
R170 Y.n1 Y.t6 26.5955
R171 Y.n16 Y.t3 24.9236
R172 Y.n16 Y.t1 24.9236
R173 Y.n15 Y.t5 24.9236
R174 Y.n15 Y.t2 24.9236
R175 Y Y.n14 24.1783
R176 Y Y.n17 19.3427
R177 Y.n14 Y.n2 5.81868
R178 VPB.t5 VPB.t15 556.386
R179 VPB.t12 VPB.t1 284.113
R180 VPB.t2 VPB.t11 248.599
R181 VPB.t0 VPB.t2 248.599
R182 VPB.t1 VPB.t0 248.599
R183 VPB.t13 VPB.t12 248.599
R184 VPB.t14 VPB.t13 248.599
R185 VPB.t15 VPB.t14 248.599
R186 VPB.t4 VPB.t5 248.599
R187 VPB.t3 VPB.t4 248.599
R188 VPB.t6 VPB.t3 248.599
R189 VPB.t7 VPB.t6 248.599
R190 VPB.t8 VPB.t7 248.599
R191 VPB.t9 VPB.t8 248.599
R192 VPB.t10 VPB.t9 248.599
R193 VPB VPB.t10 189.409
R194 D.n2 D.t6 234.392
R195 D.n1 D.t0 221.72
R196 D.n8 D.t1 221.72
R197 D.n6 D.t2 221.72
R198 D.n2 D.t7 162.091
R199 D.n10 D.n9 152
R200 D.n7 D.n0 152
R201 D.n5 D.n4 152
R202 D.n3 D.n2 152
R203 D.n1 D.t4 149.421
R204 D.n8 D.t5 149.421
R205 D.n6 D.t3 149.421
R206 D.n9 D.n1 37.4894
R207 D.n9 D.n8 37.4894
R208 D.n8 D.n7 37.4894
R209 D.n7 D.n6 37.4894
R210 D.n6 D.n5 37.4894
R211 D.n10 D.n0 26.8805
R212 D.n4 D 24.9605
R213 D.n5 D.n2 24.1005
R214 D D.n3 21.4405
R215 D.n3 D 8.0005
R216 D.n4 D 4.4805
R217 D D.n0 1.9205
R218 D D.n10 0.6405
R219 A.n0 A.t0 234.573
R220 A.n3 A.t1 221.72
R221 A.n5 A.t2 221.72
R222 A.n4 A.t6 221.72
R223 A.n0 A.t7 162.274
R224 A A.n0 154.881
R225 A.n2 A.n1 152
R226 A.n7 A.n6 152
R227 A.n3 A.t4 149.421
R228 A.n5 A.t5 149.421
R229 A.n4 A.t3 149.421
R230 A.n5 A.n4 74.9783
R231 A.n6 A.n3 53.5561
R232 A.n2 A.n0 40.1672
R233 A.n1 A 28.8005
R234 A.n7 A 26.2405
R235 A.n3 A.n2 21.4227
R236 A.n6 A.n5 21.4227
R237 A A.n7 3.2005
R238 A.n1 A 0.6405
R239 B.n0 B.t4 221.72
R240 B.n2 B.t5 221.72
R241 B.n7 B.t6 221.72
R242 B.n3 B.t7 221.72
R243 B.n4 B.n3 194.845
R244 B B.n1 162.881
R245 B.n9 B.n8 152
R246 B.n6 B.n5 152
R247 B.n0 B.t2 149.421
R248 B.n2 B.t0 149.421
R249 B.n7 B.t3 149.421
R250 B.n3 B.t1 149.421
R251 B.n1 B.n0 37.4894
R252 B.n2 B.n1 37.4894
R253 B.n8 B.n2 37.4894
R254 B.n8 B.n7 37.4894
R255 B.n7 B.n6 37.4894
R256 B.n6 B.n3 37.4894
R257 B.n4 B 16.6405
R258 B B.n9 16.0005
R259 B.n5 B 16.0005
R260 B.n9 B 13.4405
R261 B.n5 B 13.4405
R262 B B.n4 12.8005
R263 a_803_47.n4 a_803_47.t2 305.594
R264 a_803_47.n2 a_803_47.n1 185
R265 a_803_47.n5 a_803_47.n4 185
R266 a_803_47.n2 a_803_47.t4 179.204
R267 a_803_47.n3 a_803_47.n0 97.0637
R268 a_803_47.n4 a_803_47.n3 48.6962
R269 a_803_47.n3 a_803_47.n2 48.1396
R270 a_803_47.n0 a_803_47.t1 31.3851
R271 a_803_47.n0 a_803_47.t7 29.539
R272 a_803_47.n1 a_803_47.t6 24.9236
R273 a_803_47.n1 a_803_47.t5 24.9236
R274 a_803_47.t3 a_803_47.n5 24.9236
R275 a_803_47.n5 a_803_47.t0 24.9236
R276 VGND.n2 VGND.n0 205.85
R277 VGND.n2 VGND.n1 205.812
R278 VGND.n0 VGND.t2 24.9236
R279 VGND.n0 VGND.t1 24.9236
R280 VGND.n1 VGND.t3 24.9236
R281 VGND.n1 VGND.t0 24.9236
R282 VGND VGND.n2 0.56252
C0 A Y 0.285339f
C1 B VGND 0.033063f
C2 VPB D 0.133279f
C3 VPWR Y 1.54639f
C4 A VGND 0.0344f
C5 VPB C 0.121158f
C6 VPWR VGND 0.157147f
C7 D C 0.064343f
C8 VPB B 0.137603f
C9 Y VGND 0.037539f
C10 VPB A 0.133308f
C11 VPB VPWR 0.165034f
C12 C B 0.033231f
C13 VPB Y 0.033927f
C14 D VPWR 0.095209f
C15 VPB VGND 0.010343f
C16 C VPWR 0.050251f
C17 D Y 0.176233f
C18 B A 0.042327f
C19 C Y 0.212028f
C20 D VGND 0.065788f
C21 B VPWR 0.058268f
C22 C VGND 0.030813f
C23 A VPWR 0.093918f
C24 B Y 0.24258f
C25 VGND VNB 0.836562f
C26 Y VNB 0.025935f
C27 VPWR VNB 0.790844f
C28 A VNB 0.417528f
C29 B VNB 0.397122f
C30 C VNB 0.363172f
C31 D VNB 0.417482f
C32 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_1 VPB VNB VGND VPWR Y C B D A_N
X0 Y.t1 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47.t0 D.t0 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.118125 ps=1.04 w=0.65 l=0.15
X2 VPWR.t4 C.t0 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t2 A_N.t0 a_41_93.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR.t3 a_41_93.t2 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
X5 a_316_47.t0 C.t1 a_232_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t2 a_41_93.t3 a_423_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_423_47.t0 B.t1 a_316_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.125125 ps=1.035 w=0.65 l=0.15
X8 Y.t0 D.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X9 VGND.t1 A_N.t1 a_41_93.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.1113 ps=1.37 w=0.42 l=0.15
R0 B.n0 B.t0 241.536
R1 B.n0 B.t1 169.237
R2 B B.n0 154.63
R3 VPWR.n4 VPWR.t3 354.726
R4 VPWR.n3 VPWR.n2 313.337
R5 VPWR.n8 VPWR.n1 224.139
R6 VPWR.n1 VPWR.t2 95.3969
R7 VPWR.n2 VPWR.t4 38.4155
R8 VPWR.n2 VPWR.t1 37.4305
R9 VPWR.n7 VPWR.n6 34.6358
R10 VPWR.n1 VPWR.t0 26.3637
R11 VPWR.n4 VPWR.n3 18.5848
R12 VPWR.n8 VPWR.n7 14.3064
R13 VPWR.n6 VPWR.n5 9.3005
R14 VPWR.n7 VPWR.n0 9.3005
R15 VPWR.n9 VPWR.n8 9.16498
R16 VPWR.n6 VPWR.n3 1.50638
R17 VPWR.n5 VPWR.n4 0.81264
R18 VPWR.n9 VPWR.n0 0.141672
R19 VPWR VPWR.n9 0.121778
R20 VPWR.n5 VPWR.n0 0.120292
R21 Y.n2 Y.n0 252.339
R22 Y.n2 Y.n1 205.087
R23 Y Y.n4 186.31
R24 Y.n4 Y.n3 185
R25 Y.n3 Y.n2 87.4741
R26 Y.n1 Y.t3 50.2355
R27 Y.n4 Y.t2 37.8467
R28 Y.n0 Y.t4 26.5955
R29 Y.n0 Y.t0 26.5955
R30 Y.n1 Y.t1 26.5955
R31 Y Y.n3 8.58232
R32 VPB.t1 VPB.t3 319.627
R33 VPB.t4 VPB.t1 316.668
R34 VPB.t2 VPB.t0 287.072
R35 VPB VPB.t2 269.315
R36 VPB.t0 VPB.t4 248.599
R37 D.n0 D.t1 236.18
R38 D.n0 D.t0 163.881
R39 D D.n0 154.607
R40 VGND VGND.n0 221.02
R41 VGND.n0 VGND.t1 65.7148
R42 VGND.n0 VGND.t0 29.539
R43 a_232_47.t0 a_232_47.t1 49.8467
R44 VNB.t0 VNB.t1 1537.86
R45 VNB.t3 VNB.t2 1537.86
R46 VNB.t4 VNB.t0 1523.62
R47 VNB.t2 VNB.t4 1196.12
R48 VNB VNB.t3 1139.16
R49 C.n0 C.t0 236.18
R50 C.n0 C.t1 163.881
R51 C C.n0 153.487
R52 A_N A_N.n0 155.685
R53 A_N.n0 A_N.t0 142.994
R54 A_N.n0 A_N.t1 126.927
R55 a_41_93.t0 a_41_93.n1 720.221
R56 a_41_93.n1 a_41_93.n0 346.68
R57 a_41_93.n0 a_41_93.t2 236.18
R58 a_41_93.n1 a_41_93.t1 225
R59 a_41_93.n0 a_41_93.t3 163.881
R60 a_316_47.t0 a_316_47.t1 71.0774
R61 a_423_47.t0 a_423_47.t1 72.0005
C0 D C 0.079607f
C1 D VPB 0.031831f
C2 C VPB 0.02995f
C3 C B 0.094117f
C4 D VPWR 0.022205f
C5 B VPB 0.028738f
C6 D A_N 0.065226f
C7 C VPWR 0.017889f
C8 VPWR VPB 0.095142f
C9 D Y 0.020099f
C10 C A_N 3.73e-19
C11 B VPWR 0.01496f
C12 A_N VPB 0.042324f
C13 D VGND 0.014903f
C14 C Y 0.040828f
C15 Y VPB 0.019327f
C16 B Y 0.041915f
C17 C VGND 0.012914f
C18 VPWR A_N 0.020952f
C19 VGND VPB 0.0096f
C20 B VGND 0.009795f
C21 VPWR Y 0.401971f
C22 VPWR VGND 0.064985f
C23 A_N Y 8.57e-19
C24 A_N VGND 0.010976f
C25 Y VGND 0.066946f
C26 VGND VNB 0.399267f
C27 Y VNB 0.073761f
C28 A_N VNB 0.125593f
C29 VPWR VNB 0.368796f
C30 B VNB 0.092716f
C31 C VNB 0.097487f
C32 D VNB 0.100872f
C33 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_2 VNB VPB VGND VPWR A_N Y B C D
X0 Y.t1 a_27_47.t2 a_215_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_465_47.t1 B.t0 a_215_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t1 D.t0 a_655_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X3 a_215_47.t3 B.t1 a_465_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t8 A_N.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_655_47.t1 D.t1 VGND.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_655_47.t3 C.t0 a_465_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t1 B.t2 Y.t8 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t9 B.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_465_47.t2 C.t1 a_655_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VPWR.t5 a_27_47.t3 Y.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR.t7 C.t2 Y.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR.t3 D.t2 Y.t7 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=2.8 as=0.135 ps=1.27 w=1 l=0.15
X13 Y.t5 D.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X14 a_215_47.t0 a_27_47.t4 Y.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y.t2 a_27_47.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 Y.t4 C.t3 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X17 VGND.t2 A_N.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t0 a_27_47.n2 731.396
R1 a_27_47.n2 a_27_47.t1 276.529
R2 a_27_47.n2 a_27_47.n1 227.917
R3 a_27_47.n0 a_27_47.t3 212.081
R4 a_27_47.n1 a_27_47.t5 212.081
R5 a_27_47.n0 a_27_47.t4 139.78
R6 a_27_47.n1 a_27_47.t2 139.78
R7 a_27_47.n1 a_27_47.n0 61.346
R8 a_215_47.n0 a_215_47.t3 305.068
R9 a_215_47.n0 a_215_47.t1 189.496
R10 a_215_47.n1 a_215_47.n0 185
R11 a_215_47.n1 a_215_47.t2 24.9236
R12 a_215_47.t0 a_215_47.n1 24.9236
R13 Y.n3 Y.n1 347.93
R14 Y.n7 Y.n6 206.25
R15 Y.n3 Y.n2 206.25
R16 Y.n5 Y.n4 206.25
R17 Y Y.n0 187.452
R18 Y.n5 Y.n3 57.0187
R19 Y.n7 Y.n5 29.6732
R20 Y.n6 Y.t3 26.5955
R21 Y.n6 Y.t2 26.5955
R22 Y.n1 Y.t7 26.5955
R23 Y.n1 Y.t5 26.5955
R24 Y.n2 Y.t6 26.5955
R25 Y.n2 Y.t4 26.5955
R26 Y.n4 Y.t8 26.5955
R27 Y.n4 Y.t9 26.5955
R28 Y.n0 Y.t0 24.9236
R29 Y.n0 Y.t1 24.9236
R30 Y Y.n7 4.26717
R31 VNB.t7 VNB.t1 2677.02
R32 VNB.t4 VNB.t3 2677.02
R33 VNB.t5 VNB.t0 1452.43
R34 VNB.t0 VNB.t8 1196.12
R35 VNB.t1 VNB.t5 1196.12
R36 VNB.t6 VNB.t7 1196.12
R37 VNB.t2 VNB.t6 1196.12
R38 VNB.t3 VNB.t2 1196.12
R39 VNB VNB.t4 911.327
R40 B.n1 B.t2 212.081
R41 B.n2 B.t3 212.081
R42 B.n1 B.n0 180.482
R43 B.n4 B.n3 152
R44 B.n1 B.t1 139.78
R45 B.n2 B.t0 139.78
R46 B.n3 B.n1 45.2793
R47 B.n0 B 25.2805
R48 B B.n4 22.4005
R49 B.n3 B.n2 16.0672
R50 B.n4 B 7.0405
R51 B.n0 B 4.1605
R52 a_465_47.n1 a_465_47.n0 452.896
R53 a_465_47.n0 a_465_47.t3 24.9236
R54 a_465_47.n0 a_465_47.t2 24.9236
R55 a_465_47.n1 a_465_47.t0 24.9236
R56 a_465_47.t1 a_465_47.n1 24.9236
R57 D.n2 D.t3 219.383
R58 D.n1 D.t2 212.081
R59 D.n0 D 196.507
R60 D.n4 D.n3 152
R61 D.n2 D.t0 139.78
R62 D.n0 D.t1 139.78
R63 D.n3 D.n2 35.7853
R64 D.n4 D 26.5605
R65 D.n3 D.n1 18.2581
R66 D.n1 D.n0 7.30353
R67 D D.n4 2.8805
R68 a_655_47.t0 a_655_47.n1 300.377
R69 a_655_47.n1 a_655_47.t1 182.746
R70 a_655_47.n1 a_655_47.n0 94.8398
R71 a_655_47.n0 a_655_47.t2 33.2313
R72 a_655_47.n0 a_655_47.t3 33.2313
R73 VGND.n1 VGND.t2 244.06
R74 VGND.n1 VGND.n0 218.162
R75 VGND.n0 VGND.t0 24.9236
R76 VGND.n0 VGND.t1 24.9236
R77 VGND VGND.n1 0.146938
R78 A_N.n0 A_N.t0 323.55
R79 A_N.n0 A_N.t1 195.017
R80 A_N.n1 A_N.n0 152
R81 A_N.n1 A_N 15.2005
R82 A_N A_N.n1 2.93383
R83 VPWR.n23 VPWR.t8 648.322
R84 VPWR.n17 VPWR.n3 320.976
R85 VPWR.n9 VPWR.n7 315.334
R86 VPWR.n8 VPWR.t3 261.997
R87 VPWR.n1 VPWR.t4 228.946
R88 VPWR.n5 VPWR.n4 138.554
R89 VPWR.n4 VPWR.t6 76.3123
R90 VPWR.n4 VPWR.t1 60.5526
R91 VPWR.n7 VPWR.t2 37.4305
R92 VPWR.n16 VPWR.n15 34.6358
R93 VPWR.n11 VPWR.n10 34.6358
R94 VPWR.n24 VPWR.n23 34.5993
R95 VPWR.n7 VPWR.t7 33.4905
R96 VPWR.n18 VPWR.n17 32.377
R97 VPWR.n18 VPWR.n1 27.0577
R98 VPWR.n3 VPWR.t0 26.5955
R99 VPWR.n3 VPWR.t5 26.5955
R100 VPWR.n15 VPWR.n5 19.9534
R101 VPWR.n10 VPWR.n9 14.6829
R102 VPWR.n22 VPWR.n21 10.706
R103 VPWR.n10 VPWR.n6 9.3005
R104 VPWR.n12 VPWR.n11 9.3005
R105 VPWR.n13 VPWR.n5 9.3005
R106 VPWR.n15 VPWR.n14 9.3005
R107 VPWR.n16 VPWR.n2 9.3005
R108 VPWR.n19 VPWR.n18 9.3005
R109 VPWR.n21 VPWR.n20 9.3005
R110 VPWR.n22 VPWR.n0 9.3005
R111 VPWR.n9 VPWR.n8 7.48436
R112 VPWR.n17 VPWR.n16 2.25932
R113 VPWR.n11 VPWR.n5 1.12991
R114 VPWR.n8 VPWR.n6 0.61214
R115 VPWR.n21 VPWR.n1 0.555725
R116 VPWR.n23 VPWR.n22 0.233227
R117 VPWR.n12 VPWR.n6 0.120292
R118 VPWR.n13 VPWR.n12 0.120292
R119 VPWR.n14 VPWR.n13 0.120292
R120 VPWR.n14 VPWR.n2 0.120292
R121 VPWR.n19 VPWR.n2 0.120292
R122 VPWR.n20 VPWR.n19 0.120292
R123 VPWR.n20 VPWR.n0 0.120292
R124 VPWR.n24 VPWR.n0 0.120292
R125 VPWR VPWR.n24 0.0213333
R126 VPB.t8 VPB.t4 556.386
R127 VPB.t1 VPB.t6 526.792
R128 VPB.t7 VPB.t2 301.87
R129 VPB.t2 VPB.t3 248.599
R130 VPB.t6 VPB.t7 248.599
R131 VPB.t0 VPB.t1 248.599
R132 VPB.t5 VPB.t0 248.599
R133 VPB.t4 VPB.t5 248.599
R134 VPB VPB.t8 189.409
R135 C.n3 C.t3 219.383
R136 C.n2 C.t2 212.081
R137 C.n1 C.n0 152
R138 C.n5 C.n4 152
R139 C.n1 C.t0 141.242
R140 C.n3 C.t1 139.78
R141 C.n4 C.n2 48.2005
R142 C C.n5 18.5605
R143 C.n0 C 16.6405
R144 C.n0 C 12.8005
R145 C.n5 C 10.8805
R146 C.n2 C.n1 5.84292
R147 C.n4 C.n3 5.84292
C0 D Y 0.057679f
C1 C VGND 0.021358f
C2 VPWR Y 0.820498f
C3 D VGND 0.033632f
C4 VPB A_N 0.105575f
C5 VPWR VGND 0.112306f
C6 VPB B 0.070959f
C7 Y VGND 0.018003f
C8 VPB C 0.065819f
C9 VPB D 0.078576f
C10 VPB VPWR 0.132279f
C11 B C 0.036233f
C12 VPB Y 0.019172f
C13 A_N VPWR 0.020075f
C14 B VPWR 0.034993f
C15 VPB VGND 0.010854f
C16 C D 0.069591f
C17 A_N Y 0.00283f
C18 A_N VGND 0.017122f
C19 C VPWR 0.035026f
C20 B Y 0.151748f
C21 C Y 0.133313f
C22 B VGND 0.021753f
C23 D VPWR 0.076794f
C24 VGND VNB 0.63011f
C25 Y VNB 0.015271f
C26 VPWR VNB 0.547387f
C27 D VNB 0.246043f
C28 C VNB 0.194869f
C29 B VNB 0.207633f
C30 A_N VNB 0.209286f
C31 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_4 VNB VPB VGND VPWR D C B Y A_N
X0 a_991_47.t3 C.t0 a_633_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y.t19 B.t0 VPWR.t16 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_991_47.t6 D.t0 VGND.t3 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t8 a_27_47.t2 a_215_47.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_991_47.t7 D.t1 VGND.t2 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t9 a_27_47.t3 a_215_47.t2 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_633_47.t7 B.t1 a_215_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t15 B.t2 Y.t18 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t3 C.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_633_47.t0 B.t3 a_215_47.t6 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t1 D.t2 a_991_47.t4 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t2 C.t2 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t0 D.t3 a_991_47.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_215_47.t1 a_27_47.t4 Y.t10 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t1 C.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X15 a_215_47.t5 B.t4 a_633_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_215_47.t4 B.t5 a_633_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t5 D.t4 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t17 B.t6 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y.t5 D.t5 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t9 a_27_47.t5 Y.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR.t7 D.t6 Y.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 Y.t12 a_27_47.t6 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_633_47.t5 C.t4 a_991_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_633_47.t4 C.t5 a_991_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VPWR.t11 a_27_47.t7 Y.t13 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y.t7 D.t7 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR.t0 C.t6 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_215_47.t0 a_27_47.t8 Y.t14 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t15 a_27_47.t9 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR.t4 A_N.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X31 a_991_47.t0 C.t7 a_633_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 VPWR.t13 B.t7 Y.t16 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X33 VGND.t4 A_N.t1 a_27_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C.n0 C.t6 221.72
R1 C.n2 C.t1 221.72
R2 C.n7 C.t2 221.72
R3 C.n3 C.t3 221.72
R4 C.n4 C.n3 206.448
R5 C C.n1 163.201
R6 C.n9 C.n8 152
R7 C.n6 C.n5 152
R8 C.n0 C.t0 149.421
R9 C.n2 C.t5 149.421
R10 C.n7 C.t7 149.421
R11 C.n3 C.t4 149.421
R12 C.n2 C.n1 38.382
R13 C.n8 C.n2 37.4894
R14 C.n8 C.n7 37.4894
R15 C.n7 C.n6 37.4894
R16 C.n6 C.n3 37.4894
R17 C.n1 C.n0 36.5968
R18 C C.n4 16.9605
R19 C C.n9 16.0005
R20 C.n5 C 16.0005
R21 C.n9 C 13.4405
R22 C.n5 C 13.4405
R23 C.n4 C 12.4805
R24 a_633_47.n2 a_633_47.n0 224.822
R25 a_633_47.n4 a_633_47.n3 224.822
R26 a_633_47.n2 a_633_47.n1 185
R27 a_633_47.n5 a_633_47.n4 185
R28 a_633_47.n4 a_633_47.n2 64.4746
R29 a_633_47.n3 a_633_47.t1 24.9236
R30 a_633_47.n3 a_633_47.t7 24.9236
R31 a_633_47.n1 a_633_47.t3 24.9236
R32 a_633_47.n1 a_633_47.t5 24.9236
R33 a_633_47.n0 a_633_47.t6 24.9236
R34 a_633_47.n0 a_633_47.t4 24.9236
R35 a_633_47.n5 a_633_47.t2 24.9236
R36 a_633_47.t0 a_633_47.n5 24.9236
R37 a_991_47.n1 a_991_47.t2 319.277
R38 a_991_47.n1 a_991_47.n0 185
R39 a_991_47.n3 a_991_47.t7 176.972
R40 a_991_47.n3 a_991_47.n2 99.5638
R41 a_991_47.n5 a_991_47.n4 88.3446
R42 a_991_47.n4 a_991_47.n1 55.3569
R43 a_991_47.n4 a_991_47.n3 51.8339
R44 a_991_47.n0 a_991_47.t1 24.9236
R45 a_991_47.n0 a_991_47.t0 24.9236
R46 a_991_47.n2 a_991_47.t5 24.9236
R47 a_991_47.n2 a_991_47.t6 24.9236
R48 a_991_47.n5 a_991_47.t4 24.9236
R49 a_991_47.t3 a_991_47.n5 24.9236
R50 VNB.t2 VNB.t5 2677.02
R51 VNB.t8 VNB.t11 2677.02
R52 VNB.t10 VNB.t15 1196.12
R53 VNB.t14 VNB.t10 1196.12
R54 VNB.t9 VNB.t14 1196.12
R55 VNB.t6 VNB.t9 1196.12
R56 VNB.t4 VNB.t6 1196.12
R57 VNB.t3 VNB.t4 1196.12
R58 VNB.t5 VNB.t3 1196.12
R59 VNB.t0 VNB.t2 1196.12
R60 VNB.t1 VNB.t0 1196.12
R61 VNB.t7 VNB.t1 1196.12
R62 VNB.t13 VNB.t7 1196.12
R63 VNB.t12 VNB.t13 1196.12
R64 VNB.t16 VNB.t12 1196.12
R65 VNB.t11 VNB.t16 1196.12
R66 VNB VNB.t8 911.327
R67 B.n1 B.t7 240.695
R68 B.n0 B.t0 221.72
R69 B.n6 B.t2 221.72
R70 B.n7 B.t6 221.72
R71 B.n1 B.t5 168.394
R72 B.n1 B 159.361
R73 B.n3 B.n2 152
R74 B.n5 B.n4 152
R75 B.n9 B.n8 152
R76 B.n0 B.t3 149.421
R77 B.n6 B.t4 149.421
R78 B.n7 B.t1 149.421
R79 B.n8 B.n6 69.6227
R80 B.n5 B.n0 58.9116
R81 B.n2 B.n1 44.6301
R82 B.n3 B 18.2405
R83 B.n9 B 17.2805
R84 B.n2 B.n0 16.9598
R85 B.n6 B.n5 16.0672
R86 B.n4 B 16.0005
R87 B.n4 B 13.4405
R88 B B.n9 12.1605
R89 B B.n3 11.2005
R90 B.n8 B.n7 5.35606
R91 VPWR.n41 VPWR.n2 320.976
R92 VPWR.n35 VPWR.n34 320.976
R93 VPWR.n32 VPWR.n5 320.976
R94 VPWR.n10 VPWR.n9 320.976
R95 VPWR.n20 VPWR.n12 320.976
R96 VPWR.n15 VPWR.n14 320.976
R97 VPWR.n1 VPWR.t4 318.584
R98 VPWR.n16 VPWR.t5 255.091
R99 VPWR.n1 VPWR.t12 223.463
R100 VPWR.n27 VPWR.n8 139.048
R101 VPWR.n8 VPWR.t13 73.983
R102 VPWR.n8 VPWR.t1 73.9827
R103 VPWR.n16 VPWR.n15 39.0069
R104 VPWR.n31 VPWR.n6 34.6358
R105 VPWR.n36 VPWR.n33 34.6358
R106 VPWR.n40 VPWR.n3 34.6358
R107 VPWR.n19 VPWR.n13 34.6358
R108 VPWR.n22 VPWR.n21 34.6358
R109 VPWR.n26 VPWR.n25 34.6358
R110 VPWR.n42 VPWR.n41 32.377
R111 VPWR.n20 VPWR.n19 27.8593
R112 VPWR.n2 VPWR.t10 26.5955
R113 VPWR.n2 VPWR.t11 26.5955
R114 VPWR.n34 VPWR.t14 26.5955
R115 VPWR.n34 VPWR.t9 26.5955
R116 VPWR.n5 VPWR.t16 26.5955
R117 VPWR.n5 VPWR.t15 26.5955
R118 VPWR.n9 VPWR.t3 26.5955
R119 VPWR.n9 VPWR.t2 26.5955
R120 VPWR.n12 VPWR.t8 26.5955
R121 VPWR.n12 VPWR.t0 26.5955
R122 VPWR.n14 VPWR.t6 26.5955
R123 VPWR.n14 VPWR.t7 26.5955
R124 VPWR.n35 VPWR.n3 26.3534
R125 VPWR.n43 VPWR.n42 24.4711
R126 VPWR.n22 VPWR.n10 21.8358
R127 VPWR.n33 VPWR.n32 20.3299
R128 VPWR.n32 VPWR.n31 14.3064
R129 VPWR.n25 VPWR.n10 12.8005
R130 VPWR.n27 VPWR.n26 9.41227
R131 VPWR.n17 VPWR.n13 9.3005
R132 VPWR.n19 VPWR.n18 9.3005
R133 VPWR.n21 VPWR.n11 9.3005
R134 VPWR.n23 VPWR.n22 9.3005
R135 VPWR.n25 VPWR.n24 9.3005
R136 VPWR.n26 VPWR.n7 9.3005
R137 VPWR.n28 VPWR.n27 9.3005
R138 VPWR.n29 VPWR.n6 9.3005
R139 VPWR.n31 VPWR.n30 9.3005
R140 VPWR.n33 VPWR.n4 9.3005
R141 VPWR.n37 VPWR.n36 9.3005
R142 VPWR.n38 VPWR.n3 9.3005
R143 VPWR.n40 VPWR.n39 9.3005
R144 VPWR.n42 VPWR.n0 9.3005
R145 VPWR.n43 VPWR.n1 9.12056
R146 VPWR.n36 VPWR.n35 8.28285
R147 VPWR.n27 VPWR.n6 7.90638
R148 VPWR.n21 VPWR.n20 6.77697
R149 VPWR.n44 VPWR.n43 4.0883
R150 VPWR.n41 VPWR.n40 2.25932
R151 VPWR.n17 VPWR.n16 2.22239
R152 VPWR.n15 VPWR.n13 0.753441
R153 VPWR.n44 VPWR.n0 0.200784
R154 VPWR VPWR.n44 0.18088
R155 VPWR.n18 VPWR.n17 0.120292
R156 VPWR.n18 VPWR.n11 0.120292
R157 VPWR.n23 VPWR.n11 0.120292
R158 VPWR.n24 VPWR.n23 0.120292
R159 VPWR.n24 VPWR.n7 0.120292
R160 VPWR.n28 VPWR.n7 0.120292
R161 VPWR.n29 VPWR.n28 0.120292
R162 VPWR.n30 VPWR.n29 0.120292
R163 VPWR.n30 VPWR.n4 0.120292
R164 VPWR.n37 VPWR.n4 0.120292
R165 VPWR.n38 VPWR.n37 0.120292
R166 VPWR.n39 VPWR.n38 0.120292
R167 VPWR.n39 VPWR.n0 0.120292
R168 Y.n16 Y.n15 245.524
R169 Y.n5 Y.n3 235.923
R170 Y.n2 Y.n0 224.822
R171 Y.n5 Y.n4 206.25
R172 Y.n7 Y.n6 206.25
R173 Y.n9 Y.n8 206.25
R174 Y.n11 Y.n10 206.25
R175 Y.n13 Y.n12 206.25
R176 Y.n16 Y.n14 202.095
R177 Y.n2 Y.n1 185
R178 Y.n11 Y.n9 59.9278
R179 Y.n17 Y.n13 36.655
R180 Y.n7 Y.n5 29.6732
R181 Y.n9 Y.n7 29.6732
R182 Y.n13 Y.n11 29.6732
R183 Y.n14 Y.t11 26.5955
R184 Y.n14 Y.t12 26.5955
R185 Y.n15 Y.t13 26.5955
R186 Y.n15 Y.t15 26.5955
R187 Y.n3 Y.t4 26.5955
R188 Y.n3 Y.t5 26.5955
R189 Y.n4 Y.t6 26.5955
R190 Y.n4 Y.t7 26.5955
R191 Y.n6 Y.t0 26.5955
R192 Y.n6 Y.t3 26.5955
R193 Y.n8 Y.t2 26.5955
R194 Y.n8 Y.t1 26.5955
R195 Y.n10 Y.t16 26.5955
R196 Y.n10 Y.t19 26.5955
R197 Y.n12 Y.t18 26.5955
R198 Y.n12 Y.t17 26.5955
R199 Y.n0 Y.t14 24.9236
R200 Y.n0 Y.t8 24.9236
R201 Y.n1 Y.t10 24.9236
R202 Y.n1 Y.t9 24.9236
R203 Y Y.n17 16.4231
R204 Y.n18 Y 9.66088
R205 Y Y.n18 6.76276
R206 Y.n17 Y 2.03686
R207 Y.n18 Y 1.65976
R208 Y Y.n16 0.582318
R209 Y Y.n2 0.474574
R210 VPB.t13 VPB.t1 556.386
R211 VPB.t4 VPB.t12 556.386
R212 VPB.t6 VPB.t5 248.599
R213 VPB.t7 VPB.t6 248.599
R214 VPB.t8 VPB.t7 248.599
R215 VPB.t0 VPB.t8 248.599
R216 VPB.t3 VPB.t0 248.599
R217 VPB.t2 VPB.t3 248.599
R218 VPB.t1 VPB.t2 248.599
R219 VPB.t16 VPB.t13 248.599
R220 VPB.t15 VPB.t16 248.599
R221 VPB.t14 VPB.t15 248.599
R222 VPB.t9 VPB.t14 248.599
R223 VPB.t10 VPB.t9 248.599
R224 VPB.t11 VPB.t10 248.599
R225 VPB.t12 VPB.t11 248.599
R226 VPB VPB.t4 189.409
R227 D.n0 D.t5 221.72
R228 D.n6 D.t6 221.72
R229 D.n7 D.t7 221.72
R230 D.n1 D.t4 218.507
R231 D.n1 D 194.77
R232 D.n3 D.n2 152
R233 D.n5 D.n4 152
R234 D.n9 D.n8 152
R235 D.n0 D.t3 149.421
R236 D.n6 D.t0 149.421
R237 D.n7 D.t2 149.421
R238 D.n1 D.t1 146.208
R239 D.n2 D.n0 37.4894
R240 D.n5 D.n0 37.4894
R241 D.n6 D.n5 37.4894
R242 D.n8 D.n6 37.4894
R243 D.n8 D.n7 37.4894
R244 D.n2 D.n1 36.566
R245 D.n4 D 26.2405
R246 D.n3 D 25.9205
R247 D.n9 D 23.6805
R248 D D.n9 5.7605
R249 D.n4 D 3.2005
R250 D D.n3 0.6405
R251 VGND.n32 VGND.t4 287.534
R252 VGND.n10 VGND.n9 213.507
R253 VGND.n8 VGND.n7 207.213
R254 VGND.n10 VGND.n8 36.6918
R255 VGND.n13 VGND.n12 34.6358
R256 VGND.n14 VGND.n13 34.6358
R257 VGND.n14 VGND.n5 34.6358
R258 VGND.n18 VGND.n5 34.6358
R259 VGND.n19 VGND.n18 34.6358
R260 VGND.n20 VGND.n19 34.6358
R261 VGND.n20 VGND.n3 34.6358
R262 VGND.n24 VGND.n3 34.6358
R263 VGND.n25 VGND.n24 34.6358
R264 VGND.n26 VGND.n25 34.6358
R265 VGND.n26 VGND.n1 34.6358
R266 VGND.n30 VGND.n1 34.6358
R267 VGND.n31 VGND.n30 34.6358
R268 VGND.n9 VGND.t2 24.9236
R269 VGND.n9 VGND.t0 24.9236
R270 VGND.n7 VGND.t3 24.9236
R271 VGND.n7 VGND.t1 24.9236
R272 VGND.n32 VGND.n31 22.9652
R273 VGND.n12 VGND.n11 9.3005
R274 VGND.n13 VGND.n6 9.3005
R275 VGND.n15 VGND.n14 9.3005
R276 VGND.n16 VGND.n5 9.3005
R277 VGND.n18 VGND.n17 9.3005
R278 VGND.n19 VGND.n4 9.3005
R279 VGND.n21 VGND.n20 9.3005
R280 VGND.n22 VGND.n3 9.3005
R281 VGND.n24 VGND.n23 9.3005
R282 VGND.n25 VGND.n2 9.3005
R283 VGND.n27 VGND.n26 9.3005
R284 VGND.n28 VGND.n1 9.3005
R285 VGND.n30 VGND.n29 9.3005
R286 VGND.n31 VGND.n0 9.3005
R287 VGND.n33 VGND.n32 7.4049
R288 VGND.n12 VGND.n8 3.76521
R289 VGND.n11 VGND.n10 1.9288
R290 VGND.n33 VGND.n0 0.144904
R291 VGND.n11 VGND.n6 0.120292
R292 VGND.n15 VGND.n6 0.120292
R293 VGND.n16 VGND.n15 0.120292
R294 VGND.n17 VGND.n16 0.120292
R295 VGND.n17 VGND.n4 0.120292
R296 VGND.n21 VGND.n4 0.120292
R297 VGND.n22 VGND.n21 0.120292
R298 VGND.n23 VGND.n22 0.120292
R299 VGND.n23 VGND.n2 0.120292
R300 VGND.n27 VGND.n2 0.120292
R301 VGND.n28 VGND.n27 0.120292
R302 VGND.n29 VGND.n28 0.120292
R303 VGND.n29 VGND.n0 0.120292
R304 VGND VGND.n33 0.117202
R305 a_27_47.t0 a_27_47.n8 265.675
R306 a_27_47.n1 a_27_47.t5 221.72
R307 a_27_47.n2 a_27_47.t6 221.72
R308 a_27_47.n4 a_27_47.t7 221.72
R309 a_27_47.n6 a_27_47.t9 221.72
R310 a_27_47.n7 a_27_47.n6 194.845
R311 a_27_47.n3 a_27_47.n0 178.881
R312 a_27_47.n8 a_27_47.t1 169.24
R313 a_27_47.n5 a_27_47.n0 152
R314 a_27_47.n1 a_27_47.t4 149.421
R315 a_27_47.n2 a_27_47.t3 149.421
R316 a_27_47.n4 a_27_47.t8 149.421
R317 a_27_47.n6 a_27_47.t2 149.421
R318 a_27_47.n2 a_27_47.n1 74.9783
R319 a_27_47.n3 a_27_47.n2 37.4894
R320 a_27_47.n4 a_27_47.n3 37.4894
R321 a_27_47.n5 a_27_47.n4 37.4894
R322 a_27_47.n6 a_27_47.n5 37.4894
R323 a_27_47.n8 a_27_47.n7 29.7605
R324 a_27_47.n7 a_27_47.n0 28.8005
R325 a_215_47.n1 a_215_47.t4 319.277
R326 a_215_47.n1 a_215_47.n0 185
R327 a_215_47.n3 a_215_47.n2 185
R328 a_215_47.n5 a_215_47.n4 185
R329 a_215_47.t3 a_215_47.n5 183.096
R330 a_215_47.n3 a_215_47.n1 51.2005
R331 a_215_47.n5 a_215_47.n3 51.2005
R332 a_215_47.n4 a_215_47.t2 24.9236
R333 a_215_47.n4 a_215_47.t0 24.9236
R334 a_215_47.n2 a_215_47.t7 24.9236
R335 a_215_47.n2 a_215_47.t1 24.9236
R336 a_215_47.n0 a_215_47.t6 24.9236
R337 a_215_47.n0 a_215_47.t5 24.9236
R338 A_N.n0 A_N.t0 233.989
R339 A_N.n0 A_N.t1 161.69
R340 A_N A_N.n0 160
C0 VPB C 0.13951f
C1 VPB VPWR 0.186918f
C2 VPB Y 0.033677f
C3 A_N VPWR 0.017587f
C4 B C 0.045994f
C5 B VPWR 0.055484f
C6 C D 0.060585f
C7 VPB VGND 0.012266f
C8 D VPWR 0.098527f
C9 B Y 0.23982f
C10 C VPWR 0.058942f
C11 A_N VGND 0.015275f
C12 D Y 0.175245f
C13 B VGND 0.031291f
C14 C Y 0.231566f
C15 VPWR Y 1.54678f
C16 D VGND 0.061578f
C17 C VGND 0.033908f
C18 VPWR VGND 0.175807f
C19 Y VGND 0.039329f
C20 VPB A_N 0.042776f
C21 VPB B 0.131586f
C22 VPB D 0.136371f
C23 VGND VNB 0.944727f
C24 Y VNB 0.017884f
C25 VPWR VNB 0.82419f
C26 D VNB 0.422179f
C27 C VNB 0.397228f
C28 B VNB 0.381201f
C29 A_N VNB 0.147468f
C30 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4bb_1 VNB VPB VPWR VGND A_N Y C D B_N
X0 VGND.t0 B_N.t0 a_27_93.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_496_21.t0 A_N.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1827 pd=1.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 Y.t1 a_496_21.t2 a_426_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X3 VPWR.t5 a_496_21.t3 Y.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_426_47.t1 a_27_93.t2 a_326_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11375 ps=1 w=0.65 l=0.15
X5 VPWR.t0 B_N.t1 a_27_93.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 a_496_21.t1 A_N.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1827 pd=1.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y.t2 a_27_93.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X8 a_218_47.t0 D.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11975 ps=1.045 w=0.65 l=0.15
X9 a_326_47.t1 C.t0 a_218_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.12675 ps=1.04 w=0.65 l=0.15
X10 Y.t3 D.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.17575 ps=1.395 w=1 l=0.15
X11 VPWR.t4 C.t1 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.195 ps=1.39 w=1 l=0.15
R0 B_N.n0 B_N.t1 329.007
R1 B_N B_N.n0 154.012
R2 B_N.n0 B_N.t0 126.567
R3 a_27_93.n1 a_27_93.t1 747.097
R4 a_27_93.n1 a_27_93.n0 298.863
R5 a_27_93.n0 a_27_93.t3 241.536
R6 a_27_93.t0 a_27_93.n1 231.101
R7 a_27_93.n0 a_27_93.t2 169.237
R8 VGND.n1 VGND.t2 243.274
R9 VGND.n1 VGND.n0 224.964
R10 VGND.n0 VGND.t0 67.1434
R11 VGND.n0 VGND.t1 29.539
R12 VGND VGND.n1 0.15698
R13 VNB.t5 VNB.t3 2677.02
R14 VNB.t0 VNB.t1 1552.1
R15 VNB.t1 VNB.t4 1537.86
R16 VNB.t2 VNB.t5 1423.95
R17 VNB.t4 VNB.t2 1423.95
R18 VNB VNB.t0 925.567
R19 A_N.n0 A_N.t0 336.329
R20 A_N.n0 A_N.t1 204.583
R21 A_N.n1 A_N.n0 152
R22 A_N.n1 A_N 14.8485
R23 A_N A_N.n1 2.5605
R24 VPWR.n6 VPWR.t5 853.981
R25 VPWR.n5 VPWR.t1 650.85
R26 VPWR.n13 VPWR.n1 310.574
R27 VPWR.n3 VPWR.n2 310.502
R28 VPWR.n1 VPWR.t0 105.41
R29 VPWR.n1 VPWR.t3 36.2649
R30 VPWR.n12 VPWR.n11 34.6358
R31 VPWR.n8 VPWR.n7 34.6358
R32 VPWR.n2 VPWR.t2 34.4755
R33 VPWR.n2 VPWR.t4 34.4755
R34 VPWR.n13 VPWR.n12 16.9417
R35 VPWR.n7 VPWR.n6 13.0216
R36 VPWR.n7 VPWR.n4 9.3005
R37 VPWR.n9 VPWR.n8 9.3005
R38 VPWR.n11 VPWR.n10 9.3005
R39 VPWR.n12 VPWR.n0 9.3005
R40 VPWR.n8 VPWR.n3 7.52991
R41 VPWR.n14 VPWR.n13 7.4049
R42 VPWR.n6 VPWR.n5 6.68025
R43 VPWR.n5 VPWR.n4 4.04238
R44 VPWR.n11 VPWR.n3 2.25932
R45 VPWR.n14 VPWR.n0 0.144904
R46 VPWR.n9 VPWR.n4 0.120292
R47 VPWR.n10 VPWR.n9 0.120292
R48 VPWR.n10 VPWR.n0 0.120292
R49 VPWR VPWR.n14 0.118504
R50 a_496_21.t0 a_496_21.n1 705.682
R51 a_496_21.n1 a_496_21.t1 325.557
R52 a_496_21.n1 a_496_21.n0 285.99
R53 a_496_21.n0 a_496_21.t3 212.081
R54 a_496_21.n0 a_496_21.t2 139.78
R55 VPB.t2 VPB.t1 556.386
R56 VPB.t0 VPB.t4 322.587
R57 VPB.t4 VPB.t5 319.627
R58 VPB.t3 VPB.t2 295.95
R59 VPB.t5 VPB.t3 295.95
R60 VPB VPB.t0 192.369
R61 a_426_47.t0 a_426_47.t1 64.6159
R62 Y.n2 Y.n1 269.658
R63 Y.n2 Y.n0 202.095
R64 Y.n4 Y.t1 130.138
R65 Y.n1 Y.t4 38.4155
R66 Y.n1 Y.t3 38.4155
R67 Y.n0 Y.t0 34.4755
R68 Y.n0 Y.t2 34.4755
R69 Y.n3 Y 14.3365
R70 Y Y.n2 10.9181
R71 Y.n4 Y 4.70956
R72 Y Y.n4 3.7234
R73 Y.n3 Y 3.0725
R74 Y Y.n3 1.50638
R75 a_326_47.t0 a_326_47.t1 64.6159
R76 D.n0 D.t1 236.18
R77 D.n0 D.t0 163.881
R78 D D.n0 155.328
R79 a_218_47.t0 a_218_47.t1 72.0005
R80 C.n0 C.t1 239.505
R81 C.n0 C.t0 167.204
R82 C C.n0 154.279
C0 A_N VPWR 0.015524f
C1 C Y 0.037671f
C2 D VGND 0.017182f
C3 VPWR VGND 0.082326f
C4 C A_N 7.91e-20
C5 C VGND 0.010604f
C6 A_N Y 0.013903f
C7 Y VGND 0.101326f
C8 A_N VGND 0.02761f
C9 VPB B_N 0.096045f
C10 VPB D 0.032085f
C11 VPB VPWR 0.093109f
C12 B_N D 0.064876f
C13 VPB C 0.029076f
C14 B_N VPWR 0.04603f
C15 VPB Y 0.011404f
C16 B_N C 0.001096f
C17 VPB A_N 0.09848f
C18 B_N Y 0.015056f
C19 D VPWR 0.02438f
C20 VPB VGND 0.011577f
C21 B_N A_N 0.003275f
C22 D C 0.06895f
C23 C VPWR 0.01849f
C24 D Y 0.028097f
C25 B_N VGND 0.012328f
C26 VPWR Y 0.330453f
C27 VGND VNB 0.507586f
C28 Y VNB 0.014283f
C29 VPWR VNB 0.407232f
C30 A_N VNB 0.167615f
C31 C VNB 0.094697f
C32 D VNB 0.100764f
C33 B_N VNB 0.142346f
C34 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4bb_2 VNB VPB VGND VPWR A_N B_N Y C D
X0 VPWR.t1 a_193_47.t2 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t4 D.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t7 C.t0 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 D.t1 a_781_47.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t1 a_193_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 Y.t8 C.t1 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6 a_591_47.t3 C.t2 a_781_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_781_47.t0 C.t3 a_591_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t5 B_N.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_193_47.t0 A_N.t0 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1974 pd=1.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 Y.t0 a_193_47.t4 a_341_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_591_47.t0 a_27_47.t2 a_341_47.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_341_47.t0 a_193_47.t5 Y.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_341_47.t2 a_27_47.t3 a_591_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR.t3 a_27_47.t4 Y.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X16 Y.t6 a_27_47.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_193_47.t1 A_N.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1974 pd=1.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VGND.t1 B_N.t1 a_27_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_193_47.n2 a_193_47.t1 735.87
R1 a_193_47.t0 a_193_47.n2 282.711
R2 a_193_47.n2 a_193_47.n1 231.603
R3 a_193_47.n0 a_193_47.t2 221.72
R4 a_193_47.n1 a_193_47.t3 212.081
R5 a_193_47.n0 a_193_47.t5 149.421
R6 a_193_47.n1 a_193_47.t4 139.78
R7 a_193_47.n1 a_193_47.n0 72.5439
R8 Y.n6 Y.n4 309.358
R9 Y.n1 Y.t4 262.517
R10 Y.n6 Y.n5 216.613
R11 Y.n1 Y.n0 206.25
R12 Y.n7 Y.n3 202.095
R13 Y.n2 Y.n1 51.7823
R14 Y.n7 Y.n6 39.2732
R15 Y.n3 Y.t5 26.5955
R16 Y.n3 Y.t6 26.5955
R17 Y.n4 Y.t2 26.5955
R18 Y.n4 Y.t1 26.5955
R19 Y.n0 Y.t7 26.5955
R20 Y.n0 Y.t8 26.5955
R21 Y.n5 Y.t3 24.9236
R22 Y.n5 Y.t0 24.9236
R23 Y Y.n7 16.0005
R24 Y.n2 Y 14.2694
R25 Y Y.n2 1.74595
R26 VPWR.n17 VPWR.n1 605.481
R27 VPWR.n8 VPWR.n7 329.356
R28 VPWR.n11 VPWR.n4 316.245
R29 VPWR.n2 VPWR.t0 257.474
R30 VPWR.n6 VPWR.n5 139.048
R31 VPWR.n5 VPWR.t3 73.983
R32 VPWR.n5 VPWR.t8 73.9827
R33 VPWR.n1 VPWR.t6 63.3219
R34 VPWR.n1 VPWR.t5 63.3219
R35 VPWR.n16 VPWR.n15 34.6358
R36 VPWR.n12 VPWR.n11 32.7534
R37 VPWR.n10 VPWR.n6 32.7534
R38 VPWR.n17 VPWR.n16 28.9887
R39 VPWR.n4 VPWR.t4 26.5955
R40 VPWR.n4 VPWR.t1 26.5955
R41 VPWR.n7 VPWR.t2 26.5955
R42 VPWR.n7 VPWR.t7 26.5955
R43 VPWR.n12 VPWR.n2 18.0711
R44 VPWR.n11 VPWR.n10 17.6946
R45 VPWR.n15 VPWR.n2 16.5652
R46 VPWR.n10 VPWR.n9 9.3005
R47 VPWR.n11 VPWR.n3 9.3005
R48 VPWR.n13 VPWR.n12 9.3005
R49 VPWR.n15 VPWR.n14 9.3005
R50 VPWR.n16 VPWR.n0 9.3005
R51 VPWR.n18 VPWR.n17 7.21821
R52 VPWR.n8 VPWR.n6 3.73121
R53 VPWR.n9 VPWR.n8 0.396258
R54 VPWR.n18 VPWR.n0 0.147279
R55 VPWR.n9 VPWR.n3 0.120292
R56 VPWR.n13 VPWR.n3 0.120292
R57 VPWR.n14 VPWR.n13 0.120292
R58 VPWR.n14 VPWR.n0 0.120292
R59 VPWR VPWR.n18 0.116099
R60 VPB.t6 VPB.t0 680.686
R61 VPB.t3 VPB.t8 556.386
R62 VPB.t7 VPB.t2 248.599
R63 VPB.t8 VPB.t7 248.599
R64 VPB.t4 VPB.t3 248.599
R65 VPB.t1 VPB.t4 248.599
R66 VPB.t0 VPB.t1 248.599
R67 VPB.t5 VPB.t6 248.599
R68 VPB VPB.t5 192.369
R69 D.n2 D.n0 234.038
R70 D.n3 D.t0 221.72
R71 D.n2 D.n1 161.738
R72 D D.n4 159.361
R73 D.n2 D 153.601
R74 D.n3 D.t1 149.421
R75 D.n4 D.n2 56.2338
R76 D.n4 D.n3 5.35606
R77 C.n0 C.t0 221.72
R78 C.n2 C.t1 221.72
R79 C.n3 C.n2 194.845
R80 C C.n1 161.28
R81 C.n0 C.t3 149.421
R82 C.n2 C.t2 149.421
R83 C.n1 C.n0 37.4894
R84 C.n2 C.n1 37.4894
R85 C C.n3 19.5205
R86 C.n3 C 9.9205
R87 a_781_47.n0 a_781_47.t1 399.058
R88 a_781_47.n0 a_781_47.t2 24.9236
R89 a_781_47.t0 a_781_47.n0 24.9236
R90 VGND.n1 VGND.t2 287.488
R91 VGND.n1 VGND.n0 210.393
R92 VGND.n0 VGND.t0 38.5719
R93 VGND.n0 VGND.t1 38.5719
R94 VGND VGND.n1 0.143722
R95 VNB.t4 VNB.t1 3275.08
R96 VNB.t3 VNB.t7 2677.02
R97 VNB.t6 VNB.t8 1196.12
R98 VNB.t7 VNB.t6 1196.12
R99 VNB.t2 VNB.t3 1196.12
R100 VNB.t0 VNB.t2 1196.12
R101 VNB.t1 VNB.t0 1196.12
R102 VNB.t5 VNB.t4 1196.12
R103 VNB VNB.t5 925.567
R104 a_591_47.n1 a_591_47.n0 439.632
R105 a_591_47.n0 a_591_47.t1 24.9236
R106 a_591_47.n0 a_591_47.t0 24.9236
R107 a_591_47.t2 a_591_47.n1 24.9236
R108 a_591_47.n1 a_591_47.t3 24.9236
R109 B_N.n0 B_N.t0 314.908
R110 B_N.n0 B_N.t1 234.573
R111 B_N.n1 B_N.n0 152
R112 B_N.n1 B_N 10.9719
R113 B_N B_N.n1 6.79234
R114 a_27_47.n3 a_27_47.t1 761.735
R115 a_27_47.t0 a_27_47.n3 323.12
R116 a_27_47.n0 a_27_47.t4 221.72
R117 a_27_47.n1 a_27_47.t5 221.72
R118 a_27_47.n3 a_27_47.n2 176.724
R119 a_27_47.n0 a_27_47.t3 149.421
R120 a_27_47.n1 a_27_47.t2 149.421
R121 a_27_47.n2 a_27_47.n0 69.6227
R122 a_27_47.n2 a_27_47.n1 5.35606
R123 A_N.n0 A_N.t1 295.949
R124 A_N.n0 A_N.t0 228.469
R125 A_N.n1 A_N.n0 152
R126 A_N.n1 A_N 8.68621
R127 A_N A_N.n1 6.85764
R128 a_341_47.n1 a_341_47.t2 305.594
R129 a_341_47.t1 a_341_47.n1 296.363
R130 a_341_47.n1 a_341_47.n0 185
R131 a_341_47.n0 a_341_47.t3 24.9236
R132 a_341_47.n0 a_341_47.t0 24.9236
C0 VPB Y 0.021819f
C1 VPB D 0.072712f
C2 VPB VGND 0.007695f
C3 VPB VPWR 0.133193f
C4 B_N VGND 0.016979f
C5 A_N Y 0.002125f
C6 B_N VPWR 0.016943f
C7 A_N VGND 0.016111f
C8 C Y 0.138971f
C9 C D 0.06757f
C10 A_N VPWR 0.017103f
C11 C VGND 0.019663f
C12 D Y 0.076756f
C13 C VPWR 0.037317f
C14 Y VGND 0.014344f
C15 D VGND 0.030555f
C16 VPWR Y 0.81164f
C17 D VPWR 0.064289f
C18 VPWR VGND 0.080327f
C19 VPB B_N 0.086836f
C20 VPB A_N 0.09531f
C21 VPB C 0.072699f
C22 B_N A_N 0.128745f
C23 VGND VNB 0.672214f
C24 Y VNB 0.021433f
C25 VPWR VNB 0.593314f
C26 D VNB 0.239265f
C27 C VNB 0.209309f
C28 A_N VNB 0.128579f
C29 B_N VNB 0.196942f
C30 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4bb_4 VNB VPB VGND VPWR C Y A_N B_N D
X0 Y.t9 a_27_47.t2 a_432_47.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y.t5 a_27_47.t3 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t8 a_27_47.t4 a_432_47.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t16 C.t0 Y.t18 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_850_47.t7 a_193_47.t2 a_432_47.t4 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t4 D.t0 a_1266_47.t5 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t5 a_27_47.t5 Y.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t13 C.t1 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.555 ps=2.11 w=1 l=0.15
X8 Y.t3 a_27_47.t6 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VPWR.t7 D.t1 Y.t10 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X10 a_432_47.t1 a_27_47.t7 Y.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_432_47.t5 a_193_47.t3 a_850_47.t6 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_432_47.t0 a_27_47.t8 Y.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_432_47.t6 a_193_47.t4 a_850_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t11 D.t2 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t11 a_193_47.t5 Y.t14 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.555 pd=2.11 as=0.135 ps=1.27 w=1 l=0.15
X16 a_193_47.t1 B_N.t0 VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.495 pd=2.99 as=0.135 ps=1.27 w=1 l=0.15
X17 Y.t15 a_193_47.t6 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR.t9 D.t3 Y.t12 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_193_47.t0 B_N.t1 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.32175 pd=2.29 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y.t19 D.t4 VPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_850_47.t1 C.t2 a_1266_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1885 ps=1.88 w=0.65 l=0.15
X22 a_850_47.t4 a_193_47.t7 a_432_47.t7 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_850_47.t2 C.t3 a_1266_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VPWR.t2 C.t4 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND.t3 D.t5 a_1266_47.t4 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y.t0 C.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR.t13 a_193_47.t8 Y.t16 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1266_47.t1 C.t6 a_850_47.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t17 a_193_47.t9 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_1266_47.t0 C.t7 a_850_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_1266_47.t7 D.t6 VGND.t2 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_1266_47.t6 D.t7 VGND.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VPWR.t1 A_N.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 VPWR.t3 a_27_47.t9 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 VGND.t0 A_N.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t0 a_27_47.n5 903.072
R1 a_27_47.n5 a_27_47.n4 316.318
R2 a_27_47.n5 a_27_47.t1 301.127
R3 a_27_47.n1 a_27_47.t9 221.72
R4 a_27_47.n2 a_27_47.t3 221.72
R5 a_27_47.n0 a_27_47.t5 221.72
R6 a_27_47.n4 a_27_47.t6 212.081
R7 a_27_47.n1 a_27_47.t8 149.421
R8 a_27_47.n2 a_27_47.t4 149.421
R9 a_27_47.n0 a_27_47.t7 149.421
R10 a_27_47.n4 a_27_47.t2 139.78
R11 a_27_47.n2 a_27_47.n1 74.9783
R12 a_27_47.n3 a_27_47.n2 68.3552
R13 a_27_47.n4 a_27_47.n3 65.7593
R14 a_27_47.n3 a_27_47.n0 3.35269
R15 a_432_47.n3 a_432_47.t3 334.026
R16 a_432_47.n1 a_432_47.t5 305.594
R17 a_432_47.n1 a_432_47.n0 185
R18 a_432_47.n3 a_432_47.n2 185
R19 a_432_47.n5 a_432_47.n4 185
R20 a_432_47.n4 a_432_47.n1 46.7483
R21 a_432_47.n4 a_432_47.n3 46.7483
R22 a_432_47.n2 a_432_47.t2 24.9236
R23 a_432_47.n2 a_432_47.t1 24.9236
R24 a_432_47.n0 a_432_47.t7 24.9236
R25 a_432_47.n0 a_432_47.t6 24.9236
R26 a_432_47.n5 a_432_47.t4 24.9236
R27 a_432_47.t0 a_432_47.n5 24.9236
R28 Y.n16 Y.n15 354.651
R29 Y.n5 Y.n3 235.923
R30 Y.n2 Y.n0 228.008
R31 Y.n5 Y.n4 206.25
R32 Y.n7 Y.n6 206.25
R33 Y.n9 Y.n8 206.25
R34 Y.n11 Y.n10 206.25
R35 Y.n13 Y.n12 206.25
R36 Y.n16 Y.n14 202.095
R37 Y.n2 Y.n1 185
R38 Y.n11 Y.n9 78.546
R39 Y.n7 Y.n5 29.6732
R40 Y.n9 Y.n7 29.6732
R41 Y.n13 Y.n11 29.6732
R42 Y.n18 Y.n17 29.3522
R43 Y.n14 Y.t2 26.5955
R44 Y.n14 Y.t5 26.5955
R45 Y.n15 Y.t4 26.5955
R46 Y.n15 Y.t3 26.5955
R47 Y.n3 Y.t10 26.5955
R48 Y.n3 Y.t11 26.5955
R49 Y.n4 Y.t12 26.5955
R50 Y.n4 Y.t19 26.5955
R51 Y.n6 Y.t1 26.5955
R52 Y.n6 Y.t0 26.5955
R53 Y.n8 Y.t18 26.5955
R54 Y.n8 Y.t13 26.5955
R55 Y.n10 Y.t14 26.5955
R56 Y.n10 Y.t15 26.5955
R57 Y.n12 Y.t16 26.5955
R58 Y.n12 Y.t17 26.5955
R59 Y.n0 Y.t7 24.9236
R60 Y.n0 Y.t9 24.9236
R61 Y.n1 Y.t6 24.9236
R62 Y.n1 Y.t8 24.9236
R63 Y.n17 Y.n13 21.8187
R64 Y Y.n16 16.0005
R65 Y.n18 Y.n2 7.9365
R66 Y.n17 Y 1.45505
R67 Y Y.n18 0.662569
R68 VNB.t6 VNB.t10 4570.87
R69 VNB.t12 VNB.t4 3588.35
R70 VNB.t3 VNB.t17 1196.12
R71 VNB.t16 VNB.t3 1196.12
R72 VNB.t15 VNB.t16 1196.12
R73 VNB.t1 VNB.t15 1196.12
R74 VNB.t5 VNB.t1 1196.12
R75 VNB.t0 VNB.t5 1196.12
R76 VNB.t4 VNB.t0 1196.12
R77 VNB.t14 VNB.t12 1196.12
R78 VNB.t13 VNB.t14 1196.12
R79 VNB.t11 VNB.t13 1196.12
R80 VNB.t7 VNB.t11 1196.12
R81 VNB.t9 VNB.t7 1196.12
R82 VNB.t8 VNB.t9 1196.12
R83 VNB.t10 VNB.t8 1196.12
R84 VNB.t2 VNB.t6 1196.12
R85 VNB VNB.t2 925.567
R86 VPWR.n56 VPWR.n1 605.481
R87 VPWR.n42 VPWR.n41 320.976
R88 VPWR.n40 VPWR.n7 320.976
R89 VPWR.n24 VPWR.n23 320.976
R90 VPWR.n21 VPWR.n13 320.976
R91 VPWR.n16 VPWR.n15 320.976
R92 VPWR.n48 VPWR.n4 316.245
R93 VPWR.n32 VPWR.n8 292.5
R94 VPWR.n34 VPWR.n33 292.5
R95 VPWR.n31 VPWR.n30 292.5
R96 VPWR.n49 VPWR.t4 257.474
R97 VPWR.n17 VPWR.t7 253.232
R98 VPWR.n33 VPWR.n31 81.7555
R99 VPWR.n33 VPWR.n32 67.9655
R100 VPWR.n17 VPWR.n16 37.305
R101 VPWR.n32 VPWR.t11 36.4455
R102 VPWR.n54 VPWR.n2 34.6358
R103 VPWR.n55 VPWR.n54 34.6358
R104 VPWR.n39 VPWR.n38 34.6358
R105 VPWR.n47 VPWR.n5 34.6358
R106 VPWR.n20 VPWR.n14 34.6358
R107 VPWR.n25 VPWR.n22 34.6358
R108 VPWR.n29 VPWR.n11 34.6358
R109 VPWR.n43 VPWR.n40 32.7534
R110 VPWR.n31 VPWR.t10 32.5055
R111 VPWR.n50 VPWR.n48 32.377
R112 VPWR.n43 VPWR.n42 30.4946
R113 VPWR.n56 VPWR.n55 28.9887
R114 VPWR.n1 VPWR.t15 26.5955
R115 VPWR.n1 VPWR.t1 26.5955
R116 VPWR.n4 VPWR.t6 26.5955
R117 VPWR.n4 VPWR.t5 26.5955
R118 VPWR.n41 VPWR.t14 26.5955
R119 VPWR.n41 VPWR.t3 26.5955
R120 VPWR.n7 VPWR.t12 26.5955
R121 VPWR.n7 VPWR.t13 26.5955
R122 VPWR.n23 VPWR.t0 26.5955
R123 VPWR.n23 VPWR.t16 26.5955
R124 VPWR.n13 VPWR.t17 26.5955
R125 VPWR.n13 VPWR.t2 26.5955
R126 VPWR.n15 VPWR.t8 26.5955
R127 VPWR.n15 VPWR.t9 26.5955
R128 VPWR.n21 VPWR.n20 25.977
R129 VPWR.n38 VPWR.n8 25.2163
R130 VPWR.n25 VPWR.n24 19.9534
R131 VPWR.n50 VPWR.n49 18.4476
R132 VPWR.n48 VPWR.n47 18.0711
R133 VPWR.n49 VPWR.n2 16.1887
R134 VPWR.n24 VPWR.n11 14.6829
R135 VPWR.n30 VPWR.n29 10.9104
R136 VPWR.n18 VPWR.n14 9.3005
R137 VPWR.n20 VPWR.n19 9.3005
R138 VPWR.n22 VPWR.n12 9.3005
R139 VPWR.n26 VPWR.n25 9.3005
R140 VPWR.n27 VPWR.n11 9.3005
R141 VPWR.n29 VPWR.n28 9.3005
R142 VPWR.n10 VPWR.n9 9.3005
R143 VPWR.n36 VPWR.n35 9.3005
R144 VPWR.n38 VPWR.n37 9.3005
R145 VPWR.n39 VPWR.n6 9.3005
R146 VPWR.n44 VPWR.n43 9.3005
R147 VPWR.n45 VPWR.n5 9.3005
R148 VPWR.n47 VPWR.n46 9.3005
R149 VPWR.n48 VPWR.n3 9.3005
R150 VPWR.n51 VPWR.n50 9.3005
R151 VPWR.n52 VPWR.n2 9.3005
R152 VPWR.n54 VPWR.n53 9.3005
R153 VPWR.n55 VPWR.n0 9.3005
R154 VPWR.n22 VPWR.n21 8.65932
R155 VPWR.n57 VPWR.n56 7.21821
R156 VPWR.n42 VPWR.n5 4.14168
R157 VPWR.n35 VPWR.n34 3.8273
R158 VPWR.n30 VPWR.n10 3.23349
R159 VPWR.n16 VPWR.n14 2.63579
R160 VPWR.n34 VPWR.n10 2.2438
R161 VPWR.n18 VPWR.n17 2.13159
R162 VPWR.n40 VPWR.n39 1.88285
R163 VPWR.n35 VPWR.n8 0.726273
R164 VPWR.n57 VPWR.n0 0.147279
R165 VPWR.n19 VPWR.n18 0.120292
R166 VPWR.n19 VPWR.n12 0.120292
R167 VPWR.n26 VPWR.n12 0.120292
R168 VPWR.n27 VPWR.n26 0.120292
R169 VPWR.n28 VPWR.n27 0.120292
R170 VPWR.n28 VPWR.n9 0.120292
R171 VPWR.n36 VPWR.n9 0.120292
R172 VPWR.n37 VPWR.n36 0.120292
R173 VPWR.n37 VPWR.n6 0.120292
R174 VPWR.n44 VPWR.n6 0.120292
R175 VPWR.n45 VPWR.n44 0.120292
R176 VPWR.n46 VPWR.n45 0.120292
R177 VPWR.n46 VPWR.n3 0.120292
R178 VPWR.n51 VPWR.n3 0.120292
R179 VPWR.n52 VPWR.n51 0.120292
R180 VPWR.n53 VPWR.n52 0.120292
R181 VPWR.n53 VPWR.n0 0.120292
R182 VPWR VPWR.n57 0.116099
R183 VPB.t15 VPB.t4 950
R184 VPB.t11 VPB.t10 745.794
R185 VPB.t8 VPB.t7 248.599
R186 VPB.t9 VPB.t8 248.599
R187 VPB.t17 VPB.t9 248.599
R188 VPB.t2 VPB.t17 248.599
R189 VPB.t0 VPB.t2 248.599
R190 VPB.t16 VPB.t0 248.599
R191 VPB.t10 VPB.t16 248.599
R192 VPB.t12 VPB.t11 248.599
R193 VPB.t13 VPB.t12 248.599
R194 VPB.t14 VPB.t13 248.599
R195 VPB.t3 VPB.t14 248.599
R196 VPB.t6 VPB.t3 248.599
R197 VPB.t5 VPB.t6 248.599
R198 VPB.t4 VPB.t5 248.599
R199 VPB.t1 VPB.t15 248.599
R200 VPB VPB.t1 192.369
R201 C.n0 C.t4 221.72
R202 C.n2 C.t5 221.72
R203 C.n7 C.t0 221.72
R204 C.n3 C.t1 221.72
R205 C.n4 C.n3 194.845
R206 C C.n1 167.68
R207 C.n9 C.n8 152
R208 C.n6 C.n5 152
R209 C.n0 C.t7 149.421
R210 C.n2 C.t3 149.421
R211 C.n7 C.t6 149.421
R212 C.n3 C.t2 149.421
R213 C.n1 C.n0 37.4894
R214 C.n2 C.n1 37.4894
R215 C.n8 C.n2 37.4894
R216 C.n8 C.n7 37.4894
R217 C.n7 C.n6 37.4894
R218 C.n6 C.n3 37.4894
R219 C.n4 C 21.4405
R220 C.n5 C 20.8005
R221 C.n9 C 18.2405
R222 C C.n9 11.2005
R223 C.n5 C 8.6405
R224 C C.n4 8.0005
R225 a_193_47.t1 a_193_47.n9 810.715
R226 a_193_47.n9 a_193_47.t0 302.928
R227 a_193_47.n1 a_193_47.t5 221.72
R228 a_193_47.n3 a_193_47.t6 221.72
R229 a_193_47.n5 a_193_47.t8 221.72
R230 a_193_47.n6 a_193_47.t9 221.72
R231 a_193_47.n2 a_193_47.n0 179.201
R232 a_193_47.n8 a_193_47.n7 152
R233 a_193_47.n4 a_193_47.n0 152
R234 a_193_47.n1 a_193_47.t3 149.421
R235 a_193_47.n3 a_193_47.t7 149.421
R236 a_193_47.n5 a_193_47.t4 149.421
R237 a_193_47.n6 a_193_47.t2 149.421
R238 a_193_47.n9 a_193_47.n8 41.9093
R239 a_193_47.n4 a_193_47.n3 38.382
R240 a_193_47.n7 a_193_47.n6 38.382
R241 a_193_47.n2 a_193_47.n1 37.4894
R242 a_193_47.n3 a_193_47.n2 37.4894
R243 a_193_47.n5 a_193_47.n4 36.5968
R244 a_193_47.n7 a_193_47.n5 36.5968
R245 a_193_47.n8 a_193_47.n0 26.2405
R246 a_850_47.n2 a_850_47.n0 231.749
R247 a_850_47.n4 a_850_47.n3 228.008
R248 a_850_47.n2 a_850_47.n1 185
R249 a_850_47.n5 a_850_47.n4 185
R250 a_850_47.n4 a_850_47.n2 124.844
R251 a_850_47.n3 a_850_47.t5 24.9236
R252 a_850_47.n3 a_850_47.t7 24.9236
R253 a_850_47.n1 a_850_47.t3 24.9236
R254 a_850_47.n1 a_850_47.t1 24.9236
R255 a_850_47.n0 a_850_47.t0 24.9236
R256 a_850_47.n0 a_850_47.t2 24.9236
R257 a_850_47.t6 a_850_47.n5 24.9236
R258 a_850_47.n5 a_850_47.t4 24.9236
R259 D.n1 D.t1 233.868
R260 D.n4 D.t2 221.72
R261 D.n6 D.t3 221.72
R262 D.n7 D.t4 221.72
R263 D.n1 D.t7 161.567
R264 D D.n1 154.881
R265 D.n3 D.n2 152
R266 D.n5 D.n0 152
R267 D.n9 D.n8 152
R268 D.n4 D.t0 149.421
R269 D.n6 D.t6 149.421
R270 D.n7 D.t5 149.421
R271 D.n4 D.n3 37.4894
R272 D.n5 D.n4 37.4894
R273 D.n6 D.n5 37.4894
R274 D.n8 D.n6 37.4894
R275 D.n8 D.n7 37.4894
R276 D.n3 D.n1 24.1005
R277 D.n2 D 24.0005
R278 D D.n0 21.4405
R279 D D.n9 18.8805
R280 D.n9 D 10.5605
R281 D D.n0 8.0005
R282 D.n2 D 5.4405
R283 a_1266_47.n1 a_1266_47.t6 306.553
R284 a_1266_47.t3 a_1266_47.n5 302.491
R285 a_1266_47.n1 a_1266_47.n0 185
R286 a_1266_47.n3 a_1266_47.n2 185
R287 a_1266_47.n5 a_1266_47.n4 185
R288 a_1266_47.n3 a_1266_47.n1 43.0085
R289 a_1266_47.n5 a_1266_47.n3 43.0085
R290 a_1266_47.n4 a_1266_47.t2 24.9236
R291 a_1266_47.n4 a_1266_47.t1 24.9236
R292 a_1266_47.n2 a_1266_47.t4 24.9236
R293 a_1266_47.n2 a_1266_47.t0 24.9236
R294 a_1266_47.n0 a_1266_47.t5 24.9236
R295 a_1266_47.n0 a_1266_47.t7 24.9236
R296 VGND.n9 VGND.n8 205.927
R297 VGND.n11 VGND.n10 200.516
R298 VGND.n37 VGND.n36 199.739
R299 VGND.n12 VGND.n7 34.6358
R300 VGND.n16 VGND.n7 34.6358
R301 VGND.n17 VGND.n16 34.6358
R302 VGND.n18 VGND.n17 34.6358
R303 VGND.n18 VGND.n5 34.6358
R304 VGND.n22 VGND.n5 34.6358
R305 VGND.n23 VGND.n22 34.6358
R306 VGND.n24 VGND.n23 34.6358
R307 VGND.n24 VGND.n3 34.6358
R308 VGND.n28 VGND.n3 34.6358
R309 VGND.n29 VGND.n28 34.6358
R310 VGND.n30 VGND.n29 34.6358
R311 VGND.n30 VGND.n1 34.6358
R312 VGND.n34 VGND.n1 34.6358
R313 VGND.n35 VGND.n34 34.6358
R314 VGND.n12 VGND.n11 27.8593
R315 VGND.n8 VGND.t1 24.9236
R316 VGND.n8 VGND.t4 24.9236
R317 VGND.n10 VGND.t2 24.9236
R318 VGND.n10 VGND.t3 24.9236
R319 VGND.n36 VGND.t5 24.9236
R320 VGND.n36 VGND.t0 24.9236
R321 VGND.n37 VGND.n35 22.9652
R322 VGND.n13 VGND.n12 9.3005
R323 VGND.n14 VGND.n7 9.3005
R324 VGND.n16 VGND.n15 9.3005
R325 VGND.n17 VGND.n6 9.3005
R326 VGND.n19 VGND.n18 9.3005
R327 VGND.n20 VGND.n5 9.3005
R328 VGND.n22 VGND.n21 9.3005
R329 VGND.n23 VGND.n4 9.3005
R330 VGND.n25 VGND.n24 9.3005
R331 VGND.n26 VGND.n3 9.3005
R332 VGND.n28 VGND.n27 9.3005
R333 VGND.n29 VGND.n2 9.3005
R334 VGND.n31 VGND.n30 9.3005
R335 VGND.n32 VGND.n1 9.3005
R336 VGND.n34 VGND.n33 9.3005
R337 VGND.n35 VGND.n0 9.3005
R338 VGND.n38 VGND.n37 7.12063
R339 VGND.n11 VGND.n9 6.15047
R340 VGND.n13 VGND.n9 0.653323
R341 VGND.n38 VGND.n0 0.148519
R342 VGND.n14 VGND.n13 0.120292
R343 VGND.n15 VGND.n14 0.120292
R344 VGND.n15 VGND.n6 0.120292
R345 VGND.n19 VGND.n6 0.120292
R346 VGND.n20 VGND.n19 0.120292
R347 VGND.n21 VGND.n20 0.120292
R348 VGND.n21 VGND.n4 0.120292
R349 VGND.n25 VGND.n4 0.120292
R350 VGND.n26 VGND.n25 0.120292
R351 VGND.n27 VGND.n26 0.120292
R352 VGND.n27 VGND.n2 0.120292
R353 VGND.n31 VGND.n2 0.120292
R354 VGND.n32 VGND.n31 0.120292
R355 VGND.n33 VGND.n32 0.120292
R356 VGND.n33 VGND.n0 0.120292
R357 VGND VGND.n38 0.114842
R358 B_N.n0 B_N.t0 241.536
R359 B_N.n0 B_N.t1 169.237
R360 B_N B_N.n0 157.781
R361 A_N.n0 A_N.t0 230.155
R362 A_N.n0 A_N.t1 157.856
R363 A_N A_N.n0 153.962
C0 VPB C 0.138302f
C1 A_N B_N 0.105204f
C2 Y VGND 0.032548f
C3 VPB D 0.134132f
C4 VPB VPWR 0.213645f
C5 VPB Y 0.035889f
C6 A_N VPWR 0.017822f
C7 B_N VPWR 0.018591f
C8 C D 0.060549f
C9 C VPWR 0.054172f
C10 VPB VGND 0.011395f
C11 C Y 0.23587f
C12 D VPWR 0.097213f
C13 A_N VGND 0.017141f
C14 D Y 0.175239f
C15 B_N VGND 0.018039f
C16 VPWR Y 1.55974f
C17 C VGND 0.035668f
C18 VPB A_N 0.040386f
C19 D VGND 0.068179f
C20 VPB B_N 0.034714f
C21 VPWR VGND 0.15054f
C22 VGND VNB 1.09218f
C23 Y VNB 0.024838f
C24 VPWR VNB 0.944105f
C25 D VNB 0.419124f
C26 C VNB 0.402046f
C27 B_N VNB 0.095033f
C28 A_N VNB 0.156146f
C29 VPB VNB 2.0223f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR.t0 A.t0 a_109_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297.t0 B.t0 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t0 231.835
R1 A.n0 A.t1 157.07
R2 A A.n0 154.012
R3 a_109_297.t0 a_109_297.t1 41.3705
R4 VPWR VPWR.t0 250.668
R5 VPB.t0 VPB.t1 213.084
R6 VPB VPB.t0 189.409
R7 Y Y.n0 593.34
R8 Y.n2 Y.n0 289.24
R9 Y.n2 Y.n1 176.839
R10 Y.n0 Y.t1 26.5955
R11 Y.n1 Y.t2 24.9236
R12 Y.n1 Y.t0 24.9236
R13 Y Y.n2 11.3699
R14 VGND.n0 VGND.t0 163.721
R15 VGND.n0 VGND.t1 161.042
R16 VGND VGND.n0 0.489856
R17 VNB.t0 VNB.t1 1196.12
R18 VNB VNB.t0 911.327
R19 B.n0 B.t0 230.363
R20 B B.n0 158.4
R21 B.n0 B.t1 158.064
C0 A VGND 0.048556f
C1 Y VPWR 0.099513f
C2 B VPB 0.036697f
C3 Y VGND 0.154448f
C4 A VPB 0.041461f
C5 Y VPB 0.013918f
C6 B A 0.058413f
C7 B Y 0.087653f
C8 A Y 0.047068f
C9 VPWR VGND 0.031443f
C10 VPWR VPB 0.044857f
C11 VGND VPB 0.004563f
C12 B VPWR 0.014836f
C13 A VPWR 0.052823f
C14 B VGND 0.045088f
C15 VGND VNB 0.263197f
C16 VPWR VNB 0.214143f
C17 Y VNB 0.060508f
C18 A VNB 0.14927f
C19 B VNB 0.143121f
C20 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_4 VPB VNB VGND VPWR Y B A
X0 VPWR.t3 A.t0 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t3 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t2 A.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 A.t3 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t7 B.t0 Y.t10 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t1 A.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND.t0 A.t5 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t7 B.t1 Y.t11 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND.t4 B.t2 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t5 B.t3 a_27_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t1 A.t6 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y.t8 B.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y.t9 B.t5 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297.t5 B.t6 Y.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t7 B.t7 a_27_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297.t0 A.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n2 A.t7 212.081
R1 A.n1 A.t0 212.081
R2 A.n7 A.t2 212.081
R3 A.n8 A.t6 212.081
R4 A.n4 A.n3 173.761
R5 A A.n9 152.641
R6 A.n5 A.n4 152
R7 A.n6 A.n0 152
R8 A.n2 A.t5 139.78
R9 A.n1 A.t1 139.78
R10 A.n7 A.t3 139.78
R11 A.n8 A.t4 139.78
R12 A.n6 A.n5 49.6611
R13 A.n9 A.n7 45.2793
R14 A.n3 A.n1 42.3581
R15 A.n4 A.n0 21.7605
R16 A A.n0 21.1205
R17 A.n3 A.n2 18.9884
R18 A.n9 A.n8 16.0672
R19 A.n5 A.n1 7.30353
R20 A.n7 A.n6 4.38232
R21 a_27_297.n1 a_27_297.t7 361.329
R22 a_27_297.n1 a_27_297.n0 296.538
R23 a_27_297.n3 a_27_297.t1 278.985
R24 a_27_297.n3 a_27_297.n2 207.26
R25 a_27_297.n5 a_27_297.n4 188.952
R26 a_27_297.n4 a_27_297.n3 57.3598
R27 a_27_297.n4 a_27_297.n1 53.3404
R28 a_27_297.n2 a_27_297.t3 26.5955
R29 a_27_297.n2 a_27_297.t2 26.5955
R30 a_27_297.n0 a_27_297.t4 26.5955
R31 a_27_297.n0 a_27_297.t5 26.5955
R32 a_27_297.n5 a_27_297.t6 26.5955
R33 a_27_297.t0 a_27_297.n5 26.5955
R34 VPWR.n2 VPWR.n0 321.752
R35 VPWR.n2 VPWR.n1 315.784
R36 VPWR.n1 VPWR.t2 26.5955
R37 VPWR.n1 VPWR.t1 26.5955
R38 VPWR.n0 VPWR.t0 26.5955
R39 VPWR.n0 VPWR.t3 26.5955
R40 VPWR VPWR.n2 0.57222
R41 VPB.t4 VPB.t7 248.599
R42 VPB.t5 VPB.t4 248.599
R43 VPB.t6 VPB.t5 248.599
R44 VPB.t0 VPB.t6 248.599
R45 VPB.t3 VPB.t0 248.599
R46 VPB.t2 VPB.t3 248.599
R47 VPB.t1 VPB.t2 248.599
R48 VPB VPB.t1 201.246
R49 VGND.n5 VGND.t4 287.832
R50 VGND.n6 VGND.n4 207.965
R51 VGND.n9 VGND.n8 207.965
R52 VGND.n15 VGND.n1 207.965
R53 VGND.n17 VGND.t1 150.922
R54 VGND.n10 VGND.n7 34.6358
R55 VGND.n14 VGND.n2 34.6358
R56 VGND.n16 VGND.n15 32.377
R57 VGND.n9 VGND.n2 26.3534
R58 VGND.n4 VGND.t6 24.9236
R59 VGND.n4 VGND.t7 24.9236
R60 VGND.n8 VGND.t5 24.9236
R61 VGND.n8 VGND.t0 24.9236
R62 VGND.n1 VGND.t3 24.9236
R63 VGND.n1 VGND.t2 24.9236
R64 VGND.n17 VGND.n16 24.4711
R65 VGND.n6 VGND.n5 21.0905
R66 VGND.n7 VGND.n6 20.3299
R67 VGND.n18 VGND.n17 9.3005
R68 VGND.n7 VGND.n3 9.3005
R69 VGND.n11 VGND.n10 9.3005
R70 VGND.n12 VGND.n2 9.3005
R71 VGND.n14 VGND.n13 9.3005
R72 VGND.n16 VGND.n0 9.3005
R73 VGND.n10 VGND.n9 8.28285
R74 VGND.n15 VGND.n14 2.25932
R75 VGND.n5 VGND.n3 0.929432
R76 VGND.n11 VGND.n3 0.120292
R77 VGND.n12 VGND.n11 0.120292
R78 VGND.n13 VGND.n12 0.120292
R79 VGND.n13 VGND.n0 0.120292
R80 VGND.n18 VGND.n0 0.120292
R81 VGND VGND.n18 0.0213333
R82 Y.n2 Y.n1 332.332
R83 Y.n2 Y.n0 296.493
R84 Y.n5 Y.n3 135.249
R85 Y.n5 Y.n4 98.982
R86 Y.n7 Y.n6 98.982
R87 Y.n9 Y.n8 98.982
R88 Y Y.n9 39.3605
R89 Y.n7 Y.n5 36.2672
R90 Y.n9 Y.n7 36.2672
R91 Y.n1 Y.t6 26.5955
R92 Y.n1 Y.t7 26.5955
R93 Y.n0 Y.t10 26.5955
R94 Y.n0 Y.t5 26.5955
R95 Y.n3 Y.t2 24.9236
R96 Y.n3 Y.t1 24.9236
R97 Y.n4 Y.t0 24.9236
R98 Y.n4 Y.t3 24.9236
R99 Y.n6 Y.t11 24.9236
R100 Y.n6 Y.t8 24.9236
R101 Y.n8 Y.t4 24.9236
R102 Y.n8 Y.t9 24.9236
R103 Y Y.n2 23.3605
R104 VNB.t6 VNB.t4 1196.12
R105 VNB.t7 VNB.t6 1196.12
R106 VNB.t5 VNB.t7 1196.12
R107 VNB.t0 VNB.t5 1196.12
R108 VNB.t3 VNB.t0 1196.12
R109 VNB.t2 VNB.t3 1196.12
R110 VNB.t1 VNB.t2 1196.12
R111 VNB VNB.t1 968.285
R112 B.n3 B.t0 212.081
R113 B.n5 B.t3 212.081
R114 B.n7 B.t6 212.081
R115 B.n1 B.t7 212.081
R116 B.n4 B.n0 173.761
R117 B.n9 B.n2 173.761
R118 B.n6 B.n0 152
R119 B.n9 B.n8 152
R120 B.n3 B.t2 139.78
R121 B.n5 B.t5 139.78
R122 B.n7 B.t1 139.78
R123 B.n1 B.t4 139.78
R124 B.n8 B.n6 49.6611
R125 B.n5 B.n4 44.549
R126 B.n7 B.n2 43.0884
R127 B.n2 B.n1 18.2581
R128 B B.n9 17.6005
R129 B.n4 B.n3 16.7975
R130 B.n8 B.n7 6.57323
R131 B.n6 B.n5 5.11262
R132 B B.n0 4.1605
C0 VGND A 0.086395f
C1 B Y 0.354248f
C2 B VGND 0.048539f
C3 VPWR Y 0.029873f
C4 VPWR VGND 0.08158f
C5 Y VGND 0.564035f
C6 VPB A 0.120043f
C7 B VPB 0.1207f
C8 B A 0.062515f
C9 VPWR VPB 0.081483f
C10 VPWR A 0.079468f
C11 Y VPB 0.018966f
C12 Y A 0.165354f
C13 VGND VPB 0.007434f
C14 B VPWR 0.02936f
C15 VGND VNB 0.530513f
C16 Y VNB 0.083073f
C17 VPWR VNB 0.400525f
C18 B VNB 0.378897f
C19 A VNB 0.391512f
C20 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_8 VPB VNB VGND VPWR A B Y
X0 VPWR.t7 A.t0 a_27_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t15 B.t0 a_27_297.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297.t12 B.t1 Y.t14 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y.t7 A.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t6 A.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t23 B.t2 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_297.t11 B.t3 Y.t13 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t12 B.t4 a_27_297.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t6 A.t3 Y.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297.t5 A.t4 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y.t5 A.t5 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11 VGND.t4 A.t6 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t3 A.t7 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t2 A.t8 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t4 A.t9 a_27_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297.t8 B.t5 Y.t11 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X16 Y.t10 B.t6 a_27_297.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR.t3 A.t10 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X18 Y.t1 A.t11 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297.t14 B.t7 Y.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 Y.t0 A.t12 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t22 B.t8 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t21 B.t9 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y.t20 B.t10 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 Y.t8 B.t11 a_27_297.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_27_297.t2 A.t13 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND.t11 B.t12 Y.t19 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR.t1 A.t14 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND.t10 B.t13 Y.t18 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VGND.t9 B.t14 Y.t17 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VGND.t8 B.t15 Y.t16 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_27_297.t0 A.t15 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n5 A.t4 212.081
R1 A.n7 A.t9 212.081
R2 A.n3 A.t13 212.081
R3 A.n13 A.t14 212.081
R4 A.n15 A.t15 212.081
R5 A.n1 A.t0 212.081
R6 A.n21 A.t2 212.081
R7 A.n22 A.t10 212.081
R8 A.n6 A.n4 173.761
R9 A A.n23 152.321
R10 A.n8 A.n4 152
R11 A.n10 A.n9 152
R12 A.n12 A.n11 152
R13 A.n14 A.n2 152
R14 A.n17 A.n16 152
R15 A.n19 A.n18 152
R16 A.n20 A.n0 152
R17 A.n5 A.t8 139.78
R18 A.n7 A.t12 139.78
R19 A.n3 A.t7 139.78
R20 A.n13 A.t11 139.78
R21 A.n15 A.t6 139.78
R22 A.n1 A.t1 139.78
R23 A.n21 A.t3 139.78
R24 A.n22 A.t5 139.78
R25 A.n9 A.n8 49.6611
R26 A.n20 A.n19 49.6611
R27 A.n7 A.n6 45.2793
R28 A.n23 A.n21 45.2793
R29 A.n12 A.n3 42.3581
R30 A.n16 A.n1 42.3581
R31 A.n14 A.n13 30.6732
R32 A.n15 A.n14 30.6732
R33 A.n10 A.n4 21.7605
R34 A.n11 A.n10 21.7605
R35 A.n11 A.n2 21.7605
R36 A.n17 A.n2 21.7605
R37 A.n18 A.n17 21.7605
R38 A.n18 A.n0 21.7605
R39 A A.n0 21.4405
R40 A.n13 A.n12 18.9884
R41 A.n16 A.n15 18.9884
R42 A.n6 A.n5 16.0672
R43 A.n23 A.n22 16.0672
R44 A.n9 A.n3 7.30353
R45 A.n19 A.n1 7.30353
R46 A.n8 A.n7 4.38232
R47 A.n21 A.n20 4.38232
R48 a_27_297.n4 a_27_297.t8 371.904
R49 a_27_297.n4 a_27_297.n3 300.885
R50 a_27_297.n6 a_27_297.n5 300.885
R51 a_27_297.n8 a_27_297.n7 300.885
R52 a_27_297.n1 a_27_297.t3 267.507
R53 a_27_297.n11 a_27_297.n10 207.483
R54 a_27_297.n1 a_27_297.n0 207.483
R55 a_27_297.n13 a_27_297.n12 207.482
R56 a_27_297.n9 a_27_297.n2 187.506
R57 a_27_297.n9 a_27_297.n8 65.4258
R58 a_27_297.n11 a_27_297.n9 55.9405
R59 a_27_297.n6 a_27_297.n4 44.424
R60 a_27_297.n8 a_27_297.n6 44.424
R61 a_27_297.n12 a_27_297.n1 35.9624
R62 a_27_297.n12 a_27_297.n11 35.9624
R63 a_27_297.n2 a_27_297.t9 26.5955
R64 a_27_297.n2 a_27_297.t5 26.5955
R65 a_27_297.n3 a_27_297.t13 26.5955
R66 a_27_297.n3 a_27_297.t14 26.5955
R67 a_27_297.n5 a_27_297.t15 26.5955
R68 a_27_297.n5 a_27_297.t12 26.5955
R69 a_27_297.n7 a_27_297.t10 26.5955
R70 a_27_297.n7 a_27_297.t11 26.5955
R71 a_27_297.n10 a_27_297.t4 26.5955
R72 a_27_297.n10 a_27_297.t2 26.5955
R73 a_27_297.n0 a_27_297.t7 26.5955
R74 a_27_297.n0 a_27_297.t6 26.5955
R75 a_27_297.n13 a_27_297.t1 26.5955
R76 a_27_297.t0 a_27_297.n13 26.5955
R77 VPWR.n7 VPWR.n6 323.32
R78 VPWR.n10 VPWR.n3 316.245
R79 VPWR.n5 VPWR.n4 316.245
R80 VPWR.n12 VPWR.n1 316.245
R81 VPWR.n10 VPWR.n9 30.4946
R82 VPWR.n1 VPWR.t6 26.5955
R83 VPWR.n1 VPWR.t3 26.5955
R84 VPWR.n3 VPWR.t0 26.5955
R85 VPWR.n3 VPWR.t7 26.5955
R86 VPWR.n4 VPWR.t2 26.5955
R87 VPWR.n4 VPWR.t1 26.5955
R88 VPWR.n6 VPWR.t5 26.5955
R89 VPWR.n6 VPWR.t4 26.5955
R90 VPWR.n12 VPWR.n11 24.4711
R91 VPWR.n11 VPWR.n10 19.9534
R92 VPWR.n9 VPWR.n5 13.9299
R93 VPWR.n9 VPWR.n8 9.3005
R94 VPWR.n10 VPWR.n2 9.3005
R95 VPWR.n11 VPWR.n0 9.3005
R96 VPWR.n7 VPWR.n5 8.64394
R97 VPWR.n13 VPWR.n12 7.34101
R98 VPWR.n8 VPWR.n7 0.95509
R99 VPWR.n13 VPWR.n0 0.145717
R100 VPWR.n8 VPWR.n2 0.120292
R101 VPWR.n2 VPWR.n0 0.120292
R102 VPWR VPWR.n13 0.117681
R103 VPB.t13 VPB.t8 248.599
R104 VPB.t14 VPB.t13 248.599
R105 VPB.t15 VPB.t14 248.599
R106 VPB.t12 VPB.t15 248.599
R107 VPB.t10 VPB.t12 248.599
R108 VPB.t11 VPB.t10 248.599
R109 VPB.t9 VPB.t11 248.599
R110 VPB.t5 VPB.t9 248.599
R111 VPB.t4 VPB.t5 248.599
R112 VPB.t2 VPB.t4 248.599
R113 VPB.t1 VPB.t2 248.599
R114 VPB.t0 VPB.t1 248.599
R115 VPB.t7 VPB.t0 248.599
R116 VPB.t6 VPB.t7 248.599
R117 VPB.t3 VPB.t6 248.599
R118 VPB VPB.t3 204.207
R119 B.n3 B.t5 212.081
R120 B.n4 B.t6 212.081
R121 B.n6 B.t7 212.081
R122 B.n2 B.t11 212.081
R123 B.n11 B.t1 212.081
R124 B.n13 B.t0 212.081
R125 B.n16 B.t3 212.081
R126 B.n14 B.t4 212.081
R127 B.n15 B.n1 173.761
R128 B.n8 B.n7 152
R129 B.n10 B.n9 152
R130 B.n12 B.n0 152
R131 B.n19 B.n18 152
R132 B.n17 B.n1 152
R133 B.n3 B.t15 139.78
R134 B.n4 B.t2 139.78
R135 B.n6 B.t14 139.78
R136 B.n2 B.t9 139.78
R137 B.n11 B.t12 139.78
R138 B.n13 B.t10 139.78
R139 B.n16 B.t13 139.78
R140 B.n14 B.t8 139.78
R141 B.n8 B.n5 92.1128
R142 B.n4 B.n3 61.346
R143 B.n18 B.n17 49.6611
R144 B.n13 B.n12 44.549
R145 B.n16 B.n15 43.0884
R146 B.n7 B.n6 40.1672
R147 B.n11 B.n10 32.8641
R148 B.n6 B.n5 29.6015
R149 B.n10 B.n2 28.4823
R150 B.n5 B.n4 25.1769
R151 B.n9 B.n8 21.7605
R152 B.n9 B.n0 21.7605
R153 B.n19 B.n1 21.7605
R154 B.n7 B.n2 21.1793
R155 B.n15 B.n14 18.2581
R156 B.n12 B.n11 16.7975
R157 B B.n0 16.0005
R158 B.n17 B.n16 6.57323
R159 B B.n19 5.7605
R160 B.n18 B.n13 5.11262
R161 Y.n2 Y.n0 345.822
R162 Y.n2 Y.n1 301.397
R163 Y.n4 Y.n3 301.397
R164 Y.n6 Y.n5 301.397
R165 Y.n10 Y.n8 135.249
R166 Y.n10 Y.n9 98.982
R167 Y.n12 Y.n11 98.982
R168 Y.n14 Y.n13 98.982
R169 Y.n16 Y.n15 98.982
R170 Y.n18 Y.n17 98.982
R171 Y.n20 Y.n19 98.982
R172 Y.n21 Y.n7 95.6388
R173 Y.n21 Y.n20 48.0005
R174 Y.n4 Y.n2 44.424
R175 Y.n6 Y.n4 44.424
R176 Y Y.n21 41.3897
R177 Y.n12 Y.n10 36.2672
R178 Y.n14 Y.n12 36.2672
R179 Y.n16 Y.n14 36.2672
R180 Y.n18 Y.n16 36.2672
R181 Y.n20 Y.n18 36.2672
R182 Y.n0 Y.t13 26.5955
R183 Y.n0 Y.t12 26.5955
R184 Y.n1 Y.t14 26.5955
R185 Y.n1 Y.t15 26.5955
R186 Y.n3 Y.t9 26.5955
R187 Y.n3 Y.t8 26.5955
R188 Y.n5 Y.t11 26.5955
R189 Y.n5 Y.t10 26.5955
R190 Y.n7 Y.t16 24.9236
R191 Y.n7 Y.t23 24.9236
R192 Y.n8 Y.t6 24.9236
R193 Y.n8 Y.t5 24.9236
R194 Y.n9 Y.t4 24.9236
R195 Y.n9 Y.t7 24.9236
R196 Y.n11 Y.t3 24.9236
R197 Y.n11 Y.t1 24.9236
R198 Y.n13 Y.t2 24.9236
R199 Y.n13 Y.t0 24.9236
R200 Y.n15 Y.t18 24.9236
R201 Y.n15 Y.t22 24.9236
R202 Y.n17 Y.t19 24.9236
R203 Y.n17 Y.t20 24.9236
R204 Y.n19 Y.t17 24.9236
R205 Y.n19 Y.t21 24.9236
R206 Y Y.n6 2.30263
R207 VGND.n9 VGND.t8 287.257
R208 VGND.n11 VGND.n10 207.965
R209 VGND.n13 VGND.n12 207.965
R210 VGND.n19 VGND.n7 207.965
R211 VGND.n22 VGND.n21 207.965
R212 VGND.n28 VGND.n4 207.965
R213 VGND.n31 VGND.n30 207.965
R214 VGND.n37 VGND.n1 207.965
R215 VGND.n39 VGND.t5 150.922
R216 VGND.n18 VGND.n8 34.6358
R217 VGND.n23 VGND.n20 34.6358
R218 VGND.n27 VGND.n5 34.6358
R219 VGND.n32 VGND.n29 34.6358
R220 VGND.n36 VGND.n2 34.6358
R221 VGND.n14 VGND.n13 32.377
R222 VGND.n38 VGND.n37 32.377
R223 VGND.n14 VGND.n11 30.8711
R224 VGND.n19 VGND.n18 26.3534
R225 VGND.n31 VGND.n2 26.3534
R226 VGND.n10 VGND.t15 24.9236
R227 VGND.n10 VGND.t9 24.9236
R228 VGND.n12 VGND.t13 24.9236
R229 VGND.n12 VGND.t11 24.9236
R230 VGND.n7 VGND.t12 24.9236
R231 VGND.n7 VGND.t10 24.9236
R232 VGND.n21 VGND.t14 24.9236
R233 VGND.n21 VGND.t2 24.9236
R234 VGND.n4 VGND.t0 24.9236
R235 VGND.n4 VGND.t3 24.9236
R236 VGND.n30 VGND.t1 24.9236
R237 VGND.n30 VGND.t4 24.9236
R238 VGND.n1 VGND.t7 24.9236
R239 VGND.n1 VGND.t6 24.9236
R240 VGND.n39 VGND.n38 24.4711
R241 VGND.n23 VGND.n22 20.3299
R242 VGND.n29 VGND.n28 20.3299
R243 VGND.n22 VGND.n5 14.3064
R244 VGND.n28 VGND.n27 14.3064
R245 VGND.n11 VGND.n9 10.9193
R246 VGND.n40 VGND.n39 9.3005
R247 VGND.n15 VGND.n14 9.3005
R248 VGND.n16 VGND.n8 9.3005
R249 VGND.n18 VGND.n17 9.3005
R250 VGND.n20 VGND.n6 9.3005
R251 VGND.n24 VGND.n23 9.3005
R252 VGND.n25 VGND.n5 9.3005
R253 VGND.n27 VGND.n26 9.3005
R254 VGND.n29 VGND.n3 9.3005
R255 VGND.n33 VGND.n32 9.3005
R256 VGND.n34 VGND.n2 9.3005
R257 VGND.n36 VGND.n35 9.3005
R258 VGND.n38 VGND.n0 9.3005
R259 VGND.n20 VGND.n19 8.28285
R260 VGND.n32 VGND.n31 8.28285
R261 VGND.n13 VGND.n8 2.25932
R262 VGND.n37 VGND.n36 2.25932
R263 VGND.n15 VGND.n9 0.572285
R264 VGND.n16 VGND.n15 0.120292
R265 VGND.n17 VGND.n16 0.120292
R266 VGND.n17 VGND.n6 0.120292
R267 VGND.n24 VGND.n6 0.120292
R268 VGND.n25 VGND.n24 0.120292
R269 VGND.n26 VGND.n25 0.120292
R270 VGND.n26 VGND.n3 0.120292
R271 VGND.n33 VGND.n3 0.120292
R272 VGND.n34 VGND.n33 0.120292
R273 VGND.n35 VGND.n34 0.120292
R274 VGND.n35 VGND.n0 0.120292
R275 VGND.n40 VGND.n0 0.120292
R276 VGND VGND.n40 0.0226354
R277 VNB.t15 VNB.t8 1196.12
R278 VNB.t9 VNB.t15 1196.12
R279 VNB.t13 VNB.t9 1196.12
R280 VNB.t11 VNB.t13 1196.12
R281 VNB.t12 VNB.t11 1196.12
R282 VNB.t10 VNB.t12 1196.12
R283 VNB.t14 VNB.t10 1196.12
R284 VNB.t2 VNB.t14 1196.12
R285 VNB.t0 VNB.t2 1196.12
R286 VNB.t3 VNB.t0 1196.12
R287 VNB.t1 VNB.t3 1196.12
R288 VNB.t4 VNB.t1 1196.12
R289 VNB.t7 VNB.t4 1196.12
R290 VNB.t6 VNB.t7 1196.12
R291 VNB.t5 VNB.t6 1196.12
R292 VNB VNB.t5 982.524
C0 Y VGND 1.07787f
C1 VPB A 0.247191f
C2 VPB B 0.246859f
C3 A B 0.063776f
C4 VPB VPWR 0.132293f
C5 A VPWR 0.15961f
C6 VPB Y 0.019684f
C7 B VPWR 0.067937f
C8 A Y 0.375704f
C9 VPB VGND 0.010296f
C10 B Y 0.745396f
C11 A VGND 0.120249f
C12 B VGND 0.116971f
C13 VPWR Y 0.047801f
C14 VPWR VGND 0.143561f
C15 VGND VNB 0.850474f
C16 Y VNB 0.077644f
C17 VPWR VNB 0.662671f
C18 B VNB 0.745716f
C19 A VNB 0.756478f
C20 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2b_1 VPB VNB VGND VPWR B_N A Y
X0 Y.t1 a_74_47.t2 a_265_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR.t1 B_N.t0 a_74_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1573 pd=1.39 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_265_297.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.1573 ps=1.39 w=1 l=0.15
X3 Y.t0 A.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VGND.t0 B_N.t1 a_74_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t1 a_74_47.t3 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_74_47.n1 a_74_47.t1 654.968
R1 a_74_47.t0 a_74_47.n1 302.779
R2 a_74_47.n1 a_74_47.n0 246.404
R3 a_74_47.n0 a_74_47.t2 236.18
R4 a_74_47.n0 a_74_47.t3 163.881
R5 a_265_297.t0 a_265_297.t1 41.3705
R6 Y Y.n0 589.914
R7 Y.n2 Y.n0 585
R8 Y.n2 Y.n1 211.56
R9 Y.n0 Y.t1 26.5955
R10 Y.n1 Y.t2 24.9236
R11 Y.n1 Y.t0 24.9236
R12 Y Y.n2 2.85764
R13 VPB VPB.t1 334.425
R14 VPB.t1 VPB.t0 319.627
R15 VPB.t0 VPB.t2 213.084
R16 B_N B_N.n0 221.946
R17 B_N.n0 B_N.t1 176.733
R18 B_N.n0 B_N.t0 119.624
R19 VPWR VPWR.n0 317.954
R20 VPWR.n0 VPWR.t1 121.953
R21 VPWR.n0 VPWR.t0 25.6105
R22 A.n0 A.t0 236.18
R23 A.n0 A.t1 163.881
R24 A A.n0 156.678
R25 VGND.n1 VGND.t1 282.298
R26 VGND.n1 VGND.n0 129.262
R27 VGND.n0 VGND.t0 57.8133
R28 VGND.n0 VGND.t2 24.7549
R29 VGND VGND.n1 0.55669
R30 VNB VNB.t0 1594.82
R31 VNB.t0 VNB.t2 1381.23
R32 VNB.t2 VNB.t1 1196.12
C0 VPWR VGND 0.046161f
C1 VPB VPWR 0.075008f
C2 B_N VGND 0.027194f
C3 VPB B_N 0.061515f
C4 A VPWR 0.020882f
C5 A B_N 0.044907f
C6 VPWR B_N 0.012306f
C7 Y VGND 0.175424f
C8 VPB Y 0.02233f
C9 A Y 0.019983f
C10 VPWR Y 0.102774f
C11 VPB VGND 0.010151f
C12 B_N Y 0.002335f
C13 A VGND 0.027938f
C14 VPB A 0.031643f
C15 VGND VNB 0.329149f
C16 Y VNB 0.085029f
C17 B_N VNB 0.21207f
C18 VPWR VNB 0.268516f
C19 A VNB 0.09622f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2b_2 VPB VNB VGND VPWR Y A B_N
X0 Y.t3 a_251_21.t2 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t5 a_251_21.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t0 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t0 A.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t1 A.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X5 VGND.t2 a_251_21.t4 Y.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t3 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR.t2 B_N.t0 a_251_21.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND.t4 B_N.t1 a_251_21.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_27_297.t1 a_251_21.t5 Y.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 a_251_21.n2 a_251_21.t1 725.646
R1 a_251_21.t0 a_251_21.n2 248.954
R2 a_251_21.n1 a_251_21.t5 212.081
R3 a_251_21.n0 a_251_21.t2 212.081
R4 a_251_21.n2 a_251_21.n1 207.535
R5 a_251_21.n1 a_251_21.t4 139.78
R6 a_251_21.n0 a_251_21.t3 139.78
R7 a_251_21.n1 a_251_21.n0 61.346
R8 a_27_297.n0 a_27_297.t1 298.418
R9 a_27_297.n0 a_27_297.t3 288.243
R10 a_27_297.n1 a_27_297.n0 187.506
R11 a_27_297.n1 a_27_297.t2 26.5955
R12 a_27_297.t0 a_27_297.n1 26.5955
R13 Y.n2 Y.n1 337.207
R14 Y Y.n4 186.358
R15 Y.n4 Y.n3 185
R16 Y.n2 Y.n0 137.189
R17 Y.n1 Y.t2 26.5955
R18 Y.n1 Y.t3 26.5955
R19 Y.n4 Y.t4 24.9236
R20 Y.n4 Y.t5 24.9236
R21 Y.n0 Y.t0 24.9236
R22 Y.n0 Y.t1 24.9236
R23 Y Y.n3 11.8308
R24 Y.n3 Y.n2 3.10353
R25 VPB.t1 VPB.t4 556.386
R26 VPB.t2 VPB.t1 248.599
R27 VPB.t0 VPB.t2 248.599
R28 VPB.t3 VPB.t0 248.599
R29 VPB VPB.t3 201.246
R30 VGND.n4 VGND.t4 264.288
R31 VGND.n8 VGND.n1 207.965
R32 VGND.n3 VGND.t2 160.8
R33 VGND.n10 VGND.t1 151.194
R34 VGND.n7 VGND.n2 34.6358
R35 VGND.n9 VGND.n8 32.377
R36 VGND.n3 VGND.n2 26.3534
R37 VGND.n1 VGND.t3 24.9236
R38 VGND.n1 VGND.t0 24.9236
R39 VGND.n10 VGND.n9 24.4711
R40 VGND.n4 VGND.n3 15.4369
R41 VGND.n11 VGND.n10 9.3005
R42 VGND.n5 VGND.n2 9.3005
R43 VGND.n7 VGND.n6 9.3005
R44 VGND.n9 VGND.n0 9.3005
R45 VGND.n8 VGND.n7 2.25932
R46 VGND.n5 VGND.n4 0.572285
R47 VGND.n6 VGND.n5 0.120292
R48 VGND.n6 VGND.n0 0.120292
R49 VGND.n11 VGND.n0 0.120292
R50 VGND VGND.n11 0.0213333
R51 VNB.t2 VNB.t4 2677.02
R52 VNB.t3 VNB.t2 1196.12
R53 VNB.t0 VNB.t3 1196.12
R54 VNB.t1 VNB.t0 1196.12
R55 VNB VNB.t1 968.285
R56 A.n0 A.t0 212.081
R57 A.n1 A.t3 212.081
R58 A A.n2 153.601
R59 A.n0 A.t1 139.78
R60 A.n1 A.t2 139.78
R61 A.n2 A.n0 38.7066
R62 A.n2 A.n1 22.6399
R63 VPWR.n1 VPWR.t2 676.692
R64 VPWR.n1 VPWR.n0 322.19
R65 VPWR.n0 VPWR.t1 26.5955
R66 VPWR.n0 VPWR.t0 26.5955
R67 VPWR VPWR.n1 0.151166
R68 B_N.n0 B_N.t0 333.173
R69 B_N B_N.n0 164.708
R70 B_N.n0 B_N.t1 130.732
C0 VPB VPWR 0.080685f
C1 A VPWR 0.04237f
C2 VPB Y 0.005224f
C3 B_N VPWR 0.043028f
C4 A Y 0.069669f
C5 B_N Y 0.00143f
C6 VGND VPB 0.009577f
C7 VPWR Y 0.009649f
C8 VGND A 0.033005f
C9 VGND B_N 0.053975f
C10 VGND VPWR 0.064184f
C11 VGND Y 0.281397f
C12 VPB A 0.055356f
C13 VPB B_N 0.10759f
C14 VGND VNB 0.466325f
C15 Y VNB 0.016372f
C16 VPWR VNB 0.34094f
C17 B_N VNB 0.206554f
C18 A VNB 0.203992f
C19 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2b_4 VNB VPB VGND VPWR Y B_N A
X0 VPWR.t4 A.t0 a_27_297.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t11 A.t1 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t6 A.t2 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t7 A.t3 Y.t10 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t0 a_419_21.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t9 A.t4 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND.t5 A.t5 Y.t8 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t0 a_419_21.t3 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND.t1 a_419_21.t4 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t3 a_419_21.t5 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t2 A.t6 a_27_297.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y.t4 a_419_21.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t4 B_N.t0 a_419_21.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.182 ps=1.86 w=0.65 l=0.15
X13 Y.t5 a_419_21.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t0 B_N.t1 a_419_21.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.27 ps=2.54 w=1 l=0.15
X15 a_27_297.t2 a_419_21.t8 Y.t6 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y.t7 a_419_21.t9 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297.t4 A.t7 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n2 A.t7 212.081
R1 A.n1 A.t0 212.081
R2 A.n7 A.t2 212.081
R3 A.n8 A.t6 212.081
R4 A.n4 A.n3 173.761
R5 A A.n9 152.641
R6 A.n5 A.n4 152
R7 A.n6 A.n0 152
R8 A.n2 A.t5 139.78
R9 A.n1 A.t1 139.78
R10 A.n7 A.t3 139.78
R11 A.n8 A.t4 139.78
R12 A.n6 A.n5 49.6611
R13 A.n9 A.n7 45.2793
R14 A.n3 A.n1 42.3581
R15 A.n4 A.n0 21.7605
R16 A A.n0 21.1205
R17 A.n3 A.n2 18.9884
R18 A.n9 A.n8 16.0672
R19 A.n5 A.n1 7.30353
R20 A.n7 A.n6 4.38232
R21 a_27_297.n5 a_27_297.n4 296.538
R22 a_27_297.n1 a_27_297.t5 278.786
R23 a_27_297.t0 a_27_297.n5 267.592
R24 a_27_297.n1 a_27_297.n0 207.26
R25 a_27_297.n3 a_27_297.n2 188.952
R26 a_27_297.n3 a_27_297.n1 57.3601
R27 a_27_297.n5 a_27_297.n3 53.34
R28 a_27_297.n2 a_27_297.t3 26.5955
R29 a_27_297.n2 a_27_297.t4 26.5955
R30 a_27_297.n0 a_27_297.t7 26.5955
R31 a_27_297.n0 a_27_297.t6 26.5955
R32 a_27_297.n4 a_27_297.t1 26.5955
R33 a_27_297.n4 a_27_297.t2 26.5955
R34 VPWR.n4 VPWR.n3 316.245
R35 VPWR.n6 VPWR.n1 310.5
R36 VPWR.n2 VPWR.t0 246.484
R37 VPWR.n1 VPWR.t3 26.5955
R38 VPWR.n1 VPWR.t2 26.5955
R39 VPWR.n3 VPWR.t1 26.5955
R40 VPWR.n3 VPWR.t4 26.5955
R41 VPWR.n6 VPWR.n5 21.4593
R42 VPWR.n5 VPWR.n4 16.9417
R43 VPWR.n5 VPWR.n0 9.3005
R44 VPWR.n4 VPWR.n2 7.56304
R45 VPWR.n7 VPWR.n6 7.1994
R46 VPWR.n2 VPWR.n0 0.147879
R47 VPWR.n7 VPWR.n0 0.147518
R48 VPWR VPWR.n7 0.114555
R49 VPB.t0 VPB.t4 574.144
R50 VPB.t1 VPB.t0 248.599
R51 VPB.t2 VPB.t1 248.599
R52 VPB.t3 VPB.t2 248.599
R53 VPB.t5 VPB.t3 248.599
R54 VPB.t8 VPB.t5 248.599
R55 VPB.t7 VPB.t8 248.599
R56 VPB.t6 VPB.t7 248.599
R57 VPB VPB.t6 201.246
R58 VGND.n11 VGND.n4 207.965
R59 VGND.n14 VGND.n13 207.965
R60 VGND.n20 VGND.n1 207.965
R61 VGND.n7 VGND.t4 157.48
R62 VGND.n6 VGND.t1 152.594
R63 VGND.n22 VGND.t6 150.53
R64 VGND.n10 VGND.n5 34.6358
R65 VGND.n15 VGND.n12 34.6358
R66 VGND.n19 VGND.n2 34.6358
R67 VGND.n21 VGND.n20 32.377
R68 VGND.n14 VGND.n2 26.3534
R69 VGND.n4 VGND.t3 24.9236
R70 VGND.n4 VGND.t0 24.9236
R71 VGND.n13 VGND.t2 24.9236
R72 VGND.n13 VGND.t5 24.9236
R73 VGND.n1 VGND.t8 24.9236
R74 VGND.n1 VGND.t7 24.9236
R75 VGND.n22 VGND.n21 24.4711
R76 VGND.n12 VGND.n11 20.3299
R77 VGND.n11 VGND.n10 14.3064
R78 VGND.n7 VGND.n6 11.8922
R79 VGND.n23 VGND.n22 9.3005
R80 VGND.n8 VGND.n5 9.3005
R81 VGND.n10 VGND.n9 9.3005
R82 VGND.n12 VGND.n3 9.3005
R83 VGND.n16 VGND.n15 9.3005
R84 VGND.n17 VGND.n2 9.3005
R85 VGND.n19 VGND.n18 9.3005
R86 VGND.n21 VGND.n0 9.3005
R87 VGND.n15 VGND.n14 8.28285
R88 VGND.n6 VGND.n5 7.90638
R89 VGND.n20 VGND.n19 2.25932
R90 VGND.n8 VGND.n7 0.714832
R91 VGND.n9 VGND.n8 0.120292
R92 VGND.n9 VGND.n3 0.120292
R93 VGND.n16 VGND.n3 0.120292
R94 VGND.n17 VGND.n16 0.120292
R95 VGND.n18 VGND.n17 0.120292
R96 VGND.n18 VGND.n0 0.120292
R97 VGND.n23 VGND.n0 0.120292
R98 VGND VGND.n23 0.0213333
R99 Y Y.n0 309.719
R100 Y.n9 Y.n1 298.637
R101 Y.n8 Y.n2 141.293
R102 Y.n6 Y.n4 135.249
R103 Y.n6 Y.n5 98.982
R104 Y.n7 Y.n3 95.6388
R105 Y.n7 Y.n6 48.0005
R106 Y.n9 Y.n8 26.7641
R107 Y.n0 Y.t0 26.5955
R108 Y.n0 Y.t3 26.5955
R109 Y.n1 Y.t6 26.5955
R110 Y.n1 Y.t7 26.5955
R111 Y.n3 Y.t1 24.9236
R112 Y.n3 Y.t4 24.9236
R113 Y.n4 Y.t10 24.9236
R114 Y.n4 Y.t9 24.9236
R115 Y.n5 Y.t8 24.9236
R116 Y.n5 Y.t11 24.9236
R117 Y.n2 Y.t2 24.9236
R118 Y.n2 Y.t5 24.9236
R119 Y Y.n9 12.1605
R120 Y.n8 Y.n7 5.68939
R121 VNB.t1 VNB.t4 2762.46
R122 VNB.t3 VNB.t1 1196.12
R123 VNB.t0 VNB.t3 1196.12
R124 VNB.t2 VNB.t0 1196.12
R125 VNB.t5 VNB.t2 1196.12
R126 VNB.t8 VNB.t5 1196.12
R127 VNB.t7 VNB.t8 1196.12
R128 VNB.t6 VNB.t7 1196.12
R129 VNB VNB.t6 968.285
R130 a_419_21.t1 a_419_21.n8 252.549
R131 a_419_21.n6 a_419_21.t2 212.081
R132 a_419_21.n4 a_419_21.t5 212.081
R133 a_419_21.n2 a_419_21.t8 212.081
R134 a_419_21.n1 a_419_21.t9 212.081
R135 a_419_21.n3 a_419_21.n0 173.761
R136 a_419_21.n8 a_419_21.t0 153.874
R137 a_419_21.n5 a_419_21.n0 152
R138 a_419_21.n6 a_419_21.t4 139.78
R139 a_419_21.n4 a_419_21.t7 139.78
R140 a_419_21.n2 a_419_21.t3 139.78
R141 a_419_21.n1 a_419_21.t6 139.78
R142 a_419_21.n7 a_419_21.n6 112.322
R143 a_419_21.n2 a_419_21.n1 61.346
R144 a_419_21.n3 a_419_21.n2 54.0429
R145 a_419_21.n5 a_419_21.n4 42.3581
R146 a_419_21.n7 a_419_21.n0 30.5712
R147 a_419_21.n6 a_419_21.n5 18.9884
R148 a_419_21.n8 a_419_21.n7 14.5696
R149 a_419_21.n4 a_419_21.n3 7.30353
R150 B_N.n0 B_N.t1 229.754
R151 B_N B_N.n0 159.315
R152 B_N.n0 B_N.t0 157.453
C0 A VGND 0.067619f
C1 B_N VGND 0.051879f
C2 VPB A 0.119415f
C3 VPB B_N 0.04669f
C4 VPWR Y 0.020844f
C5 VPWR VGND 0.102679f
C6 Y VGND 0.544571f
C7 VPB VPWR 0.116357f
C8 A VPWR 0.07913f
C9 VPB Y 0.009206f
C10 A Y 0.176949f
C11 B_N VPWR 0.055498f
C12 VPB VGND 0.009839f
C13 VGND VNB 0.651371f
C14 Y VNB 0.025042f
C15 VPWR VNB 0.516619f
C16 B_N VNB 0.150465f
C17 A VNB 0.389045f
C18 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_1 VPB VNB VGND VPWR C B A Y
X0 VPWR.t0 A.t0 a_193_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297.t1 B.t0 a_109_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t2 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t2 A.t1 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297.t0 C.t0 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND.t0 C.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t0 229.001
R1 A A.n0 170.726
R2 A.n0 A.t1 156.702
R3 a_193_297.t0 a_193_297.t1 53.1905
R4 VPWR VPWR.t0 345.317
R5 VPB.t2 VPB.t1 248.599
R6 VPB.t0 VPB.t2 248.599
R7 VPB VPB.t0 189.409
R8 B.n0 B.t0 241.536
R9 B.n0 B.t1 169.237
R10 B B.n0 165.518
R11 a_109_297.t0 a_109_297.t1 53.1905
R12 VGND.n1 VGND.t2 284.839
R13 VGND.n1 VGND.n0 205.357
R14 VGND.n0 VGND.t1 24.9236
R15 VGND.n0 VGND.t0 24.9236
R16 VGND VGND.n1 0.636176
R17 Y.n1 Y.t0 276.308
R18 Y.n2 Y.t1 223.29
R19 Y.n1 Y.n0 192.906
R20 Y.n2 Y.n1 169.476
R21 Y.n0 Y.t3 24.9236
R22 Y.n0 Y.t2 24.9236
R23 Y Y.n2 2.7631
R24 VNB.t1 VNB.t2 1196.12
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 911.327
R27 C.n0 C.t0 231.017
R28 C.n0 C.t1 158.716
R29 C C.n0 156.268
C0 C B 0.093635f
C1 VPB A 0.043587f
C2 VPB Y 0.013918f
C3 C Y 0.091882f
C4 B A 0.05655f
C5 VPB VPWR 0.04706f
C6 C VPWR 0.009396f
C7 B Y 0.201894f
C8 VPB VGND 0.004665f
C9 A Y 0.111098f
C10 B VPWR 0.012958f
C11 C VGND 0.016667f
C12 B VGND 0.019155f
C13 A VPWR 0.047669f
C14 Y VPWR 0.170502f
C15 A VGND 0.048255f
C16 Y VGND 0.131904f
C17 VPWR VGND 0.040648f
C18 VPB C 0.036858f
C19 VPB B 0.028594f
C20 VGND VNB 0.26567f
C21 VPWR VNB 0.236658f
C22 Y VNB 0.080649f
C23 A VNB 0.176956f
C24 B VNB 0.093371f
C25 C VNB 0.143786f
C26 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_2 VPB VNB VGND VPWR A B C Y
X0 Y.t5 C.t0 a_281_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297.t1 B.t0 a_27_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t2 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297.t3 A.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t3 A.t1 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t0 A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X6 VGND.t0 B.t2 Y.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t5 C.t1 Y.t7 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t6 C.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR.t0 A.t3 a_27_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297.t2 C.t3 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297.t0 B.t3 a_281_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
R0 C.n0 C.t3 212.081
R1 C.n1 C.t0 212.081
R2 C C.n2 165.709
R3 C.n0 C.t1 139.78
R4 C.n1 C.t2 139.78
R5 C.n2 C.n0 48.2005
R6 C.n2 C.n1 13.146
R7 a_281_297.n0 a_281_297.t2 371.904
R8 a_281_297.n1 a_281_297.n0 357.356
R9 a_281_297.n0 a_281_297.t3 329.063
R10 a_281_297.t0 a_281_297.n1 26.5955
R11 a_281_297.n1 a_281_297.t1 26.5955
R12 Y Y.n0 311.889
R13 Y.n3 Y.n1 135.249
R14 Y.n3 Y.n2 98.982
R15 Y.n5 Y.n4 98.982
R16 Y.n5 Y.n3 74.6672
R17 Y.n0 Y.t4 26.5955
R18 Y.n0 Y.t5 26.5955
R19 Y.n1 Y.t1 24.9236
R20 Y.n1 Y.t0 24.9236
R21 Y.n2 Y.t3 24.9236
R22 Y.n2 Y.t2 24.9236
R23 Y.n4 Y.t7 24.9236
R24 Y.n4 Y.t6 24.9236
R25 Y Y.n5 21.0865
R26 VPB.t1 VPB.t5 568.225
R27 VPB.t5 VPB.t4 248.599
R28 VPB.t3 VPB.t1 248.599
R29 VPB.t2 VPB.t3 248.599
R30 VPB.t0 VPB.t2 248.599
R31 VPB VPB.t0 201.246
R32 B.n0 B.t3 212.081
R33 B.n1 B.t0 212.081
R34 B B.n2 152.671
R35 B.n0 B.t2 139.78
R36 B.n1 B.t1 139.78
R37 B.n2 B.n0 32.8641
R38 B.n2 B.n1 28.4823
R39 a_27_297.n0 a_27_297.t0 371.904
R40 a_27_297.n0 a_27_297.t2 279.267
R41 a_27_297.n1 a_27_297.n0 208.506
R42 a_27_297.t1 a_27_297.n1 26.5955
R43 a_27_297.n1 a_27_297.t3 26.5955
R44 VGND.n3 VGND.t5 287.342
R45 VGND.n5 VGND.t0 263.462
R46 VGND.n4 VGND.t4 263.462
R47 VGND.n11 VGND.n1 207.965
R48 VGND.n13 VGND.t2 151.584
R49 VGND.n10 VGND.n2 34.6358
R50 VGND.n12 VGND.n11 32.377
R51 VGND.n1 VGND.t1 24.9236
R52 VGND.n1 VGND.t3 24.9236
R53 VGND.n13 VGND.n12 24.4711
R54 VGND.n5 VGND.n2 21.6534
R55 VGND.n14 VGND.n13 9.3005
R56 VGND.n7 VGND.n6 9.3005
R57 VGND.n8 VGND.n2 9.3005
R58 VGND.n10 VGND.n9 9.3005
R59 VGND.n12 VGND.n0 9.3005
R60 VGND.n6 VGND.n4 8.6005
R61 VGND.n4 VGND.n3 7.64062
R62 VGND.n11 VGND.n10 2.25932
R63 VGND.n6 VGND.n5 2.2005
R64 VGND.n7 VGND.n3 0.582239
R65 VGND.n8 VGND.n7 0.120292
R66 VGND.n9 VGND.n8 0.120292
R67 VGND.n9 VGND.n0 0.120292
R68 VGND.n14 VGND.n0 0.120292
R69 VGND VGND.n14 0.0213333
R70 VNB.t0 VNB.t4 2733.98
R71 VNB.t4 VNB.t5 1196.12
R72 VNB.t1 VNB.t0 1196.12
R73 VNB.t3 VNB.t1 1196.12
R74 VNB.t2 VNB.t3 1196.12
R75 VNB VNB.t2 968.285
R76 A.n0 A.t0 212.081
R77 A.n1 A.t3 212.081
R78 A A.n2 152.849
R79 A.n0 A.t1 139.78
R80 A.n1 A.t2 139.78
R81 A.n2 A.n0 38.7066
R82 A.n2 A.n1 22.6399
R83 VPWR VPWR.n0 324.387
R84 VPWR.n0 VPWR.t1 26.5955
R85 VPWR.n0 VPWR.t0 26.5955
C0 VPB B 0.059332f
C1 A B 0.069132f
C2 VPB C 0.067833f
C3 A C 3.63e-19
C4 VPB VPWR 0.077026f
C5 A VPWR 0.04397f
C6 B C 0.036601f
C7 VPB Y 0.013147f
C8 A Y 0.061458f
C9 B VPWR 0.022934f
C10 VPB VGND 0.009613f
C11 C VPWR 0.018605f
C12 B Y 0.118347f
C13 A VGND 0.056318f
C14 C Y 0.167791f
C15 B VGND 0.030998f
C16 C VGND 0.031166f
C17 VPWR Y 0.017335f
C18 VPWR VGND 0.072894f
C19 Y VGND 0.477898f
C20 VPB A 0.056239f
C21 VGND VNB 0.483019f
C22 Y VNB 0.075161f
C23 VPWR VNB 0.363175f
C24 C VNB 0.210714f
C25 B VNB 0.184258f
C26 A VNB 0.207334f
C27 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_4 VPB VNB VGND VPWR B A Y C
X0 VPWR.t3 A.t0 a_27_297.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_449_297.t7 C.t0 Y.t15 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297.t2 B.t0 a_449_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 Y.t7 A.t1 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t6 A.t2 VPWR.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t14 C.t1 a_449_297.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_449_297.t5 C.t2 Y.t13 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t6 A.t3 Y.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t12 C.t3 a_449_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t5 A.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND.t4 A.t5 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t3 B.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t11 C.t4 Y.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_449_297.t3 B.t2 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t1 A.t6 a_27_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y.t0 B.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y.t1 B.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y.t10 C.t5 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t9 C.t6 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297.t0 B.t5 a_449_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t0 B.t6 Y.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_449_297.t1 B.t7 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND.t8 C.t7 Y.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_27_297.t4 A.t7 VPWR.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n2 A.t7 212.081
R1 A.n1 A.t0 212.081
R2 A.n7 A.t2 212.081
R3 A.n8 A.t6 212.081
R4 A.n4 A.n3 172.725
R5 A A.n9 153.829
R6 A.n5 A.n4 152
R7 A.n6 A.n0 152
R8 A.n2 A.t5 139.78
R9 A.n1 A.t1 139.78
R10 A.n7 A.t3 139.78
R11 A.n8 A.t4 139.78
R12 A.n6 A.n5 49.6611
R13 A.n9 A.n7 48.2005
R14 A.n3 A.n1 39.4369
R15 A.n3 A.n2 21.9096
R16 A.n4 A.n0 20.7243
R17 A A.n0 18.8957
R18 A.n9 A.n8 13.146
R19 A.n5 A.n1 10.2247
R20 A.n7 A.n6 1.46111
R21 a_27_297.n4 a_27_297.t2 849.22
R22 a_27_297.n5 a_27_297.n4 303.188
R23 a_27_297.n2 a_27_297.t5 279.267
R24 a_27_297.n2 a_27_297.n1 208.507
R25 a_27_297.n3 a_27_297.n0 189.831
R26 a_27_297.n3 a_27_297.n2 61.957
R27 a_27_297.n4 a_27_297.n3 29.0658
R28 a_27_297.n0 a_27_297.t1 26.5955
R29 a_27_297.n0 a_27_297.t4 26.5955
R30 a_27_297.n1 a_27_297.t7 26.5955
R31 a_27_297.n1 a_27_297.t6 26.5955
R32 a_27_297.n5 a_27_297.t3 26.5955
R33 a_27_297.t0 a_27_297.n5 26.5955
R34 VPWR.n2 VPWR.n0 323.974
R35 VPWR.n2 VPWR.n1 323.86
R36 VPWR.n1 VPWR.t2 26.5955
R37 VPWR.n1 VPWR.t1 26.5955
R38 VPWR.n0 VPWR.t0 26.5955
R39 VPWR.n0 VPWR.t3 26.5955
R40 VPWR VPWR.n2 0.505993
R41 VPB.t6 VPB.t2 248.599
R42 VPB.t7 VPB.t6 248.599
R43 VPB.t4 VPB.t7 248.599
R44 VPB.t5 VPB.t4 248.599
R45 VPB.t3 VPB.t5 248.599
R46 VPB.t0 VPB.t3 248.599
R47 VPB.t1 VPB.t0 248.599
R48 VPB.t8 VPB.t1 248.599
R49 VPB.t11 VPB.t8 248.599
R50 VPB.t10 VPB.t11 248.599
R51 VPB.t9 VPB.t10 248.599
R52 VPB VPB.t9 201.246
R53 C.n0 C.t0 212.081
R54 C.n2 C.t1 212.081
R55 C.n4 C.t2 212.081
R56 C.n3 C.t3 212.081
R57 C C.n1 168
R58 C C.n5 157.761
R59 C.n0 C.t6 139.78
R60 C.n2 C.t7 139.78
R61 C.n4 C.t5 139.78
R62 C.n3 C.t4 139.78
R63 C.n4 C.n3 61.346
R64 C.n5 C.n4 51.1217
R65 C.n2 C.n1 39.4369
R66 C.n1 C.n0 21.9096
R67 C.n5 C.n2 10.2247
R68 Y.n2 Y.n0 636.367
R69 Y.n2 Y.n1 585
R70 Y.n5 Y.n3 135.249
R71 Y.n5 Y.n4 98.982
R72 Y.n7 Y.n6 98.982
R73 Y.n9 Y.n8 98.982
R74 Y.n11 Y.n10 98.982
R75 Y.n13 Y.n12 98.982
R76 Y Y.n2 98.7591
R77 Y Y.n13 66.2074
R78 Y.n7 Y.n5 36.2672
R79 Y.n9 Y.n7 36.2672
R80 Y.n11 Y.n9 36.2672
R81 Y.n13 Y.n11 36.2672
R82 Y.n1 Y.t15 26.5955
R83 Y.n1 Y.t14 26.5955
R84 Y.n0 Y.t13 26.5955
R85 Y.n0 Y.t12 26.5955
R86 Y.n3 Y.t6 24.9236
R87 Y.n3 Y.t5 24.9236
R88 Y.n4 Y.t4 24.9236
R89 Y.n4 Y.t7 24.9236
R90 Y.n6 Y.t3 24.9236
R91 Y.n6 Y.t0 24.9236
R92 Y.n8 Y.t11 24.9236
R93 Y.n8 Y.t1 24.9236
R94 Y.n10 Y.t8 24.9236
R95 Y.n10 Y.t10 24.9236
R96 Y.n12 Y.t2 24.9236
R97 Y.n12 Y.t9 24.9236
R98 a_449_297.n3 a_449_297.n1 653.904
R99 a_449_297.n4 a_449_297.n0 639.12
R100 a_449_297.n5 a_449_297.n4 585
R101 a_449_297.n3 a_449_297.n2 187.506
R102 a_449_297.n4 a_449_297.n3 70.2743
R103 a_449_297.n2 a_449_297.t4 26.5955
R104 a_449_297.n2 a_449_297.t3 26.5955
R105 a_449_297.n1 a_449_297.t0 26.5955
R106 a_449_297.n1 a_449_297.t1 26.5955
R107 a_449_297.n0 a_449_297.t2 26.5955
R108 a_449_297.n0 a_449_297.t7 26.5955
R109 a_449_297.t6 a_449_297.n5 26.5955
R110 a_449_297.n5 a_449_297.t5 26.5955
R111 B.n1 B.n0 352.291
R112 B.n0 B.t0 236.18
R113 B.n2 B.t2 212.081
R114 B.n4 B.t5 212.081
R115 B.n5 B.t7 212.081
R116 B.n0 B.t6 163.881
R117 B B.n6 163.582
R118 B.n3 B.n1 152
R119 B.n2 B.t4 139.78
R120 B.n4 B.t1 139.78
R121 B.n5 B.t3 139.78
R122 B.n3 B.n2 59.8853
R123 B.n6 B.n4 48.2005
R124 B.n6 B.n5 13.146
R125 B B.n1 9.14336
R126 B.n4 B.n3 1.46111
R127 VGND.n8 VGND.t0 293.212
R128 VGND.n9 VGND.n7 207.965
R129 VGND.n12 VGND.n11 207.965
R130 VGND.n18 VGND.n4 207.965
R131 VGND.n21 VGND.n20 207.965
R132 VGND.n27 VGND.n1 207.965
R133 VGND.n29 VGND.t5 150.922
R134 VGND.n13 VGND.n10 34.6358
R135 VGND.n17 VGND.n5 34.6358
R136 VGND.n22 VGND.n19 34.6358
R137 VGND.n26 VGND.n2 34.6358
R138 VGND.n9 VGND.n8 32.6509
R139 VGND.n28 VGND.n27 32.377
R140 VGND.n21 VGND.n2 26.3534
R141 VGND.n7 VGND.t9 24.9236
R142 VGND.n7 VGND.t8 24.9236
R143 VGND.n11 VGND.t10 24.9236
R144 VGND.n11 VGND.t11 24.9236
R145 VGND.n4 VGND.t1 24.9236
R146 VGND.n4 VGND.t3 24.9236
R147 VGND.n20 VGND.t2 24.9236
R148 VGND.n20 VGND.t4 24.9236
R149 VGND.n1 VGND.t7 24.9236
R150 VGND.n1 VGND.t6 24.9236
R151 VGND.n29 VGND.n28 24.4711
R152 VGND.n13 VGND.n12 20.3299
R153 VGND.n19 VGND.n18 20.3299
R154 VGND.n12 VGND.n5 14.3064
R155 VGND.n18 VGND.n17 14.3064
R156 VGND.n30 VGND.n29 9.3005
R157 VGND.n10 VGND.n6 9.3005
R158 VGND.n14 VGND.n13 9.3005
R159 VGND.n15 VGND.n5 9.3005
R160 VGND.n17 VGND.n16 9.3005
R161 VGND.n19 VGND.n3 9.3005
R162 VGND.n23 VGND.n22 9.3005
R163 VGND.n24 VGND.n2 9.3005
R164 VGND.n26 VGND.n25 9.3005
R165 VGND.n28 VGND.n0 9.3005
R166 VGND.n10 VGND.n9 8.28285
R167 VGND.n22 VGND.n21 8.28285
R168 VGND.n27 VGND.n26 2.25932
R169 VGND.n8 VGND.n6 1.45203
R170 VGND.n14 VGND.n6 0.120292
R171 VGND.n15 VGND.n14 0.120292
R172 VGND.n16 VGND.n15 0.120292
R173 VGND.n16 VGND.n3 0.120292
R174 VGND.n23 VGND.n3 0.120292
R175 VGND.n24 VGND.n23 0.120292
R176 VGND.n25 VGND.n24 0.120292
R177 VGND.n25 VGND.n0 0.120292
R178 VGND.n30 VGND.n0 0.120292
R179 VGND VGND.n30 0.0213333
R180 VNB.t9 VNB.t0 1196.12
R181 VNB.t8 VNB.t9 1196.12
R182 VNB.t10 VNB.t8 1196.12
R183 VNB.t11 VNB.t10 1196.12
R184 VNB.t1 VNB.t11 1196.12
R185 VNB.t3 VNB.t1 1196.12
R186 VNB.t2 VNB.t3 1196.12
R187 VNB.t4 VNB.t2 1196.12
R188 VNB.t7 VNB.t4 1196.12
R189 VNB.t6 VNB.t7 1196.12
R190 VNB.t5 VNB.t6 1196.12
R191 VNB VNB.t5 968.285
C0 VPWR VGND 0.058535f
C1 Y VGND 0.869307f
C2 VPB A 0.12099f
C3 VPB B 0.131222f
C4 VPB C 0.114202f
C5 A B 0.064455f
C6 VPB VPWR 0.109781f
C7 B C 0.266547f
C8 VPB Y 0.031564f
C9 A VPWR 0.089804f
C10 A Y 0.166186f
C11 B VPWR 0.02432f
C12 VPB VGND 0.009386f
C13 B Y 0.443998f
C14 C VPWR 0.014894f
C15 A VGND 0.091482f
C16 C Y 0.176307f
C17 B VGND 0.056808f
C18 C VGND 0.050592f
C19 VPWR Y 0.056209f
C20 VGND VNB 0.702973f
C21 Y VNB 0.126464f
C22 VPWR VNB 0.548794f
C23 C VNB 0.350113f
C24 B VNB 0.388866f
C25 A VNB 0.392851f
C26 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_1 VPB VNB VGND VPWR C_N B Y A
X0 VGND.t0 a_91_199.t2 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y.t2 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t1 A.t0 a_245_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199.t0 C_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND.t3 A.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297.t0 B.t1 a_161_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199.t1 C_N.t1 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297.t0 a_91_199.t3 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
R0 a_91_199.n1 a_91_199.t1 648.322
R1 a_91_199.t0 a_91_199.n1 344.796
R2 a_91_199.n1 a_91_199.n0 318.776
R3 a_91_199.n0 a_91_199.t3 234.804
R4 a_91_199.n0 a_91_199.t2 162.504
R5 Y.n2 Y.t0 393.575
R6 Y.n1 Y.n0 257.599
R7 Y.n1 Y.t1 132.192
R8 Y.n2 Y.n1 60.3299
R9 Y.n0 Y.t3 24.9236
R10 Y.n0 Y.t2 24.9236
R11 Y Y.n2 1.86956
R12 VGND.n2 VGND.n0 205.625
R13 VGND.n2 VGND.n1 116.099
R14 VGND.n1 VGND.t1 57.875
R15 VGND.n0 VGND.t2 24.9236
R16 VGND.n0 VGND.t0 24.9236
R17 VGND.n1 VGND.t3 24.6931
R18 VGND VGND.n2 0.830774
R19 VNB VNB.t0 1666.02
R20 VNB.t3 VNB.t1 1381.23
R21 VNB.t2 VNB.t3 1196.12
R22 VNB.t0 VNB.t2 1196.12
R23 B.n0 B.t1 241.536
R24 B.n0 B.t0 169.237
R25 B B.n0 153.756
R26 A.n0 A.t0 241.536
R27 A.n0 A.t1 169.237
R28 A A.n0 154.168
R29 a_245_297.t0 a_245_297.t1 53.1905
R30 VPWR VPWR.n0 612.967
R31 VPWR.n0 VPWR.t0 96.1553
R32 VPWR.n0 VPWR.t1 27.3647
R33 VPB VPB.t0 346.262
R34 VPB.t3 VPB.t2 287.072
R35 VPB.t1 VPB.t3 248.599
R36 VPB.t0 VPB.t1 248.599
R37 C_N.n0 C_N.t1 201.369
R38 C_N C_N.n0 154.582
R39 C_N.n0 C_N.t0 132.282
R40 a_161_297.t0 a_161_297.t1 53.1905
C0 VPB Y 0.021749f
C1 B A 0.108301f
C2 B Y 0.034729f
C3 A Y 0.003603f
C4 VPWR VPB 0.072582f
C5 VPWR B 0.010174f
C6 C_N VPB 0.057935f
C7 VGND VPB 0.008114f
C8 VPWR A 0.018159f
C9 C_N B 2.93e-19
C10 C_N A 0.091376f
C11 VGND B 0.013535f
C12 VPWR Y 0.074972f
C13 VGND A 0.041088f
C14 C_N Y 0.001167f
C15 VGND Y 0.221777f
C16 VPWR C_N 0.007204f
C17 VPB B 0.026494f
C18 VPWR VGND 0.054345f
C19 VPB A 0.031044f
C20 C_N VGND 0.017997f
C21 VGND VNB 0.359992f
C22 C_N VNB 0.124851f
C23 VPWR VNB 0.303327f
C24 Y VNB 0.111033f
C25 A VNB 0.095278f
C26 B VNB 0.087995f
C27 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_1 VPWR VGND VPB VNB TE Z A
X0 a_276_297.t0 a_27_47.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1 Z.t0 A.t0 a_204_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2 VPWR.t0 TE.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 Z.t1 A.t1 a_276_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4 a_204_47.t1 TE.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5 VGND.t0 TE.t2 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t0 a_27_47.n0 704.985
R1 a_27_47.n0 a_27_47.t2 393.536
R2 a_27_47.n0 a_27_47.t1 273.269
R3 VPWR VPWR.n0 322.656
R4 VPWR.n0 VPWR.t1 93.6562
R5 VPWR.n0 VPWR.t0 35.1791
R6 a_276_297.t0 a_276_297.t1 71.9055
R7 VPB.t0 VPB.t1 494.238
R8 VPB.t1 VPB.t2 304.829
R9 VPB VPB.t0 189.409
R10 A.n0 A.t1 229.754
R11 A.n0 A.t0 157.453
R12 A.n1 A.n0 152
R13 A.n1 A 15.2005
R14 A A.n1 2.93383
R15 a_204_47.t0 a_204_47.t1 133.846
R16 Z Z.t1 816.716
R17 Z.n0 Z.t0 128.907
R18 Z.n0 Z 112.183
R19 Z Z.n0 3.19519
R20 VNB.t1 VNB.t0 2491.91
R21 VNB.t2 VNB.t1 1352.75
R22 VNB VNB.t2 911.327
R23 TE.n1 TE.t0 358.288
R24 TE.n0 TE.t1 257.067
R25 TE.n0 TE.t2 189.588
R26 TE.n2 TE.n1 171.946
R27 TE.n1 TE.n0 40.1672
R28 TE.n2 TE 7.93093
R29 TE TE.n2 1.53093
R30 VGND VGND.n0 190.419
R31 VGND.n0 VGND.t1 41.6488
R32 VGND.n0 VGND.t0 38.5719
C0 VPB TE 0.120084f
C1 VPB A 0.044798f
C2 VPB Z 0.00678f
C3 VPB VPWR 0.04882f
C4 TE A 0.005655f
C5 TE Z 0.002295f
C6 VPB VGND 0.004742f
C7 TE VPWR 0.02085f
C8 TE VGND 0.032026f
C9 A Z 0.171086f
C10 A VPWR 0.01187f
C11 A VGND 0.011538f
C12 VPWR Z 0.096503f
C13 Z VGND 0.09789f
C14 VPWR VGND 0.047226f
C15 VGND VNB 0.295665f
C16 Z VNB 0.052382f
C17 VPWR VNB 0.247074f
C18 A VNB 0.174637f
C19 TE VNB 0.288109f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_2 VGND VPWR VPB VNB TE Z A
X0 VPWR.t1 a_27_47.t2 a_215_309.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.2444 ps=2.4 w=0.94 l=0.15
X1 a_204_47.t3 A.t0 Z.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t2 TE.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 Z.t3 A.t1 a_204_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_215_309.t0 A.t2 Z.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Z.t0 A.t3 a_215_309.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16025 ps=1.325 w=1 l=0.15
X6 a_204_47.t1 TE.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7 VGND.t0 TE.t2 a_204_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_215_309.t2 a_27_47.t3 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.16025 pd=1.325 as=0.1269 ps=1.21 w=0.94 l=0.15
X9 VGND.t2 TE.t3 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t1 a_27_47.n1 676.984
R1 a_27_47.n1 a_27_47.t0 264.101
R2 a_27_47.n0 a_27_47.t2 253.853
R3 a_27_47.n1 a_27_47.n0 232.799
R4 a_27_47.n0 a_27_47.t3 189.588
R5 a_215_309.n1 a_215_309.t3 431.471
R6 a_215_309.t0 a_215_309.n1 397.534
R7 a_215_309.n1 a_215_309.n0 286.329
R8 a_215_309.n0 a_215_309.t2 34.5803
R9 a_215_309.n0 a_215_309.t1 31.6921
R10 VPWR.n1 VPWR.t2 736.409
R11 VPWR.n1 VPWR.n0 315.274
R12 VPWR.n0 VPWR.t0 28.2931
R13 VPWR.n0 VPWR.t1 28.2931
R14 VPWR VPWR.n1 0.487289
R15 VPB.t4 VPB.t3 556.386
R16 VPB.t2 VPB.t1 281.154
R17 VPB.t1 VPB.t0 248.599
R18 VPB.t3 VPB.t2 248.599
R19 VPB VPB.t4 189.409
R20 A.n1 A.t2 212.081
R21 A.n0 A.t3 212.081
R22 A.n2 A.n1 189.245
R23 A.n1 A.t0 139.78
R24 A.n0 A.t1 139.78
R25 A.n1 A.n0 61.346
R26 A.n2 A 12.8005
R27 A A.n2 2.47068
R28 Z Z.n0 591.4
R29 Z.n2 Z.n0 585
R30 Z Z.n1 185.195
R31 Z.n0 Z.t1 26.5955
R32 Z.n0 Z.t0 26.5955
R33 Z.n1 Z.t2 24.9236
R34 Z.n1 Z.t3 24.9236
R35 Z Z.n2 6.78838
R36 Z.n2 Z 6.4005
R37 a_204_47.n1 a_204_47.t3 313.663
R38 a_204_47.n1 a_204_47.n0 262.096
R39 a_204_47.t2 a_204_47.n1 209.923
R40 a_204_47.n0 a_204_47.t0 24.9236
R41 a_204_47.n0 a_204_47.t1 24.9236
R42 VNB.t0 VNB.t3 2677.02
R43 VNB.t1 VNB.t2 1352.75
R44 VNB.t3 VNB.t4 1196.12
R45 VNB.t2 VNB.t0 1196.12
R46 VNB VNB.t1 911.327
R47 TE.n2 TE.t0 322.94
R48 TE.n0 TE.t2 263.493
R49 TE.n1 TE.t3 189.588
R50 TE.n3 TE.n2 173.91
R51 TE.n0 TE.t1 128.534
R52 TE.n1 TE.n0 128.534
R53 TE.n2 TE.n1 40.1672
R54 TE.n3 TE 14.8903
R55 TE TE.n3 2.87397
R56 VGND.n1 VGND.t0 287.022
R57 VGND.n1 VGND.n0 190.831
R58 VGND.n0 VGND.t2 47.1434
R59 VGND.n0 VGND.t1 33.0774
R60 VGND VGND.n1 0.514329
C0 VGND TE 0.048679f
C1 Z A 0.122693f
C2 A VPWR 0.019617f
C3 VGND A 0.022759f
C4 Z VPWR 0.009749f
C5 Z VGND 0.009975f
C6 VGND VPWR 0.062104f
C7 VPB TE 0.107428f
C8 VPB A 0.07437f
C9 Z VPB 0.005146f
C10 VPB VPWR 0.07323f
C11 TE A 0.004934f
C12 Z TE 0.001007f
C13 VGND VPB 0.006901f
C14 TE VPWR 0.021524f
C15 VGND VNB 0.386303f
C16 Z VNB 0.013872f
C17 VPWR VNB 0.321877f
C18 A VNB 0.265273f
C19 TE VNB 0.343821f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_4 VPWR VGND VPB VNB TE Z A
X0 VPWR.t4 a_27_47.t2 a_215_309.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.2444 ps=2.4 w=0.94 l=0.15
X1 a_215_309.t3 A.t0 Z.t6 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t3 TE.t0 a_193_47.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X3 Z.t2 A.t1 a_193_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Z.t1 A.t2 a_193_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_193_47.t6 TE.t1 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Z.t5 A.t3 a_215_309.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16025 ps=1.325 w=1 l=0.15
X7 a_193_47.t5 TE.t2 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_193_47.t1 A.t4 Z.t7 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_193_47.t0 A.t5 Z.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t0 TE.t3 a_193_47.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_215_309.t6 a_27_47.t3 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.16025 pd=1.325 as=0.1269 ps=1.21 w=0.94 l=0.15
X12 VPWR.t2 a_27_47.t4 a_215_309.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X13 a_215_309.t4 a_27_47.t5 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X14 a_215_309.t1 A.t6 Z.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t0 TE.t4 a_27_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X16 Z.t3 A.t7 a_215_309.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t4 TE.t5 a_27_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t0 a_27_47.n3 771.813
R1 a_27_47.n0 a_27_47.t2 310.087
R2 a_27_47.n3 a_27_47.n2 261.25
R3 a_27_47.n3 a_27_47.t1 258.488
R4 a_27_47.n2 a_27_47.t3 188.517
R5 a_27_47.n1 a_27_47.t4 175.127
R6 a_27_47.n0 a_27_47.t5 175.127
R7 a_27_47.n1 a_27_47.n0 134.96
R8 a_27_47.n2 a_27_47.n1 72.3005
R9 a_215_309.n1 a_215_309.t7 848.899
R10 a_215_309.n3 a_215_309.t1 380.67
R11 a_215_309.n1 a_215_309.n0 316.457
R12 a_215_309.n3 a_215_309.n2 298.673
R13 a_215_309.n5 a_215_309.n4 286.329
R14 a_215_309.n4 a_215_309.n1 95.5466
R15 a_215_309.n4 a_215_309.n3 77.476
R16 a_215_309.n5 a_215_309.t6 34.5803
R17 a_215_309.n0 a_215_309.t5 28.2931
R18 a_215_309.n0 a_215_309.t4 28.2931
R19 a_215_309.n2 a_215_309.t2 26.5955
R20 a_215_309.n2 a_215_309.t3 26.5955
R21 a_215_309.n6 a_215_309.t0 24.357
R22 a_215_309.n7 a_215_309.n6 23.6405
R23 a_215_309.n6 a_215_309.n5 7.33561
R24 VPWR.n6 VPWR.t0 867.492
R25 VPWR.n2 VPWR.n1 313.512
R26 VPWR.n4 VPWR.n3 309.726
R27 VPWR.n3 VPWR.t1 28.2931
R28 VPWR.n3 VPWR.t4 28.2931
R29 VPWR.n1 VPWR.t3 28.2931
R30 VPWR.n1 VPWR.t2 28.2931
R31 VPWR.n5 VPWR.n4 22.9652
R32 VPWR.n6 VPWR.n5 20.7064
R33 VPWR.n5 VPWR.n0 9.3005
R34 VPWR.n7 VPWR.n6 7.12063
R35 VPWR.n4 VPWR.n2 6.4669
R36 VPWR.n2 VPWR.n0 0.65503
R37 VPWR.n7 VPWR.n0 0.148519
R38 VPWR VPWR.n7 0.11354
R39 VPB.t4 VPB.t8 556.386
R40 VPB.t7 VPB.t0 281.154
R41 VPB.t2 VPB.t1 248.599
R42 VPB.t3 VPB.t2 248.599
R43 VPB.t0 VPB.t3 248.599
R44 VPB.t6 VPB.t7 248.599
R45 VPB.t5 VPB.t6 248.599
R46 VPB.t8 VPB.t5 248.599
R47 VPB VPB.t4 189.409
R48 A.n2 A.t6 235.148
R49 A.n4 A.t7 221.72
R50 A.n6 A.t0 212.081
R51 A.n5 A.t3 212.081
R52 A.n2 A.t5 162.847
R53 A.n2 A.n1 152
R54 A.n3 A.n0 152
R55 A.n8 A.n7 152
R56 A.n4 A.t2 149.421
R57 A.n6 A.t4 139.78
R58 A.n5 A.t1 139.78
R59 A.n6 A.n5 61.346
R60 A.n7 A.n6 58.2625
R61 A.n4 A.n3 46.4153
R62 A.n8 A.n0 17.0672
R63 A.n3 A.n2 15.1746
R64 A.n7 A.n4 14.282
R65 A.n1 A 13.8044
R66 A.n1 A 9.28677
R67 A A.n0 3.26325
R68 A A.n8 2.76128
R69 Z Z.n1 312.416
R70 Z.n2 Z.n0 298.45
R71 Z.n5 Z.n3 222.883
R72 Z.n5 Z.n4 185
R73 Z.n0 Z.t6 26.5955
R74 Z.n0 Z.t5 26.5955
R75 Z.n1 Z.t4 26.5955
R76 Z.n1 Z.t3 26.5955
R77 Z.n4 Z.t7 24.9236
R78 Z.n4 Z.t2 24.9236
R79 Z.n3 Z.t0 24.9236
R80 Z.n3 Z.t1 24.9236
R81 Z.n2 Z 21.0829
R82 Z Z.n2 2.86366
R83 Z Z.n5 0.168921
R84 TE.n4 TE.t4 265.101
R85 TE.n0 TE.t3 263.493
R86 TE.n5 TE.n4 173.91
R87 TE.n3 TE.t5 152.633
R88 TE.n2 TE.n1 141.387
R89 TE.n1 TE.n0 134.96
R90 TE.n2 TE.t2 128.534
R91 TE.n1 TE.t0 128.534
R92 TE.n0 TE.t1 128.534
R93 TE.n3 TE.n2 110.861
R94 TE.n4 TE.n3 40.1672
R95 TE.n5 TE 14.8903
R96 TE TE.n5 2.87397
R97 a_193_47.n4 a_193_47.t0 321.914
R98 a_193_47.n2 a_193_47.n1 257.283
R99 a_193_47.t3 a_193_47.n5 209.923
R100 a_193_47.n2 a_193_47.n0 194.036
R101 a_193_47.n4 a_193_47.n3 185
R102 a_193_47.n5 a_193_47.n2 67.5605
R103 a_193_47.n5 a_193_47.n4 53.8792
R104 a_193_47.n1 a_193_47.t5 28.6159
R105 a_193_47.n1 a_193_47.t7 24.9236
R106 a_193_47.n0 a_193_47.t4 24.9236
R107 a_193_47.n0 a_193_47.t6 24.9236
R108 a_193_47.n3 a_193_47.t2 24.9236
R109 a_193_47.n3 a_193_47.t1 24.9236
R110 VGND.n1 VGND.t0 289.212
R111 VGND.n3 VGND.n2 198.964
R112 VGND.n6 VGND.n5 198.964
R113 VGND.n2 VGND.t2 24.9236
R114 VGND.n2 VGND.t3 24.9236
R115 VGND.n5 VGND.t1 24.9236
R116 VGND.n5 VGND.t4 24.9236
R117 VGND.n6 VGND.n4 22.9652
R118 VGND.n4 VGND.n3 16.9417
R119 VGND.n4 VGND.n0 9.3005
R120 VGND.n7 VGND.n6 7.12063
R121 VGND.n3 VGND.n1 6.71591
R122 VGND.n1 VGND.n0 0.699298
R123 VGND.n7 VGND.n0 0.148519
R124 VGND VGND.n7 0.11354
R125 VNB.t5 VNB.t3 2776.7
R126 VNB.t6 VNB.t8 1253.07
R127 VNB.t2 VNB.t0 1196.12
R128 VNB.t1 VNB.t2 1196.12
R129 VNB.t3 VNB.t1 1196.12
R130 VNB.t7 VNB.t5 1196.12
R131 VNB.t8 VNB.t7 1196.12
R132 VNB.t4 VNB.t6 1196.12
R133 VNB VNB.t4 911.327
C0 VGND A 0.034434f
C1 VGND VPWR 0.096829f
C2 VGND Z 0.025679f
C3 VPB TE 0.072689f
C4 VPB A 0.134147f
C5 VPB VPWR 0.104071f
C6 TE A 0.004655f
C7 TE VPWR 0.022881f
C8 VPB Z 0.008834f
C9 A VPWR 0.031926f
C10 TE Z 9.28e-19
C11 A Z 0.287773f
C12 VPWR Z 0.020604f
C13 VGND VPB 0.00831f
C14 VGND TE 0.075224f
C15 VGND VNB 0.567203f
C16 Z VNB 0.026655f
C17 VPWR VNB 0.470273f
C18 A VNB 0.422286f
C19 TE VNB 0.428395f
C20 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_8 VPWR VGND VPB VNB A Z TE
X0 VPWR.t7 a_27_47.t2 a_215_309.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.2444 ps=2.4 w=0.94 l=0.15
X1 a_215_309.t15 A.t0 Z.t7 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_47.t7 A.t1 Z.t15 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_215_309.t13 a_27_47.t3 VPWR.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.16025 pd=1.325 as=0.1269 ps=1.21 w=0.94 l=0.15
X4 Z.t6 A.t2 a_215_309.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t7 TE.t0 a_193_47.t12 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X6 a_215_309.t1 A.t3 Z.t5 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t5 a_27_47.t4 a_215_309.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X8 a_215_309.t11 a_27_47.t5 VPWR.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X9 Z.t4 A.t4 a_215_309.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_193_47.t13 TE.t1 VGND.t6 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Z.t14 A.t5 a_193_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_193_47.t14 TE.t2 VGND.t5 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_193_47.t15 TE.t3 VGND.t4 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_193_47.t11 TE.t4 VGND.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_193_47.t5 A.t6 Z.t13 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_193_47.t4 A.t7 Z.t12 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_193_47.t3 A.t8 Z.t11 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_215_309.t3 A.t9 Z.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t2 TE.t5 a_193_47.t10 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VPWR.t3 a_27_47.t6 a_215_309.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X21 VGND.t1 TE.t6 a_193_47.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND.t0 TE.t7 a_193_47.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Z.t2 A.t10 a_215_309.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Z.t10 A.t11 a_193_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_215_309.t9 a_27_47.t7 VPWR.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X26 Z.t1 A.t12 a_215_309.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16025 ps=1.325 w=1 l=0.15
X27 a_215_309.t6 A.t13 Z.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Z.t9 A.t14 a_193_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VPWR.t1 a_27_47.t8 a_215_309.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X30 Z.t8 A.t15 a_193_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_215_309.t7 a_27_47.t9 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X32 VPWR.t8 TE.t8 a_27_47.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X33 VGND.t8 TE.t9 a_27_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t0 a_27_47.n7 771.813
R1 a_27_47.n7 a_27_47.n6 326.413
R2 a_27_47.n0 a_27_47.t2 310.087
R3 a_27_47.n7 a_27_47.t1 258.488
R4 a_27_47.n6 a_27_47.t3 188.517
R5 a_27_47.n5 a_27_47.t4 175.127
R6 a_27_47.n4 a_27_47.t5 175.127
R7 a_27_47.n3 a_27_47.t6 175.127
R8 a_27_47.n2 a_27_47.t7 175.127
R9 a_27_47.n1 a_27_47.t8 175.127
R10 a_27_47.n0 a_27_47.t9 175.127
R11 a_27_47.n5 a_27_47.n4 134.96
R12 a_27_47.n4 a_27_47.n3 134.96
R13 a_27_47.n3 a_27_47.n2 134.96
R14 a_27_47.n2 a_27_47.n1 134.96
R15 a_27_47.n1 a_27_47.n0 134.96
R16 a_27_47.n6 a_27_47.n5 72.3005
R17 a_215_309.n5 a_215_309.t14 848.899
R18 a_215_309.n12 a_215_309.t15 382.825
R19 a_215_309.n7 a_215_309.n2 316.457
R20 a_215_309.n6 a_215_309.n3 316.457
R21 a_215_309.n5 a_215_309.n4 316.457
R22 a_215_309.n13 a_215_309.n12 298.675
R23 a_215_309.n10 a_215_309.n1 298.673
R24 a_215_309.n11 a_215_309.n0 298.673
R25 a_215_309.n9 a_215_309.n8 287.745
R26 a_215_309.n9 a_215_309.n7 84.5663
R27 a_215_309.n10 a_215_309.n9 70.913
R28 a_215_309.n7 a_215_309.n6 63.2476
R29 a_215_309.n6 a_215_309.n5 63.2476
R30 a_215_309.n12 a_215_309.n11 63.2476
R31 a_215_309.n11 a_215_309.n10 63.2476
R32 a_215_309.n8 a_215_309.t13 34.5803
R33 a_215_309.n8 a_215_309.t5 31.6921
R34 a_215_309.n2 a_215_309.t12 28.2931
R35 a_215_309.n2 a_215_309.t11 28.2931
R36 a_215_309.n3 a_215_309.t10 28.2931
R37 a_215_309.n3 a_215_309.t9 28.2931
R38 a_215_309.n4 a_215_309.t8 28.2931
R39 a_215_309.n4 a_215_309.t7 28.2931
R40 a_215_309.n1 a_215_309.t4 26.5955
R41 a_215_309.n1 a_215_309.t6 26.5955
R42 a_215_309.n0 a_215_309.t2 26.5955
R43 a_215_309.n0 a_215_309.t3 26.5955
R44 a_215_309.t0 a_215_309.n13 26.5955
R45 a_215_309.n13 a_215_309.t1 26.5955
R46 VPWR.n16 VPWR.t8 867.492
R47 VPWR.n6 VPWR.n5 315.265
R48 VPWR.n14 VPWR.n2 309.726
R49 VPWR.n4 VPWR.n3 309.726
R50 VPWR.n8 VPWR.n7 309.726
R51 VPWR.n2 VPWR.t0 28.2931
R52 VPWR.n2 VPWR.t7 28.2931
R53 VPWR.n3 VPWR.t2 28.2931
R54 VPWR.n3 VPWR.t1 28.2931
R55 VPWR.n7 VPWR.t4 28.2931
R56 VPWR.n7 VPWR.t3 28.2931
R57 VPWR.n5 VPWR.t6 28.2931
R58 VPWR.n5 VPWR.t5 28.2931
R59 VPWR.n9 VPWR.n4 27.4829
R60 VPWR.n15 VPWR.n14 22.9652
R61 VPWR.n14 VPWR.n13 21.4593
R62 VPWR.n16 VPWR.n15 20.7064
R63 VPWR.n13 VPWR.n4 16.9417
R64 VPWR.n9 VPWR.n8 10.9181
R65 VPWR.n10 VPWR.n9 9.3005
R66 VPWR.n11 VPWR.n4 9.3005
R67 VPWR.n13 VPWR.n12 9.3005
R68 VPWR.n14 VPWR.n1 9.3005
R69 VPWR.n15 VPWR.n0 9.3005
R70 VPWR.n17 VPWR.n16 7.12063
R71 VPWR.n8 VPWR.n6 6.68181
R72 VPWR.n10 VPWR.n6 0.975011
R73 VPWR.n17 VPWR.n0 0.148519
R74 VPWR.n11 VPWR.n10 0.120292
R75 VPWR.n12 VPWR.n11 0.120292
R76 VPWR.n12 VPWR.n1 0.120292
R77 VPWR.n1 VPWR.n0 0.120292
R78 VPWR VPWR.n17 0.11354
R79 VPB.t15 VPB.t14 556.386
R80 VPB.t13 VPB.t5 281.154
R81 VPB.t0 VPB.t16 248.599
R82 VPB.t1 VPB.t0 248.599
R83 VPB.t2 VPB.t1 248.599
R84 VPB.t3 VPB.t2 248.599
R85 VPB.t4 VPB.t3 248.599
R86 VPB.t6 VPB.t4 248.599
R87 VPB.t5 VPB.t6 248.599
R88 VPB.t12 VPB.t13 248.599
R89 VPB.t11 VPB.t12 248.599
R90 VPB.t10 VPB.t11 248.599
R91 VPB.t9 VPB.t10 248.599
R92 VPB.t8 VPB.t9 248.599
R93 VPB.t7 VPB.t8 248.599
R94 VPB.t14 VPB.t7 248.599
R95 VPB VPB.t15 189.409
R96 A.n1 A.t0 234.392
R97 A.n14 A.t9 221.72
R98 A.n8 A.t10 221.72
R99 A.n5 A.t2 221.72
R100 A.n10 A.t13 212.081
R101 A.n9 A.t12 212.081
R102 A.n19 A.t3 212.081
R103 A.n7 A.t4 212.081
R104 A.n1 A.t1 162.091
R105 A A.n11 157.272
R106 A.n2 A.n1 152
R107 A.n4 A.n3 152
R108 A.n6 A.n0 152
R109 A.n21 A.n20 152
R110 A.n18 A.n17 152
R111 A.n16 A.n15 152
R112 A.n13 A.n12 152
R113 A.n14 A.t7 149.421
R114 A.n8 A.t11 149.421
R115 A.n5 A.t15 149.421
R116 A.n10 A.t6 139.78
R117 A.n9 A.t5 139.78
R118 A.n19 A.t8 139.78
R119 A.n7 A.t14 139.78
R120 A.n10 A.n9 61.346
R121 A.n20 A.n6 58.9116
R122 A.n11 A.n10 58.2625
R123 A.n5 A.n4 49.9857
R124 A.n19 A.n18 46.7399
R125 A.n13 A.n8 46.4153
R126 A.n15 A.n7 40.4106
R127 A.n15 A.n14 32.1338
R128 A.n14 A.n13 28.5635
R129 A.n3 A.n2 17.0672
R130 A.n17 A.n16 17.0672
R131 A.n21 A 16.8162
R132 A.n18 A.n7 14.6066
R133 A.n11 A.n8 14.282
R134 A A.n0 12.2985
R135 A.n12 A 11.7966
R136 A.n4 A.n1 11.6042
R137 A.n12 A 11.2946
R138 A A.n0 10.7927
R139 A.n6 A.n5 10.7116
R140 A A.n21 6.27501
R141 A.n16 A 5.77305
R142 A.n3 A 4.76913
R143 A.n20 A.n19 2.92171
R144 A.n2 A 1.2554
R145 A.n17 A 0.25148
R146 Z.n10 Z.n9 298.863
R147 Z.n8 Z.n0 298.45
R148 Z.n12 Z.n11 292.406
R149 Z.n15 Z.n14 292.406
R150 Z.n3 Z.n1 235.01
R151 Z.n3 Z.n2 185
R152 Z.n5 Z.n4 185
R153 Z.n7 Z.n6 185
R154 Z.n5 Z.n3 50.0098
R155 Z.n7 Z.n5 37.8835
R156 Z Z.n8 33.1299
R157 Z.n13 Z 30.1181
R158 Z.n14 Z.t7 26.5955
R159 Z.n14 Z.t6 26.5955
R160 Z.n0 Z.t0 26.5955
R161 Z.n0 Z.t1 26.5955
R162 Z.n9 Z.t3 26.5955
R163 Z.n9 Z.t2 26.5955
R164 Z.n11 Z.t5 26.5955
R165 Z.n11 Z.t4 26.5955
R166 Z.n6 Z.t13 24.9236
R167 Z.n6 Z.t14 24.9236
R168 Z.n4 Z.t12 24.9236
R169 Z.n4 Z.t10 24.9236
R170 Z.n2 Z.t11 24.9236
R171 Z.n2 Z.t9 24.9236
R172 Z.n1 Z.t15 24.9236
R173 Z.n1 Z.t8 24.9236
R174 Z.n16 Z 24.0946
R175 Z Z.n7 23.0742
R176 Z Z.n13 14.3064
R177 Z Z.n10 8.28285
R178 Z.n13 Z.n12 6.46014
R179 Z.n16 Z.n15 6.46014
R180 Z.n12 Z 3.39383
R181 Z.n15 Z 3.39383
R182 Z.n10 Z 3.29747
R183 Z.n13 Z 3.29747
R184 Z Z.n16 3.29747
R185 Z.n8 Z 2.86366
R186 Z.n10 Z 1.50638
R187 Z.n8 Z 1.50638
R188 a_193_47.t7 a_193_47.n13 321.914
R189 a_193_47.n4 a_193_47.n3 257.283
R190 a_193_47.n7 a_193_47.t6 209.923
R191 a_193_47.n4 a_193_47.n2 194.036
R192 a_193_47.n5 a_193_47.n1 194.036
R193 a_193_47.n6 a_193_47.n0 194.036
R194 a_193_47.n13 a_193_47.n12 185
R195 a_193_47.n11 a_193_47.n10 185
R196 a_193_47.n9 a_193_47.n8 185
R197 a_193_47.n7 a_193_47.n6 66.4954
R198 a_193_47.n6 a_193_47.n5 63.2476
R199 a_193_47.n5 a_193_47.n4 63.2476
R200 a_193_47.n9 a_193_47.n7 53.6128
R201 a_193_47.n13 a_193_47.n11 51.2005
R202 a_193_47.n11 a_193_47.n9 51.2005
R203 a_193_47.n3 a_193_47.t11 28.6159
R204 a_193_47.n8 a_193_47.t2 24.9236
R205 a_193_47.n8 a_193_47.t5 24.9236
R206 a_193_47.n10 a_193_47.t1 24.9236
R207 a_193_47.n10 a_193_47.t4 24.9236
R208 a_193_47.n12 a_193_47.t0 24.9236
R209 a_193_47.n12 a_193_47.t3 24.9236
R210 a_193_47.n3 a_193_47.t12 24.9236
R211 a_193_47.n2 a_193_47.t10 24.9236
R212 a_193_47.n2 a_193_47.t13 24.9236
R213 a_193_47.n1 a_193_47.t8 24.9236
R214 a_193_47.n1 a_193_47.t14 24.9236
R215 a_193_47.n0 a_193_47.t9 24.9236
R216 a_193_47.n0 a_193_47.t15 24.9236
R217 VNB.t9 VNB.t6 2776.7
R218 VNB.t12 VNB.t13 1253.07
R219 VNB.t0 VNB.t7 1196.12
R220 VNB.t3 VNB.t0 1196.12
R221 VNB.t1 VNB.t3 1196.12
R222 VNB.t4 VNB.t1 1196.12
R223 VNB.t2 VNB.t4 1196.12
R224 VNB.t5 VNB.t2 1196.12
R225 VNB.t6 VNB.t5 1196.12
R226 VNB.t16 VNB.t9 1196.12
R227 VNB.t8 VNB.t16 1196.12
R228 VNB.t15 VNB.t8 1196.12
R229 VNB.t11 VNB.t15 1196.12
R230 VNB.t14 VNB.t11 1196.12
R231 VNB.t13 VNB.t14 1196.12
R232 VNB.t10 VNB.t12 1196.12
R233 VNB VNB.t10 911.327
R234 TE.n8 TE.t8 265.101
R235 TE.n0 TE.t7 263.493
R236 TE.n9 TE.n8 173.91
R237 TE.n7 TE.t9 152.633
R238 TE.n6 TE.n5 141.387
R239 TE.n1 TE.n0 134.96
R240 TE.n2 TE.n1 134.96
R241 TE.n3 TE.n2 134.96
R242 TE.n4 TE.n3 134.96
R243 TE.n5 TE.n4 134.96
R244 TE.n6 TE.t4 128.534
R245 TE.n5 TE.t0 128.534
R246 TE.n4 TE.t1 128.534
R247 TE.n3 TE.t5 128.534
R248 TE.n2 TE.t2 128.534
R249 TE.n1 TE.t6 128.534
R250 TE.n0 TE.t3 128.534
R251 TE.n7 TE.n6 110.861
R252 TE.n8 TE.n7 40.1672
R253 TE.n9 TE 14.8903
R254 TE TE.n9 2.87397
R255 VGND.n4 VGND.t0 288.531
R256 VGND.n6 VGND.n5 198.964
R257 VGND.n9 VGND.n8 198.964
R258 VGND.n13 VGND.n2 198.964
R259 VGND.n16 VGND.n15 198.964
R260 VGND.n9 VGND.n7 33.5064
R261 VGND.n13 VGND.n1 27.4829
R262 VGND.n5 VGND.t4 24.9236
R263 VGND.n5 VGND.t1 24.9236
R264 VGND.n8 VGND.t5 24.9236
R265 VGND.n8 VGND.t2 24.9236
R266 VGND.n2 VGND.t6 24.9236
R267 VGND.n2 VGND.t7 24.9236
R268 VGND.n15 VGND.t3 24.9236
R269 VGND.n15 VGND.t8 24.9236
R270 VGND.n16 VGND.n14 22.9652
R271 VGND.n14 VGND.n13 16.9417
R272 VGND.n6 VGND.n4 11.2483
R273 VGND.n9 VGND.n1 10.9181
R274 VGND.n7 VGND.n3 9.3005
R275 VGND.n10 VGND.n9 9.3005
R276 VGND.n11 VGND.n1 9.3005
R277 VGND.n13 VGND.n12 9.3005
R278 VGND.n14 VGND.n0 9.3005
R279 VGND.n17 VGND.n16 7.12063
R280 VGND.n7 VGND.n6 4.89462
R281 VGND.n4 VGND.n3 1.30422
R282 VGND.n17 VGND.n0 0.148519
R283 VGND.n10 VGND.n3 0.120292
R284 VGND.n11 VGND.n10 0.120292
R285 VGND.n12 VGND.n11 0.120292
R286 VGND.n12 VGND.n0 0.120292
R287 VGND VGND.n17 0.11354
C0 VPB TE 0.074108f
C1 VPB A 0.261492f
C2 TE A 0.004655f
C3 VPB VPWR 0.155017f
C4 TE VPWR 0.025519f
C5 VPB Z 0.013586f
C6 VPB VGND 0.010304f
C7 TE Z 0.001157f
C8 A VPWR 0.062992f
C9 A Z 0.652786f
C10 TE VGND 0.122603f
C11 VPWR Z 0.040111f
C12 A VGND 0.067918f
C13 VPWR VGND 0.157639f
C14 Z VGND 0.045821f
C15 VGND VNB 0.880714f
C16 Z VNB 0.025406f
C17 VPWR VNB 0.734487f
C18 A VNB 0.791088f
C19 TE VNB 0.68091f
C20 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fa_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_1 VPB VNB VGND VPWR B COUT A CIN SUM
X0 a_76_199.t1 B.t0 a_208_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X1 VGND.t5 A.t0 a_382_47.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_738_413.t2 A.t1 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_1091_47.t0 CIN.t0 a_995_47.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 VPWR.t7 CIN.t1 a_738_413.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_382_413.t1 B.t1 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR.t4 A.t2 a_382_413.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_995_47.t0 a_76_199.t4 a_738_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X8 a_382_413.t0 CIN.t2 a_76_199.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 SUM.t1 a_995_47.t4 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10235 ps=0.995 w=0.65 l=0.15
X10 a_208_47.t0 A.t3 VGND.t4 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.10235 ps=0.995 w=0.42 l=0.15
X11 VGND.t7 CIN.t3 a_738_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_76_199.t2 B.t2 a_208_413.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X13 a_208_413.t1 A.t4 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.14785 ps=1.345 w=0.42 l=0.15
X14 a_738_413.t1 B.t3 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VGND A a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10235 pd=0.995 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_738_47.t2 B.t4 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 a_738_47.t3 A.t5 VGND.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR A a_1163_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14785 pd=1.345 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_382_47.t0 CIN.t4 a_76_199.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_382_47.t1 B.t5 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 SUM.t0 a_995_47.t5 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14785 ps=1.345 w=1 l=0.15
X22 a_995_47.t1 a_76_199.t5 a_738_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X23 VPWR.t0 a_76_199.t6 COUT.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14785 pd=1.345 as=0.26 ps=2.52 w=1 l=0.15
X24 a_1091_413.t0 CIN.t5 a_995_47.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 VGND.t0 a_76_199.t7 COUT.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10235 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n0 B.t0 384.529
R1 B.n3 B.n2 373.283
R2 B.n5 B.t5 351.861
R3 B.n4 B.t1 297.233
R4 B.n6 B.n5 214.362
R5 B.n7 B.n3 167.825
R6 B.n3 B.n1 167.63
R7 B.n7 B.n6 163.79
R8 B.n8 B.n0 157.921
R9 B.n0 B.t2 156.382
R10 B.n5 B.t4 109.215
R11 B.n4 B.t3 102.659
R12 B.n6 B.n4 47.4474
R13 B.n8 B.n7 10.8599
R14 B B.n8 2.7205
R15 a_208_47.t0 a_208_47.t1 85.7148
R16 a_76_199.n3 a_76_199.n1 661.067
R17 a_76_199.n0 a_76_199.t5 373.283
R18 a_76_199.n2 a_76_199.t6 241.536
R19 a_76_199.n4 a_76_199.n0 189.024
R20 a_76_199.n5 a_76_199.n4 185.815
R21 a_76_199.n2 a_76_199.t7 169.237
R22 a_76_199.n0 a_76_199.t4 167.63
R23 a_76_199.n3 a_76_199.n2 152
R24 a_76_199.n4 a_76_199.n3 72.1596
R25 a_76_199.n1 a_76_199.t3 63.3219
R26 a_76_199.n1 a_76_199.t2 63.3219
R27 a_76_199.t0 a_76_199.n5 38.5719
R28 a_76_199.n5 a_76_199.t1 38.5719
R29 VNB.t10 VNB.t4 3801.94
R30 VNB.t6 VNB.t7 2677.02
R31 VNB.t2 VNB.t0 1409.71
R32 VNB.t3 VNB.t10 1366.99
R33 VNB.t0 VNB.t8 1281.55
R34 VNB.t5 VNB.t3 1267.31
R35 VNB.t11 VNB.t5 1196.12
R36 VNB.t7 VNB.t11 1196.12
R37 VNB.t9 VNB.t6 1196.12
R38 VNB.t1 VNB.t9 1196.12
R39 VNB.t8 VNB.t1 1196.12
R40 VNB VNB.t2 911.327
R41 A.n3 A.t1 373.283
R42 A.n2 A.n0 347.577
R43 A.n7 A.t4 334.723
R44 A.n5 A.t2 323.476
R45 A.n5 A.t0 217.436
R46 A.n7 A.t3 206.19
R47 A.n2 A.n1 193.337
R48 A.n6 A.n5 169.833
R49 A.n3 A.t5 167.63
R50 A.n4 A.n2 166.843
R51 A.n4 A.n3 166.421
R52 A.n8 A.n7 152
R53 A.n8 A.n6 11.595
R54 A A.n8 2.13383
R55 A.n6 A.n4 1.55989
R56 a_382_47.n0 a_382_47.t1 497.418
R57 a_382_47.n0 a_382_47.t2 38.5719
R58 a_382_47.t0 a_382_47.n0 38.5719
R59 VGND.n6 VGND.t1 252.518
R60 VGND.n9 VGND.t3 239.281
R61 VGND.n19 VGND.n18 199.739
R62 VGND.n5 VGND.n4 198.964
R63 VGND.n12 VGND.n11 198.964
R64 VGND.n18 VGND.t4 60.0005
R65 VGND.n4 VGND.t6 38.5719
R66 VGND.n4 VGND.t7 38.5719
R67 VGND.n11 VGND.t2 38.5719
R68 VGND.n11 VGND.t5 38.5719
R69 VGND.n16 VGND.n1 34.6358
R70 VGND.n17 VGND.n16 34.6358
R71 VGND.n12 VGND.n10 27.1064
R72 VGND.n9 VGND.n3 25.6005
R73 VGND.n18 VGND.t0 25.4291
R74 VGND.n19 VGND.n17 22.9652
R75 VGND.n10 VGND.n9 18.824
R76 VGND.n12 VGND.n1 17.3181
R77 VGND.n5 VGND.n3 12.8005
R78 VGND.n7 VGND.n3 9.3005
R79 VGND.n9 VGND.n8 9.3005
R80 VGND.n10 VGND.n2 9.3005
R81 VGND.n13 VGND.n12 9.3005
R82 VGND.n14 VGND.n1 9.3005
R83 VGND.n16 VGND.n15 9.3005
R84 VGND.n17 VGND.n0 9.3005
R85 VGND.n6 VGND.n5 7.49061
R86 VGND.n20 VGND.n19 7.12063
R87 VGND.n7 VGND.n6 0.154139
R88 VGND.n20 VGND.n0 0.148519
R89 VGND.n8 VGND.n7 0.120292
R90 VGND.n8 VGND.n2 0.120292
R91 VGND.n13 VGND.n2 0.120292
R92 VGND.n14 VGND.n13 0.120292
R93 VGND.n15 VGND.n14 0.120292
R94 VGND.n15 VGND.n0 0.120292
R95 VGND VGND.n20 0.11354
R96 VPWR.n11 VPWR.t3 663.062
R97 VPWR.n8 VPWR.t1 632.74
R98 VPWR.n19 VPWR.n1 605.481
R99 VPWR.n13 VPWR.n4 598.965
R100 VPWR.n7 VPWR.n6 598.965
R101 VPWR.n1 VPWR.t6 98.5005
R102 VPWR.n4 VPWR.t2 63.3219
R103 VPWR.n4 VPWR.t4 63.3219
R104 VPWR.n6 VPWR.t5 63.3219
R105 VPWR.n6 VPWR.t7 63.3219
R106 VPWR.n17 VPWR.n2 34.6358
R107 VPWR.n18 VPWR.n17 34.6358
R108 VPWR.n19 VPWR.n18 28.9887
R109 VPWR.n1 VPWR.t0 27.9557
R110 VPWR.n13 VPWR.n12 27.1064
R111 VPWR.n11 VPWR.n10 25.6005
R112 VPWR.n12 VPWR.n11 18.824
R113 VPWR.n13 VPWR.n2 17.3181
R114 VPWR.n10 VPWR.n7 12.8005
R115 VPWR.n10 VPWR.n9 9.3005
R116 VPWR.n11 VPWR.n5 9.3005
R117 VPWR.n12 VPWR.n3 9.3005
R118 VPWR.n14 VPWR.n13 9.3005
R119 VPWR.n15 VPWR.n2 9.3005
R120 VPWR.n17 VPWR.n16 9.3005
R121 VPWR.n18 VPWR.n0 9.3005
R122 VPWR.n8 VPWR.n7 7.49285
R123 VPWR.n20 VPWR.n19 7.12063
R124 VPWR.n9 VPWR.n8 0.151895
R125 VPWR.n20 VPWR.n0 0.148519
R126 VPWR.n9 VPWR.n5 0.120292
R127 VPWR.n5 VPWR.n3 0.120292
R128 VPWR.n14 VPWR.n3 0.120292
R129 VPWR.n15 VPWR.n14 0.120292
R130 VPWR.n16 VPWR.n15 0.120292
R131 VPWR.n16 VPWR.n0 0.120292
R132 VPWR VPWR.n20 0.11354
R133 a_738_413.n1 a_738_413.n0 1258.85
R134 a_738_413.t0 a_738_413.n1 75.0481
R135 a_738_413.n0 a_738_413.t3 63.3219
R136 a_738_413.n0 a_738_413.t1 63.3219
R137 a_738_413.n1 a_738_413.t2 63.3219
R138 VPB.t0 VPB.t3 790.188
R139 VPB.t6 VPB.t4 556.386
R140 VPB.t1 VPB.t7 292.991
R141 VPB.t2 VPB.t0 284.113
R142 VPB.t7 VPB.t5 266.356
R143 VPB.t9 VPB.t2 263.397
R144 VPB.t10 VPB.t9 248.599
R145 VPB.t4 VPB.t10 248.599
R146 VPB.t8 VPB.t6 248.599
R147 VPB.t11 VPB.t8 248.599
R148 VPB.t5 VPB.t11 248.599
R149 VPB VPB.t1 189.409
R150 CIN.n3 CIN.t0 373.283
R151 CIN.n2 CIN.n0 357.442
R152 CIN.n1 CIN.t3 346.022
R153 CIN.n0 CIN.t2 325.082
R154 CIN.n0 CIN.t4 215.829
R155 CIN.n1 CIN.t1 193.337
R156 CIN.n3 CIN.t5 167.63
R157 CIN.n2 CIN.n1 152
R158 CIN.n4 CIN.n3 152
R159 CIN.n4 CIN.n2 88.4259
R160 CIN CIN.n4 5.3765
R161 a_995_47.n2 a_995_47.n0 712.774
R162 a_995_47.n3 a_995_47.n2 303.64
R163 a_995_47.n1 a_995_47.t5 241.536
R164 a_995_47.n1 a_995_47.t4 169.237
R165 a_995_47.n2 a_995_47.n1 152
R166 a_995_47.n0 a_995_47.t1 91.4648
R167 a_995_47.n0 a_995_47.t2 63.3219
R168 a_995_47.t0 a_995_47.n3 55.7148
R169 a_995_47.n3 a_995_47.t3 38.5719
R170 a_382_413.n0 a_382_413.t1 1316.86
R171 a_382_413.n0 a_382_413.t2 63.3219
R172 a_382_413.t0 a_382_413.n0 63.3219
R173 a_738_47.n1 a_738_47.n0 458.848
R174 a_738_47.t0 a_738_47.n1 45.7148
R175 a_738_47.n0 a_738_47.t1 38.5719
R176 a_738_47.n0 a_738_47.t2 38.5719
R177 a_738_47.n1 a_738_47.t3 38.5719
R178 SUM.t0 SUM 758.202
R179 SUM.n1 SUM.t0 755.481
R180 SUM.n0 SUM.t1 209.923
R181 SUM.n3 SUM 11.4429
R182 SUM.n2 SUM.n1 8.8005
R183 SUM SUM.n0 6.5605
R184 SUM.n0 SUM 4.3205
R185 SUM SUM.n3 1.74595
R186 SUM SUM.n2 1.55202
R187 SUM.n3 SUM 1.4405
R188 SUM.n2 SUM 1.2805
R189 SUM.n1 SUM 0.8005
R190 a_208_413.t0 a_208_413.t1 140.714
R191 COUT COUT.t0 787.909
R192 COUT.n1 COUT.t0 744.115
R193 COUT.n0 COUT.t1 209.923
R194 COUT.n1 COUT.n0 75.4783
R195 COUT.n0 COUT 6.64665
R196 COUT COUT.n1 0.492808
C0 VPWR SUM 0.07457f
C1 VGND SUM 0.071274f
C2 A B 0.772692f
C3 VPB A 0.275133f
C4 a_1163_47# VGND 0.001753f
C5 A CIN 0.455174f
C6 VPB B 0.337167f
C7 a_1163_413# A 1.05e-19
C8 a_1163_47# SUM 2.86e-20
C9 A COUT 0.00345f
C10 B CIN 0.612022f
C11 VPB CIN 0.231534f
C12 a_1163_413# B 3.18e-19
C13 A VPWR 0.070501f
C14 B COUT 5.98e-19
C15 VPB COUT 0.010944f
C16 B VPWR 0.252869f
C17 A VGND 0.102674f
C18 VPB VPWR 0.156127f
C19 B VGND 0.045605f
C20 CIN VPWR 0.057695f
C21 A SUM 0.005403f
C22 VPB VGND 0.005193f
C23 a_1163_413# VPWR 7.42e-19
C24 B SUM 0.001114f
C25 CIN VGND 0.060425f
C26 COUT VPWR 0.066634f
C27 VPB SUM 0.017933f
C28 a_1163_47# A 7.66e-19
C29 COUT VGND 0.055667f
C30 a_1163_47# B 6.11e-20
C31 VPWR VGND 0.042632f
C32 SUM VNB 0.100307f
C33 VGND VNB 0.812356f
C34 VPWR VNB 0.669221f
C35 COUT VNB 0.094108f
C36 CIN VNB 0.325368f
C37 B VNB 0.471308f
C38 A VNB 0.495819f
C39 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fa_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_2 VPB VNB VGND VPWR A COUT B CIN SUM
X0 a_1171_369# CIN a_1086_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.103625 pd=0.965 as=0.088 ps=0.915 w=0.64 l=0.15
X1 VGND.t3 CIN.t0 a_829_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND.t1 a_1086_47# SUM.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X3 COUT.t1 a_80_21.t4 VPWR.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_829_369.t2 A.t0 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0944 pd=0.935 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VPWR.t5 CIN.t1 a_829_369.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 a_473_371.t1 B.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1638 pd=1.78 as=0.08505 ps=0.9 w=0.63 l=0.15
X7 a_294_47.t1 A.t1 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1034 ps=1 w=0.42 l=0.15
X8 VPWR.t8 A.t2 a_473_371.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.08505 pd=0.9 as=0.08505 ps=0.9 w=0.63 l=0.15
X9 a_829_369.t3 B.t1 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 a_829_47.t3 B.t2 VGND.t10 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_829_47.t1 A.t3 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_473_371.t0 CIN.t2 a_80_21.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.08505 pd=0.9 as=0.102375 ps=0.955 w=0.63 l=0.15
X13 a_473_47.t0 CIN.t3 a_80_21.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_473_47.t1 B.t3 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VPWR.t3 a_1086_47# SUM.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t9 a_80_21.t5 COUT.t3 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 COUT.t2 a_80_21.t6 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X18 SUM.t0 a_1086_47# VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148625 ps=1.325 w=1 l=0.15
X19 a_80_21.t3 B.t4 a_289_371.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.102375 pd=0.955 as=0.092925 ps=0.925 w=0.63 l=0.15
X20 a_80_21.t2 B.t5 a_294_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X21 VGND.t6 A.t4 a_473_47.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 SUM.t2 a_1086_47# VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10235 ps=0.995 w=0.65 l=0.15
X23 VPWR.t6 a_80_21.t7 COUT.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.148625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X24 a_289_371.t1 A.t5 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.092925 pd=0.925 as=0.148625 ps=1.325 w=0.63 l=0.15
X25 a_1194_47.t0 CIN.t4 a_1086_47# VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X26 a_1086_47# a_80_21.t8 a_829_47.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.06195 ps=0.715 w=0.42 l=0.15
X27 VGND.t2 A.t6 a_1266_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10235 pd=0.995 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1266_371.t0 B.t6 a_1171_369# VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.02 as=0.103625 ps=0.965 w=0.63 l=0.15
X29 VPWR.t0 A.t7 a_1266_371.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.148625 pd=1.325 as=0.12285 ps=1.02 w=0.63 l=0.15
X30 a_1266_47.t0 B.t7 a_1194_47.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 a_1086_47# a_80_21.t9 a_829_369.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.088 pd=0.915 as=0.0944 ps=0.935 w=0.64 l=0.15
R0 CIN.n2 CIN.n0 343.332
R1 CIN.n4 CIN.t4 321.87
R2 CIN.n1 CIN.t0 320.315
R3 CIN.n0 CIN.t2 291.342
R4 CIN.n0 CIN.t3 215.829
R5 CIN.n4 CIN.n3 183.696
R6 CIN.n1 CIN.t1 183.696
R7 CIN.n5 CIN.n4 156.096
R8 CIN.n2 CIN.n1 152
R9 CIN.n5 CIN.n2 84.872
R10 CIN CIN.n5 9.4725
R11 VPB.t2 VPB.t14 556.386
R12 VPB.t11 VPB.t9 532.711
R13 VPB.t9 VPB.t0 319.627
R14 VPB.t0 VPB.t3 281.154
R15 VPB.t10 VPB.t7 281.154
R16 VPB.t1 VPB.t6 281.154
R17 VPB.t13 VPB.t11 263.397
R18 VPB.t6 VPB.t10 263.397
R19 VPB.t3 VPB.t4 248.599
R20 VPB.t8 VPB.t13 248.599
R21 VPB.t14 VPB.t8 248.599
R22 VPB.t12 VPB.t2 248.599
R23 VPB.t7 VPB.t12 248.599
R24 VPB.t5 VPB.t1 248.599
R25 VPB VPB.t5 195.327
R26 a_829_47.n1 a_829_47.n0 458.848
R27 a_829_47.n0 a_829_47.t2 45.7148
R28 a_829_47.n0 a_829_47.t1 38.5719
R29 a_829_47.t0 a_829_47.n1 38.5719
R30 a_829_47.n1 a_829_47.t3 38.5719
R31 VGND.n12 VGND.t1 292.711
R32 VGND.n34 VGND.t8 282.565
R33 VGND.n22 VGND.t10 239.281
R34 VGND.n32 VGND.n2 199.739
R35 VGND.n11 VGND.n10 198.964
R36 VGND.n20 VGND.n8 198.964
R37 VGND.n26 VGND.n5 198.964
R38 VGND.n2 VGND.t9 48.2862
R39 VGND.n10 VGND.t0 46.8576
R40 VGND.n10 VGND.t2 38.5719
R41 VGND.n8 VGND.t5 38.5719
R42 VGND.n8 VGND.t3 38.5719
R43 VGND.n5 VGND.t4 38.5719
R44 VGND.n5 VGND.t6 38.5719
R45 VGND.n2 VGND.t7 38.5719
R46 VGND.n15 VGND.n14 34.6358
R47 VGND.n16 VGND.n15 34.6358
R48 VGND.n16 VGND.n7 34.6358
R49 VGND.n28 VGND.n27 34.6358
R50 VGND.n28 VGND.n1 34.6358
R51 VGND.n20 VGND.n7 32.0005
R52 VGND.n34 VGND.n33 32.0005
R53 VGND.n26 VGND.n4 27.4829
R54 VGND.n22 VGND.n21 25.977
R55 VGND.n33 VGND.n32 24.8476
R56 VGND.n32 VGND.n1 19.577
R57 VGND.n22 VGND.n4 18.4476
R58 VGND.n27 VGND.n26 16.9417
R59 VGND.n21 VGND.n20 12.424
R60 VGND.n35 VGND.n34 11.9358
R61 VGND.n14 VGND.n13 9.3005
R62 VGND.n15 VGND.n9 9.3005
R63 VGND.n17 VGND.n16 9.3005
R64 VGND.n18 VGND.n7 9.3005
R65 VGND.n20 VGND.n19 9.3005
R66 VGND.n21 VGND.n6 9.3005
R67 VGND.n23 VGND.n22 9.3005
R68 VGND.n24 VGND.n4 9.3005
R69 VGND.n26 VGND.n25 9.3005
R70 VGND.n27 VGND.n3 9.3005
R71 VGND.n29 VGND.n28 9.3005
R72 VGND.n30 VGND.n1 9.3005
R73 VGND.n32 VGND.n31 9.3005
R74 VGND.n33 VGND.n0 9.3005
R75 VGND.n12 VGND.n11 8.65317
R76 VGND.n14 VGND.n11 8.28285
R77 VGND.n13 VGND.n12 0.602713
R78 VGND.n13 VGND.n9 0.120292
R79 VGND.n17 VGND.n9 0.120292
R80 VGND.n18 VGND.n17 0.120292
R81 VGND.n19 VGND.n18 0.120292
R82 VGND.n19 VGND.n6 0.120292
R83 VGND.n23 VGND.n6 0.120292
R84 VGND.n24 VGND.n23 0.120292
R85 VGND.n25 VGND.n24 0.120292
R86 VGND.n25 VGND.n3 0.120292
R87 VGND.n29 VGND.n3 0.120292
R88 VGND.n30 VGND.n29 0.120292
R89 VGND.n31 VGND.n30 0.120292
R90 VGND.n31 VGND.n0 0.120292
R91 VGND.n35 VGND.n0 0.120292
R92 VGND VGND.n35 0.0226354
R93 VNB.t7 VNB.t15 2677.02
R94 VNB.t0 VNB.t1 1537.86
R95 VNB.t10 VNB.t3 1537.86
R96 VNB.t14 VNB.t11 1423.95
R97 VNB.t2 VNB.t0 1409.71
R98 VNB.t12 VNB.t2 1366.99
R99 VNB.t11 VNB.t6 1352.75
R100 VNB.t8 VNB.t10 1267.31
R101 VNB.t5 VNB.t8 1196.12
R102 VNB.t15 VNB.t5 1196.12
R103 VNB.t9 VNB.t7 1196.12
R104 VNB.t4 VNB.t9 1196.12
R105 VNB.t6 VNB.t4 1196.12
R106 VNB.t13 VNB.t14 1196.12
R107 VNB.t3 VNB.t12 1025.24
R108 VNB VNB.t13 939.807
R109 SUM SUM.n0 376.337
R110 SUM SUM.n1 135.415
R111 SUM.n1 SUM.t2 47.0774
R112 SUM.n0 SUM.t1 26.5955
R113 SUM.n0 SUM.t0 26.5955
R114 SUM.n1 SUM.t3 24.9236
R115 a_80_21.n7 a_80_21.n6 394.661
R116 a_80_21.n0 a_80_21.t9 337.937
R117 a_80_21.n3 a_80_21.t7 212.081
R118 a_80_21.n4 a_80_21.t4 212.081
R119 a_80_21.n2 a_80_21.n0 189.532
R120 a_80_21.n2 a_80_21.n1 185.786
R121 a_80_21.n6 a_80_21.n5 173.459
R122 a_80_21.n0 a_80_21.t8 167.63
R123 a_80_21.n3 a_80_21.t5 139.78
R124 a_80_21.n4 a_80_21.t6 139.78
R125 a_80_21.n6 a_80_21.n2 71.312
R126 a_80_21.n7 a_80_21.t3 59.4132
R127 a_80_21.t1 a_80_21.n7 42.2148
R128 a_80_21.n1 a_80_21.t0 38.5719
R129 a_80_21.n1 a_80_21.t2 38.5719
R130 a_80_21.n5 a_80_21.n4 33.5944
R131 a_80_21.n5 a_80_21.n3 27.752
R132 VPWR.n32 VPWR.n2 598.965
R133 VPWR.n26 VPWR.n5 598.965
R134 VPWR.n20 VPWR.n8 598.965
R135 VPWR.n13 VPWR.n11 598.965
R136 VPWR.n6 VPWR.t10 374.937
R137 VPWR.n12 VPWR.t3 362.296
R138 VPWR.n34 VPWR.t7 350.582
R139 VPWR.n11 VPWR.t0 57.8497
R140 VPWR.n2 VPWR.t4 46.9053
R141 VPWR.n2 VPWR.t6 43.9275
R142 VPWR.n5 VPWR.t1 42.2148
R143 VPWR.n5 VPWR.t8 42.2148
R144 VPWR.n8 VPWR.t9 41.5552
R145 VPWR.n8 VPWR.t5 41.5552
R146 VPWR.n27 VPWR.n3 34.6358
R147 VPWR.n31 VPWR.n3 34.6358
R148 VPWR.n15 VPWR.n14 34.6358
R149 VPWR.n15 VPWR.n9 34.6358
R150 VPWR.n19 VPWR.n9 34.6358
R151 VPWR.n11 VPWR.t2 32.9831
R152 VPWR.n34 VPWR.n33 32.0005
R153 VPWR.n20 VPWR.n19 32.0005
R154 VPWR.n26 VPWR.n25 27.4829
R155 VPWR.n21 VPWR.n6 25.977
R156 VPWR.n32 VPWR.n31 22.5887
R157 VPWR.n33 VPWR.n32 21.8358
R158 VPWR.n25 VPWR.n6 18.4476
R159 VPWR.n27 VPWR.n26 16.9417
R160 VPWR.n14 VPWR.n13 16.5652
R161 VPWR.n21 VPWR.n20 12.424
R162 VPWR.n35 VPWR.n34 11.9358
R163 VPWR.n14 VPWR.n10 9.3005
R164 VPWR.n16 VPWR.n15 9.3005
R165 VPWR.n17 VPWR.n9 9.3005
R166 VPWR.n19 VPWR.n18 9.3005
R167 VPWR.n20 VPWR.n7 9.3005
R168 VPWR.n22 VPWR.n21 9.3005
R169 VPWR.n23 VPWR.n6 9.3005
R170 VPWR.n25 VPWR.n24 9.3005
R171 VPWR.n26 VPWR.n4 9.3005
R172 VPWR.n28 VPWR.n27 9.3005
R173 VPWR.n29 VPWR.n3 9.3005
R174 VPWR.n31 VPWR.n30 9.3005
R175 VPWR.n32 VPWR.n1 9.3005
R176 VPWR.n33 VPWR.n0 9.3005
R177 VPWR.n13 VPWR.n12 6.60549
R178 VPWR.n12 VPWR.n10 0.892535
R179 VPWR.n16 VPWR.n10 0.120292
R180 VPWR.n17 VPWR.n16 0.120292
R181 VPWR.n18 VPWR.n17 0.120292
R182 VPWR.n18 VPWR.n7 0.120292
R183 VPWR.n22 VPWR.n7 0.120292
R184 VPWR.n23 VPWR.n22 0.120292
R185 VPWR.n24 VPWR.n23 0.120292
R186 VPWR.n24 VPWR.n4 0.120292
R187 VPWR.n28 VPWR.n4 0.120292
R188 VPWR.n29 VPWR.n28 0.120292
R189 VPWR.n30 VPWR.n29 0.120292
R190 VPWR.n30 VPWR.n1 0.120292
R191 VPWR.n1 VPWR.n0 0.120292
R192 VPWR.n35 VPWR.n0 0.120292
R193 VPWR VPWR.n35 0.0226354
R194 COUT.n1 COUT 595.668
R195 COUT.n2 COUT.n1 585
R196 COUT COUT.n0 291.382
R197 COUT.n1 COUT.t0 26.5955
R198 COUT.n1 COUT.t1 26.5955
R199 COUT.n0 COUT.t3 24.9236
R200 COUT.n0 COUT.t2 24.9236
R201 COUT.n2 COUT 10.0576
R202 COUT COUT.n3 10.0576
R203 COUT.n3 COUT 8.62091
R204 COUT.n3 COUT.n2 0.610024
R205 A.n1 A.t0 337.937
R206 A.n5 A.t5 300.983
R207 A.n0 A.t7 300.983
R208 A.n3 A.t2 289.736
R209 A.n3 A.t4 217.436
R210 A.n0 A.t6 206.19
R211 A.n5 A.t1 205.702
R212 A.n2 A.n0 188.26
R213 A.n4 A.n3 169.833
R214 A.n1 A.t3 167.63
R215 A.n2 A.n1 166.633
R216 A A.n5 160.915
R217 A A.n4 14.317
R218 A.n4 A.n2 1.55989
R219 a_829_369.n1 a_829_369.n0 1258.85
R220 a_829_369.n0 a_829_369.t1 49.2505
R221 a_829_369.n0 a_829_369.t2 41.5552
R222 a_829_369.t0 a_829_369.n1 41.5552
R223 a_829_369.n1 a_829_369.t3 41.5552
R224 B.n2 B.t3 393.634
R225 B.n1 B.t0 334.188
R226 B.n5 B.t5 325.082
R227 B.n0 B.t7 325.082
R228 B.n5 B.t4 182.089
R229 B.n0 B.t6 182.089
R230 B.n4 B.n0 180.215
R231 B.n3 B.n2 173.841
R232 B.n4 B.n3 162.333
R233 B B.n5 161.143
R234 B.n1 B.t1 136.567
R235 B.n2 B.t2 91.5805
R236 B.n3 B.n1 22.4938
R237 B B.n4 15.3007
R238 a_473_371.n0 a_473_371.t1 1285.37
R239 a_473_371.n0 a_473_371.t2 42.2148
R240 a_473_371.t0 a_473_371.n0 42.2148
R241 a_294_47.t0 a_294_47.t1 92.8576
R242 a_473_47.n0 a_473_47.t1 497.418
R243 a_473_47.n0 a_473_47.t2 38.5719
R244 a_473_47.t0 a_473_47.n0 38.5719
R245 a_289_371.t0 a_289_371.t1 92.2465
R246 a_1194_47.t0 a_1194_47.t1 60.0005
R247 a_1266_47.t0 a_1266_47.t1 94.2862
R248 a_1266_371.t0 a_1266_371.t1 121.953
C0 VPWR COUT 0.127521f
C1 CIN VGND 0.061194f
C2 B SUM 0.002429f
C3 a_1171_369# A 2.08e-19
C4 VPWR VGND 0.061913f
C5 a_1171_369# B 0.001729f
C6 a_1086_47# VGND 0.216712f
C7 COUT VGND 0.105281f
C8 VPWR SUM 0.124724f
C9 a_1171_369# CIN 0.001582f
C10 a_1086_47# SUM 0.224673f
C11 VPB A 0.217587f
C12 a_1171_369# VPWR 0.001873f
C13 a_1086_47# a_1171_369# 0.011019f
C14 VPB B 0.28077f
C15 VGND SUM 0.120969f
C16 A B 0.79112f
C17 VPB CIN 0.190565f
C18 A CIN 0.437816f
C19 VPB VPWR 0.175432f
C20 a_1086_47# VPB 0.07657f
C21 VPB COUT 0.008598f
C22 A VPWR 0.064029f
C23 B CIN 0.568663f
C24 a_1086_47# A 0.175657f
C25 B VPWR 0.295003f
C26 VPB VGND 0.00696f
C27 A COUT 0.004355f
C28 a_1086_47# B 0.113389f
C29 CIN VPWR 0.053148f
C30 B COUT 0.001424f
C31 VPB SUM 0.011848f
C32 A VGND 0.089193f
C33 a_1086_47# CIN 0.059656f
C34 A SUM 0.003473f
C35 B VGND 0.059878f
C36 a_1086_47# VPWR 0.246294f
C37 SUM VNB 0.058389f
C38 VGND VNB 0.931146f
C39 COUT VNB 0.055034f
C40 VPWR VNB 0.795994f
C41 CIN VNB 0.327197f
C42 B VNB 0.476923f
C43 A VNB 0.491159f
C44 VPB VNB 1.66792f
C45 a_1086_47# VNB 0.234165f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fa_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_4 VPB VNB VGND VPWR B CIN SUM COUT A
X0 a_1014_369# B.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 VPWR.t3 CIN.t0 a_1014_369# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 VPWR.t0 A.t0 a_658_369.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND.t2 A.t1 a_658_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_79_21.t1 B.t1 a_456_371.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1322 pd=1.055 as=0.092925 ps=0.925 w=0.63 l=0.15
X5 a_658_369.t2 CIN.t1 a_79_21.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1322 ps=1.055 w=0.64 l=0.15
X6 VPWR.t7 a_1271_47# SUM.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X7 a_461_47.t1 A.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1034 ps=1 w=0.42 l=0.15
X8 VPWR.t10 a_79_21.t4 COUT.t7 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.148625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X9 SUM.t6 a_1271_47# VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148625 ps=1.325 w=1 l=0.15
X10 a_658_47.t2 CIN.t2 a_79_21.t2 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0756 ps=0.78 w=0.42 l=0.15
X11 a_658_47.t0 B.t2 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 COUT.t6 a_79_21.t5 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_456_371.t1 A.t3 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.092925 pd=0.925 as=0.148625 ps=1.325 w=0.63 l=0.15
X14 a_1451_47# B a_1379_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 VPWR.t12 a_79_21.t6 COUT.t5 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t9 a_79_21.t7 COUT.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t10 a_79_21.t8 COUT.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t9 a_1271_47# SUM.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t6 a_1271_47# SUM.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X20 VGND.t5 a_1271_47# SUM.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_79_21.t0 B.t3 a_461_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.06825 ps=0.745 w=0.42 l=0.15
X22 a_1014_47# A.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 COUT.t1 a_79_21.t9 VGND.t11 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_658_369.t0 B.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 VPWR A a_1451_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148625 pd=1.325 as=0.12285 ps=1.02 w=0.63 l=0.15
X26 a_1014_47# B.t5 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_1379_47# CIN a_1271_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X28 VGND A a_1451_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11535 pd=1.035 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 SUM.t1 a_1271_47# VGND.t8 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_1356_369.t0 CIN.t3 a_1271_47# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.103625 pd=0.965 as=0.088 ps=0.915 w=0.64 l=0.15
X31 SUM.t0 a_1271_47# VGND.t7 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11535 ps=1.035 w=0.65 l=0.15
X32 SUM.t4 a_1271_47# VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X33 VGND.t13 CIN.t4 a_1014_47# VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X34 a_1014_369# A.t5 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0944 pd=0.935 as=0.0864 ps=0.91 w=0.64 l=0.15
X35 COUT.t4 a_79_21.t10 VPWR.t13 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 COUT.t0 a_79_21.t11 VGND.t12 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B.n4 B.t2 393.634
R1 B.n3 B.t4 332.58
R2 B.n7 B.t3 325.082
R3 B.n2 B.n1 325.082
R4 B.n7 B.t1 182.089
R5 B.n2 B.n0 182.089
R6 B.n6 B.n2 180.215
R7 B.n5 B.n4 173.841
R8 B B.n7 165.845
R9 B.n6 B.n5 162.333
R10 B.n3 B.t0 136.567
R11 B.n4 B.t5 91.5805
R12 B.n5 B.n3 22.4938
R13 B B.n6 15.3007
R14 VPWR.n18 VPWR.t6 826.271
R15 VPWR.n37 VPWR.n4 598.965
R16 VPWR.n31 VPWR.n7 598.965
R17 VPWR.n10 VPWR.n9 598.965
R18 VPWR.n29 VPWR.t2 374.937
R19 VPWR.n15 VPWR.t9 362.372
R20 VPWR.n44 VPWR.t13 350.582
R21 VPWR.n42 VPWR.n1 323.988
R22 VPWR.n16 VPWR.n14 323.988
R23 VPWR.n4 VPWR.t5 46.9053
R24 VPWR.n4 VPWR.t10 43.9275
R25 VPWR.n14 VPWR.t8 42.3555
R26 VPWR.n7 VPWR.t1 41.5552
R27 VPWR.n7 VPWR.t0 41.5552
R28 VPWR.n9 VPWR.t4 41.5552
R29 VPWR.n9 VPWR.t3 41.5552
R30 VPWR.n41 VPWR.n2 34.6358
R31 VPWR.n35 VPWR.n5 34.6358
R32 VPWR.n36 VPWR.n35 34.6358
R33 VPWR.n22 VPWR.n12 34.6358
R34 VPWR.n23 VPWR.n22 34.6358
R35 VPWR.n24 VPWR.n23 34.6358
R36 VPWR.n44 VPWR.n43 32.377
R37 VPWR.n24 VPWR.n10 31.624
R38 VPWR.n43 VPWR.n42 30.8711
R39 VPWR.n37 VPWR.n36 28.9887
R40 VPWR.n18 VPWR.n17 27.4829
R41 VPWR.n31 VPWR.n30 27.1064
R42 VPWR.n1 VPWR.t11 26.5955
R43 VPWR.n1 VPWR.t12 26.5955
R44 VPWR.n14 VPWR.t7 26.5955
R45 VPWR.n29 VPWR.n28 25.6005
R46 VPWR.n17 VPWR.n16 23.7181
R47 VPWR.n30 VPWR.n29 18.824
R48 VPWR.n16 VPWR.n15 17.888
R49 VPWR.n31 VPWR.n5 17.3181
R50 VPWR.n18 VPWR.n12 16.9417
R51 VPWR.n37 VPWR.n2 15.4358
R52 VPWR.n28 VPWR.n10 12.8005
R53 VPWR.n45 VPWR.n44 11.5593
R54 VPWR.n17 VPWR.n13 9.3005
R55 VPWR.n19 VPWR.n18 9.3005
R56 VPWR.n20 VPWR.n12 9.3005
R57 VPWR.n22 VPWR.n21 9.3005
R58 VPWR.n23 VPWR.n11 9.3005
R59 VPWR.n25 VPWR.n24 9.3005
R60 VPWR.n26 VPWR.n10 9.3005
R61 VPWR.n28 VPWR.n27 9.3005
R62 VPWR.n29 VPWR.n8 9.3005
R63 VPWR.n30 VPWR.n6 9.3005
R64 VPWR.n32 VPWR.n31 9.3005
R65 VPWR.n33 VPWR.n5 9.3005
R66 VPWR.n35 VPWR.n34 9.3005
R67 VPWR.n36 VPWR.n3 9.3005
R68 VPWR.n38 VPWR.n37 9.3005
R69 VPWR.n39 VPWR.n2 9.3005
R70 VPWR.n41 VPWR.n40 9.3005
R71 VPWR.n43 VPWR.n0 9.3005
R72 VPWR.n42 VPWR.n41 3.76521
R73 VPWR.n15 VPWR.n13 0.779653
R74 VPWR.n19 VPWR.n13 0.120292
R75 VPWR.n20 VPWR.n19 0.120292
R76 VPWR.n21 VPWR.n20 0.120292
R77 VPWR.n21 VPWR.n11 0.120292
R78 VPWR.n25 VPWR.n11 0.120292
R79 VPWR.n26 VPWR.n25 0.120292
R80 VPWR.n27 VPWR.n26 0.120292
R81 VPWR.n27 VPWR.n8 0.120292
R82 VPWR.n8 VPWR.n6 0.120292
R83 VPWR.n32 VPWR.n6 0.120292
R84 VPWR.n33 VPWR.n32 0.120292
R85 VPWR.n34 VPWR.n33 0.120292
R86 VPWR.n34 VPWR.n3 0.120292
R87 VPWR.n38 VPWR.n3 0.120292
R88 VPWR.n39 VPWR.n38 0.120292
R89 VPWR.n40 VPWR.n39 0.120292
R90 VPWR.n40 VPWR.n0 0.120292
R91 VPWR.n45 VPWR.n0 0.120292
R92 VPWR VPWR.n45 0.0213333
R93 VPB.t1 VPB.t11 881.932
R94 VPB.t2 VPB.t4 556.386
R95 VPB.t7 VPB.t1 514.953
R96 VPB.t3 VPB.t6 334.425
R97 VPB.t12 VPB.t9 295.95
R98 VPB.t13 VPB.t8 281.154
R99 VPB.t8 VPB.t3 263.397
R100 VPB.t9 VPB.t10 248.599
R101 VPB.t11 VPB.t12 248.599
R102 VPB.t5 VPB.t7 248.599
R103 VPB.t4 VPB.t5 248.599
R104 VPB.t0 VPB.t2 248.599
R105 VPB.t6 VPB.t0 248.599
R106 VPB.t14 VPB.t13 248.599
R107 VPB.t15 VPB.t14 248.599
R108 VPB.t16 VPB.t15 248.599
R109 VPB VPB.t16 189.409
R110 CIN.n2 CIN.n0 343.332
R111 CIN.n4 CIN.n3 321.87
R112 CIN.n1 CIN.t4 320.315
R113 CIN.n0 CIN.t1 289.736
R114 CIN.n0 CIN.t2 215.829
R115 CIN.n4 CIN.t3 183.696
R116 CIN.n1 CIN.t0 183.696
R117 CIN.n5 CIN.n4 156.096
R118 CIN.n2 CIN.n1 152
R119 CIN.n5 CIN.n2 84.872
R120 CIN CIN.n5 9.4725
R121 A.n3 A.t5 337.937
R122 A.n7 A.t3 300.983
R123 A.n2 A.n0 300.983
R124 A.n5 A.t0 288.13
R125 A.n5 A.t1 217.436
R126 A.n2 A.n1 206.19
R127 A.n7 A.t2 205.702
R128 A.n4 A.n2 188.26
R129 A.n6 A.n5 169.833
R130 A.n3 A.t4 167.63
R131 A.n4 A.n3 166.633
R132 A A.n7 165.03
R133 A A.n6 14.317
R134 A.n6 A.n4 1.55989
R135 a_658_369.t0 a_658_369.n0 1284.71
R136 a_658_369.n0 a_658_369.t1 41.5552
R137 a_658_369.n0 a_658_369.t2 41.5552
R138 a_658_47.t0 a_658_47.n0 497.418
R139 a_658_47.n0 a_658_47.t1 38.5719
R140 a_658_47.n0 a_658_47.t2 38.5719
R141 VGND.n12 VGND.t5 286.714
R142 VGND.n45 VGND.t12 282.565
R143 VGND.n16 VGND.t7 255.227
R144 VGND.n28 VGND.t1 239.281
R145 VGND.n11 VGND.n10 208.719
R146 VGND.n43 VGND.n1 208.719
R147 VGND.n38 VGND.n37 199.739
R148 VGND.n24 VGND.n23 198.964
R149 VGND.n31 VGND.n30 198.964
R150 VGND.n37 VGND.t10 48.2862
R151 VGND.n23 VGND.t3 38.5719
R152 VGND.n23 VGND.t13 38.5719
R153 VGND.n30 VGND.t0 38.5719
R154 VGND.n30 VGND.t2 38.5719
R155 VGND.n37 VGND.t4 38.5719
R156 VGND.n15 VGND.n14 34.6358
R157 VGND.n17 VGND.n8 34.6358
R158 VGND.n21 VGND.n8 34.6358
R159 VGND.n22 VGND.n21 34.6358
R160 VGND.n35 VGND.n4 34.6358
R161 VGND.n36 VGND.n35 34.6358
R162 VGND.n42 VGND.n2 34.6358
R163 VGND.n45 VGND.n44 32.377
R164 VGND.n24 VGND.n22 31.624
R165 VGND.n44 VGND.n43 30.8711
R166 VGND.n14 VGND.n11 29.7417
R167 VGND.n31 VGND.n29 27.1064
R168 VGND.n38 VGND.n36 25.977
R169 VGND.n28 VGND.n6 25.6005
R170 VGND.n10 VGND.t8 24.9236
R171 VGND.n10 VGND.t6 24.9236
R172 VGND.n1 VGND.t11 24.9236
R173 VGND.n1 VGND.t9 24.9236
R174 VGND.n29 VGND.n28 18.824
R175 VGND.n38 VGND.n2 18.4476
R176 VGND.n31 VGND.n4 17.3181
R177 VGND.n24 VGND.n6 12.8005
R178 VGND.n12 VGND.n11 11.8645
R179 VGND.n46 VGND.n45 11.5593
R180 VGND.n14 VGND.n13 9.3005
R181 VGND.n15 VGND.n9 9.3005
R182 VGND.n18 VGND.n17 9.3005
R183 VGND.n19 VGND.n8 9.3005
R184 VGND.n21 VGND.n20 9.3005
R185 VGND.n22 VGND.n7 9.3005
R186 VGND.n25 VGND.n24 9.3005
R187 VGND.n26 VGND.n6 9.3005
R188 VGND.n28 VGND.n27 9.3005
R189 VGND.n29 VGND.n5 9.3005
R190 VGND.n32 VGND.n31 9.3005
R191 VGND.n33 VGND.n4 9.3005
R192 VGND.n35 VGND.n34 9.3005
R193 VGND.n36 VGND.n3 9.3005
R194 VGND.n39 VGND.n38 9.3005
R195 VGND.n40 VGND.n2 9.3005
R196 VGND.n42 VGND.n41 9.3005
R197 VGND.n44 VGND.n0 9.3005
R198 VGND.n17 VGND.n16 8.65932
R199 VGND.n43 VGND.n42 3.76521
R200 VGND.n16 VGND.n15 1.12991
R201 VGND.n13 VGND.n12 0.779653
R202 VGND.n13 VGND.n9 0.120292
R203 VGND.n18 VGND.n9 0.120292
R204 VGND.n19 VGND.n18 0.120292
R205 VGND.n20 VGND.n19 0.120292
R206 VGND.n20 VGND.n7 0.120292
R207 VGND.n25 VGND.n7 0.120292
R208 VGND.n26 VGND.n25 0.120292
R209 VGND.n27 VGND.n26 0.120292
R210 VGND.n27 VGND.n5 0.120292
R211 VGND.n32 VGND.n5 0.120292
R212 VGND.n33 VGND.n32 0.120292
R213 VGND.n34 VGND.n33 0.120292
R214 VGND.n34 VGND.n3 0.120292
R215 VGND.n39 VGND.n3 0.120292
R216 VGND.n40 VGND.n39 0.120292
R217 VGND.n41 VGND.n40 0.120292
R218 VGND.n41 VGND.n0 0.120292
R219 VGND.n46 VGND.n0 0.120292
R220 VGND VGND.n46 0.0213333
R221 VNB.t3 VNB.t6 6721.04
R222 VNB.t2 VNB.t0 2677.02
R223 VNB.t1 VNB.t15 1452.43
R224 VNB.t6 VNB.t9 1423.95
R225 VNB.t11 VNB.t4 1423.95
R226 VNB.t4 VNB.t1 1352.75
R227 VNB.t7 VNB.t8 1196.12
R228 VNB.t9 VNB.t7 1196.12
R229 VNB.t14 VNB.t3 1196.12
R230 VNB.t0 VNB.t14 1196.12
R231 VNB.t5 VNB.t2 1196.12
R232 VNB.t15 VNB.t5 1196.12
R233 VNB.t12 VNB.t11 1196.12
R234 VNB.t10 VNB.t12 1196.12
R235 VNB.t13 VNB.t10 1196.12
R236 VNB VNB.t13 911.327
R237 a_456_371.t0 a_456_371.t1 92.2465
R238 a_79_21.n15 a_79_21.n14 394.021
R239 a_79_21.n2 a_79_21.n0 337.937
R240 a_79_21.n6 a_79_21.t4 212.081
R241 a_79_21.n11 a_79_21.t5 212.081
R242 a_79_21.n9 a_79_21.t6 212.081
R243 a_79_21.n7 a_79_21.t10 212.081
R244 a_79_21.n4 a_79_21.n2 189.532
R245 a_79_21.n4 a_79_21.n3 185.786
R246 a_79_21.n8 a_79_21.n5 177.601
R247 a_79_21.n2 a_79_21.n1 167.63
R248 a_79_21.n10 a_79_21.n5 152
R249 a_79_21.n13 a_79_21.n12 152
R250 a_79_21.n6 a_79_21.t8 139.78
R251 a_79_21.n11 a_79_21.t9 139.78
R252 a_79_21.n9 a_79_21.t7 139.78
R253 a_79_21.n7 a_79_21.t11 139.78
R254 a_79_21.n14 a_79_21.n4 73.333
R255 a_79_21.n15 a_79_21.t1 67.2307
R256 a_79_21.n3 a_79_21.t0 64.2862
R257 a_79_21.n8 a_79_21.n7 43.8187
R258 a_79_21.n12 a_79_21.n6 40.8975
R259 a_79_21.n3 a_79_21.t2 38.5719
R260 a_79_21.n16 a_79_21.t3 38.2409
R261 a_79_21.n10 a_79_21.n9 32.1338
R262 a_79_21.n11 a_79_21.n10 29.2126
R263 a_79_21.n14 a_79_21.n13 28.2358
R264 a_79_21.n13 a_79_21.n5 25.6005
R265 a_79_21.n12 a_79_21.n11 20.449
R266 a_79_21.n9 a_79_21.n8 17.5278
R267 a_79_21.n16 a_79_21.n15 15.6354
R268 a_79_21.n17 a_79_21.n16 3.33948
R269 SUM.n2 SUM.n0 373.817
R270 SUM.n2 SUM.n1 206.832
R271 SUM.n5 SUM.n3 139.154
R272 SUM.n5 SUM.n4 98.788
R273 SUM.n3 SUM.t0 39.6928
R274 SUM SUM.n2 30.9048
R275 SUM SUM.n5 26.7018
R276 SUM.n0 SUM.t7 26.5955
R277 SUM.n0 SUM.t6 26.5955
R278 SUM.n1 SUM.t5 26.5955
R279 SUM.n1 SUM.t4 26.5955
R280 SUM.n3 SUM.t3 24.9236
R281 SUM.n4 SUM.t2 24.9236
R282 SUM.n4 SUM.t1 24.9236
R283 a_461_47.t0 a_461_47.t1 92.8576
R284 COUT.n6 COUT.n0 585
R285 COUT.n5 COUT.n4 369.954
R286 COUT COUT.n0 302.55
R287 COUT.n3 COUT.n1 251.922
R288 COUT.n3 COUT.n2 98.788
R289 COUT.n5 COUT.n3 36.9161
R290 COUT.n0 COUT.t5 26.5955
R291 COUT.n0 COUT.t4 26.5955
R292 COUT.n4 COUT.t7 26.5955
R293 COUT.n4 COUT.t6 26.5955
R294 COUT.n1 COUT.t2 24.9236
R295 COUT.n1 COUT.t1 24.9236
R296 COUT.n2 COUT.t3 24.9236
R297 COUT.n2 COUT.t0 24.9236
R298 COUT COUT.n6 6.4005
R299 COUT.n6 COUT.n5 4.65505
R300 a_1356_369.n0 a_1356_369.t0 3.03127
C0 a_1451_47# a_1271_47# 0.00786f
C1 VPWR a_1451_371# 0.002106f
C2 VPB A 0.220437f
C3 a_1014_369# a_1451_371# 3.49e-19
C4 VPB B 0.284057f
C5 a_1014_47# VGND 0.146711f
C6 VGND SUM 0.253862f
C7 VPB a_1271_47# 0.140539f
C8 A B 0.801163f
C9 a_1379_47# VGND 8.64e-19
C10 VPB CIN 0.193074f
C11 A a_1271_47# 0.172418f
C12 SUM a_1451_371# 7.56e-20
C13 a_1014_47# a_1379_47# 2.04e-19
C14 A CIN 0.437174f
C15 a_1451_47# VGND 0.0024f
C16 VPB VPWR 0.206836f
C17 B a_1271_47# 0.113521f
C18 a_1014_47# a_1451_47# 3.57e-20
C19 VPB COUT 0.012538f
C20 B CIN 0.544917f
C21 A VPWR 0.064277f
C22 a_1451_47# SUM 3.81e-19
C23 CIN a_1271_47# 0.059656f
C24 VPB a_1014_369# 0.004107f
C25 VPB VGND 0.007971f
C26 A COUT 0.005042f
C27 B VPWR 0.294776f
C28 A a_1014_369# 0.010031f
C29 VPWR a_1271_47# 0.279642f
C30 a_1014_47# VPB 7.38e-19
C31 CIN VPWR 0.053466f
C32 A VGND 0.089911f
C33 B COUT 0.001816f
C34 VPB SUM 0.015402f
C35 B a_1014_369# 0.016831f
C36 a_1271_47# a_1014_369# 0.025789f
C37 a_1014_47# A 0.043259f
C38 A SUM 0.004329f
C39 B VGND 0.059993f
C40 CIN a_1014_369# 0.078088f
C41 VGND a_1271_47# 0.249725f
C42 a_1014_47# B 0.005347f
C43 a_1379_47# A 8.51e-19
C44 CIN VGND 0.061421f
C45 VPWR COUT 0.309908f
C46 B SUM 0.003336f
C47 a_1014_47# a_1271_47# 0.023091f
C48 B a_1451_371# 0.003361f
C49 SUM a_1271_47# 0.42318f
C50 VPWR a_1014_369# 0.174928f
C51 a_1271_47# a_1451_371# 0.013654f
C52 a_1451_47# A 3.14e-19
C53 a_1014_47# CIN 0.047968f
C54 VPWR VGND 0.100004f
C55 a_1379_47# a_1271_47# 0.005553f
C56 CIN a_1451_371# 7.61e-19
C57 a_1451_47# B 6.31e-19
C58 COUT VGND 0.238414f
C59 VPWR SUM 0.29959f
C60 SUM VNB 0.063014f
C61 VGND VNB 1.11447f
C62 COUT VNB 0.058002f
C63 VPWR VNB 0.951779f
C64 CIN VNB 0.331216f
C65 B VNB 0.47835f
C66 A VNB 0.487539f
C67 VPB VNB 2.0223f
C68 a_1014_47# VNB 0.015892f
C69 a_1014_369# VNB 0.004114f
C70 a_1271_47# VNB 0.416727f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fah_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fah_1 VPWR VGND VNB VPB B CI COUT SUM A
X0 a_508_297.t2 B.t0 VGND.t4 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.17 pd=1.86 as=0.171275 ps=1.18 w=0.65 l=0.15
X1 a_1332_297.t1 a_719_47.t4 a_1262_49.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.088 pd=0.915 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 a_27_47.t3 a_508_297.t4 a_719_47.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.2176 pd=1.96 as=0.088 ps=0.915 w=0.64 l=0.15
X3 a_67_199.t0 A.t0 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X4 a_508_297.t3 B.t1 VPWR.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X5 VPWR.t3 A.t1 a_310_49.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.275 ps=2.55 w=1 l=0.15
X6 a_310_49.t2 B.t2 a_1008_47.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.15225 ps=1.3 w=0.84 l=0.15
X7 a_508_297.t1 a_1008_47.t4 a_1332_297.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.088 ps=0.915 w=0.64 l=0.15
X8 a_1332_297.t2 a_719_47.t5 a_508_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2562 ps=2.29 w=0.84 l=0.15
X9 a_719_47.t0 B.t3 a_310_49.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.088 pd=0.915 as=0.16285 ps=1.8 w=0.64 l=0.15
X10 a_1640_380.t0 a_719_47.t6 a_1617_49.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1792 pd=1.84 as=0.0928 ps=0.93 w=0.64 l=0.15
X11 a_1008_47.t2 a_508_297.t5 a_310_49.t5 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.189675 pd=1.24 as=0.1664 ps=1.8 w=0.64 l=0.15
X12 VGND.t0 a_1332_297.t4 COUT.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1755 ps=1.84 w=0.65 l=0.15
X13 a_719_47.t1 B.t4 a_27_47.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.115 as=0.3594 ps=2.8 w=0.84 l=0.15
X14 a_1262_49.t2 a_719_47.t7 a_1617_49.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.340275 pd=1.73 as=0.1134 ps=1.11 w=0.84 l=0.15
X15 SUM.t0 a_1617_49.t4 VPWR.t6 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1640_380.t2 a_1262_49.t5 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_1617_49.t2 a_1008_47.t5 a_1640_380.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.21515 ps=2.2 w=0.84 l=0.15
X18 VPWR.t1 a_1332_297.t5 COUT.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VPWR.t7 a_67_199.t2 a_27_47.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.28 ps=2.56 w=1 l=0.15
X20 a_310_49.t4 a_508_297.t6 a_719_47.t2 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.1155 ps=1.115 w=0.84 l=0.15
X21 a_67_199.t1 A.t2 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.10525 ps=0.975 w=0.64 l=0.15
X22 VGND.t2 A.t3 a_310_49.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.171275 pd=1.18 as=0.1664 ps=1.8 w=0.64 l=0.15
X23 a_27_47.t1 B.t5 a_1008_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.189675 ps=1.24 w=0.64 l=0.15
X24 a_1617_49.t3 a_1008_47.t6 a_1262_49.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X25 SUM.t1 a_1617_49.t5 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t0 CI.t0 a_1262_49.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.340275 ps=1.73 w=1 l=0.15
X27 a_1008_47.t3 a_508_297.t7 a_27_47.t2 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.3 as=0.323 ps=2.73 w=0.84 l=0.15
X28 VGND.t5 a_67_199.t3 a_27_47.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X29 a_1262_49.t0 a_1008_47.t7 a_1332_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.711425 pd=3.4 as=0.1134 ps=1.11 w=0.84 l=0.15
R0 B.n3 B.t2 242.607
R1 B.n2 B.t1 212.081
R2 B.n4 B.n2 188.038
R3 B.n0 B.t4 186.374
R4 B B.n3 166.03
R5 B.n3 B.t5 154.24
R6 B.n0 B.t3 141.387
R7 B.n1 B.t0 139.78
R8 B.n1 B.n0 139.488
R9 B.n2 B.n1 14.6066
R10 B.n4 B 9.3005
R11 B B.n4 5.4405
R12 VGND.n6 VGND.n5 207.213
R13 VGND.n13 VGND.n1 207.213
R14 VGND.n4 VGND.n3 118.794
R15 VGND.n5 VGND.t4 67.042
R16 VGND.n14 VGND.n13 43.1829
R17 VGND.n6 VGND.n4 40.3541
R18 VGND.n1 VGND.t1 35.6255
R19 VGND.n7 VGND.n2 34.6358
R20 VGND.n11 VGND.n2 34.6358
R21 VGND.n12 VGND.n11 34.6358
R22 VGND.n5 VGND.t2 25.313
R23 VGND.n3 VGND.t3 24.9236
R24 VGND.n3 VGND.t0 24.9236
R25 VGND.n1 VGND.t5 22.1675
R26 VGND.n12 VGND.n0 9.3005
R27 VGND.n11 VGND.n10 9.3005
R28 VGND.n9 VGND.n2 9.3005
R29 VGND.n8 VGND.n7 9.3005
R30 VGND.n7 VGND.n6 1.88285
R31 VGND.n13 VGND.n12 0.753441
R32 VGND.n8 VGND.n4 0.147187
R33 VGND.n9 VGND.n8 0.120292
R34 VGND.n10 VGND.n9 0.120292
R35 VGND.n10 VGND.n0 0.120292
R36 VGND.n14 VGND.n0 0.120292
R37 VGND VGND.n14 0.0226354
R38 a_508_297.t3 a_508_297.n5 853.981
R39 a_508_297.n0 a_508_297.t0 769.082
R40 a_508_297.n0 a_508_297.t1 398.344
R41 a_508_297.n5 a_508_297.t2 269.195
R42 a_508_297.n1 a_508_297.t7 191.486
R43 a_508_297.n2 a_508_297.t6 186.374
R44 a_508_297.n4 a_508_297.n3 171.486
R45 a_508_297.n2 a_508_297.t4 141.387
R46 a_508_297.n1 a_508_297.t5 141.387
R47 a_508_297.n3 a_508_297.n1 106.624
R48 a_508_297.n3 a_508_297.n2 42.3581
R49 a_508_297.n4 a_508_297.n0 21.7106
R50 a_508_297.n5 a_508_297.n4 17.546
R51 VNB.t1 VNB.t2 8500.97
R52 VNB.t12 VNB.t11 2904.85
R53 VNB.t10 VNB.t9 2719.74
R54 VNB.t3 VNB.t7 2677.02
R55 VNB.t8 VNB.t0 2677.02
R56 VNB.t4 VNB.t5 2677.02
R57 VNB.t11 VNB.t8 2107.44
R58 VNB.t5 VNB.t10 1936.57
R59 VNB.t13 VNB.t4 1352.75
R60 VNB.t7 VNB.t1 1253.07
R61 VNB.t0 VNB.t3 1210.36
R62 VNB.t9 VNB.t12 1210.36
R63 VNB.t2 VNB.t6 1196.12
R64 VNB VNB.t13 925.567
R65 a_719_47.n5 a_719_47.n4 641.221
R66 a_719_47.n1 a_719_47.t6 289.2
R67 a_719_47.n1 a_719_47.t7 284.38
R68 a_719_47.n3 a_719_47.n1 234.447
R69 a_719_47.n3 a_719_47.n2 219.333
R70 a_719_47.n4 a_719_47.n0 209.471
R71 a_719_47.n2 a_719_47.t5 186.374
R72 a_719_47.n2 a_719_47.t4 146.938
R73 a_719_47.n5 a_719_47.t2 32.8338
R74 a_719_47.t1 a_719_47.n5 31.6612
R75 a_719_47.n0 a_719_47.t0 26.2505
R76 a_719_47.n0 a_719_47.t3 25.313
R77 a_719_47.n4 a_719_47.n3 11.6813
R78 a_1262_49.n5 a_1262_49.t0 757.375
R79 a_1262_49.n3 a_1262_49.n0 587.121
R80 a_1262_49.n7 a_1262_49.n6 585
R81 a_1262_49.n4 a_1262_49.t3 316.281
R82 a_1262_49.n2 a_1262_49.t5 238.155
R83 a_1262_49.n3 a_1262_49.n2 215.494
R84 a_1262_49.n4 a_1262_49.t4 210.312
R85 a_1262_49.n2 a_1262_49.n1 164.25
R86 a_1262_49.n6 a_1262_49.n5 146.905
R87 a_1262_49.n8 a_1262_49.t1 137.74
R88 a_1262_49.n7 a_1262_49.t2 84.4291
R89 a_1262_49.n5 a_1262_49.n4 69.0419
R90 a_1262_49.n6 a_1262_49.n3 43.6551
R91 a_1262_49.t1 a_1262_49.n0 25.4508
R92 a_1262_49.n9 a_1262_49.n8 24.6255
R93 a_1262_49.n10 a_1262_49.n9 21.6225
R94 a_1262_49.n9 a_1262_49.n0 13.1972
R95 a_1262_49.n8 a_1262_49.n7 4.69098
R96 a_1332_297.n3 a_1332_297.n2 615.006
R97 a_1332_297.n1 a_1332_297.t5 233.576
R98 a_1332_297.n2 a_1332_297.n0 203.964
R99 a_1332_297.n2 a_1332_297.n1 176.151
R100 a_1332_297.n1 a_1332_297.t4 161.275
R101 a_1332_297.t0 a_1332_297.n3 31.6612
R102 a_1332_297.n3 a_1332_297.t2 31.6612
R103 a_1332_297.n0 a_1332_297.t3 26.2505
R104 a_1332_297.n0 a_1332_297.t1 25.313
R105 a_27_47.n12 a_27_47.t0 852.851
R106 a_27_47.n11 a_27_47.t2 394.389
R107 a_27_47.n3 a_27_47.t1 291.488
R108 a_27_47.n10 a_27_47.t3 266.661
R109 a_27_47.n13 a_27_47.n12 231.488
R110 a_27_47.t4 a_27_47.n13 220.177
R111 a_27_47.n13 a_27_47.t5 202.655
R112 a_27_47.n12 a_27_47.n11 141.565
R113 a_27_47.n2 a_27_47.n1 115.201
R114 a_27_47.n8 a_27_47.n1 98.9872
R115 a_27_47.n4 a_27_47.n3 80.0837
R116 a_27_47.n11 a_27_47.n10 77.2186
R117 a_27_47.n7 a_27_47.n0 54.4005
R118 a_27_47.n8 a_27_47.n7 44.8005
R119 a_27_47.n6 a_27_47.n2 38.4005
R120 a_27_47.n6 a_27_47.n5 38.4005
R121 a_27_47.n3 a_27_47.n1 32.7848
R122 a_27_47.n7 a_27_47.n6 32.0005
R123 a_27_47.n4 a_27_47.n2 25.6005
R124 a_27_47.n9 a_27_47.n8 19.5373
R125 a_27_47.n10 a_27_47.n9 18.2494
R126 a_27_47.n9 a_27_47.n0 9.6005
R127 a_27_47.n5 a_27_47.n0 5.1205
R128 a_27_47.n5 a_27_47.n4 1.82907
R129 CI.n1 CI.t0 233.869
R130 CI CI.n1 175.952
R131 CI.n1 CI.n0 159.963
R132 A.n0 A.t1 214.272
R133 A.n1 A.t0 212.81
R134 A A.n2 159.041
R135 A.n1 A.t2 141.387
R136 A.n0 A.t3 138.173
R137 A.n2 A.n0 103.704
R138 A.n2 A.n1 33.5944
R139 VPWR.n3 VPWR.n2 600.515
R140 VPWR.n14 VPWR.n13 598.755
R141 VPWR.n44 VPWR.n1 598.152
R142 VPWR.n15 VPWR.n12 324.606
R143 VPWR.n2 VPWR.t3 50.2355
R144 VPWR.n43 VPWR.n42 34.6358
R145 VPWR.n18 VPWR.n11 34.6358
R146 VPWR.n19 VPWR.n18 34.6358
R147 VPWR.n20 VPWR.n19 34.6358
R148 VPWR.n20 VPWR.n9 34.6358
R149 VPWR.n24 VPWR.n9 34.6358
R150 VPWR.n25 VPWR.n24 34.6358
R151 VPWR.n26 VPWR.n25 34.6358
R152 VPWR.n26 VPWR.n7 34.6358
R153 VPWR.n30 VPWR.n7 34.6358
R154 VPWR.n31 VPWR.n30 34.6358
R155 VPWR.n32 VPWR.n31 34.6358
R156 VPWR.n32 VPWR.n5 34.6358
R157 VPWR.n36 VPWR.n5 34.6358
R158 VPWR.n37 VPWR.n36 34.6358
R159 VPWR.n38 VPWR.n37 34.6358
R160 VPWR.n42 VPWR.n3 34.2593
R161 VPWR.n1 VPWR.t7 32.5055
R162 VPWR.n2 VPWR.t5 31.5205
R163 VPWR.n14 VPWR.n11 30.8711
R164 VPWR.n1 VPWR.t2 26.5955
R165 VPWR.n13 VPWR.t4 26.5955
R166 VPWR.n13 VPWR.t0 26.5955
R167 VPWR.n12 VPWR.t6 26.5955
R168 VPWR.n12 VPWR.t1 26.5955
R169 VPWR.n44 VPWR.n43 16.5652
R170 VPWR.n38 VPWR.n3 10.1652
R171 VPWR.n16 VPWR.n11 9.3005
R172 VPWR.n18 VPWR.n17 9.3005
R173 VPWR.n19 VPWR.n10 9.3005
R174 VPWR.n21 VPWR.n20 9.3005
R175 VPWR.n22 VPWR.n9 9.3005
R176 VPWR.n24 VPWR.n23 9.3005
R177 VPWR.n25 VPWR.n8 9.3005
R178 VPWR.n27 VPWR.n26 9.3005
R179 VPWR.n28 VPWR.n7 9.3005
R180 VPWR.n30 VPWR.n29 9.3005
R181 VPWR.n31 VPWR.n6 9.3005
R182 VPWR.n33 VPWR.n32 9.3005
R183 VPWR.n34 VPWR.n5 9.3005
R184 VPWR.n36 VPWR.n35 9.3005
R185 VPWR.n37 VPWR.n4 9.3005
R186 VPWR.n39 VPWR.n38 9.3005
R187 VPWR.n40 VPWR.n3 9.3005
R188 VPWR.n42 VPWR.n41 9.3005
R189 VPWR.n43 VPWR.n0 9.3005
R190 VPWR.n45 VPWR.n44 7.30743
R191 VPWR.n15 VPWR.n14 6.37606
R192 VPWR.n16 VPWR.n15 0.184025
R193 VPWR.n45 VPWR.n0 0.146144
R194 VPWR.n17 VPWR.n16 0.120292
R195 VPWR.n17 VPWR.n10 0.120292
R196 VPWR.n21 VPWR.n10 0.120292
R197 VPWR.n22 VPWR.n21 0.120292
R198 VPWR.n23 VPWR.n22 0.120292
R199 VPWR.n23 VPWR.n8 0.120292
R200 VPWR.n27 VPWR.n8 0.120292
R201 VPWR.n28 VPWR.n27 0.120292
R202 VPWR.n29 VPWR.n28 0.120292
R203 VPWR.n29 VPWR.n6 0.120292
R204 VPWR.n33 VPWR.n6 0.120292
R205 VPWR.n34 VPWR.n33 0.120292
R206 VPWR.n35 VPWR.n34 0.120292
R207 VPWR.n35 VPWR.n4 0.120292
R208 VPWR.n39 VPWR.n4 0.120292
R209 VPWR.n40 VPWR.n39 0.120292
R210 VPWR.n41 VPWR.n40 0.120292
R211 VPWR.n41 VPWR.n0 0.120292
R212 VPWR VPWR.n45 0.117248
R213 a_67_199.t0 a_67_199.n1 893.554
R214 a_67_199.n0 a_67_199.t2 236.934
R215 a_67_199.n1 a_67_199.t1 172.631
R216 a_67_199.n0 a_67_199.t3 164.633
R217 a_67_199.n1 a_67_199.n0 152
R218 VPB.t0 VPB.t4 905.607
R219 VPB.t9 VPB.t6 722.119
R220 VPB.t11 VPB.t2 651.091
R221 VPB.t14 VPB.t13 624.456
R222 VPB.t12 VPB.t10 624.456
R223 VPB.t8 VPB.t7 568.225
R224 VPB.t1 VPB.t5 497.197
R225 VPB.t7 VPB.t12 334.425
R226 VPB.t13 VPB.t11 287.072
R227 VPB.t3 VPB.t8 266.356
R228 VPB.t10 VPB.t14 251.559
R229 VPB.t6 VPB.t15 248.599
R230 VPB.t5 VPB.t9 248.599
R231 VPB.t4 VPB.t1 248.599
R232 VPB.t2 VPB.t0 248.599
R233 VPB VPB.t3 204.207
R234 a_310_49.t0 a_310_49.n3 911.827
R235 a_310_49.n0 a_310_49.t2 731.486
R236 a_310_49.n0 a_310_49.t4 619.861
R237 a_310_49.n1 a_310_49.t5 298.389
R238 a_310_49.n1 a_310_49.t3 212.649
R239 a_310_49.n2 a_310_49.n0 180.894
R240 a_310_49.n3 a_310_49.t1 137.428
R241 a_310_49.n3 a_310_49.n2 116.617
R242 a_310_49.n2 a_310_49.n1 11.8862
R243 a_1008_47.n5 a_1008_47.n4 585
R244 a_1008_47.n4 a_1008_47.n2 416.856
R245 a_1008_47.n0 a_1008_47.t5 319.034
R246 a_1008_47.n4 a_1008_47.n3 288.983
R247 a_1008_47.n1 a_1008_47.t7 195.868
R248 a_1008_47.n1 a_1008_47.t4 138.173
R249 a_1008_47.n0 a_1008_47.t6 138.173
R250 a_1008_47.n2 a_1008_47.n0 69.3793
R251 a_1008_47.n2 a_1008_47.n1 67.9187
R252 a_1008_47.n3 a_1008_47.t2 66.1291
R253 a_1008_47.t0 a_1008_47.n5 50.1584
R254 a_1008_47.n5 a_1008_47.t3 32.2493
R255 a_1008_47.n3 a_1008_47.t1 26.0641
R256 a_1617_49.n3 a_1617_49.n2 592.529
R257 a_1617_49.n1 a_1617_49.t4 241.536
R258 a_1617_49.n2 a_1617_49.n0 239.085
R259 a_1617_49.n2 a_1617_49.n1 188.651
R260 a_1617_49.n1 a_1617_49.t5 169.237
R261 a_1617_49.t1 a_1617_49.n3 31.6612
R262 a_1617_49.n3 a_1617_49.t2 31.6612
R263 a_1617_49.n0 a_1617_49.t3 29.063
R264 a_1617_49.n0 a_1617_49.t0 25.313
R265 a_1640_380.n0 a_1640_380.t1 687.788
R266 a_1640_380.t2 a_1640_380.n0 639.976
R267 a_1640_380.n0 a_1640_380.t0 377.372
R268 COUT.n1 COUT.n0 585
R269 COUT COUT.n0 299.255
R270 COUT.n1 COUT.t1 271.817
R271 COUT.n0 COUT.t0 26.5955
R272 COUT COUT.n1 3.69281
R273 SUM SUM.t0 368.241
R274 SUM SUM.t1 154.514
C0 VGND COUT 0.102007f
C1 VPB A 0.091048f
C2 VGND SUM 0.099144f
C3 VPB B 0.17852f
C4 COUT SUM 0.00968f
C5 VPB VPWR 0.246285f
C6 A B 0.055195f
C7 VPB CI 0.036811f
C8 A VPWR 0.033037f
C9 B VPWR 0.050297f
C10 VPB VGND 0.007665f
C11 B CI 2.13e-19
C12 VPB COUT 0.017767f
C13 A VGND 0.034436f
C14 VPWR CI 0.013446f
C15 B VGND 0.079275f
C16 VPB SUM 0.01427f
C17 B COUT 4.95e-21
C18 VPWR VGND 0.053433f
C19 VPWR COUT 0.126934f
C20 CI VGND 0.031502f
C21 B SUM 1.5e-21
C22 VPWR SUM 0.109351f
C23 SUM VNB 0.094881f
C24 COUT VNB 0.01721f
C25 VGND VNB 1.32517f
C26 CI VNB 0.111457f
C27 VPWR VNB 1.09047f
C28 B VNB 0.392095f
C29 A VNB 0.234314f
C30 VPB VNB 2.46528f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fahcin_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fahcin_1 VPWR VGND VNB VPB SUM CIN COUT B A
X0 a_721_47.t2 a_489_21.t2 a_27_47.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.3 as=0.3398 ps=2.77 w=0.84 l=0.15
X1 VGND.t1 a_1636_315.t3 a_1565_49.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.1728 ps=1.82 w=0.64 l=0.15
X2 SUM.t0 a_1647_49.t2 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t4 CIN.t0 a_1251_49.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VPWR.t0 a_67_199.t6 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X5 a_67_199.t1 B.t0 a_721_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.2814 pd=2.35 as=0.15225 ps=1.3 w=0.84 l=0.15
X6 VPWR.t5 CIN.t1 a_1251_49.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_67_199.t4 a_489_21.t3 a_434_49.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.1155 ps=1.115 w=0.84 l=0.15
X8 COUT.t1 a_434_49.t4 a_1251_49.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.088 pd=0.915 as=0.192 ps=1.88 w=0.64 l=0.15
X9 a_434_49.t3 B.t1 a_67_199.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.088 pd=0.915 as=0.321225 ps=1.645 w=0.64 l=0.15
X10 a_434_49.t2 B.t2 a_27_47.t4 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.115 as=0.2629 ps=2.64 w=0.84 l=0.15
X11 VPWR.t3 a_1636_315.t4 a_1565_49.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4492 ps=1.98 w=1 l=0.15
X12 VGND.t5 B.t3 a_489_21.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.11645 pd=1.01 as=0.165325 ps=1.82 w=0.65 l=0.15
X13 a_67_199.t0 A.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.31175 pd=2.88 as=0.175 ps=1.35 w=1 l=0.15
X14 a_1142_49.t3 a_721_47.t4 COUT.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1792 pd=1.84 as=0.088 ps=0.915 w=0.64 l=0.15
X15 VGND.t3 a_67_199.t7 a_27_47.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.1696 ps=1.81 w=0.64 l=0.15
X16 a_27_47.t1 a_489_21.t4 a_434_49.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.199825 pd=1.91 as=0.088 ps=0.915 w=0.64 l=0.15
X17 a_67_199.t3 A.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.321225 pd=1.645 as=0.10525 ps=0.975 w=0.65 l=0.15
X18 VPWR.t7 B.t4 a_489_21.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47.t5 B.t5 a_721_47.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.162825 pd=1.8 as=0.165675 ps=1.165 w=0.64 l=0.15
X20 a_1251_49.t3 a_721_47.t5 COUT.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.7033 pd=3.36 as=0.1134 ps=1.11 w=0.84 l=0.15
X21 a_1142_49.t1 a_489_21.t5 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.11645 ps=1.01 w=0.64 l=0.15
X22 a_1142_49.t2 a_489_21.t6 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.3826 pd=1.79 as=0.18 ps=1.36 w=1 l=0.15
X23 a_1565_49.t0 a_434_49.t5 a_1647_49.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.4492 pd=1.98 as=0.1134 ps=1.11 w=0.84 l=0.15
X24 a_721_47.t1 a_489_21.t7 a_67_199.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.165675 pd=1.165 as=0.168125 ps=1.83 w=0.64 l=0.15
X25 a_1647_49.t1 a_721_47.t6 a_1636_315.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2184 ps=2.2 w=0.84 l=0.15
X26 a_1636_315.t1 CIN.t2 VPWR.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X27 COUT.t0 a_434_49.t6 a_1142_49.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.3826 ps=1.79 w=0.84 l=0.15
X28 a_1636_315.t2 CIN.t3 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10525 ps=0.975 w=0.65 l=0.15
R0 a_489_21.t1 a_489_21.n5 849.337
R1 a_489_21.n1 a_489_21.t0 253.917
R2 a_489_21.n0 a_489_21.t6 238.59
R3 a_489_21.n5 a_489_21.n4 208.85
R4 a_489_21.n2 a_489_21.t2 194.407
R5 a_489_21.n3 a_489_21.t3 186.374
R6 a_489_21.n1 a_489_21.n0 166.546
R7 a_489_21.n0 a_489_21.t5 164.684
R8 a_489_21.n2 a_489_21.t7 141.387
R9 a_489_21.n3 a_489_21.t4 138.173
R10 a_489_21.n4 a_489_21.n2 105.894
R11 a_489_21.n4 a_489_21.n3 41.6278
R12 a_489_21.n5 a_489_21.n1 12.3378
R13 a_27_47.n2 a_27_47.t4 745.086
R14 a_27_47.n1 a_27_47.t2 388.983
R15 a_27_47.n0 a_27_47.t5 312.3
R16 a_27_47.n0 a_27_47.t1 258.632
R17 a_27_47.t0 a_27_47.n3 221.34
R18 a_27_47.n3 a_27_47.t3 216.083
R19 a_27_47.n2 a_27_47.n1 132.004
R20 a_27_47.n3 a_27_47.n2 119.585
R21 a_27_47.n1 a_27_47.n0 76.063
R22 a_721_47.n6 a_721_47.n5 585
R23 a_721_47.n5 a_721_47.n3 580.947
R24 a_721_47.n1 a_721_47.t6 282.086
R25 a_721_47.n5 a_721_47.n4 280.137
R26 a_721_47.n2 a_721_47.t5 195.137
R27 a_721_47.n1 a_721_47.n0 144.746
R28 a_721_47.n2 a_721_47.t4 138.173
R29 a_721_47.n3 a_721_47.n2 130.725
R30 a_721_47.n4 a_721_47.t1 62.5944
R31 a_721_47.t0 a_721_47.n6 50.1584
R32 a_721_47.n6 a_721_47.t2 32.2493
R33 a_721_47.n3 a_721_47.n1 24.1005
R34 a_721_47.n4 a_721_47.t3 20.1091
R35 VPB.t11 VPB.t10 899.688
R36 VPB.t2 VPB.t6 668.847
R37 VPB.t3 VPB.t14 662.928
R38 VPB.t8 VPB.t9 630.375
R39 VPB.t4 VPB.t15 624.456
R40 VPB.t13 VPB.t12 571.184
R41 VPB.t7 VPB.t5 556.386
R42 VPB.t15 VPB.t7 301.87
R43 VPB.t1 VPB.t3 295.95
R44 VPB.t9 VPB.t4 287.072
R45 VPB.t14 VPB.t8 251.559
R46 VPB.t12 VPB.t0 248.599
R47 VPB.t6 VPB.t13 248.599
R48 VPB.t10 VPB.t2 248.599
R49 VPB.t5 VPB.t11 248.599
R50 VPB VPB.t1 195.327
R51 a_1636_315.n2 a_1636_315.t0 798.064
R52 a_1636_315.n0 a_1636_315.t4 241.536
R53 a_1636_315.t1 a_1636_315.n2 222.827
R54 a_1636_315.n1 a_1636_315.t2 169.726
R55 a_1636_315.n0 a_1636_315.t3 167.63
R56 a_1636_315.n1 a_1636_315.n0 152
R57 a_1636_315.n2 a_1636_315.n1 21.8174
R58 a_1565_49.n0 a_1565_49.t2 789.159
R59 a_1565_49.n1 a_1565_49.t0 174.72
R60 a_1565_49.n0 a_1565_49.t1 20.9089
R61 a_1565_49.n2 a_1565_49.n1 18.8622
R62 a_1565_49.n1 a_1565_49.n0 12.9785
R63 VGND.n14 VGND.t4 270.652
R64 VGND.n13 VGND.n12 208.719
R65 VGND.n1 VGND.n0 207.213
R66 VGND.n31 VGND.n30 110.424
R67 VGND.n30 VGND.t2 40.313
R68 VGND.n17 VGND.n11 34.6358
R69 VGND.n18 VGND.n17 34.6358
R70 VGND.n19 VGND.n18 34.6358
R71 VGND.n19 VGND.n9 34.6358
R72 VGND.n23 VGND.n9 34.6358
R73 VGND.n24 VGND.n23 34.6358
R74 VGND.n25 VGND.n24 34.6358
R75 VGND.n25 VGND.n7 34.6358
R76 VGND.n29 VGND.n7 34.6358
R77 VGND.n32 VGND.n5 34.6358
R78 VGND.n36 VGND.n5 34.6358
R79 VGND.n37 VGND.n36 34.6358
R80 VGND.n38 VGND.n37 34.6358
R81 VGND.n38 VGND.n3 34.6358
R82 VGND.n42 VGND.n3 34.6358
R83 VGND.n43 VGND.n42 34.6358
R84 VGND.n44 VGND.n43 34.6358
R85 VGND.n44 VGND.n1 32.7534
R86 VGND.n0 VGND.t3 30.938
R87 VGND.n12 VGND.t1 29.063
R88 VGND.n12 VGND.t6 28.73
R89 VGND.n13 VGND.n11 28.2358
R90 VGND.n0 VGND.t0 26.855
R91 VGND.n32 VGND.n31 26.3534
R92 VGND.n30 VGND.t5 24.0425
R93 VGND.n31 VGND.n29 18.0711
R94 VGND.n14 VGND.n13 13.9325
R95 VGND.n46 VGND.n1 9.54145
R96 VGND.n45 VGND.n44 9.3005
R97 VGND.n43 VGND.n2 9.3005
R98 VGND.n42 VGND.n41 9.3005
R99 VGND.n40 VGND.n3 9.3005
R100 VGND.n39 VGND.n38 9.3005
R101 VGND.n37 VGND.n4 9.3005
R102 VGND.n36 VGND.n35 9.3005
R103 VGND.n34 VGND.n5 9.3005
R104 VGND.n33 VGND.n32 9.3005
R105 VGND.n31 VGND.n6 9.3005
R106 VGND.n15 VGND.n11 9.3005
R107 VGND.n17 VGND.n16 9.3005
R108 VGND.n18 VGND.n10 9.3005
R109 VGND.n20 VGND.n19 9.3005
R110 VGND.n21 VGND.n9 9.3005
R111 VGND.n23 VGND.n22 9.3005
R112 VGND.n24 VGND.n8 9.3005
R113 VGND.n26 VGND.n25 9.3005
R114 VGND.n27 VGND.n7 9.3005
R115 VGND.n29 VGND.n28 9.3005
R116 VGND.n15 VGND.n14 0.214895
R117 VGND.n46 VGND.n45 0.141672
R118 VGND VGND.n46 0.121778
R119 VGND.n16 VGND.n15 0.120292
R120 VGND.n16 VGND.n10 0.120292
R121 VGND.n20 VGND.n10 0.120292
R122 VGND.n21 VGND.n20 0.120292
R123 VGND.n22 VGND.n21 0.120292
R124 VGND.n22 VGND.n8 0.120292
R125 VGND.n26 VGND.n8 0.120292
R126 VGND.n27 VGND.n26 0.120292
R127 VGND.n28 VGND.n27 0.120292
R128 VGND.n28 VGND.n6 0.120292
R129 VGND.n33 VGND.n6 0.120292
R130 VGND.n34 VGND.n33 0.120292
R131 VGND.n35 VGND.n34 0.120292
R132 VGND.n35 VGND.n4 0.120292
R133 VGND.n39 VGND.n4 0.120292
R134 VGND.n40 VGND.n39 0.120292
R135 VGND.n41 VGND.n40 0.120292
R136 VGND.n41 VGND.n2 0.120292
R137 VGND.n45 VGND.n2 0.120292
R138 VNB.t7 VNB.t3 8486.73
R139 VNB.t2 VNB.t1 3260.84
R140 VNB.t6 VNB.t4 2876.38
R141 VNB.t5 VNB.t0 2833.66
R142 VNB.t11 VNB.t9 2677.02
R143 VNB.t12 VNB.t10 2648.54
R144 VNB.t4 VNB.t12 1893.85
R145 VNB.t10 VNB.t5 1452.43
R146 VNB.t3 VNB.t11 1352.75
R147 VNB.t8 VNB.t2 1352.75
R148 VNB.t0 VNB.t7 1210.36
R149 VNB.t1 VNB.t6 1210.36
R150 VNB VNB.t8 939.807
R151 a_1647_49.n2 a_1647_49.n1 488.366
R152 a_1647_49.n1 a_1647_49.t2 241.536
R153 a_1647_49.n1 a_1647_49.n0 169.237
R154 a_1647_49.t0 a_1647_49.n2 31.6612
R155 a_1647_49.n2 a_1647_49.t1 31.6612
R156 VPWR.n48 VPWR.n1 606.836
R157 VPWR.n16 VPWR.n13 605.707
R158 VPWR.n7 VPWR.n6 600.515
R159 VPWR.n15 VPWR.n14 324.483
R160 VPWR.n6 VPWR.t7 44.3255
R161 VPWR.n49 VPWR.n48 43.5593
R162 VPWR.n1 VPWR.t2 42.3555
R163 VPWR.n35 VPWR.n34 34.6358
R164 VPWR.n36 VPWR.n35 34.6358
R165 VPWR.n36 VPWR.n4 34.6358
R166 VPWR.n40 VPWR.n4 34.6358
R167 VPWR.n41 VPWR.n40 34.6358
R168 VPWR.n42 VPWR.n41 34.6358
R169 VPWR.n42 VPWR.n2 34.6358
R170 VPWR.n46 VPWR.n2 34.6358
R171 VPWR.n47 VPWR.n46 34.6358
R172 VPWR.n18 VPWR.n17 34.6358
R173 VPWR.n18 VPWR.n11 34.6358
R174 VPWR.n22 VPWR.n11 34.6358
R175 VPWR.n23 VPWR.n22 34.6358
R176 VPWR.n24 VPWR.n23 34.6358
R177 VPWR.n24 VPWR.n9 34.6358
R178 VPWR.n28 VPWR.n9 34.6358
R179 VPWR.n29 VPWR.n28 34.6358
R180 VPWR.n30 VPWR.n29 34.6358
R181 VPWR.n34 VPWR.n7 32.377
R182 VPWR.n17 VPWR.n16 28.9887
R183 VPWR.n1 VPWR.t0 26.5955
R184 VPWR.n6 VPWR.t4 26.5955
R185 VPWR.n13 VPWR.t6 26.5955
R186 VPWR.n13 VPWR.t3 26.5955
R187 VPWR.n14 VPWR.t1 26.5955
R188 VPWR.n14 VPWR.t5 26.5955
R189 VPWR.n16 VPWR.n15 13.1909
R190 VPWR.n30 VPWR.n7 12.0476
R191 VPWR.n17 VPWR.n12 9.3005
R192 VPWR.n19 VPWR.n18 9.3005
R193 VPWR.n20 VPWR.n11 9.3005
R194 VPWR.n22 VPWR.n21 9.3005
R195 VPWR.n23 VPWR.n10 9.3005
R196 VPWR.n25 VPWR.n24 9.3005
R197 VPWR.n26 VPWR.n9 9.3005
R198 VPWR.n28 VPWR.n27 9.3005
R199 VPWR.n29 VPWR.n8 9.3005
R200 VPWR.n31 VPWR.n30 9.3005
R201 VPWR.n32 VPWR.n7 9.3005
R202 VPWR.n34 VPWR.n33 9.3005
R203 VPWR.n35 VPWR.n5 9.3005
R204 VPWR.n37 VPWR.n36 9.3005
R205 VPWR.n38 VPWR.n4 9.3005
R206 VPWR.n40 VPWR.n39 9.3005
R207 VPWR.n41 VPWR.n3 9.3005
R208 VPWR.n43 VPWR.n42 9.3005
R209 VPWR.n44 VPWR.n2 9.3005
R210 VPWR.n46 VPWR.n45 9.3005
R211 VPWR.n47 VPWR.n0 9.3005
R212 VPWR.n48 VPWR.n47 0.376971
R213 VPWR.n15 VPWR.n12 0.203949
R214 VPWR.n19 VPWR.n12 0.120292
R215 VPWR.n20 VPWR.n19 0.120292
R216 VPWR.n21 VPWR.n20 0.120292
R217 VPWR.n21 VPWR.n10 0.120292
R218 VPWR.n25 VPWR.n10 0.120292
R219 VPWR.n26 VPWR.n25 0.120292
R220 VPWR.n27 VPWR.n26 0.120292
R221 VPWR.n27 VPWR.n8 0.120292
R222 VPWR.n31 VPWR.n8 0.120292
R223 VPWR.n32 VPWR.n31 0.120292
R224 VPWR.n33 VPWR.n32 0.120292
R225 VPWR.n33 VPWR.n5 0.120292
R226 VPWR.n37 VPWR.n5 0.120292
R227 VPWR.n38 VPWR.n37 0.120292
R228 VPWR.n39 VPWR.n38 0.120292
R229 VPWR.n39 VPWR.n3 0.120292
R230 VPWR.n43 VPWR.n3 0.120292
R231 VPWR.n44 VPWR.n43 0.120292
R232 VPWR.n45 VPWR.n44 0.120292
R233 VPWR.n45 VPWR.n0 0.120292
R234 VPWR.n49 VPWR.n0 0.120292
R235 VPWR VPWR.n49 0.0226354
R236 SUM SUM.t0 371.428
R237 CIN.n1 CIN.t2 215.732
R238 CIN.n0 CIN.t1 212.081
R239 CIN CIN.n2 153.583
R240 CIN.n1 CIN.t3 139.78
R241 CIN.n0 CIN.t0 138.173
R242 CIN.n2 CIN.n0 100.052
R243 CIN.n2 CIN.n1 37.246
R244 a_1251_49.n0 a_1251_49.t3 440.846
R245 a_1251_49.n0 a_1251_49.t0 324.721
R246 a_1251_49.t2 a_1251_49.n1 266.731
R247 a_1251_49.n1 a_1251_49.t1 228.805
R248 a_1251_49.n1 a_1251_49.n0 21.8028
R249 a_67_199.t0 a_67_199.n7 699.885
R250 a_67_199.n0 a_67_199.t1 631.12
R251 a_67_199.n0 a_67_199.t4 629.452
R252 a_67_199.n1 a_67_199.t5 310.173
R253 a_67_199.n5 a_67_199.t6 236.18
R254 a_67_199.n2 a_67_199.n1 185
R255 a_67_199.n5 a_67_199.t7 165.488
R256 a_67_199.n6 a_67_199.n5 152
R257 a_67_199.n8 a_67_199.t0 126.081
R258 a_67_199.n3 a_67_199.n2 123.984
R259 a_67_199.n4 a_67_199.n3 95.0816
R260 a_67_199.n7 a_67_199.n6 69.5733
R261 a_67_199.n7 a_67_199.n0 63.6505
R262 a_67_199.n6 a_67_199.n4 45.5608
R263 a_67_199.n4 a_67_199.n1 41.2771
R264 a_67_199.n2 a_67_199.t2 25.313
R265 a_67_199.n3 a_67_199.t3 14.1839
R266 B.n2 B.t0 244.798
R267 B.n4 B.n0 233.519
R268 B.n1 B.t4 212.081
R269 B.n0 B.t2 186.374
R270 B B.n3 179.536
R271 B.n1 B.t3 139.78
R272 B.n0 B.t1 138.173
R273 B.n2 B.t5 138.173
R274 B.n3 B.n1 116.849
R275 B.n3 B.n2 18.9884
R276 B.n4 B 9.3005
R277 B B.n4 4.73093
R278 a_434_49.n6 a_434_49.n5 610.386
R279 a_434_49.n2 a_434_49.t5 246.482
R280 a_434_49.n2 a_434_49.n1 214.821
R281 a_434_49.n3 a_434_49.t6 202.28
R282 a_434_49.n5 a_434_49.n0 198.59
R283 a_434_49.n4 a_434_49.n2 165.602
R284 a_434_49.n4 a_434_49.n3 163.816
R285 a_434_49.n3 a_434_49.t4 154.079
R286 a_434_49.t1 a_434_49.n6 32.8338
R287 a_434_49.n6 a_434_49.t2 31.6612
R288 a_434_49.n0 a_434_49.t0 26.2505
R289 a_434_49.n0 a_434_49.t3 25.313
R290 a_434_49.n5 a_434_49.n4 12.909
R291 COUT COUT.n0 593.297
R292 COUT COUT.n1 216.15
R293 COUT.n0 COUT.t3 31.6612
R294 COUT.n0 COUT.t0 31.6612
R295 COUT.n1 COUT.t2 26.2505
R296 COUT.n1 COUT.t1 25.313
R297 A.n0 A.t0 230.363
R298 A A.n0 159.041
R299 A.n0 A.t1 158.064
R300 a_1142_49.n3 a_1142_49.n2 595.465
R301 a_1142_49.n1 a_1142_49.n0 585
R302 a_1142_49.n1 a_1142_49.t3 405.216
R303 a_1142_49.n2 a_1142_49.t1 276.404
R304 a_1142_49.n4 a_1142_49.n0 79.7386
R305 a_1142_49.n2 a_1142_49.n1 47.3703
R306 a_1142_49.n0 a_1142_49.t0 31.6612
R307 a_1142_49.n4 a_1142_49.n3 24.8276
R308 a_1142_49.n5 a_1142_49.n4 24.8194
R309 a_1142_49.n3 a_1142_49.t2 18.6209
C0 VPB A 0.042156f
C1 COUT VGND 0.005343f
C2 VPB VPWR 0.251728f
C3 SUM VGND 0.071984f
C4 VPB B 0.1721f
C5 A VPWR 0.012725f
C6 VPB CIN 0.089133f
C7 A B 0.052221f
C8 VPWR B 0.033833f
C9 VPB COUT 0.003252f
C10 VPWR CIN 0.028875f
C11 VPB SUM 0.013578f
C12 VPB VGND 0.008044f
C13 VPWR COUT 0.003816f
C14 A VGND 0.01514f
C15 B COUT 3.09e-19
C16 VPWR SUM 0.106873f
C17 VPWR VGND 0.044946f
C18 B SUM 9.28e-23
C19 B VGND 0.208167f
C20 CIN SUM 0.002316f
C21 CIN VGND 0.031418f
C22 VGND VNB 1.33068f
C23 SUM VNB 0.093722f
C24 COUT VNB 0.006405f
C25 CIN VNB 0.230607f
C26 B VNB 0.390988f
C27 VPWR VNB 1.08951f
C28 A VNB 0.109448f
C29 VPB VNB 2.46528f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fahcon_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fahcon_1 VPWR VGND VNB VPB SUM CI COUT_N B A
X0 a_1144_49.t2 B.t0 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.3826 pd=1.79 as=0.18 ps=1.36 w=1 l=0.15
X1 VPWR.t6 a_67_199.t6 a_28_47.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.26 ps=2.52 w=1 l=0.15
X2 VGND.t4 B.t1 a_488_21.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.11005 pd=0.99 as=0.16715 ps=1.82 w=0.65 l=0.15
X3 a_1589_49.t0 a_434_49.t4 a_1710_49.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.3024 pd=2.4 as=0.1134 ps=1.11 w=0.84 l=0.15
X4 SUM.t0 a_1710_49.t4 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10525 ps=0.975 w=0.65 l=0.15
X5 a_1710_49.t3 a_726_47.t4 a_1634_315.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2352 ps=2.24 w=0.84 l=0.15
X6 a_434_49.t1 B.t2 a_67_199.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.321225 ps=1.645 w=0.64 l=0.15
X7 a_434_49.t0 B.t3 a_28_47.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2629 ps=2.64 w=0.84 l=0.15
X8 a_1589_49.t3 CI.t0 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X9 COUT_N.t1 a_434_49.t5 a_1144_49.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.3826 ps=1.79 w=0.84 l=0.15
X10 a_1144_49.t3 a_726_47.t5 COUT_N.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1952 pd=1.89 as=0.088 ps=0.915 w=0.64 l=0.15
X11 SUM.t1 a_1710_49.t5 VPWR.t5 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X12 a_67_199.t0 A.t0 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.3184 pd=2.88 as=0.175 ps=1.35 w=1 l=0.15
X13 a_28_47.t2 B.t4 a_726_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.16285 pd=1.8 as=0.165675 ps=1.165 w=0.64 l=0.15
X14 VPWR.t4 CI.t1 a_1261_49.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t7 a_67_199.t7 a_28_47.t4 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 a_28_47.t0 a_488_21.t2 a_434_49.t2 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.2176 pd=1.96 as=0.0864 ps=0.91 w=0.64 l=0.15
X17 a_1144_49.t1 B.t5 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.11005 ps=0.99 w=0.64 l=0.15
X18 a_726_47.t2 a_488_21.t3 a_28_47.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.151625 pd=1.3 as=0.3314 ps=2.75 w=0.84 l=0.15
X19 a_67_199.t1 A.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.321225 pd=1.645 as=0.10525 ps=0.975 w=0.65 l=0.15
X20 VPWR.t1 a_1589_49.t4 a_1634_315.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.35 ps=2.7 w=1 l=0.15
X21 a_726_47.t3 a_488_21.t4 a_67_199.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.165675 pd=1.165 as=0.1792 ps=1.84 w=0.64 l=0.15
X22 a_1710_49.t2 a_726_47.t6 a_1589_49.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0928 pd=0.93 as=0.2912 ps=2.19 w=0.64 l=0.15
X23 a_1634_315.t1 a_434_49.t6 a_1710_49.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.3136 pd=1.62 as=0.0928 ps=0.93 w=0.64 l=0.15
X24 a_67_199.t3 B.t6 a_726_47.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=2.24 as=0.151625 ps=1.3 w=0.84 l=0.15
X25 a_1589_49.t2 CI.t2 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10525 ps=0.975 w=0.65 l=0.15
X26 a_67_199.t4 a_488_21.t5 a_434_49.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.1134 ps=1.11 w=0.84 l=0.15
X27 VPWR.t3 B.t7 a_488_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.26 ps=2.52 w=1 l=0.15
X28 VGND.t0 a_1589_49.t5 a_1634_315.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.3136 ps=1.62 w=0.64 l=0.15
X29 a_1261_49.t0 a_726_47.t7 COUT_N.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.4536 pd=2.76 as=0.1134 ps=1.11 w=0.84 l=0.15
X30 VGND.t1 CI.t3 a_1261_49.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10525 pd=0.975 as=0.1664 ps=1.8 w=0.64 l=0.15
R0 B.n4 B.t6 246.258
R1 B.n6 B.n0 230.964
R2 B.n1 B.t0 212.081
R3 B.n3 B.t7 212.081
R4 B.n0 B.t3 186.374
R5 B B.n5 179.558
R6 B.n2 B.t1 139.78
R7 B.n0 B.t2 138.173
R8 B.n1 B.t5 138.173
R9 B.n4 B.t4 138.173
R10 B.n5 B.n3 114.659
R11 B.n2 B.n1 71.5702
R12 B.n5 B.n4 18.9884
R13 B.n6 B 9.3005
R14 B B.n6 4.03013
R15 B.n3 B.n2 2.92171
R16 VPWR.n48 VPWR.n1 606.836
R17 VPWR.n7 VPWR.n6 600.515
R18 VPWR.n16 VPWR.n15 598.755
R19 VPWR.n14 VPWR.n13 324.478
R20 VPWR.n6 VPWR.t3 44.3255
R21 VPWR.n49 VPWR.n48 43.5593
R22 VPWR.n1 VPWR.t0 42.3555
R23 VPWR.n35 VPWR.n34 34.6358
R24 VPWR.n36 VPWR.n35 34.6358
R25 VPWR.n36 VPWR.n4 34.6358
R26 VPWR.n40 VPWR.n4 34.6358
R27 VPWR.n41 VPWR.n40 34.6358
R28 VPWR.n42 VPWR.n41 34.6358
R29 VPWR.n42 VPWR.n2 34.6358
R30 VPWR.n46 VPWR.n2 34.6358
R31 VPWR.n47 VPWR.n46 34.6358
R32 VPWR.n18 VPWR.n17 34.6358
R33 VPWR.n18 VPWR.n11 34.6358
R34 VPWR.n22 VPWR.n11 34.6358
R35 VPWR.n23 VPWR.n22 34.6358
R36 VPWR.n24 VPWR.n23 34.6358
R37 VPWR.n24 VPWR.n9 34.6358
R38 VPWR.n28 VPWR.n9 34.6358
R39 VPWR.n29 VPWR.n28 34.6358
R40 VPWR.n30 VPWR.n29 34.6358
R41 VPWR.n34 VPWR.n7 33.1299
R42 VPWR.n1 VPWR.t6 26.5955
R43 VPWR.n6 VPWR.t2 26.5955
R44 VPWR.n15 VPWR.t7 26.5955
R45 VPWR.n15 VPWR.t1 26.5955
R46 VPWR.n13 VPWR.t5 26.5955
R47 VPWR.n13 VPWR.t4 26.5955
R48 VPWR.n17 VPWR.n16 17.3181
R49 VPWR.n30 VPWR.n7 11.2946
R50 VPWR.n17 VPWR.n12 9.3005
R51 VPWR.n19 VPWR.n18 9.3005
R52 VPWR.n20 VPWR.n11 9.3005
R53 VPWR.n22 VPWR.n21 9.3005
R54 VPWR.n23 VPWR.n10 9.3005
R55 VPWR.n25 VPWR.n24 9.3005
R56 VPWR.n26 VPWR.n9 9.3005
R57 VPWR.n28 VPWR.n27 9.3005
R58 VPWR.n29 VPWR.n8 9.3005
R59 VPWR.n31 VPWR.n30 9.3005
R60 VPWR.n32 VPWR.n7 9.3005
R61 VPWR.n34 VPWR.n33 9.3005
R62 VPWR.n35 VPWR.n5 9.3005
R63 VPWR.n37 VPWR.n36 9.3005
R64 VPWR.n38 VPWR.n4 9.3005
R65 VPWR.n40 VPWR.n39 9.3005
R66 VPWR.n41 VPWR.n3 9.3005
R67 VPWR.n43 VPWR.n42 9.3005
R68 VPWR.n44 VPWR.n2 9.3005
R69 VPWR.n46 VPWR.n45 9.3005
R70 VPWR.n47 VPWR.n0 9.3005
R71 VPWR.n16 VPWR.n14 7.22798
R72 VPWR.n48 VPWR.n47 0.376971
R73 VPWR.n14 VPWR.n12 0.217427
R74 VPWR.n19 VPWR.n12 0.120292
R75 VPWR.n20 VPWR.n19 0.120292
R76 VPWR.n21 VPWR.n20 0.120292
R77 VPWR.n21 VPWR.n10 0.120292
R78 VPWR.n25 VPWR.n10 0.120292
R79 VPWR.n26 VPWR.n25 0.120292
R80 VPWR.n27 VPWR.n26 0.120292
R81 VPWR.n27 VPWR.n8 0.120292
R82 VPWR.n31 VPWR.n8 0.120292
R83 VPWR.n32 VPWR.n31 0.120292
R84 VPWR.n33 VPWR.n32 0.120292
R85 VPWR.n33 VPWR.n5 0.120292
R86 VPWR.n37 VPWR.n5 0.120292
R87 VPWR.n38 VPWR.n37 0.120292
R88 VPWR.n39 VPWR.n38 0.120292
R89 VPWR.n39 VPWR.n3 0.120292
R90 VPWR.n43 VPWR.n3 0.120292
R91 VPWR.n44 VPWR.n43 0.120292
R92 VPWR.n45 VPWR.n44 0.120292
R93 VPWR.n45 VPWR.n0 0.120292
R94 VPWR.n49 VPWR.n0 0.120292
R95 VPWR VPWR.n49 0.0226354
R96 a_1144_49.n3 a_1144_49.n2 595.465
R97 a_1144_49.n1 a_1144_49.n0 585
R98 a_1144_49.n1 a_1144_49.t3 398.366
R99 a_1144_49.n2 a_1144_49.t1 276.774
R100 a_1144_49.n4 a_1144_49.n0 79.7386
R101 a_1144_49.n2 a_1144_49.n1 47.3703
R102 a_1144_49.n0 a_1144_49.t0 31.6612
R103 a_1144_49.n4 a_1144_49.n3 24.8276
R104 a_1144_49.n5 a_1144_49.n4 24.8194
R105 a_1144_49.n3 a_1144_49.t2 18.6209
R106 VPB.t0 VPB.t14 899.688
R107 VPB.t1 VPB.t4 668.847
R108 VPB.t3 VPB.t7 662.928
R109 VPB.t10 VPB.t13 642.212
R110 VPB.t6 VPB.t5 621.495
R111 VPB.t15 VPB.t9 571.184
R112 VPB.t8 VPB.t2 556.386
R113 VPB.t5 VPB.t8 301.87
R114 VPB.t12 VPB.t3 295.95
R115 VPB.t13 VPB.t6 287.072
R116 VPB.t9 VPB.t11 248.599
R117 VPB.t4 VPB.t15 248.599
R118 VPB.t14 VPB.t1 248.599
R119 VPB.t2 VPB.t0 248.599
R120 VPB.t7 VPB.t10 248.599
R121 VPB VPB.t12 195.327
R122 a_67_199.n0 a_67_199.t4 719.438
R123 a_67_199.t0 a_67_199.n7 705.562
R124 a_67_199.n0 a_67_199.t3 642.293
R125 a_67_199.n1 a_67_199.t5 301.834
R126 a_67_199.n5 a_67_199.t6 236.18
R127 a_67_199.n2 a_67_199.n1 185
R128 a_67_199.n5 a_67_199.t7 165.488
R129 a_67_199.n6 a_67_199.n5 152
R130 a_67_199.n8 a_67_199.t0 141.84
R131 a_67_199.n3 a_67_199.n2 123.984
R132 a_67_199.n4 a_67_199.n3 95.0816
R133 a_67_199.n7 a_67_199.n6 69.5733
R134 a_67_199.n6 a_67_199.n4 45.5608
R135 a_67_199.n4 a_67_199.n1 41.2771
R136 a_67_199.n2 a_67_199.t2 25.313
R137 a_67_199.n7 a_67_199.n0 15.0593
R138 a_67_199.n3 a_67_199.t1 14.1839
R139 a_28_47.n2 a_28_47.t1 745.086
R140 a_28_47.n1 a_28_47.t3 391.714
R141 a_28_47.n0 a_28_47.t2 315.613
R142 a_28_47.n0 a_28_47.t0 260.591
R143 a_28_47.t5 a_28_47.n3 221.34
R144 a_28_47.n3 a_28_47.t4 216.822
R145 a_28_47.n2 a_28_47.n1 137.619
R146 a_28_47.n3 a_28_47.n2 121.754
R147 a_28_47.n1 a_28_47.n0 76.422
R148 a_488_21.t1 a_488_21.n3 849.337
R149 a_488_21.n3 a_488_21.t0 247.546
R150 a_488_21.n0 a_488_21.t3 192.946
R151 a_488_21.n1 a_488_21.t5 186.374
R152 a_488_21.n3 a_488_21.n2 182.438
R153 a_488_21.n0 a_488_21.t4 141.387
R154 a_488_21.n1 a_488_21.t2 138.173
R155 a_488_21.n2 a_488_21.n0 108.816
R156 a_488_21.n2 a_488_21.n1 43.0884
R157 VGND.n14 VGND.n13 208.719
R158 VGND.n15 VGND.n12 208.282
R159 VGND.n1 VGND.n0 207.213
R160 VGND.n32 VGND.n31 110.424
R161 VGND.n31 VGND.t3 38.438
R162 VGND.n18 VGND.n11 34.6358
R163 VGND.n19 VGND.n18 34.6358
R164 VGND.n20 VGND.n19 34.6358
R165 VGND.n20 VGND.n9 34.6358
R166 VGND.n24 VGND.n9 34.6358
R167 VGND.n25 VGND.n24 34.6358
R168 VGND.n26 VGND.n25 34.6358
R169 VGND.n26 VGND.n7 34.6358
R170 VGND.n30 VGND.n7 34.6358
R171 VGND.n33 VGND.n5 34.6358
R172 VGND.n37 VGND.n5 34.6358
R173 VGND.n38 VGND.n37 34.6358
R174 VGND.n39 VGND.n38 34.6358
R175 VGND.n39 VGND.n3 34.6358
R176 VGND.n43 VGND.n3 34.6358
R177 VGND.n44 VGND.n43 34.6358
R178 VGND.n45 VGND.n44 34.6358
R179 VGND.n45 VGND.n1 32.7534
R180 VGND.n12 VGND.t6 32.48
R181 VGND.n13 VGND.t0 30.938
R182 VGND.n0 VGND.t7 30.938
R183 VGND.n14 VGND.n11 29.7417
R184 VGND.n33 VGND.n32 27.8593
R185 VGND.n13 VGND.t5 26.855
R186 VGND.n0 VGND.t2 26.855
R187 VGND.n12 VGND.t1 25.313
R188 VGND.n31 VGND.t4 22.1675
R189 VGND.n32 VGND.n30 16.5652
R190 VGND.n15 VGND.n14 12.4327
R191 VGND.n47 VGND.n1 9.54145
R192 VGND.n46 VGND.n45 9.3005
R193 VGND.n44 VGND.n2 9.3005
R194 VGND.n43 VGND.n42 9.3005
R195 VGND.n41 VGND.n3 9.3005
R196 VGND.n40 VGND.n39 9.3005
R197 VGND.n38 VGND.n4 9.3005
R198 VGND.n37 VGND.n36 9.3005
R199 VGND.n35 VGND.n5 9.3005
R200 VGND.n34 VGND.n33 9.3005
R201 VGND.n32 VGND.n6 9.3005
R202 VGND.n16 VGND.n11 9.3005
R203 VGND.n18 VGND.n17 9.3005
R204 VGND.n19 VGND.n10 9.3005
R205 VGND.n21 VGND.n20 9.3005
R206 VGND.n22 VGND.n9 9.3005
R207 VGND.n24 VGND.n23 9.3005
R208 VGND.n25 VGND.n8 9.3005
R209 VGND.n27 VGND.n26 9.3005
R210 VGND.n28 VGND.n7 9.3005
R211 VGND.n30 VGND.n29 9.3005
R212 VGND.n16 VGND.n15 0.209004
R213 VGND.n47 VGND.n46 0.141672
R214 VGND VGND.n47 0.121778
R215 VGND.n17 VGND.n16 0.120292
R216 VGND.n17 VGND.n10 0.120292
R217 VGND.n21 VGND.n10 0.120292
R218 VGND.n22 VGND.n21 0.120292
R219 VGND.n23 VGND.n22 0.120292
R220 VGND.n23 VGND.n8 0.120292
R221 VGND.n27 VGND.n8 0.120292
R222 VGND.n28 VGND.n27 0.120292
R223 VGND.n29 VGND.n28 0.120292
R224 VGND.n29 VGND.n6 0.120292
R225 VGND.n34 VGND.n6 0.120292
R226 VGND.n35 VGND.n34 0.120292
R227 VGND.n36 VGND.n35 0.120292
R228 VGND.n36 VGND.n4 0.120292
R229 VGND.n40 VGND.n4 0.120292
R230 VGND.n41 VGND.n40 0.120292
R231 VGND.n42 VGND.n41 0.120292
R232 VGND.n42 VGND.n2 0.120292
R233 VGND.n46 VGND.n2 0.120292
R234 VNB.t4 VNB.t8 4044.01
R235 VNB.t8 VNB.t9 4015.53
R236 VNB.t3 VNB.t6 3260.84
R237 VNB.t0 VNB.t1 3218.12
R238 VNB.t14 VNB.t13 2961.81
R239 VNB.t10 VNB.t2 2677.02
R240 VNB.t5 VNB.t7 2662.78
R241 VNB.t13 VNB.t5 1893.85
R242 VNB.t7 VNB.t4 1395.47
R243 VNB.t2 VNB.t11 1352.75
R244 VNB.t1 VNB.t10 1352.75
R245 VNB.t12 VNB.t3 1352.75
R246 VNB.t9 VNB.t0 1253.07
R247 VNB.t6 VNB.t14 1196.12
R248 VNB VNB.t12 939.807
R249 a_434_49.n6 a_434_49.n5 595.899
R250 a_434_49.n1 a_434_49.t4 241.804
R251 a_434_49.n3 a_434_49.t5 202.28
R252 a_434_49.n5 a_434_49.n0 196.913
R253 a_434_49.n4 a_434_49.n1 165.95
R254 a_434_49.n1 a_434_49.t6 164.684
R255 a_434_49.n4 a_434_49.n3 163.816
R256 a_434_49.n3 a_434_49.n2 154.079
R257 a_434_49.n6 a_434_49.t3 31.6612
R258 a_434_49.t0 a_434_49.n6 31.6612
R259 a_434_49.n0 a_434_49.t2 25.313
R260 a_434_49.n0 a_434_49.t1 25.313
R261 a_434_49.n5 a_434_49.n4 12.9179
R262 a_1261_49.n0 a_1261_49.t0 463.384
R263 a_1261_49.t2 a_1261_49.n0 266.731
R264 a_1261_49.n0 a_1261_49.t1 228.805
R265 COUT_N COUT_N.n0 593.297
R266 COUT_N COUT_N.t2 301.241
R267 COUT_N.n0 COUT_N.t0 31.6612
R268 COUT_N.n0 COUT_N.t1 31.6612
R269 a_1710_49.n3 a_1710_49.n2 320.894
R270 a_1710_49.n2 a_1710_49.n0 253.381
R271 a_1710_49.n1 a_1710_49.t5 241.536
R272 a_1710_49.n2 a_1710_49.n1 196.952
R273 a_1710_49.n1 a_1710_49.t4 169.237
R274 a_1710_49.t0 a_1710_49.n3 31.6612
R275 a_1710_49.n3 a_1710_49.t3 31.6612
R276 a_1710_49.n0 a_1710_49.t2 29.063
R277 a_1710_49.n0 a_1710_49.t1 25.313
R278 a_1589_49.n2 a_1589_49.t0 342.923
R279 a_1589_49.n2 a_1589_49.t1 326.688
R280 a_1589_49.n0 a_1589_49.t4 241.536
R281 a_1589_49.t3 a_1589_49.n3 224.139
R282 a_1589_49.n1 a_1589_49.t2 169.726
R283 a_1589_49.n0 a_1589_49.t5 167.63
R284 a_1589_49.n1 a_1589_49.n0 152
R285 a_1589_49.n3 a_1589_49.n2 23.8428
R286 a_1589_49.n3 a_1589_49.n1 22.0383
R287 SUM SUM.t1 373.803
R288 SUM SUM.t0 154.212
R289 a_726_47.n4 a_726_47.n2 607.196
R290 a_726_47.n5 a_726_47.n4 585
R291 a_726_47.n4 a_726_47.n3 259.055
R292 a_726_47.n1 a_726_47.t7 195.137
R293 a_726_47.n0 a_726_47.t4 164.843
R294 a_726_47.n0 a_726_47.t6 138.173
R295 a_726_47.n1 a_726_47.t5 138.173
R296 a_726_47.n2 a_726_47.n1 130.725
R297 a_726_47.n3 a_726_47.t3 62.5944
R298 a_726_47.n2 a_726_47.n0 51.4326
R299 a_726_47.t1 a_726_47.n5 50.6612
R300 a_726_47.n5 a_726_47.t2 32.2493
R301 a_726_47.n3 a_726_47.t0 20.1091
R302 a_1634_315.n1 a_1634_315.t0 457.182
R303 a_1634_315.t3 a_1634_315.n1 319.853
R304 a_1634_315.n1 a_1634_315.n0 174.75
R305 a_1634_315.n0 a_1634_315.t1 156.562
R306 a_1634_315.n0 a_1634_315.t2 27.188
R307 CI.n1 CI.t0 215.732
R308 CI.n0 CI.t1 212.081
R309 CI CI.n2 153.583
R310 CI.n1 CI.t2 139.78
R311 CI.n0 CI.t3 138.173
R312 CI.n2 CI.n0 100.052
R313 CI.n2 CI.n1 37.246
R314 A.n0 A.t0 230.363
R315 A A.n0 159.041
R316 A.n0 A.t1 158.064
C0 SUM VGND 0.075174f
C1 A VPWR 0.012308f
C2 VPB A 0.042159f
C3 A B 0.052246f
C4 VPB VPWR 0.253651f
C5 VPWR B 0.037492f
C6 VPB B 0.215961f
C7 VPWR CI 0.032067f
C8 VPB CI 0.089916f
C9 VPWR COUT_N 0.003816f
C10 VPB COUT_N 0.003252f
C11 B COUT_N 3.12e-19
C12 A VGND 0.01514f
C13 VPWR SUM 0.10562f
C14 VPB SUM 0.013153f
C15 B SUM 1.16e-22
C16 VPWR VGND 0.041004f
C17 VPB VGND 0.009617f
C18 B VGND 0.232174f
C19 CI SUM 0.002133f
C20 CI VGND 0.031783f
C21 COUT_N VGND 0.005346f
C22 VGND VNB 1.3356f
C23 SUM VNB 0.093542f
C24 COUT_N VNB 0.006459f
C25 CI VNB 0.230588f
C26 B VNB 0.497319f
C27 VPWR VNB 1.08652f
C28 A VNB 0.109448f
C29 VPB VNB 2.46528f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_1 VPWR VGND VPB VNB
C0 VGND VPWR 0.012627f
C1 VGND VPB 0.006841f
C2 VPWR VPB 0.022269f
C3 VGND VNB 0.112285f
C4 VPWR VNB 0.096857f
C5 VPB VNB 0.161784f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_2 VGND VPWR VPB VNB
C0 VGND VPB 0.013682f
C1 VPB VPWR 0.041139f
C2 VGND VPWR 0.025254f
C3 VGND VNB 0.171784f
C4 VPWR VNB 0.144327f
C5 VPB VNB 0.25038f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_4 VGND VPWR VPB VNB
C0 VGND VPB 0.027364f
C1 VGND VPWR 0.050509f
C2 VPB VPWR 0.078879f
C3 VGND VNB 0.290784f
C4 VPWR VNB 0.239269f
C5 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_8 VGND VPWR VPB VNB
C0 VPB VGND 0.054729f
C1 VPB VPWR 0.15436f
C2 VPWR VGND 0.101017f
C3 VGND VNB 0.528782f
C4 VPWR VNB 0.429151f
C5 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ha_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ha_1 VNB VPB VGND VPWR SUM B A COUT
X0 a_297_47.t2 a_250_199.t3 a_79_21.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_297_47.t0 A.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 COUT.t0 a_250_199.t4 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 a_250_199.t0 B.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X4 a_376_413.t1 B.t1 a_79_21.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_79_21.t1 a_250_199.t5 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X6 a_674_47.t1 B.t2 a_250_199.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR.t0 A.t1 a_376_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X8 VGND.t3 B.t3 a_297_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 COUT.t1 a_250_199.t6 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR.t2 a_79_21.t3 SUM.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X11 VPWR.t1 A.t2 a_250_199.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X12 VGND.t1 A.t3 a_674_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 VGND.t2 a_79_21.t4 SUM.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_250_199.n4 a_250_199.n3 680.346
R1 a_250_199.n0 a_250_199.t5 334.723
R2 a_250_199.n1 a_250_199.n0 287.906
R3 a_250_199.n2 a_250_199.t4 241.536
R4 a_250_199.n1 a_250_199.t2 239.007
R5 a_250_199.n0 a_250_199.t3 206.19
R6 a_250_199.n2 a_250_199.t6 169.237
R7 a_250_199.n3 a_250_199.n2 152
R8 a_250_199.n3 a_250_199.n1 77.6519
R9 a_250_199.n4 a_250_199.t1 68.0124
R10 a_250_199.t0 a_250_199.n4 68.0124
R11 a_79_21.n2 a_79_21.n1 684.765
R12 a_79_21.n1 a_79_21.t2 260.188
R13 a_79_21.n0 a_79_21.t3 232.214
R14 a_79_21.n1 a_79_21.n0 181.365
R15 a_79_21.n0 a_79_21.t4 159.915
R16 a_79_21.t0 a_79_21.n2 63.3219
R17 a_79_21.n2 a_79_21.t1 63.3219
R18 a_297_47.t0 a_297_47.n0 490.642
R19 a_297_47.n0 a_297_47.t1 38.5719
R20 a_297_47.n0 a_297_47.t2 38.5719
R21 VNB.t1 VNB.t4 2976.05
R22 VNB.t2 VNB.t6 2677.02
R23 VNB.t0 VNB.t5 1352.75
R24 VNB.t3 VNB.t1 1196.12
R25 VNB.t6 VNB.t3 1196.12
R26 VNB.t4 VNB.t0 1025.24
R27 VNB VNB.t2 911.327
R28 A.n0 A.t0 405.293
R29 A.n1 A.t2 274.51
R30 A.n0 A.t1 250.549
R31 A.n1 A.t3 248.804
R32 A.n3 A.n0 216.754
R33 A.n2 A.n1 152
R34 A.n2 A 12.2316
R35 A.n3 A.n2 4.55161
R36 A A.n3 2.5605
R37 VGND.n4 VGND.n3 210.816
R38 VGND.n2 VGND.n1 199.739
R39 VGND.n8 VGND.t2 162.178
R40 VGND.n3 VGND.t1 54.2862
R41 VGND.n1 VGND.t0 38.5719
R42 VGND.n1 VGND.t3 38.5719
R43 VGND.n7 VGND.n6 34.6358
R44 VGND.n8 VGND.n7 27.1064
R45 VGND.n3 VGND.t4 25.9346
R46 VGND.n6 VGND.n2 19.9534
R47 VGND.n6 VGND.n5 9.3005
R48 VGND.n7 VGND.n0 9.3005
R49 VGND.n9 VGND.n8 7.4049
R50 VGND.n4 VGND.n2 7.17218
R51 VGND.n5 VGND.n4 0.166386
R52 VGND.n9 VGND.n0 0.144904
R53 VGND.n5 VGND.n0 0.120292
R54 VGND VGND.n9 0.117202
R55 VPWR.n5 VPWR.n4 612.782
R56 VPWR.n17 VPWR.n16 585
R57 VPWR.n20 VPWR.n19 585
R58 VPWR.n9 VPWR.n8 585
R59 VPWR.n7 VPWR.n6 585
R60 VPWR.n18 VPWR.n1 316.413
R61 VPWR.n19 VPWR.n17 194.655
R62 VPWR.n8 VPWR.n7 159.476
R63 VPWR.n17 VPWR.t5 100.846
R64 VPWR.n4 VPWR.t1 89.1195
R65 VPWR.n7 VPWR.t3 86.7743
R66 VPWR.n8 VPWR.t0 86.7743
R67 VPWR.n21 VPWR.n20 38.8357
R68 VPWR.n11 VPWR.n2 34.6358
R69 VPWR.n11 VPWR.n10 30.5443
R70 VPWR.n4 VPWR.t4 29.316
R71 VPWR.n15 VPWR.n2 29.01
R72 VPWR.n18 VPWR.t2 25.6105
R73 VPWR.n16 VPWR.n1 9.78163
R74 VPWR.n10 VPWR.n3 9.3005
R75 VPWR.n12 VPWR.n11 9.3005
R76 VPWR.n13 VPWR.n2 9.3005
R77 VPWR.n15 VPWR.n14 9.3005
R78 VPWR.n1 VPWR.n0 9.3005
R79 VPWR.n9 VPWR.n6 8.21182
R80 VPWR.n6 VPWR.n5 7.81091
R81 VPWR.n19 VPWR.n18 2.34574
R82 VPWR.n10 VPWR.n9 2.05333
R83 VPWR.n16 VPWR.n15 1.3288
R84 VPWR.n5 VPWR.n3 0.514096
R85 VPWR.n20 VPWR.n1 0.242009
R86 VPWR.n12 VPWR.n3 0.120292
R87 VPWR.n13 VPWR.n12 0.120292
R88 VPWR.n14 VPWR.n13 0.120292
R89 VPWR.n14 VPWR.n0 0.120292
R90 VPWR.n21 VPWR.n0 0.120292
R91 VPWR VPWR.n21 0.0213333
R92 COUT COUT.n0 592.718
R93 COUT.n3 COUT.n0 585
R94 COUT.n2 COUT.n0 585
R95 COUT.n1 COUT.t1 129.036
R96 COUT.n2 COUT.n1 63.4912
R97 COUT.n0 COUT.t0 26.5955
R98 COUT.n3 COUT 7.71815
R99 COUT.n1 COUT 5.70906
R100 COUT COUT.n3 5.08285
R101 COUT COUT.n2 5.08285
R102 VPB.t2 VPB.t5 541.59
R103 VPB.t1 VPB.t3 509.034
R104 VPB.t4 VPB.t1 325.546
R105 VPB.t0 VPB.t6 281.154
R106 VPB.t3 VPB.t0 260.437
R107 VPB.t5 VPB.t4 248.599
R108 VPB VPB.t2 189.409
R109 B.n0 B.t2 419.877
R110 B.n2 B.t3 360.791
R111 B.n1 B.n0 215.625
R112 B.n2 B.t1 167.992
R113 B.n0 B.t0 154.23
R114 B.n3 B.n2 152
R115 B B.n3 9.02345
R116 B.n3 B.n1 3.35788
R117 B.n1 B 1.88902
R118 a_376_413.t0 a_376_413.t1 187.619
R119 a_674_47.t0 a_674_47.t1 60.0005
R120 SUM SUM.n0 592.833
R121 SUM.n5 SUM.n0 585
R122 SUM.n4 SUM.n0 585
R123 SUM.n1 SUM.t1 128.996
R124 SUM.n0 SUM.t0 26.5955
R125 SUM SUM.n2 15.5831
R126 SUM.n5 SUM 7.83334
R127 SUM SUM.n1 6.93222
R128 SUM.n3 SUM 6.67876
R129 SUM.n1 SUM 5.79252
R130 SUM SUM.n5 5.15871
R131 SUM SUM.n4 5.15871
R132 SUM.n3 SUM 4.58557
R133 SUM.n2 SUM 3.33963
R134 SUM.n4 SUM.n3 3.24826
R135 SUM.n2 SUM 2.29304
C0 VPB VPWR 0.105209f
C1 VPB VGND 0.011728f
C2 B VPWR 0.122694f
C3 A VPWR 0.043268f
C4 B VGND 0.032029f
C5 VPB COUT 0.010336f
C6 B COUT 4.25e-19
C7 A VGND 0.035082f
C8 SUM VPWR 0.115405f
C9 SUM VGND 0.086113f
C10 A COUT 0.004901f
C11 VPWR VGND 0.09142f
C12 VPWR COUT 0.067632f
C13 VGND COUT 0.060529f
C14 VPB B 0.181716f
C15 VPB A 0.171249f
C16 B A 0.366423f
C17 VPB SUM 0.011264f
C18 COUT VNB 0.089579f
C19 VGND VNB 0.554977f
C20 VPWR VNB 0.448883f
C21 SUM VNB 0.089208f
C22 A VNB 0.255924f
C23 B VNB 0.236166f
C24 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ha_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ha_2 VNB VPB VGND VPWR COUT A B SUM
X0 VPWR.t0 A.t0 a_342_199.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.0928 ps=0.93 w=0.64 l=0.15
X1 a_766_47.t1 B.t0 a_342_199.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND.t5 B.t1 a_389_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 COUT.t1 a_342_199.t3 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND.t1 A.t1 a_766_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_342_199.t2 B.t2 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.2272 ps=1.35 w=0.64 l=0.15
X6 a_468_369.t1 B.t3 a_79_21.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.04 as=0.0864 ps=0.91 w=0.64 l=0.15
X7 a_79_21.t1 a_342_199.t4 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.2916 ps=1.765 w=0.64 l=0.15
X8 a_389_47.t1 a_342_199.t5 a_79_21.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_389_47.t0 A.t2 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 COUT.t3 a_342_199.t6 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.149 ps=1.325 w=1 l=0.15
X11 VPWR.t2 a_342_199.t7 COUT.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X12 VGND.t6 a_79_21.t3 SUM.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13 VPWR.t6 a_79_21.t4 SUM.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.2916 pd=1.765 as=0.155 ps=1.31 w=1 l=0.15
X14 VGND.t3 a_342_199.t8 COUT.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X15 SUM.t2 a_79_21.t5 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR.t1 A.t3 a_468_369.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2272 pd=1.35 as=0.128 ps=1.04 w=0.64 l=0.15
X17 SUM.t0 a_79_21.t6 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n0 A.t3 299.07
R1 A.n2 A.t0 272.747
R2 A.n2 A.t1 224.547
R3 A.n1 A.n0 217.13
R4 A.n0 A.t2 166.52
R5 A.n3 A.n2 152
R6 A A.n3 12.2316
R7 A.n3 A.n1 5.1205
R8 A.n1 A 1.99161
R9 a_342_199.n5 a_342_199.n4 597.424
R10 a_342_199.n4 a_342_199.n3 358.683
R11 a_342_199.n2 a_342_199.t1 316.659
R12 a_342_199.n3 a_342_199.t4 299.377
R13 a_342_199.n0 a_342_199.t7 212.081
R14 a_342_199.n1 a_342_199.t6 212.081
R15 a_342_199.n3 a_342_199.t5 206.19
R16 a_342_199.n2 a_342_199.n1 160.034
R17 a_342_199.n0 a_342_199.t8 139.78
R18 a_342_199.n1 a_342_199.t3 139.78
R19 a_342_199.n4 a_342_199.n2 82.9225
R20 a_342_199.n1 a_342_199.n0 67.1884
R21 a_342_199.t0 a_342_199.n5 44.6333
R22 a_342_199.n5 a_342_199.t2 44.6333
R23 VPWR.n7 VPWR.n6 601.679
R24 VPWR.n15 VPWR.n14 585
R25 VPWR.n13 VPWR.n12 585
R26 VPWR.n8 VPWR.t2 258.447
R27 VPWR.n24 VPWR.t7 251.655
R28 VPWR.n22 VPWR.n2 241.339
R29 VPWR.n2 VPWR.t4 194.351
R30 VPWR.n14 VPWR.n13 104.656
R31 VPWR.n6 VPWR.t0 58.4849
R32 VPWR.n13 VPWR.t5 56.9458
R33 VPWR.n14 VPWR.t1 56.9458
R34 VPWR.n17 VPWR.n3 34.6358
R35 VPWR.n21 VPWR.n3 34.6358
R36 VPWR.n6 VPWR.t3 31.6057
R37 VPWR.n2 VPWR.t6 30.1648
R38 VPWR.n23 VPWR.n22 27.4829
R39 VPWR.n22 VPWR.n21 27.1064
R40 VPWR.n17 VPWR.n16 27.0813
R41 VPWR.n11 VPWR.n5 24.3832
R42 VPWR.n24 VPWR.n23 23.7181
R43 VPWR.n7 VPWR.n5 22.9652
R44 VPWR.n9 VPWR.n5 9.3005
R45 VPWR.n11 VPWR.n10 9.3005
R46 VPWR.n16 VPWR.n4 9.3005
R47 VPWR.n18 VPWR.n17 9.3005
R48 VPWR.n19 VPWR.n3 9.3005
R49 VPWR.n21 VPWR.n20 9.3005
R50 VPWR.n22 VPWR.n1 9.3005
R51 VPWR.n23 VPWR.n0 9.3005
R52 VPWR.n25 VPWR.n24 9.3005
R53 VPWR.n15 VPWR.n12 7.25383
R54 VPWR.n8 VPWR.n7 6.50073
R55 VPWR.n16 VPWR.n15 1.81383
R56 VPWR.n12 VPWR.n11 0.747167
R57 VPWR.n9 VPWR.n8 0.65346
R58 VPWR.n10 VPWR.n9 0.120292
R59 VPWR.n10 VPWR.n4 0.120292
R60 VPWR.n18 VPWR.n4 0.120292
R61 VPWR.n19 VPWR.n18 0.120292
R62 VPWR.n20 VPWR.n19 0.120292
R63 VPWR.n20 VPWR.n1 0.120292
R64 VPWR.n1 VPWR.n0 0.120292
R65 VPWR.n25 VPWR.n0 0.120292
R66 VPWR VPWR.n25 0.0213333
R67 VPB.t7 VPB.t4 541.59
R68 VPB.t0 VPB.t5 509.034
R69 VPB.t6 VPB.t0 325.546
R70 VPB.t1 VPB.t3 281.154
R71 VPB.t3 VPB.t2 272.274
R72 VPB.t8 VPB.t7 272.274
R73 VPB.t5 VPB.t1 260.437
R74 VPB.t4 VPB.t6 248.599
R75 VPB VPB.t8 189.409
R76 B.n0 B.t0 382.387
R77 B.n1 B.t3 261.178
R78 B.n1 B.t1 232.258
R79 B.n0 B.t2 218.507
R80 B B.n0 193.035
R81 B.n2 B.n1 152
R82 B.n2 B 7.76443
R83 B B.n2 6.50542
R84 a_766_47.t0 a_766_47.t1 60.0005
R85 VNB.t1 VNB.t7 2976.05
R86 VNB.t8 VNB.t4 2677.02
R87 VNB.t2 VNB.t5 1352.75
R88 VNB.t5 VNB.t3 1310.03
R89 VNB.t0 VNB.t8 1310.03
R90 VNB.t6 VNB.t1 1196.12
R91 VNB.t4 VNB.t6 1196.12
R92 VNB.t7 VNB.t2 1025.24
R93 VNB VNB.t0 911.327
R94 a_389_47.t0 a_389_47.n0 490.642
R95 a_389_47.n0 a_389_47.t2 38.5719
R96 a_389_47.n0 a_389_47.t1 38.5719
R97 VGND.n6 VGND.n5 204.457
R98 VGND.n13 VGND.n12 199.739
R99 VGND.n4 VGND.t3 163.379
R100 VGND.n18 VGND.t6 162.178
R101 VGND.n20 VGND.t0 156.495
R102 VGND.n5 VGND.t1 54.2862
R103 VGND.n12 VGND.t2 38.5719
R104 VGND.n12 VGND.t5 38.5719
R105 VGND.n7 VGND.n3 34.6358
R106 VGND.n11 VGND.n3 34.6358
R107 VGND.n14 VGND.n1 34.6358
R108 VGND.n19 VGND.n18 27.4829
R109 VGND.n18 VGND.n1 27.1064
R110 VGND.n5 VGND.t4 25.9346
R111 VGND.n13 VGND.n11 24.4711
R112 VGND.n20 VGND.n19 23.7181
R113 VGND.n7 VGND.n6 22.9652
R114 VGND.n14 VGND.n13 19.9534
R115 VGND.n21 VGND.n20 9.3005
R116 VGND.n8 VGND.n7 9.3005
R117 VGND.n9 VGND.n3 9.3005
R118 VGND.n11 VGND.n10 9.3005
R119 VGND.n13 VGND.n2 9.3005
R120 VGND.n15 VGND.n14 9.3005
R121 VGND.n16 VGND.n1 9.3005
R122 VGND.n18 VGND.n17 9.3005
R123 VGND.n19 VGND.n0 9.3005
R124 VGND.n6 VGND.n4 6.88265
R125 VGND.n8 VGND.n4 0.580811
R126 VGND.n9 VGND.n8 0.120292
R127 VGND.n10 VGND.n9 0.120292
R128 VGND.n10 VGND.n2 0.120292
R129 VGND.n15 VGND.n2 0.120292
R130 VGND.n16 VGND.n15 0.120292
R131 VGND.n17 VGND.n16 0.120292
R132 VGND.n17 VGND.n0 0.120292
R133 VGND.n21 VGND.n0 0.120292
R134 VGND VGND.n21 0.0213333
R135 COUT.n2 COUT 591.4
R136 COUT.n3 COUT.n2 585
R137 COUT.n0 COUT 185.97
R138 COUT.n1 COUT.n0 185
R139 COUT.n3 COUT.n1 64.4083
R140 COUT.n2 COUT.t2 34.4755
R141 COUT.n0 COUT.t0 32.3082
R142 COUT.n2 COUT.t3 26.5955
R143 COUT.n0 COUT.t1 24.9236
R144 COUT.n1 COUT 12.2187
R145 COUT COUT.n3 3.8405
R146 a_79_21.n3 a_79_21.n2 698.694
R147 a_79_21.n2 a_79_21.t0 260.188
R148 a_79_21.n1 a_79_21.t4 212.081
R149 a_79_21.n0 a_79_21.t5 212.081
R150 a_79_21.n2 a_79_21.n1 208.387
R151 a_79_21.n1 a_79_21.t3 139.78
R152 a_79_21.n0 a_79_21.t6 139.78
R153 a_79_21.n1 a_79_21.n0 67.1884
R154 a_79_21.n3 a_79_21.t2 41.5552
R155 a_79_21.t1 a_79_21.n3 41.5552
R156 a_468_369.t0 a_468_369.t1 123.126
R157 SUM SUM.n0 592.952
R158 SUM.n6 SUM.n0 585
R159 SUM.n5 SUM.n0 585
R160 SUM.n1 SUM 185.97
R161 SUM.n2 SUM.n1 185
R162 SUM.n0 SUM.t2 34.4755
R163 SUM.n1 SUM.t0 32.3082
R164 SUM.n0 SUM.t3 26.5955
R165 SUM.n1 SUM.t1 24.9236
R166 SUM SUM.n3 15.9294
R167 SUM.n2 SUM 12.2187
R168 SUM.n6 SUM 7.95202
R169 SUM.n4 SUM 6.82717
R170 SUM SUM.n6 5.23686
R171 SUM SUM.n5 5.23686
R172 SUM.n4 SUM 4.65505
R173 SUM.n3 SUM 3.41383
R174 SUM.n5 SUM.n4 3.29747
R175 SUM.n3 SUM 2.32777
R176 SUM SUM.n2 0.970197
C0 VPB A 0.13222f
C1 VPB VGND 0.014925f
C2 B A 0.354587f
C3 VPB VPWR 0.132502f
C4 B VGND 0.034776f
C5 B VPWR 0.037622f
C6 VPB SUM 0.005386f
C7 A VGND 0.048022f
C8 VPB COUT 0.004572f
C9 A VPWR 0.037216f
C10 VPWR VGND 0.134091f
C11 B COUT 4.25e-19
C12 SUM VGND 0.13278f
C13 A COUT 0.003281f
C14 VPWR SUM 0.19025f
C15 COUT VGND 0.106554f
C16 VPWR COUT 0.129675f
C17 VPB B 0.14275f
C18 VGND VNB 0.700869f
C19 COUT VNB 0.026521f
C20 SUM VNB 0.026013f
C21 VPWR VNB 0.587299f
C22 A VNB 0.263973f
C23 B VNB 0.245429f
C24 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ha_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ha_4 VNB VPB VGND VPWR COUT A B SUM
X0 a_467_47.t5 B.t0 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.095875 ps=0.945 w=0.65 l=0.15
X1 a_1325_47.t0 B.t1 a_514_199.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 COUT.t3 a_514_199.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X3 COUT.t2 a_514_199.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_467_47.t2 a_514_199.t8 a_79_21.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_717_297.t1 A.t0 VPWR.t15 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.1475 ps=1.295 w=1 l=0.15
X6 VPWR.t11 B.t2 a_514_199.t4 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t3 a_514_199.t9 COUT.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t9 a_79_21.t6 SUM.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t11 A.t1 a_1325_47.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_514_199.t5 A.t2 VPWR.t13 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.23 ps=1.46 w=1 l=0.15
X11 COUT.t6 a_514_199.t10 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_79_21.t0 a_514_199.t11 a_467_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VPWR.t1 a_514_199.t12 COUT.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 SUM.t2 a_79_21.t7 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t5 a_514_199.t13 a_79_21.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t1 A.t3 a_467_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t7 a_79_21.t8 SUM.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 COUT.t4 a_514_199.t14 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X19 VGND.t8 a_79_21.t9 SUM.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND.t9 a_79_21.t10 SUM.t6 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 SUM.t5 a_79_21.t11 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_79_21.t2 a_514_199.t15 VPWR.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3825 ps=1.765 w=1 l=0.15
X23 a_514_199.t2 B.t3 a_1167_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0715 ps=0.87 w=0.65 l=0.15
X24 VPWR.t14 A.t4 a_890_297.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.23 pd=1.46 as=0.2875 ps=1.575 w=1 l=0.15
X25 VPWR.t12 A.t5 a_514_199.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND.t6 B.t4 a_467_47.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VGND.t4 a_514_199.t16 COUT.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VGND.t5 a_514_199.t17 COUT.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_890_297.t0 B.t5 a_79_21.t5 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.2875 pd=1.575 as=0.135 ps=1.27 w=1 l=0.15
X30 a_514_199.t3 B.t6 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VGND.t0 A.t6 a_467_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X32 SUM.t0 a_79_21.t12 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_79_21.t4 B.t7 a_717_297.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1475 ps=1.295 w=1 l=0.15
X34 SUM.t4 a_79_21.t13 VGND.t12 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B B.n4 450.856
R1 B.n0 B.t6 212.081
R2 B.n1 B.t2 212.081
R3 B.n4 B.t5 212.081
R4 B.n3 B.t7 212.081
R5 B B.n2 155.061
R6 B.n0 B.t1 139.78
R7 B.n1 B.t3 139.78
R8 B.n4 B.t4 139.78
R9 B.n3 B.t0 139.78
R10 B.n4 B.n3 61.346
R11 B.n2 B.n0 46.7399
R12 B.n2 B.n1 14.6066
R13 VGND.n25 VGND.t6 282.817
R14 VGND.n19 VGND.t0 279.74
R15 VGND.n12 VGND.n11 209.381
R16 VGND.n9 VGND.n8 199.739
R17 VGND.n28 VGND.n27 198.702
R18 VGND.n10 VGND.t5 166.952
R19 VGND.n41 VGND.t12 160.014
R20 VGND.n34 VGND.t9 156.495
R21 VGND.n39 VGND.n1 120.698
R22 VGND.n18 VGND.n17 34.6358
R23 VGND.n20 VGND.n18 34.6358
R24 VGND.n24 VGND.n6 34.6358
R25 VGND.n28 VGND.n26 34.6358
R26 VGND.n32 VGND.n4 34.6358
R27 VGND.n33 VGND.n32 34.6358
R28 VGND.n38 VGND.n2 34.6358
R29 VGND.n34 VGND.n33 32.7534
R30 VGND.n8 VGND.t2 32.3082
R31 VGND.n8 VGND.t11 32.3082
R32 VGND.n13 VGND.n12 32.0005
R33 VGND.n40 VGND.n39 30.8711
R34 VGND.n17 VGND.n9 28.9887
R35 VGND.n27 VGND.t7 27.6928
R36 VGND.n27 VGND.t1 26.7697
R37 VGND.n41 VGND.n40 25.977
R38 VGND.n11 VGND.t3 24.9236
R39 VGND.n11 VGND.t4 24.9236
R40 VGND.n1 VGND.t10 24.9236
R41 VGND.n1 VGND.t8 24.9236
R42 VGND.n34 VGND.n2 18.4476
R43 VGND.n13 VGND.n9 15.4358
R44 VGND.n42 VGND.n41 9.3005
R45 VGND.n14 VGND.n13 9.3005
R46 VGND.n15 VGND.n9 9.3005
R47 VGND.n17 VGND.n16 9.3005
R48 VGND.n18 VGND.n7 9.3005
R49 VGND.n21 VGND.n20 9.3005
R50 VGND.n22 VGND.n6 9.3005
R51 VGND.n24 VGND.n23 9.3005
R52 VGND.n26 VGND.n5 9.3005
R53 VGND.n29 VGND.n28 9.3005
R54 VGND.n30 VGND.n4 9.3005
R55 VGND.n32 VGND.n31 9.3005
R56 VGND.n33 VGND.n3 9.3005
R57 VGND.n35 VGND.n34 9.3005
R58 VGND.n36 VGND.n2 9.3005
R59 VGND.n38 VGND.n37 9.3005
R60 VGND.n40 VGND.n0 9.3005
R61 VGND.n28 VGND.n4 7.90638
R62 VGND.n19 VGND.n6 7.15344
R63 VGND.n12 VGND.n10 6.53364
R64 VGND.n25 VGND.n24 6.02403
R65 VGND.n26 VGND.n25 3.76521
R66 VGND.n39 VGND.n38 3.76521
R67 VGND.n20 VGND.n19 2.63579
R68 VGND.n14 VGND.n10 0.626657
R69 VGND.n15 VGND.n14 0.120292
R70 VGND.n16 VGND.n15 0.120292
R71 VGND.n16 VGND.n7 0.120292
R72 VGND.n21 VGND.n7 0.120292
R73 VGND.n22 VGND.n21 0.120292
R74 VGND.n23 VGND.n22 0.120292
R75 VGND.n23 VGND.n5 0.120292
R76 VGND.n29 VGND.n5 0.120292
R77 VGND.n30 VGND.n29 0.120292
R78 VGND.n31 VGND.n30 0.120292
R79 VGND.n31 VGND.n3 0.120292
R80 VGND.n35 VGND.n3 0.120292
R81 VGND.n36 VGND.n35 0.120292
R82 VGND.n37 VGND.n36 0.120292
R83 VGND.n37 VGND.n0 0.120292
R84 VGND.n42 VGND.n0 0.120292
R85 VGND VGND.n42 0.0213333
R86 a_467_47.n1 a_467_47.t3 329.344
R87 a_467_47.n2 a_467_47.t0 288.726
R88 a_467_47.n3 a_467_47.n2 195.166
R89 a_467_47.n1 a_467_47.n0 185
R90 a_467_47.n2 a_467_47.n1 75.2946
R91 a_467_47.n0 a_467_47.t1 24.9236
R92 a_467_47.n0 a_467_47.t2 24.9236
R93 a_467_47.t4 a_467_47.n3 24.9236
R94 a_467_47.n3 a_467_47.t5 24.9236
R95 VNB.t8 VNB.t0 2748.22
R96 VNB.t13 VNB.t5 2677.02
R97 VNB.t0 VNB.t9 2249.84
R98 VNB.t15 VNB.t2 1423.95
R99 VNB.t1 VNB.t11 1267.31
R100 VNB.t3 VNB.t7 1196.12
R101 VNB.t6 VNB.t3 1196.12
R102 VNB.t2 VNB.t6 1196.12
R103 VNB.t10 VNB.t15 1196.12
R104 VNB.t9 VNB.t10 1196.12
R105 VNB.t11 VNB.t8 1196.12
R106 VNB.t4 VNB.t1 1196.12
R107 VNB.t5 VNB.t4 1196.12
R108 VNB.t14 VNB.t13 1196.12
R109 VNB.t12 VNB.t14 1196.12
R110 VNB.t16 VNB.t12 1196.12
R111 VNB VNB.t16 911.327
R112 a_514_199.n13 a_514_199.n9 597.424
R113 a_514_199.n15 a_514_199.n14 597.424
R114 a_514_199.n13 a_514_199.n12 411.012
R115 a_514_199.n8 a_514_199.n0 291.166
R116 a_514_199.n11 a_514_199.t15 215.732
R117 a_514_199.n10 a_514_199.t13 212.081
R118 a_514_199.n1 a_514_199.t9 212.081
R119 a_514_199.n2 a_514_199.t10 212.081
R120 a_514_199.n4 a_514_199.t12 212.081
R121 a_514_199.n5 a_514_199.t14 212.081
R122 a_514_199.n7 a_514_199.n3 177.601
R123 a_514_199.n7 a_514_199.n6 152
R124 a_514_199.n10 a_514_199.t8 143.433
R125 a_514_199.n11 a_514_199.t11 139.78
R126 a_514_199.n1 a_514_199.t17 139.78
R127 a_514_199.n2 a_514_199.t7 139.78
R128 a_514_199.n4 a_514_199.t16 139.78
R129 a_514_199.n5 a_514_199.t6 139.78
R130 a_514_199.n14 a_514_199.n8 87.3417
R131 a_514_199.n14 a_514_199.n13 63.2476
R132 a_514_199.n2 a_514_199.n1 61.346
R133 a_514_199.n12 a_514_199.n11 48.9308
R134 a_514_199.n3 a_514_199.n2 36.5157
R135 a_514_199.n6 a_514_199.n5 36.5157
R136 a_514_199.n8 a_514_199.n7 30.8711
R137 a_514_199.n9 a_514_199.t4 26.5955
R138 a_514_199.n9 a_514_199.t5 26.5955
R139 a_514_199.t0 a_514_199.n15 26.5955
R140 a_514_199.n15 a_514_199.t3 26.5955
R141 a_514_199.n0 a_514_199.t1 24.9236
R142 a_514_199.n0 a_514_199.t2 24.9236
R143 a_514_199.n4 a_514_199.n3 24.8308
R144 a_514_199.n6 a_514_199.n4 24.8308
R145 a_514_199.n12 a_514_199.n10 8.76414
R146 a_1325_47.t0 a_1325_47.t1 49.8467
R147 COUT.n1 COUT 590.715
R148 COUT.n2 COUT.n1 585
R149 COUT.n3 COUT.n0 366.325
R150 COUT.n7 COUT.n4 239.965
R151 COUT.n6 COUT.n5 185
R152 COUT.n1 COUT.t7 26.5955
R153 COUT.n1 COUT.t6 26.5955
R154 COUT.n0 COUT.t5 26.5955
R155 COUT.n0 COUT.t4 26.5955
R156 COUT.n5 COUT.t0 24.9236
R157 COUT.n5 COUT.t2 24.9236
R158 COUT.n4 COUT.t1 24.9236
R159 COUT.n4 COUT.t3 24.9236
R160 COUT COUT.n7 13.0291
R161 COUT.n3 COUT.n2 9.6005
R162 COUT COUT.n6 8.91479
R163 COUT.n6 COUT 6.62907
R164 COUT.n2 COUT 3.42907
R165 COUT COUT.n3 2.51479
R166 COUT.n7 COUT 2.51479
R167 a_79_21.n2 a_79_21.n1 703.966
R168 a_79_21.n2 a_79_21.n0 297.224
R169 a_79_21.n8 a_79_21.n7 220.766
R170 a_79_21.n6 a_79_21.t6 212.081
R171 a_79_21.n5 a_79_21.t7 212.081
R172 a_79_21.n4 a_79_21.t8 212.081
R173 a_79_21.n3 a_79_21.t12 212.081
R174 a_79_21.n7 a_79_21.n6 150.203
R175 a_79_21.n6 a_79_21.t10 139.78
R176 a_79_21.n5 a_79_21.t11 139.78
R177 a_79_21.n4 a_79_21.t9 139.78
R178 a_79_21.n3 a_79_21.t13 139.78
R179 a_79_21.n6 a_79_21.n5 61.346
R180 a_79_21.n5 a_79_21.n4 61.346
R181 a_79_21.n4 a_79_21.n3 61.346
R182 a_79_21.n7 a_79_21.n2 53.4593
R183 a_79_21.n0 a_79_21.t3 26.5955
R184 a_79_21.n0 a_79_21.t2 26.5955
R185 a_79_21.n1 a_79_21.t5 26.5955
R186 a_79_21.n1 a_79_21.t4 26.5955
R187 a_79_21.t1 a_79_21.n8 24.9236
R188 a_79_21.n8 a_79_21.t0 24.9236
R189 A.n4 A.n3 337.224
R190 A.n1 A.t4 267.291
R191 A.n5 A.t5 241.536
R192 A.n3 A.t0 241.536
R193 A.n2 A.t2 212.081
R194 A.n4 A.n2 177.976
R195 A.n5 A.t1 169.237
R196 A.n3 A.t3 169.237
R197 A.n6 A.n5 162.667
R198 A.n2 A.n0 147.083
R199 A.n1 A.t6 139.78
R200 A A.n4 73.5759
R201 A.n2 A.n1 54.0429
R202 A A.n6 6.67876
R203 A.n6 A 4.46111
R204 VPWR.n6 VPWR.n5 612.482
R205 VPWR.n25 VPWR.n10 601.679
R206 VPWR.n23 VPWR.n12 601.679
R207 VPWR.n14 VPWR.n13 601.679
R208 VPWR.n17 VPWR.n16 313.837
R209 VPWR.n15 VPWR.t3 262.841
R210 VPWR.n43 VPWR.t6 255.904
R211 VPWR.n41 VPWR.n1 229.373
R212 VPWR.n36 VPWR.n4 115.572
R213 VPWR.n4 VPWR.t4 90.6205
R214 VPWR.n4 VPWR.t9 60.0855
R215 VPWR.n10 VPWR.t13 45.3105
R216 VPWR.n10 VPWR.t14 45.3105
R217 VPWR.n40 VPWR.n2 34.6358
R218 VPWR.n29 VPWR.n8 34.6358
R219 VPWR.n30 VPWR.n29 34.6358
R220 VPWR.n31 VPWR.n30 34.6358
R221 VPWR.n35 VPWR.n34 34.6358
R222 VPWR.n13 VPWR.t0 34.4755
R223 VPWR.n13 VPWR.t12 34.4755
R224 VPWR.n24 VPWR.n23 32.0005
R225 VPWR.n5 VPWR.t15 31.5205
R226 VPWR.n42 VPWR.n41 30.8711
R227 VPWR.n25 VPWR.n8 30.8711
R228 VPWR.n22 VPWR.n14 28.9887
R229 VPWR.n1 VPWR.t8 26.5955
R230 VPWR.n1 VPWR.t7 26.5955
R231 VPWR.n5 VPWR.t5 26.5955
R232 VPWR.n12 VPWR.t10 26.5955
R233 VPWR.n12 VPWR.t11 26.5955
R234 VPWR.n16 VPWR.t2 26.5955
R235 VPWR.n16 VPWR.t1 26.5955
R236 VPWR.n43 VPWR.n42 25.977
R237 VPWR.n18 VPWR.n17 25.977
R238 VPWR.n34 VPWR.n6 21.4593
R239 VPWR.n36 VPWR.n2 18.4476
R240 VPWR.n18 VPWR.n14 15.4358
R241 VPWR.n25 VPWR.n24 13.5534
R242 VPWR.n31 VPWR.n6 13.177
R243 VPWR.n36 VPWR.n35 12.424
R244 VPWR.n23 VPWR.n22 12.424
R245 VPWR.n19 VPWR.n18 9.3005
R246 VPWR.n20 VPWR.n14 9.3005
R247 VPWR.n22 VPWR.n21 9.3005
R248 VPWR.n23 VPWR.n11 9.3005
R249 VPWR.n24 VPWR.n9 9.3005
R250 VPWR.n26 VPWR.n25 9.3005
R251 VPWR.n27 VPWR.n8 9.3005
R252 VPWR.n29 VPWR.n28 9.3005
R253 VPWR.n30 VPWR.n7 9.3005
R254 VPWR.n32 VPWR.n31 9.3005
R255 VPWR.n34 VPWR.n33 9.3005
R256 VPWR.n35 VPWR.n3 9.3005
R257 VPWR.n37 VPWR.n36 9.3005
R258 VPWR.n38 VPWR.n2 9.3005
R259 VPWR.n40 VPWR.n39 9.3005
R260 VPWR.n42 VPWR.n0 9.3005
R261 VPWR.n44 VPWR.n43 9.3005
R262 VPWR.n17 VPWR.n15 6.53364
R263 VPWR.n41 VPWR.n40 3.76521
R264 VPWR.n19 VPWR.n15 0.626657
R265 VPWR.n20 VPWR.n19 0.120292
R266 VPWR.n21 VPWR.n20 0.120292
R267 VPWR.n21 VPWR.n11 0.120292
R268 VPWR.n11 VPWR.n9 0.120292
R269 VPWR.n26 VPWR.n9 0.120292
R270 VPWR.n27 VPWR.n26 0.120292
R271 VPWR.n28 VPWR.n27 0.120292
R272 VPWR.n28 VPWR.n7 0.120292
R273 VPWR.n32 VPWR.n7 0.120292
R274 VPWR.n33 VPWR.n32 0.120292
R275 VPWR.n33 VPWR.n3 0.120292
R276 VPWR.n37 VPWR.n3 0.120292
R277 VPWR.n38 VPWR.n37 0.120292
R278 VPWR.n39 VPWR.n38 0.120292
R279 VPWR.n39 VPWR.n0 0.120292
R280 VPWR.n44 VPWR.n0 0.120292
R281 VPWR VPWR.n44 0.0213333
R282 a_717_297.t0 a_717_297.t1 58.1155
R283 VPB.t9 VPB.t0 541.59
R284 VPB.t12 VPB.t15 429.128
R285 VPB.t15 VPB.t16 361.06
R286 VPB.t14 VPB.t1 295.95
R287 VPB.t17 VPB.t10 263.397
R288 VPB.t2 VPB.t17 263.397
R289 VPB.t4 VPB.t5 248.599
R290 VPB.t3 VPB.t4 248.599
R291 VPB.t1 VPB.t3 248.599
R292 VPB.t11 VPB.t14 248.599
R293 VPB.t13 VPB.t11 248.599
R294 VPB.t16 VPB.t13 248.599
R295 VPB.t10 VPB.t12 248.599
R296 VPB.t0 VPB.t2 248.599
R297 VPB.t8 VPB.t9 248.599
R298 VPB.t7 VPB.t8 248.599
R299 VPB.t6 VPB.t7 248.599
R300 VPB VPB.t6 189.409
R301 SUM SUM.n0 592.952
R302 SUM.n8 SUM.n0 585
R303 SUM.n7 SUM.n0 585
R304 SUM.n3 SUM.n1 220.571
R305 SUM.n4 SUM 185.97
R306 SUM.n5 SUM.n4 185
R307 SUM.n3 SUM.n2 114.736
R308 SUM.n6 SUM.n3 28.682
R309 SUM.n0 SUM.t1 26.5955
R310 SUM.n0 SUM.t0 26.5955
R311 SUM.n1 SUM.t3 26.5955
R312 SUM.n1 SUM.t2 26.5955
R313 SUM.n4 SUM.t7 24.9236
R314 SUM.n4 SUM.t4 24.9236
R315 SUM.n2 SUM.t6 24.9236
R316 SUM.n2 SUM.t5 24.9236
R317 SUM.n5 SUM 12.2187
R318 SUM SUM.n6 9.50353
R319 SUM.n8 SUM 7.95202
R320 SUM.n7 SUM 7.95202
R321 SUM SUM.n8 5.23686
R322 SUM SUM.n7 5.23686
R323 SUM.n6 SUM 3.68535
R324 SUM SUM.n5 0.970197
R325 a_890_297.t0 a_890_297.t1 113.275
C0 VPB B 0.126111f
C1 VPB VPWR 0.190961f
C2 A B 0.486152f
C3 A VPWR 0.081667f
C4 VPB SUM 0.010208f
C5 VPB COUT 0.007933f
C6 B VPWR 0.048697f
C7 A COUT 6.28e-19
C8 VPB VGND 0.013885f
C9 A VGND 0.064168f
C10 VPWR SUM 0.409225f
C11 VPWR COUT 0.303208f
C12 B VGND 0.116322f
C13 VPWR VGND 0.208698f
C14 SUM VGND 0.294788f
C15 COUT VGND 0.207901f
C16 VPB A 0.141726f
C17 VGND VNB 1.06298f
C18 COUT VNB 0.032236f
C19 SUM VNB 0.032255f
C20 VPWR VNB 0.903239f
C21 B VNB 0.389723f
C22 A VNB 0.381077f
C23 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
X0 VPWR.t11 A.t0 Y.t17 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t16 A.t1 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t15 A.t2 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t8 A.t3 Y.t14 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.515 pd=3.03 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t23 A.t4 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y.t3 A.t5 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t7 A.t6 Y.t13 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t6 A.t7 Y.t12 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y.t2 A.t8 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t1 A.t9 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t11 A.t10 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t7 A.t11 Y.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.33475 pd=2.33 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t6 A.t12 Y.t7 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t10 A.t13 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Y.t6 A.t14 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR.t3 A.t15 Y.t9 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y.t5 A.t16 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y.t8 A.t17 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR.t1 A.t18 Y.t22 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND.t3 A.t19 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND.t2 A.t20 Y.t20 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t1 A.t21 Y.t19 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t21 A.t22 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND.t0 A.t23 Y.t18 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n2 A.t3 212.081
R1 A.n1 A.t2 212.081
R2 A.n6 A.t7 212.081
R3 A.n28 A.t10 212.081
R4 A.n26 A.t15 212.081
R5 A.n7 A.t17 212.081
R6 A.n22 A.t18 212.081
R7 A.n8 A.t22 212.081
R8 A.n17 A.t0 212.081
R9 A.n9 A.t1 212.081
R10 A.n12 A.t6 212.081
R11 A.n10 A.t13 212.081
R12 A.n11 A 163.264
R13 A A.n3 154.048
R14 A.n5 A.n4 152
R15 A A.n29 152
R16 A.n27 A.n0 152
R17 A.n25 A 152
R18 A.n24 A.n23 152
R19 A.n21 A.n20 152
R20 A.n19 A.n18 152
R21 A.n16 A.n15 152
R22 A.n14 A.n13 152
R23 A.n2 A.t11 139.78
R24 A.n1 A.t9 139.78
R25 A.n6 A.t12 139.78
R26 A.n28 A.t8 139.78
R27 A.n26 A.t23 139.78
R28 A.n7 A.t5 139.78
R29 A.n22 A.t21 139.78
R30 A.n8 A.t4 139.78
R31 A.n17 A.t20 139.78
R32 A.n9 A.t16 139.78
R33 A.n12 A.t19 139.78
R34 A.n10 A.t14 139.78
R35 A.n3 A.n2 30.6732
R36 A.n3 A.n1 30.6732
R37 A.n5 A.n1 30.6732
R38 A.n6 A.n5 30.6732
R39 A.n29 A.n6 30.6732
R40 A.n29 A.n28 30.6732
R41 A.n28 A.n27 30.6732
R42 A.n27 A.n26 30.6732
R43 A.n26 A.n25 30.6732
R44 A.n25 A.n7 30.6732
R45 A.n23 A.n7 30.6732
R46 A.n23 A.n22 30.6732
R47 A.n22 A.n21 30.6732
R48 A.n21 A.n8 30.6732
R49 A.n18 A.n8 30.6732
R50 A.n18 A.n17 30.6732
R51 A.n17 A.n16 30.6732
R52 A.n16 A.n9 30.6732
R53 A.n13 A.n9 30.6732
R54 A.n13 A.n12 30.6732
R55 A.n12 A.n11 30.6732
R56 A.n11 A.n10 30.6732
R57 A A.n0 21.5045
R58 A A.n24 21.5045
R59 A.n4 A 19.4565
R60 A.n20 A 19.4565
R61 A A.n19 17.4085
R62 A.n15 A 15.3605
R63 A A.n14 13.3125
R64 A.n14 A 10.2405
R65 A.n15 A 8.1925
R66 A.n19 A 6.1445
R67 A.n20 A 4.0965
R68 A.n4 A 2.0485
R69 A A.n0 2.0485
R70 A.n24 A 2.0485
R71 Y.n1 Y.n0 205.28
R72 Y.n3 Y.n2 205.28
R73 Y.n5 Y.n4 205.28
R74 Y.n7 Y.n6 205.28
R75 Y.n9 Y.n8 205.28
R76 Y.n11 Y.n10 205.28
R77 Y.n13 Y.n12 99.1759
R78 Y.n15 Y.n14 99.1759
R79 Y.n17 Y.n16 99.1759
R80 Y.n19 Y.n18 99.1759
R81 Y.n21 Y.n20 99.1759
R82 Y.n23 Y.n22 99.1759
R83 Y Y.n11 42.5955
R84 Y.n3 Y.n1 38.4005
R85 Y.n5 Y.n3 38.4005
R86 Y.n7 Y.n5 38.4005
R87 Y.n9 Y.n7 38.4005
R88 Y.n11 Y.n9 38.4005
R89 Y.n15 Y.n13 34.3584
R90 Y.n17 Y.n15 34.3584
R91 Y.n19 Y.n17 34.3584
R92 Y.n21 Y.n19 34.3584
R93 Y.n23 Y.n21 34.3584
R94 Y.n13 Y 33.3575
R95 Y Y.n1 27.1064
R96 Y.n0 Y.t13 26.5955
R97 Y.n0 Y.t10 26.5955
R98 Y.n2 Y.t17 26.5955
R99 Y.n2 Y.t16 26.5955
R100 Y.n4 Y.t22 26.5955
R101 Y.n4 Y.t21 26.5955
R102 Y.n6 Y.t9 26.5955
R103 Y.n6 Y.t8 26.5955
R104 Y.n8 Y.t12 26.5955
R105 Y.n8 Y.t11 26.5955
R106 Y.n10 Y.t14 26.5955
R107 Y.n10 Y.t15 26.5955
R108 Y.n12 Y.t0 24.9236
R109 Y.n12 Y.t1 24.9236
R110 Y.n14 Y.t7 24.9236
R111 Y.n14 Y.t2 24.9236
R112 Y.n16 Y.t18 24.9236
R113 Y.n16 Y.t3 24.9236
R114 Y.n18 Y.t19 24.9236
R115 Y.n18 Y.t23 24.9236
R116 Y.n20 Y.t20 24.9236
R117 Y.n20 Y.t5 24.9236
R118 Y.n22 Y.t4 24.9236
R119 Y.n22 Y.t6 24.9236
R120 Y Y.n23 20.3378
R121 VPWR.n12 VPWR.t8 393.505
R122 VPWR.n29 VPWR.t4 342.375
R123 VPWR.n2 VPWR.n1 320.976
R124 VPWR.n22 VPWR.n4 320.976
R125 VPWR.n6 VPWR.n5 320.976
R126 VPWR.n16 VPWR.n8 320.976
R127 VPWR.n11 VPWR.n10 320.976
R128 VPWR.n15 VPWR.n9 34.6358
R129 VPWR.n18 VPWR.n17 34.6358
R130 VPWR.n24 VPWR.n23 34.6358
R131 VPWR.n28 VPWR.n27 34.6358
R132 VPWR.n22 VPWR.n21 32.0005
R133 VPWR.n21 VPWR.n6 31.2476
R134 VPWR.n1 VPWR.t10 26.5955
R135 VPWR.n1 VPWR.t7 26.5955
R136 VPWR.n4 VPWR.t0 26.5955
R137 VPWR.n4 VPWR.t11 26.5955
R138 VPWR.n5 VPWR.t2 26.5955
R139 VPWR.n5 VPWR.t1 26.5955
R140 VPWR.n8 VPWR.t5 26.5955
R141 VPWR.n8 VPWR.t3 26.5955
R142 VPWR.n10 VPWR.t9 26.5955
R143 VPWR.n10 VPWR.t6 26.5955
R144 VPWR.n24 VPWR.n2 25.977
R145 VPWR.n17 VPWR.n16 25.224
R146 VPWR.n12 VPWR.n11 22.6104
R147 VPWR.n11 VPWR.n9 19.2005
R148 VPWR.n29 VPWR.n28 13.5534
R149 VPWR.n30 VPWR.n29 11.1829
R150 VPWR.n16 VPWR.n15 9.41227
R151 VPWR.n13 VPWR.n9 9.3005
R152 VPWR.n15 VPWR.n14 9.3005
R153 VPWR.n17 VPWR.n7 9.3005
R154 VPWR.n19 VPWR.n18 9.3005
R155 VPWR.n21 VPWR.n20 9.3005
R156 VPWR.n23 VPWR.n3 9.3005
R157 VPWR.n25 VPWR.n24 9.3005
R158 VPWR.n27 VPWR.n26 9.3005
R159 VPWR.n28 VPWR.n0 9.3005
R160 VPWR.n27 VPWR.n2 8.65932
R161 VPWR.n18 VPWR.n6 3.38874
R162 VPWR.n23 VPWR.n22 2.63579
R163 VPWR.n13 VPWR.n12 0.554787
R164 VPWR.n14 VPWR.n13 0.120292
R165 VPWR.n14 VPWR.n7 0.120292
R166 VPWR.n19 VPWR.n7 0.120292
R167 VPWR.n20 VPWR.n19 0.120292
R168 VPWR.n20 VPWR.n3 0.120292
R169 VPWR.n25 VPWR.n3 0.120292
R170 VPWR.n26 VPWR.n25 0.120292
R171 VPWR.n26 VPWR.n0 0.120292
R172 VPWR.n30 VPWR.n0 0.120292
R173 VPWR VPWR.n30 0.0226354
R174 VPB VPB.t4 290.031
R175 VPB.t9 VPB.t8 248.599
R176 VPB.t6 VPB.t9 248.599
R177 VPB.t5 VPB.t6 248.599
R178 VPB.t3 VPB.t5 248.599
R179 VPB.t2 VPB.t3 248.599
R180 VPB.t1 VPB.t2 248.599
R181 VPB.t0 VPB.t1 248.599
R182 VPB.t11 VPB.t0 248.599
R183 VPB.t10 VPB.t11 248.599
R184 VPB.t7 VPB.t10 248.599
R185 VPB.t4 VPB.t7 248.599
R186 VGND.n29 VGND.t5 287.151
R187 VGND.n12 VGND.t7 278.007
R188 VGND.n11 VGND.n10 207.213
R189 VGND.n16 VGND.n8 207.213
R190 VGND.n6 VGND.n5 207.213
R191 VGND.n22 VGND.n4 207.213
R192 VGND.n2 VGND.n1 207.213
R193 VGND.n15 VGND.n9 34.6358
R194 VGND.n18 VGND.n17 34.6358
R195 VGND.n24 VGND.n23 34.6358
R196 VGND.n28 VGND.n27 34.6358
R197 VGND.n22 VGND.n21 32.0005
R198 VGND.n21 VGND.n6 31.2476
R199 VGND.n24 VGND.n2 25.977
R200 VGND.n17 VGND.n16 25.224
R201 VGND.n10 VGND.t8 24.9236
R202 VGND.n10 VGND.t6 24.9236
R203 VGND.n8 VGND.t9 24.9236
R204 VGND.n8 VGND.t0 24.9236
R205 VGND.n5 VGND.t10 24.9236
R206 VGND.n5 VGND.t1 24.9236
R207 VGND.n4 VGND.t11 24.9236
R208 VGND.n4 VGND.t2 24.9236
R209 VGND.n1 VGND.t4 24.9236
R210 VGND.n1 VGND.t3 24.9236
R211 VGND.n12 VGND.n11 22.6104
R212 VGND.n11 VGND.n9 19.2005
R213 VGND.n29 VGND.n28 13.5534
R214 VGND.n30 VGND.n29 11.1829
R215 VGND.n16 VGND.n15 9.41227
R216 VGND.n13 VGND.n9 9.3005
R217 VGND.n15 VGND.n14 9.3005
R218 VGND.n17 VGND.n7 9.3005
R219 VGND.n19 VGND.n18 9.3005
R220 VGND.n21 VGND.n20 9.3005
R221 VGND.n23 VGND.n3 9.3005
R222 VGND.n25 VGND.n24 9.3005
R223 VGND.n27 VGND.n26 9.3005
R224 VGND.n28 VGND.n0 9.3005
R225 VGND.n27 VGND.n2 8.65932
R226 VGND.n18 VGND.n6 3.38874
R227 VGND.n23 VGND.n22 2.63579
R228 VGND.n13 VGND.n12 0.554787
R229 VGND.n14 VGND.n13 0.120292
R230 VGND.n14 VGND.n7 0.120292
R231 VGND.n19 VGND.n7 0.120292
R232 VGND.n20 VGND.n19 0.120292
R233 VGND.n20 VGND.n3 0.120292
R234 VGND.n25 VGND.n3 0.120292
R235 VGND.n26 VGND.n25 0.120292
R236 VGND.n26 VGND.n0 0.120292
R237 VGND.n30 VGND.n0 0.120292
R238 VGND VGND.n30 0.0226354
R239 VNB VNB.t5 1395.47
R240 VNB.t8 VNB.t7 1196.12
R241 VNB.t6 VNB.t8 1196.12
R242 VNB.t9 VNB.t6 1196.12
R243 VNB.t0 VNB.t9 1196.12
R244 VNB.t10 VNB.t0 1196.12
R245 VNB.t1 VNB.t10 1196.12
R246 VNB.t11 VNB.t1 1196.12
R247 VNB.t2 VNB.t11 1196.12
R248 VNB.t4 VNB.t2 1196.12
R249 VNB.t3 VNB.t4 1196.12
R250 VNB.t5 VNB.t3 1196.12
C0 VPB A 0.383471f
C1 VPB VPWR 0.130635f
C2 A VPWR 0.181754f
C3 VPB Y 0.040341f
C4 VPB VGND 0.009331f
C5 A Y 1.26141f
C6 A VGND 0.167395f
C7 VPWR Y 1.14598f
C8 VPWR VGND 0.124118f
C9 Y VGND 0.843368f
C10 VGND VNB 0.694591f
C11 Y VNB 0.132809f
C12 VPWR VNB 0.605858f
C13 A VNB 1.13688f
C14 VPB VNB 1.22494f
.ends


* NGSPICE file created from sky130_fd_sc_hd__inv_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
X0 VPWR.t5 A.t0 Y.t8 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 Y.t7 A.t1 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t3 A.t2 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t3 A.t3 Y.t6 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t5 A.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t1 A.t5 Y.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t2 A.t6 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X7 Y.t0 A.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t1 A.t8 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X9 VGND.t2 A.t9 Y.t10 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t1 A.t10 Y.t9 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t0 A.t11 Y.t11 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n0 A.t0 212.081
R1 A.n2 A.t1 212.081
R2 A.n9 A.t3 212.081
R3 A.n3 A.t4 212.081
R4 A.n4 A.t5 212.081
R5 A.n5 A.t8 212.081
R6 A.n6 A.n5 206.042
R7 A A.n1 154.304
R8 A.n11 A.n10 152
R9 A.n8 A.n7 152
R10 A.n0 A.t11 139.78
R11 A.n2 A.t2 139.78
R12 A.n9 A.t10 139.78
R13 A.n3 A.t7 139.78
R14 A.n4 A.t9 139.78
R15 A.n5 A.t6 139.78
R16 A A.n6 62.2085
R17 A.n4 A.n3 61.346
R18 A.n5 A.n4 61.346
R19 A.n1 A.n0 42.3581
R20 A.n10 A.n2 42.3581
R21 A.n9 A.n8 42.3581
R22 A A.n11 19.2005
R23 A.n2 A.n1 18.9884
R24 A.n10 A.n9 18.9884
R25 A.n8 A.n3 18.9884
R26 A.n7 A 17.1525
R27 A.n7 A 6.4005
R28 A.n6 A 6.4005
R29 A.n11 A 4.3525
R30 Y.n3 Y.n2 267.699
R31 Y.n8 Y.n6 243.68
R32 Y.n3 Y.n1 207.965
R33 Y.n4 Y.n0 207.965
R34 Y.n8 Y.n7 205.28
R35 Y.n9 Y.n5 204.893
R36 Y.n4 Y.n3 59.7338
R37 Y.n9 Y.n8 38.7884
R38 Y.n5 Y.t8 26.5955
R39 Y.n5 Y.t7 26.5955
R40 Y.n6 Y.t4 26.5955
R41 Y.n6 Y.t1 26.5955
R42 Y.n7 Y.t6 26.5955
R43 Y.n7 Y.t5 26.5955
R44 Y.n2 Y.t10 24.9236
R45 Y.n2 Y.t2 24.9236
R46 Y.n1 Y.t9 24.9236
R47 Y.n1 Y.t0 24.9236
R48 Y.n0 Y.t11 24.9236
R49 Y.n0 Y.t3 24.9236
R50 Y.n10 Y.n4 18.1338
R51 Y Y.n9 11.3665
R52 Y.n10 Y 10.6062
R53 Y Y.n10 1.82907
R54 VPWR.n5 VPWR.t5 873.6
R55 VPWR.n2 VPWR.n1 320.976
R56 VPWR.n6 VPWR.n4 320.976
R57 VPWR.n13 VPWR.t0 279.582
R58 VPWR.n6 VPWR.n5 37.1366
R59 VPWR.n8 VPWR.n7 34.6358
R60 VPWR.n12 VPWR.n11 34.6358
R61 VPWR.n1 VPWR.t2 26.5955
R62 VPWR.n1 VPWR.t1 26.5955
R63 VPWR.n4 VPWR.t4 26.5955
R64 VPWR.n4 VPWR.t3 26.5955
R65 VPWR.n8 VPWR.n2 25.6005
R66 VPWR.n13 VPWR.n12 19.9534
R67 VPWR.n7 VPWR.n3 9.3005
R68 VPWR.n9 VPWR.n8 9.3005
R69 VPWR.n11 VPWR.n10 9.3005
R70 VPWR.n12 VPWR.n0 9.3005
R71 VPWR.n14 VPWR.n13 9.3005
R72 VPWR.n11 VPWR.n2 9.03579
R73 VPWR.n7 VPWR.n6 3.01226
R74 VPWR.n5 VPWR.n3 2.28766
R75 VPWR.n9 VPWR.n3 0.120292
R76 VPWR.n10 VPWR.n9 0.120292
R77 VPWR.n10 VPWR.n0 0.120292
R78 VPWR.n14 VPWR.n0 0.120292
R79 VPWR VPWR.n14 0.0226354
R80 VPB VPB.t0 292.991
R81 VPB.t4 VPB.t5 248.599
R82 VPB.t3 VPB.t4 248.599
R83 VPB.t2 VPB.t3 248.599
R84 VPB.t1 VPB.t2 248.599
R85 VPB.t0 VPB.t1 248.599
R86 VGND.n5 VGND.t0 287.26
R87 VGND.n13 VGND.t4 250.433
R88 VGND.n6 VGND.n4 207.213
R89 VGND.n2 VGND.n1 207.213
R90 VGND.n6 VGND.n5 36.3334
R91 VGND.n8 VGND.n7 34.6358
R92 VGND.n12 VGND.n11 34.6358
R93 VGND.n8 VGND.n2 25.6005
R94 VGND.n4 VGND.t5 24.9236
R95 VGND.n4 VGND.t1 24.9236
R96 VGND.n1 VGND.t3 24.9236
R97 VGND.n1 VGND.t2 24.9236
R98 VGND.n13 VGND.n12 22.2123
R99 VGND.n14 VGND.n13 9.3005
R100 VGND.n7 VGND.n3 9.3005
R101 VGND.n9 VGND.n8 9.3005
R102 VGND.n11 VGND.n10 9.3005
R103 VGND.n12 VGND.n0 9.3005
R104 VGND.n11 VGND.n2 9.03579
R105 VGND.n7 VGND.n6 3.01226
R106 VGND.n5 VGND.n3 2.43104
R107 VGND.n9 VGND.n3 0.120292
R108 VGND.n10 VGND.n9 0.120292
R109 VGND.n10 VGND.n0 0.120292
R110 VGND.n14 VGND.n0 0.120292
R111 VGND VGND.n14 0.0226354
R112 VNB VNB.t4 1409.71
R113 VNB.t5 VNB.t0 1196.12
R114 VNB.t1 VNB.t5 1196.12
R115 VNB.t3 VNB.t1 1196.12
R116 VNB.t2 VNB.t3 1196.12
R117 VNB.t4 VNB.t2 1196.12
C0 Y VPB 0.018383f
C1 VGND VPB 0.00676f
C2 Y A 0.543559f
C3 VGND A 0.1215f
C4 Y VPWR 0.530316f
C5 VGND VPWR 0.069534f
C6 Y VGND 0.325869f
C7 VPB A 0.212612f
C8 VPB VPWR 0.078318f
C9 A VPWR 0.136084f
C10 VGND VNB 0.421424f
C11 Y VNB 0.09005f
C12 VPWR VNB 0.373245f
C13 A VNB 0.646336f
C14 VPB VNB 0.69336f
.ends


* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_4 KAPWR VGND VPWR A X VPB VNB
X0 KAPWR.t4 A.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND.t3 a_27_47.t2 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND.t2 a_27_47.t3 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X.t7 a_27_47.t4 KAPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X.t0 a_27_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND.t4 A.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 KAPWR.t2 a_27_47.t6 X.t6 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X.t3 a_27_47.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X.t5 a_27_47.t8 KAPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 KAPWR.t0 a_27_47.t9 X.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n0 A.t0 238.59
R1 A.n0 A.t1 203.244
R2 A A.n0 154.012
R3 a_27_47.t1 a_27_47.n9 418.024
R4 a_27_47.n9 a_27_47.t0 304.587
R5 a_27_47.n6 a_27_47.t8 223.19
R6 a_27_47.n3 a_27_47.t6 221.72
R7 a_27_47.n0 a_27_47.t4 221.72
R8 a_27_47.n1 a_27_47.t9 221.72
R9 a_27_47.n3 a_27_47.t2 185.38
R10 a_27_47.n6 a_27_47.t7 184.768
R11 a_27_47.n1 a_27_47.t3 184.768
R12 a_27_47.n0 a_27_47.t5 184.768
R13 a_27_47.n4 a_27_47.n2 177.601
R14 a_27_47.n8 a_27_47.n7 152
R15 a_27_47.n5 a_27_47.n2 152
R16 a_27_47.n9 a_27_47.n8 85.4593
R17 a_27_47.n4 a_27_47.n3 56.9641
R18 a_27_47.n7 a_27_47.n6 49.0769
R19 a_27_47.n5 a_27_47.n0 41.1896
R20 a_27_47.n1 a_27_47.n5 33.3023
R21 a_27_47.n7 a_27_47.n1 26.2914
R22 a_27_47.n8 a_27_47.n2 25.6005
R23 a_27_47.n0 a_27_47.n4 18.4041
R24 KAPWR.n1 KAPWR.n0 597.986
R25 KAPWR.n1 KAPWR.t2 333.687
R26 KAPWR.n3 KAPWR.n2 305.096
R27 KAPWR.n2 KAPWR.t1 37.4305
R28 KAPWR.n2 KAPWR.t4 27.5805
R29 KAPWR.n0 KAPWR.t3 27.5805
R30 KAPWR.n0 KAPWR.t0 27.5805
R31 KAPWR.n3 KAPWR.n1 0.511798
R32 KAPWR KAPWR.n3 0.304587
R33 VPB.t4 VPB.t1 284.113
R34 VPB.t3 VPB.t2 254.518
R35 VPB.t0 VPB.t3 254.518
R36 VPB.t1 VPB.t0 254.518
R37 VPB VPB.t4 195.327
R38 X.n5 X.n3 693.095
R39 X.n2 X.n0 243.627
R40 X.n2 X.n1 200.262
R41 X.n5 X.n4 196.75
R42 X.n0 X.t1 40.0005
R43 X.n0 X.t3 40.0005
R44 X.n1 X.t2 40.0005
R45 X.n1 X.t0 40.0005
R46 X.n3 X.t4 27.5805
R47 X.n3 X.t5 27.5805
R48 X.n4 X.t6 27.5805
R49 X.n4 X.t7 27.5805
R50 X X.n6 19.2609
R51 X.n6 X.n5 13.438
R52 X.n7 X 9.00791
R53 X.n7 X.n2 6.77697
R54 X.n6 X 2.70819
R55 X X.n7 1.73877
R56 VGND.n1 VGND.t3 249.87
R57 VGND.n3 VGND.n2 205.078
R58 VGND.n6 VGND.n5 203.619
R59 VGND.n5 VGND.t0 55.7148
R60 VGND.n2 VGND.t1 40.0005
R61 VGND.n2 VGND.t2 40.0005
R62 VGND.n5 VGND.t4 40.0005
R63 VGND.n4 VGND.n3 24.4711
R64 VGND.n6 VGND.n4 24.0946
R65 VGND.n4 VGND.n0 9.3005
R66 VGND.n7 VGND.n6 7.27268
R67 VGND.n3 VGND.n1 6.71867
R68 VGND.n1 VGND.n0 0.647964
R69 VGND.n7 VGND.n0 0.146586
R70 VGND VGND.n7 0.116801
R71 VNB.t4 VNB.t0 1381.23
R72 VNB.t1 VNB.t3 1224.6
R73 VNB.t2 VNB.t1 1224.6
R74 VNB.t0 VNB.t2 1224.6
R75 VNB VNB.t4 939.807
C0 A VGND 0.042728f
C1 KAPWR X 0.300268f
C2 VPB VPWR 0.048961f
C3 X VGND 0.215037f
C4 A VPWR 0.007982f
C5 KAPWR VGND 0.059713f
C6 X VPWR 0.065438f
C7 KAPWR VPWR 0.396927f
C8 VGND VPWR 0.004316f
C9 VPB A 0.032139f
C10 VPB X 0.012134f
C11 VPB KAPWR 0.012371f
C12 A X 0.014114f
C13 VPB VGND 0.005641f
C14 A KAPWR 0.015089f
C15 VPWR VNB 0.278787f
C16 VGND VNB 0.357713f
C17 X VNB 0.06701f
C18 KAPWR VNB 0.041612f
C19 A VNB 0.147639f
C20 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_2 KAPWR VGND VPWR A X VPB VNB
X0 KAPWR.t2 A.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 KAPWR.t0 a_27_47.t2 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t2 A.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X.t0 a_27_47.t3 KAPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X.t3 a_27_47.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND.t0 a_27_47.t5 X.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 A.n0 A.t0 239.293
R1 A.n0 A.t1 171.06
R2 A A.n0 162.667
R3 a_27_47.t0 a_27_47.n3 407.61
R4 a_27_47.n3 a_27_47.t1 299.271
R5 a_27_47.n3 a_27_47.n2 215.082
R6 a_27_47.n0 a_27_47.t3 189.588
R7 a_27_47.n0 a_27_47.t2 189.588
R8 a_27_47.n1 a_27_47.t5 96.4005
R9 a_27_47.n1 a_27_47.t4 96.4005
R10 a_27_47.n2 a_27_47.n1 35.0935
R11 a_27_47.n2 a_27_47.n0 19.8724
R12 KAPWR.n1 KAPWR.t0 832.371
R13 KAPWR.n1 KAPWR.n0 305.086
R14 KAPWR.n0 KAPWR.t1 36.4455
R15 KAPWR.n0 KAPWR.t2 27.5805
R16 KAPWR KAPWR.n1 0.320212
R17 VPB.t2 VPB.t0 281.154
R18 VPB.t0 VPB.t1 248.599
R19 VPB VPB.t2 195.327
R20 X X.n0 635.053
R21 X X.n1 216.464
R22 X.n1 X.t2 38.5719
R23 X.n1 X.t3 38.5719
R24 X.n0 X.t1 26.5955
R25 X.n0 X.t0 26.5955
R26 VGND.n1 VGND.t0 245.523
R27 VGND.n1 VGND.n0 209.065
R28 VGND.n0 VGND.t1 52.8576
R29 VGND.n0 VGND.t2 40.0005
R30 VGND VGND.n1 0.549826
R31 VNB.t2 VNB.t1 1352.75
R32 VNB.t1 VNB.t0 1196.12
R33 VNB VNB.t2 939.807
C0 X VGND 0.114239f
C1 VPB VPWR 0.035289f
C2 VPB A 0.033009f
C3 A VPWR 0.008179f
C4 VPB KAPWR 0.007899f
C5 KAPWR VPWR 0.262453f
C6 A KAPWR 0.015316f
C7 VPB X 0.008051f
C8 X VPWR 0.024311f
C9 A X 0.01266f
C10 VPB VGND 0.004059f
C11 VGND VPWR 0.004216f
C12 KAPWR X 0.141577f
C13 A VGND 0.045054f
C14 KAPWR VGND 0.038723f
C15 VPWR VNB 0.203241f
C16 VGND VNB 0.262949f
C17 X VNB 0.070513f
C18 KAPWR VNB 0.031011f
C19 A VNB 0.147594f
C20 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_1 KAPWR VGND VPWR X A VPB VNB
X0 KAPWR.t0 a_75_212.t2 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212.t0 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212.t1 A.t1 KAPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND.t0 a_75_212.t3 X.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
R0 a_75_212.t1 a_75_212.n1 407.228
R1 a_75_212.n1 a_75_212.t0 294.341
R2 a_75_212.n0 a_75_212.t2 254.389
R3 a_75_212.n0 a_75_212.t3 211.01
R4 a_75_212.n1 a_75_212.n0 152
R5 X.n1 X.t0 368.521
R6 X.n0 X.t1 216.155
R7 X X.n0 82.2255
R8 X.n1 X 10.5563
R9 X X.n1 5.48477
R10 X.n0 X 5.16973
R11 KAPWR KAPWR.n0 305.26
R12 KAPWR.n0 KAPWR.t1 36.1587
R13 KAPWR.n0 KAPWR.t0 36.1587
R14 VPB.t1 VPB.t0 260.437
R15 VPB VPB.t1 91.745
R16 A.n0 A.t1 260.322
R17 A.n0 A.t0 175.169
R18 A A.n0 154.133
R19 VGND VGND.n0 205.657
R20 VGND.n0 VGND.t1 33.462
R21 VGND.n0 VGND.t0 33.462
R22 VNB.t1 VNB.t0 1253.07
R23 VNB VNB.t1 441.425
C0 VPB VGND 0.004897f
C1 KAPWR VPWR 0.1756f
C2 A KAPWR 0.013437f
C3 X KAPWR 0.075741f
C4 VPB A 0.052491f
C5 A VGND 0.018157f
C6 VPB VPWR 0.029804f
C7 VGND VPWR 0.005062f
C8 VPB X 0.012788f
C9 X VGND 0.05405f
C10 A VPWR 0.009537f
C11 X VPWR 0.028088f
C12 A X 8.48e-19
C13 KAPWR VGND 0.027221f
C14 VPB KAPWR 0.0055f
C15 VPWR VNB 0.16597f
C16 VGND VNB 0.20733f
C17 KAPWR VNB 0.020391f
C18 X VNB 0.094159f
C19 A VNB 0.164205f
C20 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_bleeder_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_bleeder_1 VPB VNB SHORT VPWR VGND
X0 a_147_105.t0 SHORT.t0 VGND.t0 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0378 pd=0.57 as=0.0936 ps=1.24 w=0.36 l=0.15
X1 VPWR.t0 SHORT.t1 a_363_105.t0 VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.0936 pd=1.24 as=0.0378 ps=0.57 w=0.36 l=0.15
X2 a_363_105.t1 SHORT.t2 a_291_105.t0 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0378 pd=0.57 as=0.0378 ps=0.57 w=0.36 l=0.15
X3 a_291_105.t1 SHORT.t3 a_219_105.t0 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0378 pd=0.57 as=0.0378 ps=0.57 w=0.36 l=0.15
X4 a_219_105.t1 SHORT.t4 a_147_105.t1 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0378 pd=0.57 as=0.0378 ps=0.57 w=0.36 l=0.15
R0 SHORT.n4 SHORT.n0 152
R1 SHORT.n7 SHORT.n6 152
R2 SHORT.n1 SHORT.t1 145.768
R3 SHORT.n6 SHORT.t0 101.951
R4 SHORT.n1 SHORT.t2 93.1872
R5 SHORT.n5 SHORT.t4 93.1872
R6 SHORT.n3 SHORT.t3 93.1872
R7 SHORT.n2 SHORT.n0 73.1551
R8 SHORT.n4 SHORT.n3 46.7399
R9 SHORT.n6 SHORT.n5 43.8187
R10 SHORT.n3 SHORT.n2 23.8919
R11 SHORT.n2 SHORT.n1 21.8408
R12 SHORT.n7 SHORT.n0 6.30775
R13 SHORT.n5 SHORT.n4 5.84292
R14 SHORT SHORT.n7 5.28746
R15 VGND VGND.t0 264.077
R16 a_147_105.t0 a_147_105.t1 70.0005
R17 VNB VNB.t4 1466.67
R18 VNB.t2 VNB.t3 1025.24
R19 VNB.t1 VNB.t2 1025.24
R20 VNB.t0 VNB.t1 1025.24
R21 VNB.t4 VNB.t0 1025.24
R22 a_363_105.t0 a_363_105.t1 70.0005
R23 VPWR VPWR.t0 315.344
R24 a_291_105.t0 a_291_105.t1 70.0005
R25 a_219_105.t0 a_219_105.t1 70.0005
C0 SHORT VGND 0.112785f
C1 VPB VPWR 0.145185f
C2 SHORT VPWR 0.143549f
C3 VGND VPWR 0.087376f
C4 VPB SHORT 0.133175f
C5 VPB VGND 0.018244f
C6 VPWR VNB 0.398527f
C7 VGND VNB 0.415639f
C8 SHORT VNB 0.386092f
C9 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_8 X A VPB VNB KAPWR VGND VPWR
X0 KAPWR.t1 A.t0 a_110_47.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 KAPWR.t2 a_110_47.t4 X.t15 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X.t14 a_110_47.t5 KAPWR.t9 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47.t2 A.t1 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X.t5 a_110_47.t6 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X.t13 a_110_47.t7 KAPWR.t8 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND.t8 a_110_47.t8 X.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 KAPWR.t7 a_110_47.t9 X.t12 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND.t1 A.t2 a_110_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND.t7 a_110_47.t10 X.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47.t0 A.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 KAPWR.t6 a_110_47.t11 X.t11 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X.t10 a_110_47.t12 KAPWR.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND.t6 a_110_47.t13 X.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND.t5 a_110_47.t14 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X.t9 a_110_47.t15 KAPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X.t0 a_110_47.t16 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 KAPWR.t3 a_110_47.t17 X.t8 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X.t7 a_110_47.t18 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X.t6 a_110_47.t19 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A.n0 A.t0 184.768
R1 A.n1 A.t1 184.768
R2 A A.n1 173.609
R3 A.n0 A.t2 146.208
R4 A.n1 A.t3 146.208
R5 A.n1 A.n0 40.6397
R6 a_110_47.n21 a_110_47.n20 316.591
R7 a_110_47.n20 a_110_47.n0 217.256
R8 a_110_47.n3 a_110_47.t17 212.081
R9 a_110_47.n4 a_110_47.t12 212.081
R10 a_110_47.n5 a_110_47.t9 212.081
R11 a_110_47.n7 a_110_47.t5 212.081
R12 a_110_47.n8 a_110_47.t4 212.081
R13 a_110_47.n14 a_110_47.t15 212.081
R14 a_110_47.n16 a_110_47.t11 212.081
R15 a_110_47.n17 a_110_47.t7 212.081
R16 a_110_47.n10 a_110_47.n6 169.409
R17 a_110_47.n3 a_110_47.t10 162.274
R18 a_110_47.n4 a_110_47.t16 162.274
R19 a_110_47.n5 a_110_47.t13 162.274
R20 a_110_47.n7 a_110_47.t18 162.274
R21 a_110_47.n8 a_110_47.t14 162.274
R22 a_110_47.n14 a_110_47.t19 162.274
R23 a_110_47.n16 a_110_47.t8 162.274
R24 a_110_47.n17 a_110_47.t6 162.274
R25 a_110_47.n19 a_110_47.n18 152
R26 a_110_47.n15 a_110_47.n1 152
R27 a_110_47.n13 a_110_47.n12 152
R28 a_110_47.n11 a_110_47.n2 152
R29 a_110_47.n10 a_110_47.n9 152
R30 a_110_47.n4 a_110_47.n3 55.2698
R31 a_110_47.n5 a_110_47.n4 55.2698
R32 a_110_47.n13 a_110_47.n2 43.7018
R33 a_110_47.n20 a_110_47.n19 43.5205
R34 a_110_47.n0 a_110_47.t1 40.0005
R35 a_110_47.n0 a_110_47.t0 40.0005
R36 a_110_47.n15 a_110_47.n14 39.8458
R37 a_110_47.n9 a_110_47.n8 35.9898
R38 a_110_47.n6 a_110_47.n5 30.8485
R39 a_110_47.n18 a_110_47.n16 28.2778
R40 a_110_47.n21 a_110_47.t3 27.5805
R41 a_110_47.t2 a_110_47.n21 27.5805
R42 a_110_47.n18 a_110_47.n17 26.9925
R43 a_110_47.n7 a_110_47.n6 24.4218
R44 a_110_47.n9 a_110_47.n7 19.2805
R45 a_110_47.n11 a_110_47.n10 17.4085
R46 a_110_47.n12 a_110_47.n11 17.4085
R47 a_110_47.n12 a_110_47.n1 17.4085
R48 a_110_47.n19 a_110_47.n1 17.4085
R49 a_110_47.n16 a_110_47.n15 15.4245
R50 a_110_47.n8 a_110_47.n2 7.7125
R51 a_110_47.n14 a_110_47.n13 3.8565
R52 KAPWR.n1 KAPWR.t3 769.928
R53 KAPWR.n5 KAPWR.n4 594.793
R54 KAPWR.n1 KAPWR.n0 594.793
R55 KAPWR.n3 KAPWR.n2 594.644
R56 KAPWR.n8 KAPWR.t0 337.877
R57 KAPWR.n7 KAPWR.n6 311.43
R58 KAPWR.n6 KAPWR.t8 27.5805
R59 KAPWR.n6 KAPWR.t1 27.5805
R60 KAPWR.n4 KAPWR.t4 27.5805
R61 KAPWR.n4 KAPWR.t6 27.5805
R62 KAPWR.n2 KAPWR.t9 27.5805
R63 KAPWR.n2 KAPWR.t2 27.5805
R64 KAPWR.n0 KAPWR.t5 27.5805
R65 KAPWR.n0 KAPWR.t7 27.5805
R66 KAPWR.n3 KAPWR.n1 0.508673
R67 KAPWR.n8 KAPWR.n7 0.496173
R68 KAPWR.n7 KAPWR.n5 0.493048
R69 KAPWR.n5 KAPWR.n3 0.489923
R70 KAPWR KAPWR.n8 0.0557885
R71 VPB.t4 VPB.t2 254.518
R72 VPB.t6 VPB.t4 254.518
R73 VPB.t8 VPB.t6 254.518
R74 VPB.t9 VPB.t8 254.518
R75 VPB.t3 VPB.t9 254.518
R76 VPB.t5 VPB.t3 254.518
R77 VPB.t7 VPB.t5 254.518
R78 VPB.t1 VPB.t7 254.518
R79 VPB.t0 VPB.t1 254.518
R80 VPB VPB.t0 195.327
R81 X.n7 X.n5 333.392
R82 X.n7 X.n6 301.392
R83 X.n9 X.n8 301.392
R84 X.n11 X.n10 298.296
R85 X.n2 X.n0 248.638
R86 X.n2 X.n1 203.463
R87 X.n4 X.n3 203.463
R88 X X.n13 199.673
R89 X.n4 X.n2 45.177
R90 X.n0 X.t4 40.0005
R91 X.n0 X.t5 40.0005
R92 X.n1 X.t1 40.0005
R93 X.n1 X.t6 40.0005
R94 X.n3 X.t2 40.0005
R95 X.n3 X.t7 40.0005
R96 X.n13 X.t3 40.0005
R97 X.n13 X.t0 40.0005
R98 X.n9 X.n7 32.0005
R99 X.n5 X.t11 27.5805
R100 X.n5 X.t13 27.5805
R101 X.n6 X.t15 27.5805
R102 X.n6 X.t9 27.5805
R103 X.n8 X.t12 27.5805
R104 X.n8 X.t14 27.5805
R105 X.n10 X.t8 27.5805
R106 X.n10 X.t10 27.5805
R107 X.n12 X.n4 27.1064
R108 X.n11 X.n9 19.2005
R109 X.n12 X 3.76132
R110 X X.n11 2.2438
R111 X X.n12 0.726273
R112 VGND.n7 VGND.t7 249.72
R113 VGND.n21 VGND.t0 244.853
R114 VGND.n19 VGND.n2 206.909
R115 VGND.n6 VGND.n5 204.692
R116 VGND.n12 VGND.n11 204.692
R117 VGND.n15 VGND.n14 204.692
R118 VGND.n5 VGND.t4 40.0005
R119 VGND.n5 VGND.t6 40.0005
R120 VGND.n11 VGND.t3 40.0005
R121 VGND.n11 VGND.t5 40.0005
R122 VGND.n14 VGND.t2 40.0005
R123 VGND.n14 VGND.t8 40.0005
R124 VGND.n2 VGND.t9 40.0005
R125 VGND.n2 VGND.t1 40.0005
R126 VGND.n10 VGND.n4 34.6358
R127 VGND.n15 VGND.n13 31.624
R128 VGND.n19 VGND.n1 27.1064
R129 VGND.n20 VGND.n19 22.5887
R130 VGND.n21 VGND.n20 22.5887
R131 VGND.n15 VGND.n1 18.0711
R132 VGND.n13 VGND.n12 13.5534
R133 VGND.n7 VGND.n6 12.6486
R134 VGND.n22 VGND.n21 9.3005
R135 VGND.n8 VGND.n4 9.3005
R136 VGND.n10 VGND.n9 9.3005
R137 VGND.n13 VGND.n3 9.3005
R138 VGND.n16 VGND.n15 9.3005
R139 VGND.n17 VGND.n1 9.3005
R140 VGND.n19 VGND.n18 9.3005
R141 VGND.n20 VGND.n0 9.3005
R142 VGND.n6 VGND.n4 9.03579
R143 VGND.n12 VGND.n10 1.50638
R144 VGND.n8 VGND.n7 1.08558
R145 VGND.n9 VGND.n8 0.120292
R146 VGND.n9 VGND.n3 0.120292
R147 VGND.n16 VGND.n3 0.120292
R148 VGND.n17 VGND.n16 0.120292
R149 VGND.n18 VGND.n17 0.120292
R150 VGND.n18 VGND.n0 0.120292
R151 VGND.n22 VGND.n0 0.120292
R152 VGND VGND.n22 0.0226354
R153 VNB.t4 VNB.t7 1224.6
R154 VNB.t6 VNB.t4 1224.6
R155 VNB.t3 VNB.t6 1224.6
R156 VNB.t5 VNB.t3 1224.6
R157 VNB.t2 VNB.t5 1224.6
R158 VNB.t8 VNB.t2 1224.6
R159 VNB.t9 VNB.t8 1224.6
R160 VNB.t1 VNB.t9 1224.6
R161 VNB.t0 VNB.t1 1224.6
R162 VNB VNB.t0 939.807
C0 A KAPWR 0.061797f
C1 VPB X 0.022318f
C2 VPB VGND 0.008825f
C3 A X 0.001679f
C4 KAPWR X 0.660006f
C5 A VGND 0.068858f
C6 VPB VPWR 0.083959f
C7 KAPWR VGND 0.111499f
C8 A VPWR 0.020216f
C9 KAPWR VPWR 0.727511f
C10 X VGND 0.490553f
C11 X VPWR 0.135811f
C12 VGND VPWR 0.008217f
C13 VPB A 0.070741f
C14 VPB KAPWR 0.029773f
C15 VPWR VNB 0.478152f
C16 VGND VNB 0.607928f
C17 X VNB 0.081251f
C18 KAPWR VNB 0.063346f
C19 A VNB 0.28981f
C20 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_16 VNB VPB KAPWR VGND VPWR A X
X0 KAPWR.t15 A.t0 a_110_47.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 KAPWR.t11 a_110_47.t8 X.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X.t10 a_110_47.t9 KAPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X.t9 a_110_47.t10 KAPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_47.t6 A.t1 KAPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 a_110_47.t3 A.t2 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 X.t12 a_110_47.t11 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 a_110_47.t5 A.t3 KAPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND.t14 A.t4 a_110_47.t2 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND.t10 a_110_47.t12 X.t23 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 KAPWR.t8 a_110_47.t13 X.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 X.t7 a_110_47.t14 KAPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND.t13 A.t5 a_110_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 KAPWR.t6 a_110_47.t15 X.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X14 VGND.t9 a_110_47.t16 X.t22 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X.t5 a_110_47.t17 KAPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X16 a_110_47.t0 A.t6 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X17 KAPWR.t12 A.t7 a_110_47.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 X.t4 a_110_47.t18 KAPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND.t8 a_110_47.t19 X.t21 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 VGND.t7 a_110_47.t20 X.t20 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 X.t19 a_110_47.t21 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 X.t3 a_110_47.t22 KAPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 X.t2 a_110_47.t23 KAPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 X.t18 a_110_47.t24 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X25 KAPWR.t1 a_110_47.t25 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 X.t0 a_110_47.t26 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 X.t17 a_110_47.t27 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 X.t16 a_110_47.t28 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X.t15 a_110_47.t29 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X.t14 a_110_47.t30 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X31 X.t13 a_110_47.t31 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
R0 A.n0 A.t7 184.768
R1 A.n1 A.t3 184.768
R2 A.n2 A.t0 184.768
R3 A.n3 A.t1 184.768
R4 A A.n3 173.609
R5 A.n0 A.t4 146.208
R6 A.n1 A.t2 146.208
R7 A.n2 A.t5 146.208
R8 A.n3 A.t6 146.208
R9 A.n1 A.n0 40.6397
R10 A.n2 A.n1 40.6397
R11 A.n3 A.n2 40.6397
R12 a_110_47.n57 a_110_47.n56 227.583
R13 a_110_47.n58 a_110_47.n2 226.815
R14 a_110_47.n57 a_110_47.n55 220.84
R15 a_110_47.n2 a_110_47.n3 217.256
R16 a_110_47.n19 a_110_47.n17 212.081
R17 a_110_47.n20 a_110_47.t26 212.081
R18 a_110_47.n21 a_110_47.n15 212.081
R19 a_110_47.n23 a_110_47.t14 212.081
R20 a_110_47.n25 a_110_47.n13 212.081
R21 a_110_47.n1 a_110_47.t22 212.081
R22 a_110_47.n30 a_110_47.n10 212.081
R23 a_110_47.n8 a_110_47.t17 212.081
R24 a_110_47.n35 a_110_47.t15 212.081
R25 a_110_47.n0 a_110_47.t10 212.081
R26 a_110_47.n40 a_110_47.t25 212.081
R27 a_110_47.n42 a_110_47.t18 212.081
R28 a_110_47.n43 a_110_47.t13 212.081
R29 a_110_47.n49 a_110_47.t9 212.081
R30 a_110_47.n51 a_110_47.t8 212.081
R31 a_110_47.n52 a_110_47.t23 212.081
R32 a_110_47.n22 a_110_47.n12 169.409
R33 a_110_47.n19 a_110_47.n18 162.274
R34 a_110_47.n20 a_110_47.t21 162.274
R35 a_110_47.n21 a_110_47.n16 162.274
R36 a_110_47.n23 a_110_47.t27 162.274
R37 a_110_47.n25 a_110_47.n14 162.274
R38 a_110_47.n1 a_110_47.t29 162.274
R39 a_110_47.n30 a_110_47.n11 162.274
R40 a_110_47.n8 a_110_47.t31 162.274
R41 a_110_47.n35 a_110_47.t12 162.274
R42 a_110_47.n0 a_110_47.t11 162.274
R43 a_110_47.n40 a_110_47.t16 162.274
R44 a_110_47.n42 a_110_47.t24 162.274
R45 a_110_47.n43 a_110_47.t19 162.274
R46 a_110_47.n49 a_110_47.t28 162.274
R47 a_110_47.n51 a_110_47.t20 162.274
R48 a_110_47.n52 a_110_47.t30 162.274
R49 a_110_47.n54 a_110_47.n53 152
R50 a_110_47.n50 a_110_47.n4 152
R51 a_110_47.n48 a_110_47.n47 152
R52 a_110_47.n46 a_110_47.n5 152
R53 a_110_47.n45 a_110_47.n44 152
R54 a_110_47.n41 a_110_47.n6 152
R55 a_110_47.n39 a_110_47.n38 152
R56 a_110_47.n37 a_110_47.n0 152
R57 a_110_47.n36 a_110_47.n7 152
R58 a_110_47.n34 a_110_47.n33 152
R59 a_110_47.n32 a_110_47.n31 152
R60 a_110_47.n29 a_110_47.n9 152
R61 a_110_47.n1 a_110_47.n28 152
R62 a_110_47.n27 a_110_47.n26 152
R63 a_110_47.n24 a_110_47.n12 152
R64 a_110_47.n20 a_110_47.n19 55.2698
R65 a_110_47.n21 a_110_47.n20 55.2698
R66 a_110_47.n26 a_110_47.n1 43.7018
R67 a_110_47.n29 a_110_47.n1 43.7018
R68 a_110_47.n0 a_110_47.n36 43.7018
R69 a_110_47.n48 a_110_47.n5 43.7018
R70 a_110_47.n39 a_110_47.n0 43.7018
R71 a_110_47.n2 a_110_47.n54 43.5205
R72 a_110_47.n2 a_110_47.n57 43.5205
R73 a_110_47.n55 a_110_47.t1 40.0005
R74 a_110_47.n55 a_110_47.t0 40.0005
R75 a_110_47.n3 a_110_47.t2 40.0005
R76 a_110_47.n3 a_110_47.t3 40.0005
R77 a_110_47.n50 a_110_47.n49 39.8458
R78 a_110_47.n44 a_110_47.n43 35.9898
R79 a_110_47.n22 a_110_47.n21 35.3472
R80 a_110_47.n35 a_110_47.n34 33.4192
R81 a_110_47.n31 a_110_47.n30 32.7765
R82 a_110_47.n25 a_110_47.n24 31.4912
R83 a_110_47.n41 a_110_47.n40 30.8485
R84 a_110_47.n53 a_110_47.n51 28.2778
R85 a_110_47.n56 a_110_47.t7 27.5805
R86 a_110_47.n56 a_110_47.t6 27.5805
R87 a_110_47.t4 a_110_47.n58 27.5805
R88 a_110_47.n58 a_110_47.t5 27.5805
R89 a_110_47.n53 a_110_47.n52 26.9925
R90 a_110_47.n42 a_110_47.n41 24.4218
R91 a_110_47.n24 a_110_47.n23 23.7792
R92 a_110_47.n31 a_110_47.n8 22.4938
R93 a_110_47.n34 a_110_47.n8 21.2085
R94 a_110_47.n23 a_110_47.n22 19.9232
R95 a_110_47.n44 a_110_47.n42 19.2805
R96 a_110_47.n27 a_110_47.n12 17.4085
R97 a_110_47.n28 a_110_47.n27 17.4085
R98 a_110_47.n28 a_110_47.n9 17.4085
R99 a_110_47.n32 a_110_47.n9 17.4085
R100 a_110_47.n33 a_110_47.n32 17.4085
R101 a_110_47.n33 a_110_47.n7 17.4085
R102 a_110_47.n37 a_110_47.n7 17.4085
R103 a_110_47.n38 a_110_47.n37 17.4085
R104 a_110_47.n38 a_110_47.n6 17.4085
R105 a_110_47.n45 a_110_47.n6 17.4085
R106 a_110_47.n46 a_110_47.n45 17.4085
R107 a_110_47.n47 a_110_47.n46 17.4085
R108 a_110_47.n47 a_110_47.n4 17.4085
R109 a_110_47.n54 a_110_47.n4 17.4085
R110 a_110_47.n51 a_110_47.n50 15.4245
R111 a_110_47.n40 a_110_47.n39 12.8538
R112 a_110_47.n26 a_110_47.n25 12.2112
R113 a_110_47.n30 a_110_47.n29 10.9258
R114 a_110_47.n36 a_110_47.n35 10.2832
R115 a_110_47.n43 a_110_47.n5 7.7125
R116 a_110_47.n49 a_110_47.n48 3.8565
R117 KAPWR.n0 KAPWR.t0 760.357
R118 KAPWR.n1 KAPWR.t3 760.163
R119 KAPWR.n0 KAPWR.t7 760.163
R120 KAPWR.n3 KAPWR.n2 594.822
R121 KAPWR.n7 KAPWR.n6 594.793
R122 KAPWR.n5 KAPWR.n4 594.793
R123 KAPWR.n9 KAPWR.n8 594.644
R124 KAPWR.n14 KAPWR.t14 237.472
R125 KAPWR.n13 KAPWR.n12 209.893
R126 KAPWR.n11 KAPWR.n10 209.893
R127 KAPWR.n12 KAPWR.t13 27.5805
R128 KAPWR.n12 KAPWR.t15 27.5805
R129 KAPWR.n10 KAPWR.t2 27.5805
R130 KAPWR.n10 KAPWR.t12 27.5805
R131 KAPWR.n8 KAPWR.t10 27.5805
R132 KAPWR.n8 KAPWR.t11 27.5805
R133 KAPWR.n6 KAPWR.t4 27.5805
R134 KAPWR.n6 KAPWR.t8 27.5805
R135 KAPWR.n4 KAPWR.t9 27.5805
R136 KAPWR.n4 KAPWR.t1 27.5805
R137 KAPWR.n2 KAPWR.t6 27.5805
R138 KAPWR.n2 KAPWR.t5 26.5955
R139 KAPWR.n9 KAPWR.n7 0.508673
R140 KAPWR.n3 KAPWR.n1 0.496173
R141 KAPWR.n7 KAPWR.n5 0.496173
R142 KAPWR.n14 KAPWR.n13 0.496173
R143 KAPWR.n1 KAPWR.n0 0.493048
R144 KAPWR.n5 KAPWR.n3 0.493048
R145 KAPWR.n13 KAPWR.n11 0.493048
R146 KAPWR.n11 KAPWR.n9 0.489923
R147 KAPWR KAPWR.n14 0.0581923
R148 VPB.t7 VPB.t0 509.034
R149 VPB.t3 VPB.t7 509.034
R150 VPB.t5 VPB.t3 509.034
R151 VPB.t9 VPB.t6 254.518
R152 VPB.t1 VPB.t9 254.518
R153 VPB.t4 VPB.t1 254.518
R154 VPB.t8 VPB.t4 254.518
R155 VPB.t10 VPB.t8 254.518
R156 VPB.t11 VPB.t10 254.518
R157 VPB.t2 VPB.t11 254.518
R158 VPB.t12 VPB.t2 254.518
R159 VPB.t13 VPB.t12 254.518
R160 VPB.t15 VPB.t13 254.518
R161 VPB.t14 VPB.t15 254.518
R162 VPB.t6 VPB.t5 251.559
R163 VPB VPB.t14 145.017
R164 X.n17 X.t5 414.159
R165 X.n18 X.t3 414.159
R166 X.n19 X.t7 414.159
R167 X.n20 X.t0 411.271
R168 X.n12 X.n10 338.599
R169 X.n12 X.n11 302.327
R170 X.n14 X.n13 302.327
R171 X.n16 X.n15 302.327
R172 X.n2 X.n0 248.638
R173 X.n7 X.t13 243.463
R174 X.n8 X.t15 243.463
R175 X.n9 X.t17 243.463
R176 X X.t19 239.607
R177 X.n2 X.n1 203.463
R178 X.n4 X.n3 203.463
R179 X.n6 X.n5 202.456
R180 X.n4 X.n2 45.177
R181 X.n8 X.n7 45.177
R182 X.n9 X.n8 45.177
R183 X.n6 X.n4 44.0476
R184 X.n7 X.n6 44.0476
R185 X.n0 X.t20 40.0005
R186 X.n0 X.t14 40.0005
R187 X.n1 X.t21 40.0005
R188 X.n1 X.t16 40.0005
R189 X.n3 X.t22 40.0005
R190 X.n3 X.t18 40.0005
R191 X.n5 X.t23 40.0005
R192 X.n5 X.t12 40.0005
R193 X.n14 X.n12 32.0005
R194 X.n16 X.n14 32.0005
R195 X.n18 X.n17 32.0005
R196 X.n19 X.n18 32.0005
R197 X.n17 X.n16 31.2005
R198 X.n10 X.t11 27.5805
R199 X.n10 X.t2 27.5805
R200 X.n11 X.t8 27.5805
R201 X.n11 X.t10 27.5805
R202 X.n13 X.t1 27.5805
R203 X.n13 X.t4 27.5805
R204 X.n15 X.t6 27.5805
R205 X.n15 X.t9 27.5805
R206 X.n21 X.n9 13.177
R207 X.n20 X.n19 10.4484
R208 X.n21 X 3.13183
R209 X X.n20 1.75844
R210 X X.n21 0.604792
R211 VGND.n10 VGND.t6 250.282
R212 VGND.n9 VGND.t4 245.481
R213 VGND.n13 VGND.t2 245.481
R214 VGND.n39 VGND.t12 240.948
R215 VGND.n33 VGND.n32 206.909
R216 VGND.n37 VGND.n2 206.909
R217 VGND.n7 VGND.n6 205.899
R218 VGND.n20 VGND.n19 205.899
R219 VGND.n23 VGND.n22 204.692
R220 VGND.n30 VGND.n29 204.692
R221 VGND.n6 VGND.t10 40.0005
R222 VGND.n19 VGND.t11 40.0005
R223 VGND.n19 VGND.t9 40.0005
R224 VGND.n22 VGND.t5 40.0005
R225 VGND.n22 VGND.t8 40.0005
R226 VGND.n29 VGND.t3 40.0005
R227 VGND.n29 VGND.t7 40.0005
R228 VGND.n32 VGND.t1 40.0005
R229 VGND.n32 VGND.t14 40.0005
R230 VGND.n2 VGND.t15 40.0005
R231 VGND.n2 VGND.t13 40.0005
R232 VGND.n6 VGND.t0 38.5719
R233 VGND.n18 VGND.n7 34.6358
R234 VGND.n24 VGND.n21 34.6358
R235 VGND.n28 VGND.n4 34.6358
R236 VGND.n33 VGND.n31 31.624
R237 VGND.n14 VGND.n13 29.7417
R238 VGND.n37 VGND.n1 27.1064
R239 VGND.n12 VGND.n9 25.224
R240 VGND.n38 VGND.n37 22.5887
R241 VGND.n39 VGND.n38 22.5887
R242 VGND.n13 VGND.n12 20.7064
R243 VGND.n33 VGND.n1 18.0711
R244 VGND.n14 VGND.n7 16.1887
R245 VGND.n31 VGND.n30 13.5534
R246 VGND.n20 VGND.n18 11.6711
R247 VGND.n40 VGND.n39 9.3005
R248 VGND.n12 VGND.n11 9.3005
R249 VGND.n13 VGND.n8 9.3005
R250 VGND.n15 VGND.n14 9.3005
R251 VGND.n16 VGND.n7 9.3005
R252 VGND.n18 VGND.n17 9.3005
R253 VGND.n21 VGND.n5 9.3005
R254 VGND.n25 VGND.n24 9.3005
R255 VGND.n26 VGND.n4 9.3005
R256 VGND.n28 VGND.n27 9.3005
R257 VGND.n31 VGND.n3 9.3005
R258 VGND.n34 VGND.n33 9.3005
R259 VGND.n35 VGND.n1 9.3005
R260 VGND.n37 VGND.n36 9.3005
R261 VGND.n38 VGND.n0 9.3005
R262 VGND.n23 VGND.n4 9.03579
R263 VGND.n10 VGND.n9 6.78128
R264 VGND.n24 VGND.n23 6.02403
R265 VGND.n21 VGND.n20 4.51815
R266 VGND.n30 VGND.n28 1.50638
R267 VGND.n11 VGND.n10 0.56336
R268 VGND.n11 VGND.n8 0.120292
R269 VGND.n15 VGND.n8 0.120292
R270 VGND.n16 VGND.n15 0.120292
R271 VGND.n17 VGND.n16 0.120292
R272 VGND.n17 VGND.n5 0.120292
R273 VGND.n25 VGND.n5 0.120292
R274 VGND.n26 VGND.n25 0.120292
R275 VGND.n27 VGND.n26 0.120292
R276 VGND.n27 VGND.n3 0.120292
R277 VGND.n34 VGND.n3 0.120292
R278 VGND.n35 VGND.n34 0.120292
R279 VGND.n36 VGND.n35 0.120292
R280 VGND.n36 VGND.n0 0.120292
R281 VGND.n40 VGND.n0 0.120292
R282 VGND VGND.n40 0.0226354
R283 VNB.t4 VNB.t6 2449.19
R284 VNB.t2 VNB.t4 2449.19
R285 VNB.t0 VNB.t2 2449.19
R286 VNB.t11 VNB.t10 1224.6
R287 VNB.t9 VNB.t11 1224.6
R288 VNB.t5 VNB.t9 1224.6
R289 VNB.t8 VNB.t5 1224.6
R290 VNB.t3 VNB.t8 1224.6
R291 VNB.t7 VNB.t3 1224.6
R292 VNB.t1 VNB.t7 1224.6
R293 VNB.t14 VNB.t1 1224.6
R294 VNB.t15 VNB.t14 1224.6
R295 VNB.t13 VNB.t15 1224.6
R296 VNB.t12 VNB.t13 1224.6
R297 VNB.t10 VNB.t0 1210.36
R298 VNB VNB.t12 697.736
C0 A VGND 0.113883f
C1 KAPWR X 1.27396f
C2 VPB VPWR 0.141271f
C3 A VPWR 0.03533f
C4 KAPWR VGND 0.20578f
C5 KAPWR VPWR 1.34584f
C6 X VGND 0.973835f
C7 X VPWR 0.277309f
C8 VGND VPWR 0.00674f
C9 VPB A 0.133144f
C10 VPB KAPWR 0.034148f
C11 VPB X 0.031597f
C12 A KAPWR 0.106184f
C13 A X 0.001281f
C14 VPB VGND 0.011113f
C15 VPWR VNB 0.818117f
C16 VGND VNB 1.01459f
C17 X VNB 0.110579f
C18 KAPWR VNB 0.057392f
C19 A VNB 0.494797f
C20 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_1 VPB VNB KAPWR VGND VPWR A Y
X0 Y.t1 A.t0 KAPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2184 ps=2.2 w=0.84 l=0.15
X1 VGND.t0 A.t1 Y.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 KAPWR.t1 A.t2 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=2.24 as=0.1134 ps=1.11 w=0.84 l=0.15
R0 A A.n1 283.014
R1 A.n0 A.t2 231.907
R2 A.n1 A.t0 231.361
R3 A.n0 A.t1 170.308
R4 A.n1 A.n0 54.0627
R5 KAPWR.n0 KAPWR.t0 403.139
R6 KAPWR.n0 KAPWR.t1 396.5
R7 KAPWR KAPWR.n0 0.0605962
R8 Y Y.n0 345.13
R9 Y.n1 Y.t2 240.419
R10 Y.n0 Y.t0 31.6612
R11 Y.n0 Y.t1 31.6612
R12 Y Y.n1 6.19224
R13 Y.n1 Y 0.0242128
R14 VPB.t1 VPB.t0 248.599
R15 VPB VPB.t1 192.369
R16 VGND VGND.t0 250.06
R17 VNB VNB.t0 2107.44
C0 VGND VPB 0.005703f
C1 VPWR Y 0.022275f
C2 VGND A 0.043271f
C3 VGND KAPWR 0.030073f
C4 VGND Y 0.10005f
C5 VPB A 0.09475f
C6 VPB KAPWR 0.022471f
C7 A KAPWR 0.047941f
C8 VPB Y 0.012263f
C9 VGND VPWR 0.005809f
C10 A Y 0.123649f
C11 KAPWR Y 0.175404f
C12 VPWR VPB 0.028996f
C13 VPWR A 0.01744f
C14 VPWR KAPWR 0.212352f
C15 VPWR VNB 0.16615f
C16 VGND VNB 0.226501f
C17 Y VNB 0.067884f
C18 KAPWR VNB 0.075678f
C19 A VNB 0.308156f
C20 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_2 VNB VPB KAPWR VPWR VGND A Y
X0 Y.t2 A.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 Y.t3 A.t1 KAPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 KAPWR.t1 A.t2 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND.t1 A.t3 Y.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 KAPWR.t0 A.t4 Y.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n1 A.t4 221.72
R1 A.n0 A.t1 221.72
R2 A.n7 A.t2 218.507
R3 A.n1 A.t3 189.052
R4 A.n2 A.t0 183.161
R5 A.n8 A.n7 181.087
R6 A.n4 A.n3 152
R7 A.n6 A.n5 152
R8 A.n3 A.n1 63.2789
R9 A.n6 A.n0 45.6184
R10 A.n7 A.n6 27.9589
R11 A.n5 A.n4 19.3427
R12 A.n8 A 16.2138
R13 A.n3 A.n2 10.3291
R14 A A.n8 9.95606
R15 A.n4 A 3.69828
R16 A.n5 A 3.12939
R17 A.n2 A.n0 2.58264
R18 VGND.n0 VGND.t0 249.679
R19 VGND.n0 VGND.t1 245.364
R20 VGND VGND.n0 0.591777
R21 Y.n2 Y.t0 445.25
R22 Y.n2 Y.n1 318.928
R23 Y.n3 Y.n0 222.707
R24 Y.n0 Y.t1 40.0005
R25 Y.n0 Y.t2 40.0005
R26 Y.n1 Y.t4 27.5805
R27 Y.n1 Y.t3 27.5805
R28 Y Y.n2 22.6425
R29 Y.n3 Y 13.4862
R30 Y Y.n3 2.05764
R31 VNB VNB.t1 2264.08
R32 VNB.t1 VNB.t0 1224.6
R33 KAPWR.n1 KAPWR.t0 333.192
R34 KAPWR.n1 KAPWR.n0 305.091
R35 KAPWR.n0 KAPWR.t2 27.5805
R36 KAPWR.n0 KAPWR.t1 27.5805
R37 KAPWR KAPWR.n1 0.317087
R38 VPB.t2 VPB.t0 254.518
R39 VPB.t1 VPB.t2 254.518
R40 VPB VPB.t1 207.166
C0 VPB Y 0.019021f
C1 VPWR VPB 0.036595f
C2 A Y 0.233176f
C3 VPB KAPWR 0.012254f
C4 VPWR A 0.025783f
C5 VPB VGND 0.004996f
C6 A KAPWR 0.043458f
C7 VPWR Y 0.052944f
C8 A VGND 0.073739f
C9 Y KAPWR 0.277661f
C10 VPWR KAPWR 0.261713f
C11 Y VGND 0.1235f
C12 VPWR VGND 0.004166f
C13 KAPWR VGND 0.038604f
C14 VPB A 0.10832f
C15 VPWR VNB 0.20334f
C16 VGND VNB 0.292563f
C17 KAPWR VNB 0.044434f
C18 Y VNB 0.109271f
C19 A VNB 0.373936f
C20 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_4 VNB VPB KAPWR VPWR VGND A Y
X0 Y.t7 A.t0 KAPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND.t3 A.t1 Y.t9 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1659 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND.t2 A.t2 Y.t8 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 KAPWR.t5 A.t3 Y.t6 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 KAPWR.t4 A.t4 Y.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y.t1 A.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y.t4 A.t6 KAPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y.t0 A.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1386 ps=1.5 w=0.42 l=0.15
X8 Y.t3 A.t8 KAPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 KAPWR.t1 A.t9 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n2 A.t4 276.168
R1 A.n8 A.t6 247.606
R2 A.n3 A.t0 221.72
R3 A.n5 A.t9 221.72
R4 A.n13 A.t8 221.72
R5 A.n7 A.t3 221.72
R6 A.n3 A.t1 186.374
R7 A.n5 A.t5 186.374
R8 A.n13 A.t2 186.374
R9 A.n7 A.t7 186.374
R10 A.n2 A.n1 152
R11 A.n4 A.n0 152
R12 A.n15 A.n14 152
R13 A.n12 A.n11 152
R14 A.n10 A.n6 152
R15 A.n9 A.n8 152
R16 A.n12 A.n6 60.6968
R17 A.n14 A.n13 54.4486
R18 A.n8 A.n7 50.8783
R19 A.n4 A.n3 38.382
R20 A.n5 A.n4 38.382
R21 A.n3 A.n2 22.3153
R22 A.n14 A.n5 22.3153
R23 A.n1 A.n0 19.3427
R24 A.n10 A.n9 19.3427
R25 A A.n15 17.3516
R26 A.n11 A 15.6449
R27 A.n11 A 10.5249
R28 A.n7 A.n6 9.81902
R29 A.n15 A 8.81828
R30 A.n13 A.n12 6.24865
R31 A.n1 A 4.83606
R32 A A.n10 3.69828
R33 A.n9 A 3.12939
R34 A A.n0 1.99161
R35 KAPWR.n1 KAPWR.t4 333.18
R36 KAPWR.n4 KAPWR.t3 332.671
R37 KAPWR.n3 KAPWR.n2 305.091
R38 KAPWR.n1 KAPWR.n0 305.091
R39 KAPWR.n2 KAPWR.t2 27.5805
R40 KAPWR.n2 KAPWR.t5 27.5805
R41 KAPWR.n0 KAPWR.t0 27.5805
R42 KAPWR.n0 KAPWR.t1 27.5805
R43 KAPWR.n3 KAPWR.n1 0.521173
R44 KAPWR.n4 KAPWR.n3 0.496173
R45 KAPWR KAPWR.n4 0.0557885
R46 Y.n7 Y.n4 315.615
R47 Y.n9 Y.n2 315.613
R48 Y.n8 Y.n3 315.613
R49 Y.n1 Y.n0 203.322
R50 Y.n6 Y.n5 202.97
R51 Y.n7 Y.n6 146.447
R52 Y.n9 Y.n8 64.7534
R53 Y.n8 Y.n7 64.7534
R54 Y.n10 Y.n1 51.9534
R55 Y.n6 Y.n1 45.177
R56 Y.n0 Y.t9 40.0005
R57 Y.n0 Y.t1 40.0005
R58 Y.n5 Y.t8 40.0005
R59 Y.n5 Y.t0 40.0005
R60 Y Y.n9 33.2554
R61 Y.n2 Y.t5 27.5805
R62 Y.n2 Y.t7 27.5805
R63 Y.n3 Y.t2 27.5805
R64 Y.n3 Y.t3 27.5805
R65 Y.n4 Y.t6 27.5805
R66 Y.n4 Y.t4 27.5805
R67 Y.n10 Y 12.5872
R68 Y Y.n10 1.9205
R69 VPB.t5 VPB.t3 254.518
R70 VPB.t0 VPB.t5 254.518
R71 VPB.t1 VPB.t0 254.518
R72 VPB.t4 VPB.t1 254.518
R73 VPB.t2 VPB.t4 254.518
R74 VPB VPB.t2 219.004
R75 VGND.n1 VGND.t3 247.148
R76 VGND.n5 VGND.t0 241.923
R77 VGND.n3 VGND.n2 204.201
R78 VGND.n2 VGND.t1 40.0005
R79 VGND.n2 VGND.t2 40.0005
R80 VGND.n4 VGND.n3 23.3417
R81 VGND.n5 VGND.n4 21.8358
R82 VGND.n4 VGND.n0 9.3005
R83 VGND.n6 VGND.n5 7.30743
R84 VGND.n3 VGND.n1 6.81041
R85 VGND.n1 VGND.n0 0.58231
R86 VGND.n6 VGND.n0 0.146144
R87 VGND VGND.n6 0.117248
R88 VNB VNB.t0 2278.32
R89 VNB.t1 VNB.t3 1224.6
R90 VNB.t2 VNB.t1 1224.6
R91 VNB.t0 VNB.t2 1224.6
C0 Y VGND 0.317378f
C1 VPB VPWR 0.056144f
C2 A VPWR 0.04747f
C3 VPB A 0.192877f
C4 KAPWR VPWR 0.486817f
C5 VPB KAPWR 0.018359f
C6 Y VPWR 0.080072f
C7 A KAPWR 0.084832f
C8 VPB Y 0.024655f
C9 VGND VPWR 0.004365f
C10 VPB VGND 0.006215f
C11 A Y 0.590483f
C12 A VGND 0.082801f
C13 KAPWR Y 0.519324f
C14 KAPWR VGND 0.070455f
C15 VPWR VNB 0.318489f
C16 VGND VNB 0.426146f
C17 Y VNB 0.154641f
C18 KAPWR VNB 0.06393f
C19 A VNB 0.602468f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_8 VNB VPB KAPWR VGND VPWR A Y
X0 Y.t7 A.t0 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 KAPWR.t11 A.t1 Y.t19 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t6 A.t2 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 Y.t5 A.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y.t18 A.t4 KAPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 KAPWR.t9 A.t5 Y.t17 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X6 KAPWR.t8 A.t6 Y.t16 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t4 A.t7 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 Y.t15 A.t8 KAPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t3 A.t9 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 Y.t14 A.t10 KAPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1375 ps=1.275 w=1 l=0.15
X11 KAPWR.t5 A.t11 Y.t13 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t2 A.t12 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 KAPWR.t4 A.t13 Y.t12 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t11 A.t14 KAPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t1 A.t15 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 KAPWR.t2 A.t16 Y.t10 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y.t9 A.t17 KAPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t8 A.t18 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND.t0 A.t19 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A.n8 A.t11 225.911
R1 A.n41 A.t18 205.375
R2 A.n7 A.t8 192.8
R3 A.n11 A.t13 192.8
R4 A.n5 A.t14 192.8
R5 A.n18 A.t16 192.8
R6 A.n23 A.t17 192.8
R7 A.n3 A.t1 192.8
R8 A.n30 A.t4 192.8
R9 A.n33 A.t6 192.8
R10 A.n1 A.t10 192.8
R11 A.n40 A.t5 192.8
R12 A.n9 A.n8 169.067
R13 A.n10 A.n9 152
R14 A.n14 A.n13 152
R15 A.n16 A.n15 152
R16 A.n20 A.n19 152
R17 A.n22 A.n21 152
R18 A.n26 A.n25 152
R19 A.n28 A.n27 152
R20 A.n31 A.n2 152
R21 A.n36 A.n35 152
R22 A.n38 A.n37 152
R23 A.n39 A.n0 152
R24 A.n42 A.n41 152
R25 A.n34 A.t0 117.287
R26 A.n32 A.t15 117.287
R27 A.n29 A.t7 117.287
R28 A.n24 A.t12 117.287
R29 A.n4 A.t3 117.287
R30 A.n17 A.t9 117.287
R31 A.n12 A.t2 117.287
R32 A.n6 A.t19 117.287
R33 A.n39 A.n38 28.5014
R34 A.n24 A.n23 24.3101
R35 A.n41 A.n40 22.6335
R36 A.n28 A.n3 21.3762
R37 A.n7 A.n6 20.957
R38 A.n13 A.n11 19.6996
R39 A.n35 A.n34 18.8614
R40 A.n19 A.n4 17.1848
R41 A.n21 A.n20 17.0672
R42 A.n36 A.n2 17.0672
R43 A.n42 A.n0 17.0672
R44 A.n27 A 16.5652
R45 A.n15 A 15.5613
R46 A.n31 A.n30 14.6701
R47 A.n14 A 13.5534
R48 A.n12 A.n5 13.4127
R49 A.n16 A.n5 12.9935
R50 A.n18 A.n17 12.5744
R51 A.n26 A 12.5495
R52 A.n37 A 11.5456
R53 A.n37 A 11.5456
R54 A.n22 A.n4 11.317
R55 A.n32 A.n31 11.317
R56 A A.n26 10.5417
R57 A.n30 A.n29 10.0596
R58 A.n17 A.n16 9.6405
R59 A A.n14 9.53776
R60 A.n33 A.n32 9.22137
R61 A.n11 A.n10 8.80224
R62 A.n34 A.n1 8.38311
R63 A.n35 A.n33 7.96398
R64 A.n15 A 7.52991
R65 A.n25 A.n3 7.12572
R66 A.n27 A 6.52599
R67 A.n19 A.n18 6.28746
R68 A.n40 A.n39 5.86833
R69 A A.n36 5.52207
R70 A A.n0 5.52207
R71 A.n10 A.n6 5.4492
R72 A.n21 A 4.51815
R73 A.n25 A.n24 3.77267
R74 A.n29 A.n28 3.77267
R75 A.n9 A 3.51423
R76 A.n8 A.n7 2.09615
R77 A.n13 A.n12 2.09615
R78 A.n20 A 1.50638
R79 A.n38 A.n1 1.25789
R80 A A.n2 0.502461
R81 A A.n42 0.502461
R82 A.n23 A.n22 0.41963
R83 VGND.n4 VGND.t0 245.494
R84 VGND.n15 VGND.t7 240.127
R85 VGND.n6 VGND.n5 200.127
R86 VGND.n9 VGND.n8 200.127
R87 VGND.n13 VGND.n2 200.127
R88 VGND.n5 VGND.t6 40.0005
R89 VGND.n5 VGND.t3 40.0005
R90 VGND.n8 VGND.t5 40.0005
R91 VGND.n8 VGND.t2 40.0005
R92 VGND.n2 VGND.t4 40.0005
R93 VGND.n2 VGND.t1 40.0005
R94 VGND.n9 VGND.n7 27.4829
R95 VGND.n13 VGND.n1 22.9652
R96 VGND.n14 VGND.n13 21.4593
R97 VGND.n15 VGND.n14 18.4476
R98 VGND.n9 VGND.n1 16.9417
R99 VGND.n7 VGND.n6 12.424
R100 VGND.n7 VGND.n3 9.3005
R101 VGND.n10 VGND.n9 9.3005
R102 VGND.n11 VGND.n1 9.3005
R103 VGND.n13 VGND.n12 9.3005
R104 VGND.n14 VGND.n0 9.3005
R105 VGND.n16 VGND.n15 7.26269
R106 VGND.n6 VGND.n4 6.80308
R107 VGND.n4 VGND.n3 0.797793
R108 VGND VGND.n16 0.231207
R109 VGND.n16 VGND.n0 0.15127
R110 VGND.n10 VGND.n3 0.120292
R111 VGND.n11 VGND.n10 0.120292
R112 VGND.n12 VGND.n11 0.120292
R113 VGND.n12 VGND.n0 0.120292
R114 Y.n14 Y.n7 321.353
R115 Y.n19 Y.n2 315.613
R116 Y.n18 Y.n3 315.613
R117 Y.n17 Y.n4 315.613
R118 Y.n16 Y.n5 315.613
R119 Y.n15 Y.n6 315.613
R120 Y.n1 Y.n0 207.569
R121 Y.n9 Y.n8 207.569
R122 Y.n11 Y.n10 207.569
R123 Y.n13 Y.n12 207.569
R124 Y.n14 Y.n13 181.459
R125 Y.n20 Y.n1 65.1299
R126 Y.n15 Y.n14 63.624
R127 Y.n19 Y.n18 63.2476
R128 Y.n18 Y.n17 63.2476
R129 Y.n17 Y.n16 63.2476
R130 Y.n16 Y.n15 63.2476
R131 Y.n9 Y.n1 50.4476
R132 Y.n11 Y.n9 50.4476
R133 Y.n13 Y.n11 50.4476
R134 Y.n0 Y.t0 40.0005
R135 Y.n0 Y.t6 40.0005
R136 Y.n8 Y.t3 40.0005
R137 Y.n8 Y.t5 40.0005
R138 Y.n10 Y.t2 40.0005
R139 Y.n10 Y.t4 40.0005
R140 Y.n12 Y.t1 40.0005
R141 Y.n12 Y.t7 40.0005
R142 Y.n2 Y.t13 26.5955
R143 Y.n2 Y.t15 26.5955
R144 Y.n3 Y.t12 26.5955
R145 Y.n3 Y.t11 26.5955
R146 Y.n4 Y.t10 26.5955
R147 Y.n4 Y.t9 26.5955
R148 Y.n5 Y.t19 26.5955
R149 Y.n5 Y.t18 26.5955
R150 Y.n6 Y.t16 26.5955
R151 Y.n6 Y.t14 26.5955
R152 Y.n7 Y.t17 26.5955
R153 Y.n7 Y.t8 26.5955
R154 Y Y.n19 26.2001
R155 Y.n20 Y 15.4079
R156 Y Y.n20 0.711611
R157 VNB VNB.t7 3602.59
R158 VNB.t6 VNB.t0 1224.6
R159 VNB.t3 VNB.t6 1224.6
R160 VNB.t5 VNB.t3 1224.6
R161 VNB.t2 VNB.t5 1224.6
R162 VNB.t4 VNB.t2 1224.6
R163 VNB.t1 VNB.t4 1224.6
R164 VNB.t7 VNB.t1 1224.6
R165 KAPWR.n1 KAPWR.t5 332.207
R166 KAPWR.n10 KAPWR.t0 331.687
R167 KAPWR.n9 KAPWR.n8 305.091
R168 KAPWR.n7 KAPWR.n6 305.091
R169 KAPWR.n5 KAPWR.n4 305.091
R170 KAPWR.n3 KAPWR.n2 305.091
R171 KAPWR.n1 KAPWR.n0 305.091
R172 KAPWR.n8 KAPWR.t9 27.5805
R173 KAPWR.n8 KAPWR.t6 26.5955
R174 KAPWR.n6 KAPWR.t10 26.5955
R175 KAPWR.n6 KAPWR.t8 26.5955
R176 KAPWR.n4 KAPWR.t1 26.5955
R177 KAPWR.n4 KAPWR.t11 26.5955
R178 KAPWR.n2 KAPWR.t3 26.5955
R179 KAPWR.n2 KAPWR.t2 26.5955
R180 KAPWR.n0 KAPWR.t7 26.5955
R181 KAPWR.n0 KAPWR.t4 26.5955
R182 KAPWR.n9 KAPWR.n7 0.521173
R183 KAPWR.n7 KAPWR.n5 0.508673
R184 KAPWR.n3 KAPWR.n1 0.496173
R185 KAPWR.n10 KAPWR.n9 0.496173
R186 KAPWR.n5 KAPWR.n3 0.411798
R187 KAPWR KAPWR.n10 0.0221346
R188 VPB.t9 VPB.t6 251.559
R189 VPB.t7 VPB.t5 248.599
R190 VPB.t4 VPB.t7 248.599
R191 VPB.t3 VPB.t4 248.599
R192 VPB.t2 VPB.t3 248.599
R193 VPB.t1 VPB.t2 248.599
R194 VPB.t11 VPB.t1 248.599
R195 VPB.t10 VPB.t11 248.599
R196 VPB.t8 VPB.t10 248.599
R197 VPB.t6 VPB.t8 248.599
R198 VPB.t0 VPB.t9 248.599
R199 VPB VPB.t0 189.409
C0 VPB A 0.371833f
C1 VPB KAPWR 0.033596f
C2 A KAPWR 0.185827f
C3 VPB Y 0.02699f
C4 VPB VGND 0.011303f
C5 A Y 1.1944f
C6 A VGND 0.173084f
C7 VPB VPWR 0.100245f
C8 KAPWR Y 1.00388f
C9 A VPWR 0.076623f
C10 KAPWR VGND 0.132214f
C11 KAPWR VPWR 0.900696f
C12 Y VGND 0.563854f
C13 Y VPWR 0.151222f
C14 VGND VPWR 0.008416f
C15 VPWR VNB 0.556555f
C16 VGND VNB 0.715601f
C17 Y VNB 0.161499f
C18 KAPWR VNB 0.059724f
C19 A VNB 1.15234f
C20 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_16 Y A KAPWR VGND VPWR VNB VPB
X0 VGND.t15 A.t0 Y.t16 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 Y.t3 A.t1 KAPWR.t23 VPB.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 KAPWR.t22 A.t2 Y.t2 VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X3 Y.t1 A.t3 KAPWR.t21 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND.t14 A.t4 Y.t15 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 KAPWR.t20 A.t5 Y.t0 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y.t14 A.t6 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND.t12 A.t7 Y.t13 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 KAPWR.t19 A.t8 Y.t39 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 KAPWR.t18 A.t9 Y.t38 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 Y.t12 A.t10 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 Y.t37 A.t11 KAPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 KAPWR.t16 A.t12 Y.t36 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2175 ps=1.435 w=1 l=0.15
X13 VGND.t10 A.t13 Y.t11 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 Y.t35 A.t14 KAPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.275 ps=2.55 w=1 l=0.15
X15 KAPWR.t14 A.t15 Y.t34 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y.t33 A.t16 KAPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 Y.t32 A.t17 KAPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 Y.t10 A.t18 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VGND.t8 A.t19 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 Y.t8 A.t20 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 VGND.t6 A.t21 Y.t7 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 Y.t31 A.t22 KAPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 KAPWR.t10 A.t23 Y.t30 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 Y.t29 A.t24 KAPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.1575 ps=1.315 w=1 l=0.15
X25 Y.t28 A.t25 KAPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 KAPWR.t7 A.t26 Y.t27 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 Y.t6 A.t27 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 Y.t26 A.t28 KAPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 KAPWR.t5 A.t29 Y.t25 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 KAPWR.t4 A.t30 Y.t24 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 Y.t5 A.t31 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 VGND.t3 A.t32 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 KAPWR.t3 A.t33 Y.t23 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 Y.t19 A.t34 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.09135 pd=0.855 as=0.06615 ps=0.735 w=0.42 l=0.15
X35 Y.t22 A.t35 KAPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 Y.t18 A.t36 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X37 KAPWR.t1 A.t37 Y.t21 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 Y.t20 A.t38 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND.t0 A.t39 Y.t17 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.09135 ps=0.855 w=0.42 l=0.15
R0 A.n5 A.t30 218.106
R1 A.n34 A.t14 218.106
R2 A.n6 A.t28 204.048
R3 A.n9 A.t29 204.048
R4 A.n2 A.t17 204.048
R5 A.n16 A.t5 204.048
R6 A.n17 A.t38 204.048
R7 A.n18 A.t26 204.048
R8 A.n19 A.t16 204.048
R9 A.n20 A.t15 204.048
R10 A.n21 A.t3 204.048
R11 A.n22 A.t37 204.048
R12 A.n23 A.t25 204.048
R13 A.n24 A.t12 204.048
R14 A.n25 A.t24 204.048
R15 A.n26 A.t2 204.048
R16 A.n27 A.t35 204.048
R17 A.n28 A.t23 204.048
R18 A.n29 A.t11 204.048
R19 A.n30 A.t9 204.048
R20 A.n31 A.t1 204.048
R21 A.n40 A.t33 204.048
R22 A.n38 A.t22 204.048
R23 A.n33 A.t8 204.048
R24 A.n16 A.t0 175.127
R25 A.n17 A.t10 175.127
R26 A.n18 A.t4 175.127
R27 A.n19 A.t18 175.127
R28 A.n20 A.t7 175.127
R29 A.n21 A.t20 175.127
R30 A.n22 A.t32 175.127
R31 A.n23 A.t27 175.127
R32 A.n24 A.t39 175.127
R33 A.n25 A.t34 175.127
R34 A.n26 A.t13 175.127
R35 A.n27 A.t6 175.127
R36 A.n28 A.t19 175.127
R37 A.n29 A.t31 175.127
R38 A.n30 A.t21 175.127
R39 A.n31 A.t36 175.127
R40 A.n5 A.n4 163.453
R41 A.n35 A.n34 163.453
R42 A.n15 A.n14 163.117
R43 A.n7 A.n4 152
R44 A.n11 A.n10 152
R45 A.n8 A.n3 152
R46 A.n42 A.n41 152
R47 A.n39 A.n1 152
R48 A.n37 A.n36 152
R49 A.n35 A.n32 152
R50 A.n25 A.n24 78.3255
R51 A.n26 A.n25 62.2588
R52 A.n17 A.n16 57.5727
R53 A.n18 A.n17 57.5727
R54 A.n19 A.n18 57.5727
R55 A.n20 A.n19 57.5727
R56 A.n21 A.n20 57.5727
R57 A.n22 A.n21 57.5727
R58 A.n23 A.n22 57.5727
R59 A.n24 A.n23 57.5727
R60 A.n27 A.n26 57.5727
R61 A.n28 A.n27 57.5727
R62 A.n29 A.n28 57.5727
R63 A.n30 A.n29 57.5727
R64 A.n31 A.n30 57.5727
R65 A.n10 A.n7 45.5227
R66 A.n37 A.n32 45.5227
R67 A.n6 A.n5 43.5144
R68 A.n34 A.n33 43.5144
R69 A.n9 A.n8 35.4811
R70 A.n39 A.n38 35.4811
R71 A.n16 A.n15 34.1422
R72 A.n41 A.n31 34.1422
R73 A.n15 A.n2 23.4311
R74 A.n41 A.n40 23.4311
R75 A.n8 A.n2 22.0922
R76 A.n40 A.n39 22.0922
R77 A A.n0 12.1637
R78 A.n11 A.n3 11.4531
R79 A.n42 A.n1 11.4531
R80 A.n36 A.n1 11.4531
R81 A.n36 A.n35 11.4531
R82 A.n10 A.n9 10.0422
R83 A.n38 A.n37 10.0422
R84 A.n13 A.n12 9.5505
R85 A.n1 A.n0 9.5505
R86 A.n14 A.n13 9.3005
R87 A.n12 A.n4 7.74787
R88 A.n13 A.n0 6.47061
R89 A.n12 A.n11 3.70576
R90 A.n7 A.n6 2.00883
R91 A.n33 A.n32 2.00883
R92 A A.n42 1.17945
R93 A.n14 A.n3 0.337342
R94 Y.n24 Y.n23 356.142
R95 Y.n11 Y.n9 308.26
R96 Y.n31 Y.n29 307.029
R97 Y.n28 Y.n15 303.724
R98 Y.n27 Y.n17 303.724
R99 Y.n26 Y.n19 303.724
R100 Y.n25 Y.n21 303.724
R101 Y.n24 Y.n22 303.724
R102 Y.n13 Y.n0 303.724
R103 Y.n7 Y.n3 303.724
R104 Y.n6 Y.n4 303.724
R105 Y.n6 Y.n5 259.678
R106 Y.n8 Y.n2 240.183
R107 Y.n11 Y.n10 239.965
R108 Y.n12 Y.n1 236.733
R109 Y.n28 Y.n14 234.665
R110 Y.n27 Y.n16 234.665
R111 Y.n26 Y.n18 234.665
R112 Y.n25 Y.n20 234.665
R113 Y Y.n30 221.571
R114 Y.n30 Y.t17 75.7148
R115 Y.n29 Y.t29 53.1905
R116 Y.n7 Y.n6 51.4931
R117 Y.n25 Y.n24 51.2005
R118 Y.n30 Y.t19 48.5719
R119 Y.n26 Y.n25 44.0325
R120 Y.n27 Y.n26 44.0325
R121 Y.n28 Y.n27 44.0325
R122 Y.n31 Y.n28 40.7045
R123 Y.n14 Y.t4 40.0005
R124 Y.n14 Y.t6 40.0005
R125 Y.n16 Y.t13 40.0005
R126 Y.n16 Y.t8 40.0005
R127 Y.n18 Y.t15 40.0005
R128 Y.n18 Y.t10 40.0005
R129 Y.n20 Y.t16 40.0005
R130 Y.n20 Y.t12 40.0005
R131 Y.n2 Y.t7 40.0005
R132 Y.n2 Y.t18 40.0005
R133 Y.n10 Y.t9 40.0005
R134 Y.n10 Y.t5 40.0005
R135 Y.n1 Y.t11 40.0005
R136 Y.n1 Y.t14 40.0005
R137 Y.n31 Y.n13 39.1685
R138 Y.n12 Y.n11 37.1205
R139 Y.n11 Y.n8 36.8645
R140 Y.n29 Y.t36 32.5055
R141 Y.n15 Y.t21 27.5805
R142 Y.n15 Y.t28 27.5805
R143 Y.n17 Y.t34 27.5805
R144 Y.n17 Y.t1 27.5805
R145 Y.n19 Y.t27 27.5805
R146 Y.n19 Y.t33 27.5805
R147 Y.n21 Y.t0 27.5805
R148 Y.n21 Y.t20 27.5805
R149 Y.n22 Y.t25 27.5805
R150 Y.n22 Y.t32 27.5805
R151 Y.n23 Y.t24 27.5805
R152 Y.n23 Y.t26 27.5805
R153 Y.n0 Y.t2 27.5805
R154 Y.n0 Y.t22 27.5805
R155 Y.n3 Y.t38 27.5805
R156 Y.n3 Y.t3 27.5805
R157 Y.n5 Y.t39 27.5805
R158 Y.n5 Y.t35 27.5805
R159 Y.n4 Y.t23 27.5805
R160 Y.n4 Y.t31 27.5805
R161 Y.n9 Y.t30 27.5805
R162 Y.n9 Y.t37 27.5805
R163 Y.n31 Y 3.47479
R164 Y Y.n31 2.5605
R165 Y.n8 Y.n7 0.7685
R166 Y.n13 Y.n12 0.2565
R167 VGND.n7 VGND.t15 251.076
R168 VGND.n40 VGND.t1 246.096
R169 VGND.n19 VGND.n18 210.316
R170 VGND.n9 VGND.n8 206.494
R171 VGND.n12 VGND.n11 206.494
R172 VGND.n22 VGND.n21 206.494
R173 VGND.n28 VGND.n27 206.494
R174 VGND.n31 VGND.n30 206.494
R175 VGND.n38 VGND.n37 206.494
R176 VGND.n27 VGND.t10 47.1434
R177 VGND.n27 VGND.t2 42.8576
R178 VGND.n8 VGND.t11 40.0005
R179 VGND.n8 VGND.t14 40.0005
R180 VGND.n11 VGND.t9 40.0005
R181 VGND.n11 VGND.t12 40.0005
R182 VGND.n18 VGND.t7 40.0005
R183 VGND.n18 VGND.t3 40.0005
R184 VGND.n21 VGND.t5 40.0005
R185 VGND.n21 VGND.t0 40.0005
R186 VGND.n30 VGND.t13 40.0005
R187 VGND.n30 VGND.t8 40.0005
R188 VGND.n37 VGND.t4 40.0005
R189 VGND.n37 VGND.t6 40.0005
R190 VGND.n13 VGND.n10 34.6358
R191 VGND.n17 VGND.n5 34.6358
R192 VGND.n26 VGND.n3 34.6358
R193 VGND.n32 VGND.n29 34.6358
R194 VGND.n36 VGND.n1 34.6358
R195 VGND.n22 VGND.n20 34.2593
R196 VGND.n40 VGND.n39 30.4946
R197 VGND.n9 VGND.n7 19.3233
R198 VGND.n22 VGND.n3 15.0593
R199 VGND.n39 VGND.n38 14.3064
R200 VGND.n20 VGND.n19 10.5417
R201 VGND.n31 VGND.n1 9.78874
R202 VGND.n10 VGND.n6 9.3005
R203 VGND.n14 VGND.n13 9.3005
R204 VGND.n15 VGND.n5 9.3005
R205 VGND.n17 VGND.n16 9.3005
R206 VGND.n20 VGND.n4 9.3005
R207 VGND.n23 VGND.n22 9.3005
R208 VGND.n24 VGND.n3 9.3005
R209 VGND.n26 VGND.n25 9.3005
R210 VGND.n29 VGND.n2 9.3005
R211 VGND.n33 VGND.n32 9.3005
R212 VGND.n34 VGND.n1 9.3005
R213 VGND.n36 VGND.n35 9.3005
R214 VGND.n39 VGND.n0 9.3005
R215 VGND.n13 VGND.n12 8.65932
R216 VGND.n28 VGND.n26 7.52991
R217 VGND.n19 VGND.n17 7.15344
R218 VGND.n29 VGND.n28 7.15344
R219 VGND.n41 VGND.n40 6.82589
R220 VGND.n12 VGND.n5 6.02403
R221 VGND.n32 VGND.n31 4.89462
R222 VGND.n10 VGND.n9 1.50638
R223 VGND.n7 VGND.n6 1.46762
R224 VGND VGND.n41 0.465247
R225 VGND.n38 VGND.n36 0.376971
R226 VGND.n41 VGND.n0 0.159177
R227 VGND.n14 VGND.n6 0.120292
R228 VGND.n15 VGND.n14 0.120292
R229 VGND.n16 VGND.n15 0.120292
R230 VGND.n16 VGND.n4 0.120292
R231 VGND.n23 VGND.n4 0.120292
R232 VGND.n24 VGND.n23 0.120292
R233 VGND.n25 VGND.n24 0.120292
R234 VGND.n25 VGND.n2 0.120292
R235 VGND.n33 VGND.n2 0.120292
R236 VGND.n34 VGND.n33 0.120292
R237 VGND.n35 VGND.n34 0.120292
R238 VGND.n35 VGND.n0 0.120292
R239 VNB VNB.t1 5866.67
R240 VNB.t2 VNB.t0 1666.02
R241 VNB.t10 VNB.t2 1324.27
R242 VNB.t11 VNB.t15 1224.6
R243 VNB.t14 VNB.t11 1224.6
R244 VNB.t9 VNB.t14 1224.6
R245 VNB.t12 VNB.t9 1224.6
R246 VNB.t7 VNB.t12 1224.6
R247 VNB.t3 VNB.t7 1224.6
R248 VNB.t5 VNB.t3 1224.6
R249 VNB.t0 VNB.t5 1224.6
R250 VNB.t13 VNB.t10 1224.6
R251 VNB.t8 VNB.t13 1224.6
R252 VNB.t4 VNB.t8 1224.6
R253 VNB.t6 VNB.t4 1224.6
R254 VNB.t1 VNB.t6 1224.6
R255 KAPWR.n1 KAPWR.t4 332.212
R256 KAPWR.n21 KAPWR.n20 305.096
R257 KAPWR.n19 KAPWR.n18 305.096
R258 KAPWR.n17 KAPWR.n16 305.096
R259 KAPWR.n15 KAPWR.n14 305.096
R260 KAPWR.n13 KAPWR.n12 305.096
R261 KAPWR.n11 KAPWR.n10 305.096
R262 KAPWR.n9 KAPWR.n8 305.096
R263 KAPWR.n7 KAPWR.n6 305.096
R264 KAPWR.n5 KAPWR.n4 305.096
R265 KAPWR.n3 KAPWR.n2 305.096
R266 KAPWR.n1 KAPWR.n0 305.096
R267 KAPWR.n22 KAPWR.t15 236.488
R268 KAPWR.n12 KAPWR.t22 31.5205
R269 KAPWR.n12 KAPWR.t9 30.5355
R270 KAPWR.n10 KAPWR.t8 28.5655
R271 KAPWR.n20 KAPWR.t11 27.5805
R272 KAPWR.n20 KAPWR.t19 27.5805
R273 KAPWR.n18 KAPWR.t23 27.5805
R274 KAPWR.n18 KAPWR.t3 27.5805
R275 KAPWR.n16 KAPWR.t17 27.5805
R276 KAPWR.n16 KAPWR.t18 27.5805
R277 KAPWR.n14 KAPWR.t2 27.5805
R278 KAPWR.n14 KAPWR.t10 27.5805
R279 KAPWR.n8 KAPWR.t21 27.5805
R280 KAPWR.n8 KAPWR.t1 27.5805
R281 KAPWR.n6 KAPWR.t13 27.5805
R282 KAPWR.n6 KAPWR.t14 27.5805
R283 KAPWR.n4 KAPWR.t0 27.5805
R284 KAPWR.n4 KAPWR.t7 27.5805
R285 KAPWR.n2 KAPWR.t12 27.5805
R286 KAPWR.n2 KAPWR.t20 27.5805
R287 KAPWR.n0 KAPWR.t6 27.5805
R288 KAPWR.n0 KAPWR.t5 27.5805
R289 KAPWR.n10 KAPWR.t16 26.5955
R290 KAPWR.n11 KAPWR.n9 0.533673
R291 KAPWR.n17 KAPWR.n15 0.533673
R292 KAPWR.n7 KAPWR.n5 0.521173
R293 KAPWR.n13 KAPWR.n11 0.521173
R294 KAPWR.n21 KAPWR.n19 0.521173
R295 KAPWR.n19 KAPWR.n17 0.508673
R296 KAPWR.n3 KAPWR.n1 0.496173
R297 KAPWR.n9 KAPWR.n7 0.496173
R298 KAPWR.n15 KAPWR.n13 0.496173
R299 KAPWR.n22 KAPWR.n21 0.496173
R300 KAPWR.n5 KAPWR.n3 0.477423
R301 KAPWR KAPWR.n22 0.0293462
R302 VPB.t9 VPB.t16 346.262
R303 VPB.t22 VPB.t9 275.235
R304 VPB.t6 VPB.t4 254.518
R305 VPB.t5 VPB.t6 254.518
R306 VPB.t12 VPB.t5 254.518
R307 VPB.t20 VPB.t12 254.518
R308 VPB.t0 VPB.t20 254.518
R309 VPB.t7 VPB.t0 254.518
R310 VPB.t13 VPB.t7 254.518
R311 VPB.t14 VPB.t13 254.518
R312 VPB.t21 VPB.t14 254.518
R313 VPB.t1 VPB.t21 254.518
R314 VPB.t8 VPB.t1 254.518
R315 VPB.t16 VPB.t8 254.518
R316 VPB.t2 VPB.t22 254.518
R317 VPB.t10 VPB.t2 254.518
R318 VPB.t17 VPB.t10 254.518
R319 VPB.t18 VPB.t17 254.518
R320 VPB.t23 VPB.t18 254.518
R321 VPB.t3 VPB.t23 254.518
R322 VPB.t11 VPB.t3 254.518
R323 VPB.t19 VPB.t11 254.518
R324 VPB.t15 VPB.t19 254.518
R325 VPB VPB.t15 201.246
C0 VPB KAPWR 0.03281f
C1 A KAPWR 0.680499f
C2 VPB Y 0.047038f
C3 VPB VGND 0.007999f
C4 A Y 1.67561f
C5 A VGND 0.795781f
C6 VPB VPWR 0.168046f
C7 KAPWR Y 1.8976f
C8 A VPWR 0.152946f
C9 KAPWR VGND 0.059235f
C10 KAPWR VPWR 1.67779f
C11 Y VGND 0.804977f
C12 Y VPWR 0.331167f
C13 VGND VPWR 0.004565f
C14 VPB A 0.7812f
C15 VPWR VNB 0.97722f
C16 VGND VNB 1.29662f
C17 Y VNB 0.137982f
C18 KAPWR VNB 0.071079f
C19 A VNB 2.36074f
C20 VPB VNB 2.19949f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_3.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_3 VPWR VGND KAPWR VPB VNB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
R0 VGND.n1 VGND.t2 259.082
R1 VGND.n0 VGND.t0 216.798
R2 VGND.n2 VGND.t1 214.456
R3 VGND.n3 VGND.n2 9.71789
R4 VGND.n1 VGND.n0 7.01592
R5 VGND.n3 VGND.n0 3.76277
R6 VGND.n2 VGND.n1 1.18311
R7 VGND VGND.n3 0.0226354
R8 KAPWR.n1 KAPWR.t0 381.443
R9 KAPWR.n4 KAPWR.t1 381.443
R10 KAPWR.n2 KAPWR.t2 242.282
R11 KAPWR.n1 KAPWR.n0 9.93905
R12 KAPWR.n5 KAPWR.n4 9.71789
R13 KAPWR.n3 KAPWR.n0 9.3005
R14 KAPWR.n4 KAPWR.n3 5.98311
R15 KAPWR.n3 KAPWR.n2 4.8005
R16 KAPWR.n2 KAPWR.n1 1.18311
R17 KAPWR.n5 KAPWR.n0 0.221654
R18 KAPWR KAPWR.n5 0.03175
R19 VPB VPB.t0 315.767
R20 VNB VNB.t0 1487.5
C0 VPB KAPWR 0.037232f
C1 VGND KAPWR 0.345679f
C2 VPB VPWR 0.027424f
C3 VGND VPWR 0.016799f
C4 KAPWR VPWR 0.261774f
C5 VPB VGND 0.079601f
C6 VPWR VNB 0.165266f
C7 KAPWR VNB 0.314272f
C8 VGND VNB 0.428813f
C9 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_4 VGND VPWR KAPWR VPB VNB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
R0 VGND.n1 VGND.t2 218.308
R1 VGND.n0 VGND.t0 218.243
R2 VGND.n2 VGND.t1 214.456
R3 VGND.n3 VGND.n2 9.70901
R4 VGND.n1 VGND.n0 6.78155
R5 VGND.n2 VGND.n1 2.7239
R6 VGND.n3 VGND.n0 1.75362
R7 VGND VGND.n3 0.0226354
R8 KAPWR.n6 KAPWR.t1 388.656
R9 KAPWR.n2 KAPWR.t0 388.656
R10 KAPWR.n1 KAPWR.t2 210.964
R11 KAPWR.n3 KAPWR.n2 9.93905
R12 KAPWR.n7 KAPWR.n6 9.71789
R13 KAPWR.n4 KAPWR.n3 9.3005
R14 KAPWR.n5 KAPWR.n0 9.3005
R15 KAPWR.n5 KAPWR.n4 6.4005
R16 KAPWR.n6 KAPWR.n5 5.98311
R17 KAPWR.n4 KAPWR.n1 3.2005
R18 KAPWR.n2 KAPWR.n1 2.78311
R19 KAPWR.n3 KAPWR.n0 0.221654
R20 KAPWR.n7 KAPWR.n0 0.221654
R21 KAPWR KAPWR.n7 0.03175
R22 VPB VPB.t0 458.724
R23 VNB VNB.t0 2207.12
C0 VPB KAPWR 0.048521f
C1 VGND KAPWR 0.535692f
C2 VPB VPWR 0.032492f
C3 VGND VPWR 0.025664f
C4 KAPWR VPWR 0.359985f
C5 VPB VGND 0.116183f
C6 VPWR VNB 0.203066f
C7 KAPWR VNB 0.425681f
C8 VGND VNB 0.556326f
C9 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_6 VPWR VGND KAPWR VPB VNB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
R0 VGND.n1 VGND.t0 219.12
R1 VGND.n0 VGND.t1 214.456
R2 VGND.n0 VGND.t2 121.927
R3 VGND.n1 VGND.n0 4.29166
R4 VGND VGND.n1 0.929743
R5 KAPWR.n3 KAPWR.t0 806.106
R6 KAPWR.t0 KAPWR.n2 751.692
R7 KAPWR.n7 KAPWR.t1 388.656
R8 KAPWR.n2 KAPWR.t2 133.512
R9 KAPWR.n8 KAPWR.n7 9.71789
R10 KAPWR.n5 KAPWR.n4 9.3005
R11 KAPWR.n6 KAPWR.n0 9.3005
R12 KAPWR.n6 KAPWR.n5 6.4005
R13 KAPWR.n7 KAPWR.n6 5.98311
R14 KAPWR.n5 KAPWR.n1 4.38311
R15 KAPWR.n4 KAPWR.n3 3.44285
R16 KAPWR.n3 KAPWR.n1 2.1691
R17 KAPWR.n2 KAPWR.n1 1.85174
R18 KAPWR.n4 KAPWR.n0 0.221654
R19 KAPWR.n8 KAPWR.n0 0.221654
R20 KAPWR KAPWR.n8 0.03175
R21 VPB VPB.t0 730.997
R22 VNB VNB.t0 3517.15
C0 VPB KAPWR 0.04586f
C1 VGND KAPWR 0.88823f
C2 VPB VPWR 0.042629f
C3 VGND VPWR 0.042169f
C4 KAPWR VPWR 0.555378f
C5 VPB VGND 0.161001f
C6 VPWR VNB 0.278668f
C7 KAPWR VNB 0.597928f
C8 VGND VNB 0.766353f
C9 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso0n_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso0n_1 VPWR VGND X SLEEP_B A VPB VNB
X0 VPWR.t1 SLEEP_B.t0 a_59_75.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X.t0 a_59_75.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND.t1 SLEEP_B.t1 a_145_75.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75.t1 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X.t1 a_59_75.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75.t1 A.t1 a_59_75.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
R0 SLEEP_B.n0 SLEEP_B.t0 261.887
R1 SLEEP_B SLEEP_B.n0 156.864
R2 SLEEP_B.n0 SLEEP_B.t1 155.847
R3 a_59_75.n2 a_59_75.n1 672.948
R4 a_59_75.n1 a_59_75.t2 314.563
R5 a_59_75.n0 a_59_75.t3 236.18
R6 a_59_75.n0 a_59_75.t4 163.881
R7 a_59_75.n1 a_59_75.n0 152
R8 a_59_75.t0 a_59_75.n2 63.3219
R9 a_59_75.n2 a_59_75.t1 63.3219
R10 VPWR.n1 VPWR.t2 682.442
R11 VPWR.n1 VPWR.n0 331.682
R12 VPWR.n0 VPWR.t1 116.341
R13 VPWR.n0 VPWR.t0 28.4453
R14 VPWR VPWR.n1 0.401673
R15 VPB.t1 VPB.t0 319.627
R16 VPB VPB.t2 298.911
R17 VPB.t2 VPB.t1 248.599
R18 X.n0 X 590.984
R19 X.n1 X.n0 585
R20 X X.t1 269.426
R21 X.n0 X.t0 46.2955
R22 X X.n3 11.2645
R23 X X.n2 6.6565
R24 X.n3 X 6.1445
R25 X.n3 X 4.63498
R26 X.n2 X 3.61789
R27 X.n1 X 3.47876
R28 X.n2 X.n1 2.36572
R29 a_145_75.t0 a_145_75.t1 77.1434
R30 VGND VGND.n0 212.421
R31 VGND.n0 VGND.t1 72.8576
R32 VGND.n0 VGND.t0 22.3257
R33 VNB.t1 VNB.t0 1537.86
R34 VNB VNB.t2 1438.19
R35 VNB.t2 VNB.t1 1196.12
R36 A.n0 A.t0 256.07
R37 A.n1 A.n0 152
R38 A.n0 A.t1 150.03
R39 A A.n1 9.22489
R40 A.n1 A 7.6805
C0 VPWR SLEEP_B 0.011747f
C1 X VGND 0.099328f
C2 A SLEEP_B 0.097088f
C3 VGND VPB 0.007995f
C4 VGND VPWR 0.046078f
C5 VGND A 0.014715f
C6 X VPB 0.012653f
C7 VGND SLEEP_B 0.011461f
C8 X VPWR 0.111215f
C9 X A 1.68e-19
C10 X SLEEP_B 0.002761f
C11 VPB VPWR 0.072934f
C12 VPB A 0.080573f
C13 VPB SLEEP_B 0.06287f
C14 VPWR A 0.036234f
C15 VGND VNB 0.311398f
C16 X VNB 0.100184f
C17 SLEEP_B VNB 0.112872f
C18 A VNB 0.173792f
C19 VPWR VNB 0.273451f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_12 VGND VPWR KAPWR VPB VNB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
R0 VGND.n6 VGND.t2 538.312
R1 VGND.n4 VGND.t0 219.992
R2 VGND.n16 VGND.n15 214.956
R3 VGND.n17 VGND.t1 214.456
R4 VGND.n6 VGND.n5 152
R5 VGND.n8 VGND.n7 152
R6 VGND.n15 VGND.n14 152
R7 VGND.t2 VGND.n2 68.6994
R8 VGND.n7 VGND.n6 62.9556
R9 VGND.n7 VGND.n2 31.4781
R10 VGND.n15 VGND.n2 31.4781
R11 VGND.n18 VGND.n17 9.56351
R12 VGND.n1 VGND.n0 9.3005
R13 VGND.n13 VGND.n12 9.3005
R14 VGND.n11 VGND.n3 9.3005
R15 VGND.n10 VGND.n9 9.3005
R16 VGND.n5 VGND.n4 5.29077
R17 VGND.n13 VGND.n1 4.03338
R18 VGND.n9 VGND.n5 3.59502
R19 VGND.n14 VGND.n3 3.59502
R20 VGND.n17 VGND.n16 2.63064
R21 VGND.n9 VGND.n8 2.01694
R22 VGND.n8 VGND.n3 2.01694
R23 VGND.n16 VGND.n1 1.14023
R24 VGND.n14 VGND.n13 0.438856
R25 VGND.n10 VGND.n4 0.283314
R26 VGND.n11 VGND.n10 0.120292
R27 VGND.n12 VGND.n11 0.120292
R28 VGND.n12 VGND.n0 0.120292
R29 VGND.n18 VGND.n0 0.120292
R30 VGND VGND.n18 0.0226354
R31 KAPWR.n15 KAPWR.t2 571.745
R32 KAPWR.n29 KAPWR.t1 388.656
R33 KAPWR.n8 KAPWR.t0 388.656
R34 KAPWR.n13 KAPWR.n6 214.956
R35 KAPWR.n15 KAPWR.n3 152
R36 KAPWR.n17 KAPWR.n16 152
R37 KAPWR.n13 KAPWR.n12 152
R38 KAPWR.t2 KAPWR.n14 107.793
R39 KAPWR.n16 KAPWR.n15 62.9556
R40 KAPWR.n16 KAPWR.n14 32.4617
R41 KAPWR.n14 KAPWR.n13 30.4944
R42 KAPWR.n9 KAPWR.n8 9.78832
R43 KAPWR.n30 KAPWR.n29 9.71789
R44 KAPWR.n9 KAPWR.n7 9.3005
R45 KAPWR.n11 KAPWR.n10 9.3005
R46 KAPWR.n5 KAPWR.n4 9.3005
R47 KAPWR.n19 KAPWR.n18 9.3005
R48 KAPWR.n21 KAPWR.n20 9.3005
R49 KAPWR.n22 KAPWR.n2 9.3005
R50 KAPWR.n24 KAPWR.n23 9.3005
R51 KAPWR.n25 KAPWR.n1 9.3005
R52 KAPWR.n27 KAPWR.n26 9.3005
R53 KAPWR.n28 KAPWR.n0 9.3005
R54 KAPWR.n23 KAPWR.n22 6.4005
R55 KAPWR.n23 KAPWR.n1 6.4005
R56 KAPWR.n27 KAPWR.n1 6.4005
R57 KAPWR.n28 KAPWR.n27 6.4005
R58 KAPWR.n29 KAPWR.n28 5.98311
R59 KAPWR.n22 KAPWR.n21 5.62176
R60 KAPWR.n11 KAPWR.n7 4.08939
R61 KAPWR.n18 KAPWR.n3 3.82272
R62 KAPWR.n12 KAPWR.n5 3.46717
R63 KAPWR.n8 KAPWR.n6 2.84494
R64 KAPWR.n17 KAPWR.n5 2.22272
R65 KAPWR.n18 KAPWR.n17 1.86717
R66 KAPWR.n7 KAPWR.n6 0.978278
R67 KAPWR.n12 KAPWR.n11 0.622722
R68 KAPWR.n21 KAPWR.n3 0.267167
R69 KAPWR.n10 KAPWR.n9 0.221654
R70 KAPWR.n10 KAPWR.n4 0.221654
R71 KAPWR.n19 KAPWR.n4 0.221654
R72 KAPWR.n20 KAPWR.n19 0.221654
R73 KAPWR.n20 KAPWR.n2 0.221654
R74 KAPWR.n24 KAPWR.n2 0.221654
R75 KAPWR.n25 KAPWR.n24 0.221654
R76 KAPWR.n26 KAPWR.n25 0.221654
R77 KAPWR.n26 KAPWR.n0 0.221654
R78 KAPWR.n30 KAPWR.n0 0.221654
R79 KAPWR KAPWR.n30 0.03175
R80 VPB VPB.t0 1547.82
R81 VNB VNB.t0 7447.25
C0 VGND KAPWR 1.97765f
C1 VPWR VPB 0.073134f
C2 VPWR VGND 0.093539f
C3 VPWR KAPWR 1.1426f
C4 VPB VGND 0.336357f
C5 VPB KAPWR 0.072947f
C6 VPWR VNB 0.505511f
C7 KAPWR VNB 1.19099f
C8 VGND VNB 1.46641f
C9 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_8 VPWR VGND KAPWR VPB VNB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
R0 VGND.n4 VGND.t0 219.518
R1 VGND.n10 VGND.t1 214.456
R2 VGND.n9 VGND.n8 200.692
R3 VGND.n3 VGND.n2 190.399
R4 VGND.n8 VGND.n7 152
R5 VGND.n2 VGND.t2 34.2973
R6 VGND.n11 VGND.n10 9.56351
R7 VGND.n1 VGND.n0 9.3005
R8 VGND.n6 VGND.n5 9.3005
R9 VGND.n4 VGND.n3 5.14426
R10 VGND.n8 VGND.n2 4.85762
R11 VGND.n6 VGND.n3 3.50735
R12 VGND.n7 VGND.n1 3.2005
R13 VGND.n10 VGND.n9 2.63064
R14 VGND.n9 VGND.n1 1.14023
R15 VGND.n7 VGND.n6 0.833377
R16 VGND.n5 VGND.n4 0.53311
R17 VGND.n5 VGND.n0 0.120292
R18 VGND.n11 VGND.n0 0.120292
R19 VGND VGND.n11 0.0226354
R20 KAPWR.n18 KAPWR.t1 388.656
R21 KAPWR.n5 KAPWR.t0 388.656
R22 KAPWR.n9 KAPWR.n4 202.66
R23 KAPWR.n11 KAPWR.n10 190.165
R24 KAPWR.n9 KAPWR.n8 152
R25 KAPWR.n10 KAPWR.t2 50.5057
R26 KAPWR.n6 KAPWR.n5 9.78832
R27 KAPWR.n19 KAPWR.n18 9.71789
R28 KAPWR.n7 KAPWR.n6 9.3005
R29 KAPWR.n3 KAPWR.n2 9.3005
R30 KAPWR.n13 KAPWR.n12 9.3005
R31 KAPWR.n14 KAPWR.n1 9.3005
R32 KAPWR.n16 KAPWR.n15 9.3005
R33 KAPWR.n17 KAPWR.n0 9.3005
R34 KAPWR.n10 KAPWR.n9 7.11866
R35 KAPWR.n16 KAPWR.n1 6.4005
R36 KAPWR.n17 KAPWR.n16 6.4005
R37 KAPWR.n18 KAPWR.n17 5.98311
R38 KAPWR.n12 KAPWR.n1 5.57151
R39 KAPWR.n11 KAPWR.n3 3.91161
R40 KAPWR.n8 KAPWR.n7 3.42272
R41 KAPWR.n5 KAPWR.n4 2.66717
R42 KAPWR.n7 KAPWR.n4 1.15606
R43 KAPWR.n8 KAPWR.n3 0.667167
R44 KAPWR.n6 KAPWR.n2 0.221654
R45 KAPWR.n13 KAPWR.n2 0.221654
R46 KAPWR.n14 KAPWR.n13 0.221654
R47 KAPWR.n15 KAPWR.n14 0.221654
R48 KAPWR.n15 KAPWR.n0 0.221654
R49 KAPWR.n19 KAPWR.n0 0.221654
R50 KAPWR.n12 KAPWR.n11 0.178278
R51 KAPWR KAPWR.n19 0.03175
R52 VPB VPB.t0 1003.27
R53 VNB VNB.t0 4827.18
C0 KAPWR VPB 0.055151f
C1 VPWR VPB 0.052767f
C2 KAPWR VGND 1.25219f
C3 VPWR VGND 0.059275f
C4 KAPWR VPWR 0.751273f
C5 VPB VGND 0.219439f
C6 VPWR VNB 0.354269f
C7 KAPWR VNB 0.796151f
C8 VGND VNB 0.998917f
C9 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputisolatch_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputisolatch_1 VGND VPWR VPB VNB SLEEP_B Q D
X0 a_381_369.t0 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_575_47.t1 a_27_47.t2 a_476_47.t3 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0486 pd=0.63 as=0.0621 ps=0.705 w=0.36 l=0.15
X2 a_476_47.t2 a_27_47.t3 a_381_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X3 a_476_47.t0 a_193_47.t2 a_381_47.t1 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.066 ps=0.745 w=0.36 l=0.15
X4 VGND.t4 a_629_21.t2 a_575_47.t0 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0936 pd=1.24 as=0.0486 ps=0.63 w=0.36 l=0.15
X5 Q.t0 a_476_47.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_193_47.t1 a_27_47.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.62 as=0.07425 ps=0.82 w=0.55 l=0.15
X7 a_193_47.t0 a_27_47.t5 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR.t5 a_629_21.t3 a_560_413.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.07245 ps=0.765 w=0.42 l=0.15
X9 VGND.t2 a_476_47.t5 a_629_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 Q.t1 a_476_47.t6 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR.t4 a_476_47.t7 a_629_21.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_381_47.t0 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 VPWR.t2 SLEEP_B.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.07425 pd=0.82 as=0.143 ps=1.62 w=0.55 l=0.15
X14 a_560_413.t1 a_193_47.t3 a_476_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND.t3 SLEEP_B.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 373.283
R1 D D.n0 155.244
R2 D.n0 D.t1 127.284
R3 VPWR.n2 VPWR.t0 717.596
R4 VPWR.n4 VPWR.t5 678.236
R5 VPWR.n15 VPWR.n1 604.394
R6 VPWR.n6 VPWR.n5 332.916
R7 VPWR.n1 VPWR.t1 48.355
R8 VPWR.n1 VPWR.t2 48.355
R9 VPWR.n9 VPWR.n8 34.6358
R10 VPWR.n10 VPWR.n9 34.6358
R11 VPWR.n8 VPWR.n4 33.8829
R12 VPWR.n5 VPWR.t3 26.5955
R13 VPWR.n5 VPWR.t4 26.5955
R14 VPWR.n14 VPWR.n13 26.5725
R15 VPWR.n15 VPWR.n14 22.9652
R16 VPWR.n10 VPWR.n2 21.9179
R17 VPWR.n8 VPWR.n7 9.3005
R18 VPWR.n9 VPWR.n3 9.3005
R19 VPWR.n11 VPWR.n10 9.3005
R20 VPWR.n13 VPWR.n12 9.3005
R21 VPWR.n14 VPWR.n0 9.3005
R22 VPWR.n6 VPWR.n4 8.11084
R23 VPWR.n16 VPWR.n15 7.12063
R24 VPWR.n7 VPWR.n6 0.390468
R25 VPWR.n13 VPWR.n2 0.233227
R26 VPWR.n16 VPWR.n0 0.148519
R27 VPWR.n7 VPWR.n3 0.120292
R28 VPWR.n11 VPWR.n3 0.120292
R29 VPWR.n12 VPWR.n11 0.120292
R30 VPWR.n12 VPWR.n0 0.120292
R31 VPWR VPWR.n16 0.114842
R32 a_381_369.t0 a_381_369.t1 132.286
R33 VPB.t7 VPB.t6 562.306
R34 VPB.t2 VPB.t0 556.386
R35 VPB.t3 VPB.t7 292.991
R36 VPB.t0 VPB.t1 281.154
R37 VPB.t6 VPB.t5 248.599
R38 VPB.t1 VPB.t3 248.599
R39 VPB.t4 VPB.t2 248.599
R40 VPB VPB.t4 142.056
R41 a_27_47.t1 a_27_47.n3 717.703
R42 a_27_47.n1 a_27_47.n0 432.644
R43 a_27_47.n0 a_27_47.t2 425.945
R44 a_27_47.n3 a_27_47.t0 300.767
R45 a_27_47.n2 a_27_47.t5 273.134
R46 a_27_47.n1 a_27_47.t4 245.821
R47 a_27_47.n0 a_27_47.t3 219.042
R48 a_27_47.n3 a_27_47.n2 165.145
R49 a_27_47.n2 a_27_47.n1 38.5605
R50 a_476_47.n4 a_476_47.n3 722.672
R51 a_476_47.n3 a_476_47.n2 280.625
R52 a_476_47.n3 a_476_47.n1 243.968
R53 a_476_47.n0 a_476_47.t6 212.081
R54 a_476_47.n1 a_476_47.t7 212.081
R55 a_476_47.n0 a_476_47.t4 139.78
R56 a_476_47.n1 a_476_47.t5 139.78
R57 a_476_47.n2 a_476_47.t0 68.3338
R58 a_476_47.t1 a_476_47.n4 63.3219
R59 a_476_47.n4 a_476_47.t2 63.3219
R60 a_476_47.n1 a_476_47.n0 61.346
R61 a_476_47.n2 a_476_47.t3 46.6672
R62 a_575_47.t0 a_575_47.t1 90.0005
R63 VNB.t4 VNB.t1 2705.5
R64 VNB.t6 VNB.t0 2677.02
R65 VNB.t5 VNB.t7 1409.71
R66 VNB.t0 VNB.t5 1352.75
R67 VNB.t1 VNB.t2 1196.12
R68 VNB.t7 VNB.t4 1196.12
R69 VNB.t3 VNB.t6 1196.12
R70 VNB VNB.t3 683.495
R71 a_193_47.t1 a_193_47.n1 646.532
R72 a_193_47.n1 a_193_47.t0 333.841
R73 a_193_47.n0 a_193_47.t2 328.108
R74 a_193_47.n0 a_193_47.t3 300.252
R75 a_193_47.n1 a_193_47.n0 109.177
R76 a_381_47.n0 a_381_47.t1 66.6672
R77 a_381_47.n0 a_381_47.t0 26.3935
R78 a_381_47.n1 a_381_47.n0 14.4005
R79 a_629_21.t1 a_629_21.n0 393.961
R80 a_629_21.n1 a_629_21.t2 375.961
R81 a_629_21.n0 a_629_21.t0 277.123
R82 a_629_21.n0 a_629_21.n1 170.424
R83 a_629_21.n1 a_629_21.t3 147.814
R84 VGND.n5 VGND.t4 247.262
R85 VGND.n11 VGND.t0 238.311
R86 VGND.n4 VGND.n3 226.88
R87 VGND.n14 VGND.n13 199.739
R88 VGND.n13 VGND.t5 38.5719
R89 VGND.n13 VGND.t3 38.5719
R90 VGND.n7 VGND.n6 34.6358
R91 VGND.n7 VGND.n1 34.6358
R92 VGND.n3 VGND.t1 24.9236
R93 VGND.n3 VGND.t2 24.9236
R94 VGND.n12 VGND.n11 22.9652
R95 VGND.n14 VGND.n12 22.9652
R96 VGND.n11 VGND.n1 21.4593
R97 VGND.n6 VGND.n5 20.7064
R98 VGND.n6 VGND.n2 9.3005
R99 VGND.n8 VGND.n7 9.3005
R100 VGND.n9 VGND.n1 9.3005
R101 VGND.n11 VGND.n10 9.3005
R102 VGND.n12 VGND.n0 9.3005
R103 VGND.n15 VGND.n14 7.12063
R104 VGND.n5 VGND.n4 6.83752
R105 VGND.n4 VGND.n2 0.462689
R106 VGND.n15 VGND.n0 0.148519
R107 VGND.n8 VGND.n2 0.120292
R108 VGND.n9 VGND.n8 0.120292
R109 VGND.n10 VGND.n9 0.120292
R110 VGND.n10 VGND.n0 0.120292
R111 VGND VGND.n15 0.114842
R112 Q.n0 Q.t1 374.774
R113 Q.n1 Q.t0 209.923
R114 Q Q.n1 82.223
R115 Q Q.n0 8.17402
R116 Q.n0 Q 6.98766
R117 Q.n1 Q 6.9619
R118 a_560_413.t0 a_560_413.t1 161.821
R119 SLEEP_B.n0 SLEEP_B.t0 284.916
R120 SLEEP_B.n0 SLEEP_B.t1 235.109
R121 SLEEP_B SLEEP_B.n0 154.101
C0 VPB VPWR 0.122469f
C1 VPB VGND 0.014191f
C2 SLEEP_B VPWR 0.019063f
C3 SLEEP_B VGND 0.018836f
C4 VPB Q 0.011685f
C5 D VPWR 0.014418f
C6 D VGND 0.033288f
C7 VPWR VGND 0.109434f
C8 VPWR Q 0.102729f
C9 VGND Q 0.052705f
C10 VPB SLEEP_B 0.075689f
C11 VPB D 0.048998f
C12 Q VNB 0.084805f
C13 VGND VNB 0.617039f
C14 VPWR VNB 0.489488f
C15 D VNB 0.127168f
C16 SLEEP_B VNB 0.197909f
C17 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso1p_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso1p_1 VPB VNB VGND VPWR X SLEEP A
X0 VGND.t1 SLEEP.t0 a_68_297.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X.t1 a_68_297.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR.t0 SLEEP.t1 a_150_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X.t0 a_68_297.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297.t0 A.t1 a_68_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 SLEEP.n0 SLEEP.t0 206.19
R1 SLEEP SLEEP.n0 154.657
R2 SLEEP.n0 SLEEP.t1 148.35
R3 a_68_297.n1 a_68_297.t1 662.71
R4 a_68_297.n2 a_68_297.n1 260.308
R5 a_68_297.n1 a_68_297.n0 241.601
R6 a_68_297.n0 a_68_297.t4 236.18
R7 a_68_297.n0 a_68_297.t3 163.881
R8 a_68_297.n2 a_68_297.t2 38.5719
R9 a_68_297.t0 a_68_297.n2 38.5719
R10 VGND.n1 VGND.t0 253.421
R11 VGND.n1 VGND.n0 217.375
R12 VGND.n0 VGND.t1 55.7148
R13 VGND.n0 VGND.t2 26.8576
R14 VGND VGND.n1 0.437652
R15 VNB.t1 VNB.t2 1381.23
R16 VNB VNB.t0 1338.51
R17 VNB.t0 VNB.t1 1196.12
R18 A.n0 A.t0 192.639
R19 A A.n0 158.172
R20 A.n0 A.t1 134.799
R21 X.n0 X.t0 340.584
R22 X X.t1 174.464
R23 X.n0 X 2.4386
R24 X X.n0 1.43601
R25 a_150_297.t0 a_150_297.t1 98.5005
R26 VPWR VPWR.n0 320.877
R27 VPWR.n0 VPWR.t0 96.1553
R28 VPWR.n0 VPWR.t1 25.6105
R29 VPB VPB.t0 313.707
R30 VPB.t1 VPB.t2 287.072
R31 VPB.t0 VPB.t1 213.084
C0 VPWR X 0.128567f
C1 A SLEEP 0.07509f
C2 A X 1.65e-19
C3 VPWR VGND 0.046447f
C4 A VGND 0.043653f
C5 SLEEP X 0.013051f
C6 SLEEP VGND 0.034653f
C7 X VGND 0.113947f
C8 VPB VPWR 0.080528f
C9 VPB A 0.046202f
C10 VPB SLEEP 0.030968f
C11 VPB X 0.020902f
C12 VPWR A 0.008552f
C13 VPB VGND 0.011204f
C14 VPWR SLEEP 0.008464f
C15 VGND VNB 0.320425f
C16 X VNB 0.100952f
C17 SLEEP VNB 0.110717f
C18 A VNB 0.182719f
C19 VPWR VNB 0.268565f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso1n_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso1n_1 VGND VPWR VNB VPB A X SLEEP_B
X0 a_219_297.t0 a_27_53.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X1 VGND.t3 SLEEP_B.t0 a_27_53.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t0 A.t0 a_301_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X.t0 a_219_297.t3 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_301_297.t1 a_27_53.t3 a_219_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X.t1 a_219_297.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6 a_27_53.t1 SLEEP_B.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND.t2 A.t1 a_219_297.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 a_27_53.n1 a_27_53.t1 672.086
R1 a_27_53.t0 a_27_53.n1 261.192
R2 a_27_53.n0 a_27_53.t2 186.03
R3 a_27_53.n1 a_27_53.n0 171.394
R4 a_27_53.n0 a_27_53.t3 137.829
R5 VGND.n3 VGND.n2 202.195
R6 VGND.n7 VGND.n6 185
R7 VGND.n9 VGND.n8 185
R8 VGND.n8 VGND.n7 137.143
R9 VGND.n2 VGND.t2 52.8576
R10 VGND.n7 VGND.t0 38.5719
R11 VGND.n8 VGND.t3 38.5719
R12 VGND.n10 VGND.n9 38.1787
R13 VGND.n6 VGND.n3 29.3949
R14 VGND.n2 VGND.t1 27.5691
R15 VGND.n1 VGND.n0 9.3005
R16 VGND.n5 VGND.n4 9.3005
R17 VGND.n5 VGND.n1 9.05896
R18 VGND.n4 VGND.n3 2.16256
R19 VGND.n6 VGND.n5 0.197423
R20 VGND.n9 VGND.n1 0.197423
R21 VGND.n4 VGND.n0 0.120292
R22 VGND.n10 VGND.n0 0.120292
R23 VGND VGND.n10 0.0213333
R24 a_219_297.n1 a_219_297.t1 731.812
R25 a_219_297.n2 a_219_297.n1 263.83
R26 a_219_297.n0 a_219_297.t4 240.484
R27 a_219_297.n0 a_219_297.t3 168.185
R28 a_219_297.n1 a_219_297.n0 152
R29 a_219_297.n2 a_219_297.t2 38.5719
R30 a_219_297.t0 a_219_297.n2 38.5719
R31 VNB.t3 VNB.t1 2563.11
R32 VNB.t2 VNB.t0 1395.47
R33 VNB.t1 VNB.t2 1196.12
R34 VNB VNB.t3 911.327
R35 SLEEP_B.n0 SLEEP_B.t0 185.376
R36 SLEEP_B SLEEP_B.n0 157.632
R37 SLEEP_B.n0 SLEEP_B.t1 137.177
R38 A A.t0 563.896
R39 A.t0 A.t1 392.027
R40 a_301_297.t0 a_301_297.t1 98.5005
R41 VPWR.n1 VPWR.t2 708.777
R42 VPWR.n1 VPWR.n0 321.704
R43 VPWR.n0 VPWR.t0 96.1553
R44 VPWR.n0 VPWR.t1 26.5955
R45 VPWR VPWR.n1 0.065704
R46 VPB.t3 VPB.t2 568.225
R47 VPB.t0 VPB.t1 290.031
R48 VPB.t2 VPB.t0 213.084
R49 VPB VPB.t3 189.409
R50 X X.t1 360.769
R51 X X.t0 287.072
C0 X VPWR 0.087835f
C1 SLEEP_B A 2.16e-19
C2 VGND VPB 0.009103f
C3 VPWR A 0.194142f
C4 SLEEP_B VGND 0.0173f
C5 X A 0.002526f
C6 VGND VPWR 0.057039f
C7 X VGND 0.035406f
C8 VGND A 0.01651f
C9 SLEEP_B VPB 0.046613f
C10 VPB VPWR 0.097059f
C11 X VPB 0.010908f
C12 SLEEP_B VPWR 0.037442f
C13 VPB A 0.160525f
C14 VGND VNB 0.353111f
C15 X VNB 0.08883f
C16 SLEEP_B VNB 0.169579f
C17 A VNB 0.135517f
C18 VPWR VNB 0.324987f
C19 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso0p_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso0p_1 X SLEEP A VGND VPWR VPB VNB
X0 VPWR.t1 A.t0 a_207_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X.t1 a_207_413.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47.t1 a_27_413.t2 a_207_413.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X.t0 a_207_413.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413.t2 a_27_413.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR.t0 SLEEP.t0 a_27_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND.t0 A.t1 a_297_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413.t1 SLEEP.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A.n0 A.t1 293.969
R1 A.n1 A.n0 152
R2 A.n0 A.t0 138.338
R3 A A.n1 14.0392
R4 A.n1 A 4.95534
R5 a_207_413.n2 a_207_413.n1 625.684
R6 a_207_413.n1 a_207_413.t1 262.252
R7 a_207_413.n0 a_207_413.t3 240.484
R8 a_207_413.n1 a_207_413.n0 174.924
R9 a_207_413.n0 a_207_413.t4 166.692
R10 a_207_413.t0 a_207_413.n2 68.0124
R11 a_207_413.n2 a_207_413.t2 68.0124
R12 VPWR.n9 VPWR.n1 602.456
R13 VPWR.n3 VPWR.n2 585
R14 VPWR.n5 VPWR.n4 585
R15 VPWR.n4 VPWR.n3 159.476
R16 VPWR.n1 VPWR.t3 96.1553
R17 VPWR.n3 VPWR.t1 86.7743
R18 VPWR.n4 VPWR.t2 66.8398
R19 VPWR.n1 VPWR.t0 63.3219
R20 VPWR.n8 VPWR.n7 27.724
R21 VPWR.n9 VPWR.n8 22.9652
R22 VPWR.n7 VPWR.n6 9.3005
R23 VPWR.n8 VPWR.n0 9.3005
R24 VPWR.n6 VPWR.n5 9.01185
R25 VPWR.n10 VPWR.n9 7.12063
R26 VPWR.n5 VPWR.n2 6.8005
R27 VPWR.n7 VPWR.n2 1.0005
R28 VPWR.n10 VPWR.n0 0.148519
R29 VPWR.n6 VPWR.n0 0.120292
R30 VPWR VPWR.n10 0.114842
R31 VPB.t1 VPB.t2 526.792
R32 VPB.t0 VPB.t3 290.031
R33 VPB.t3 VPB.t1 260.437
R34 VPB VPB.t0 192.369
R35 X.n1 X.t1 358.94
R36 X.n0 X.t0 209.923
R37 X X.n0 79.4838
R38 X.n1 X 7.91583
R39 X.n0 X 6.66717
R40 X X.n1 6.2537
R41 a_27_413.t0 a_27_413.n1 725.558
R42 a_27_413.n0 a_27_413.t3 381.656
R43 a_27_413.n1 a_27_413.t1 243.694
R44 a_27_413.n0 a_27_413.t2 197.62
R45 a_27_413.n1 a_27_413.n0 164.994
R46 a_297_47.t0 a_297_47.t1 68.5719
R47 VNB.t3 VNB.t2 2677.02
R48 VNB.t0 VNB.t1 1395.47
R49 VNB.t2 VNB.t0 1110.68
R50 VNB VNB.t3 925.567
R51 VGND.n1 VGND.t2 247.484
R52 VGND.n1 VGND.n0 206.194
R53 VGND.n0 VGND.t0 58.5719
R54 VGND.n0 VGND.t1 25.4291
R55 VGND VGND.n1 0.0759566
R56 SLEEP.n0 SLEEP.t0 327.99
R57 SLEEP.n0 SLEEP.t1 199.457
R58 SLEEP.n1 SLEEP.n0 152
R59 SLEEP.n1 SLEEP 12.1605
R60 SLEEP SLEEP.n1 2.34717
C0 VGND SLEEP 0.047311f
C1 X A 0.030307f
C2 A VPWR 0.086692f
C3 X VPWR 0.055194f
C4 VGND A 0.01869f
C5 X VGND 0.065151f
C6 VGND VPWR 0.056424f
C7 VPB SLEEP 0.080056f
C8 VPB A 0.111061f
C9 X VPB 0.012221f
C10 VPB VPWR 0.063352f
C11 VGND VPB 0.007626f
C12 SLEEP VPWR 0.018219f
C13 VGND VNB 0.368472f
C14 X VNB 0.089221f
C15 VPWR VNB 0.291542f
C16 A VNB 0.132317f
C17 SLEEP VNB 0.201458f
C18 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_4 VNB VPB VGND VPWR X A SLEEP
X0 VPWR.t4 SLEEP.t0 a_27_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t3 SLEEP.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t2 SLEEP.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t3 SLEEP.t3 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297.t4 a_419_21.t2 X.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 X.t1 SLEEP.t4 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND.t1 SLEEP.t5 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t5 a_419_21.t3 X.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND.t6 a_419_21.t4 X.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X.t7 a_419_21.t5 a_27_297.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t2 SLEEP.t6 a_27_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 X.t8 a_419_21.t6 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t0 A.t0 a_419_21.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.182 ps=1.86 w=0.65 l=0.15
X13 X.t9 a_419_21.t7 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t0 A.t1 a_419_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.27 ps=2.54 w=1 l=0.15
X15 a_27_297.t6 a_419_21.t8 X.t10 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X.t11 a_419_21.t9 a_27_297.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297.t0 SLEEP.t7 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 SLEEP.n2 SLEEP.t7 212.081
R1 SLEEP.n1 SLEEP.t0 212.081
R2 SLEEP.n7 SLEEP.t2 212.081
R3 SLEEP.n8 SLEEP.t6 212.081
R4 SLEEP.n4 SLEEP.n3 173.761
R5 SLEEP SLEEP.n9 152.641
R6 SLEEP.n5 SLEEP.n4 152
R7 SLEEP.n6 SLEEP.n0 152
R8 SLEEP.n2 SLEEP.t5 139.78
R9 SLEEP.n1 SLEEP.t1 139.78
R10 SLEEP.n7 SLEEP.t3 139.78
R11 SLEEP.n8 SLEEP.t4 139.78
R12 SLEEP.n6 SLEEP.n5 49.6611
R13 SLEEP.n9 SLEEP.n7 45.2793
R14 SLEEP.n3 SLEEP.n1 42.3581
R15 SLEEP.n4 SLEEP.n0 21.7605
R16 SLEEP SLEEP.n0 21.1205
R17 SLEEP.n3 SLEEP.n2 18.9884
R18 SLEEP.n9 SLEEP.n8 16.0672
R19 SLEEP.n5 SLEEP.n1 7.30353
R20 SLEEP.n7 SLEEP.n6 4.38232
R21 a_27_297.n1 a_27_297.n0 296.538
R22 a_27_297.n3 a_27_297.t1 278.786
R23 a_27_297.n1 a_27_297.t4 267.592
R24 a_27_297.n3 a_27_297.n2 207.26
R25 a_27_297.n5 a_27_297.n4 188.952
R26 a_27_297.n4 a_27_297.n3 57.3598
R27 a_27_297.n4 a_27_297.n1 53.3404
R28 a_27_297.n2 a_27_297.t3 26.5955
R29 a_27_297.n2 a_27_297.t2 26.5955
R30 a_27_297.n0 a_27_297.t5 26.5955
R31 a_27_297.n0 a_27_297.t6 26.5955
R32 a_27_297.n5 a_27_297.t7 26.5955
R33 a_27_297.t0 a_27_297.n5 26.5955
R34 VPWR.n4 VPWR.n3 316.245
R35 VPWR.n6 VPWR.n1 310.5
R36 VPWR.n2 VPWR.t0 246.484
R37 VPWR.n1 VPWR.t3 26.5955
R38 VPWR.n1 VPWR.t2 26.5955
R39 VPWR.n3 VPWR.t1 26.5955
R40 VPWR.n3 VPWR.t4 26.5955
R41 VPWR.n6 VPWR.n5 21.4593
R42 VPWR.n5 VPWR.n4 16.9417
R43 VPWR.n5 VPWR.n0 9.3005
R44 VPWR.n4 VPWR.n2 7.56304
R45 VPWR.n7 VPWR.n6 7.1994
R46 VPWR.n2 VPWR.n0 0.147879
R47 VPWR.n7 VPWR.n0 0.147518
R48 VPWR VPWR.n7 0.114555
R49 VPB.t5 VPB.t0 574.144
R50 VPB.t6 VPB.t5 248.599
R51 VPB.t7 VPB.t6 248.599
R52 VPB.t8 VPB.t7 248.599
R53 VPB.t1 VPB.t8 248.599
R54 VPB.t4 VPB.t1 248.599
R55 VPB.t3 VPB.t4 248.599
R56 VPB.t2 VPB.t3 248.599
R57 VPB VPB.t2 201.246
R58 VGND.n11 VGND.n4 207.965
R59 VGND.n14 VGND.n13 207.965
R60 VGND.n20 VGND.n1 207.965
R61 VGND.n7 VGND.t0 157.48
R62 VGND.n6 VGND.t6 152.594
R63 VGND.n22 VGND.t2 150.53
R64 VGND.n10 VGND.n5 34.6358
R65 VGND.n15 VGND.n12 34.6358
R66 VGND.n19 VGND.n2 34.6358
R67 VGND.n21 VGND.n20 32.377
R68 VGND.n14 VGND.n2 26.3534
R69 VGND.n4 VGND.t8 24.9236
R70 VGND.n4 VGND.t5 24.9236
R71 VGND.n13 VGND.t7 24.9236
R72 VGND.n13 VGND.t1 24.9236
R73 VGND.n1 VGND.t4 24.9236
R74 VGND.n1 VGND.t3 24.9236
R75 VGND.n22 VGND.n21 24.4711
R76 VGND.n12 VGND.n11 20.3299
R77 VGND.n11 VGND.n10 14.3064
R78 VGND.n7 VGND.n6 11.8922
R79 VGND.n23 VGND.n22 9.3005
R80 VGND.n8 VGND.n5 9.3005
R81 VGND.n10 VGND.n9 9.3005
R82 VGND.n12 VGND.n3 9.3005
R83 VGND.n16 VGND.n15 9.3005
R84 VGND.n17 VGND.n2 9.3005
R85 VGND.n19 VGND.n18 9.3005
R86 VGND.n21 VGND.n0 9.3005
R87 VGND.n15 VGND.n14 8.28285
R88 VGND.n6 VGND.n5 7.90638
R89 VGND.n20 VGND.n19 2.25932
R90 VGND.n8 VGND.n7 0.714832
R91 VGND.n9 VGND.n8 0.120292
R92 VGND.n9 VGND.n3 0.120292
R93 VGND.n16 VGND.n3 0.120292
R94 VGND.n17 VGND.n16 0.120292
R95 VGND.n18 VGND.n17 0.120292
R96 VGND.n18 VGND.n0 0.120292
R97 VGND.n23 VGND.n0 0.120292
R98 VGND VGND.n23 0.0213333
R99 X X.n0 309.719
R100 X.n9 X.n1 298.637
R101 X.n8 X.n2 141.293
R102 X.n6 X.n4 135.249
R103 X.n6 X.n5 98.982
R104 X.n7 X.n3 95.6388
R105 X.n7 X.n6 48.0005
R106 X.n9 X.n8 26.7641
R107 X.n0 X.t4 26.5955
R108 X.n0 X.t7 26.5955
R109 X.n1 X.t10 26.5955
R110 X.n1 X.t11 26.5955
R111 X.n3 X.t5 24.9236
R112 X.n3 X.t8 24.9236
R113 X.n4 X.t2 24.9236
R114 X.n4 X.t1 24.9236
R115 X.n5 X.t0 24.9236
R116 X.n5 X.t3 24.9236
R117 X.n2 X.t6 24.9236
R118 X.n2 X.t9 24.9236
R119 X X.n9 12.1605
R120 X.n8 X.n7 5.68939
R121 VNB.t6 VNB.t0 2762.46
R122 VNB.t8 VNB.t6 1196.12
R123 VNB.t5 VNB.t8 1196.12
R124 VNB.t7 VNB.t5 1196.12
R125 VNB.t1 VNB.t7 1196.12
R126 VNB.t4 VNB.t1 1196.12
R127 VNB.t3 VNB.t4 1196.12
R128 VNB.t2 VNB.t3 1196.12
R129 VNB VNB.t2 968.285
R130 a_419_21.t0 a_419_21.n8 252.549
R131 a_419_21.n6 a_419_21.t2 212.081
R132 a_419_21.n4 a_419_21.t5 212.081
R133 a_419_21.n2 a_419_21.t8 212.081
R134 a_419_21.n1 a_419_21.t9 212.081
R135 a_419_21.n3 a_419_21.n0 173.761
R136 a_419_21.n8 a_419_21.t1 153.874
R137 a_419_21.n5 a_419_21.n0 152
R138 a_419_21.n6 a_419_21.t4 139.78
R139 a_419_21.n4 a_419_21.t7 139.78
R140 a_419_21.n2 a_419_21.t3 139.78
R141 a_419_21.n1 a_419_21.t6 139.78
R142 a_419_21.n7 a_419_21.n6 112.322
R143 a_419_21.n2 a_419_21.n1 61.346
R144 a_419_21.n3 a_419_21.n2 54.0429
R145 a_419_21.n5 a_419_21.n4 42.3581
R146 a_419_21.n7 a_419_21.n0 30.5712
R147 a_419_21.n6 a_419_21.n5 18.9884
R148 a_419_21.n8 a_419_21.n7 14.5696
R149 a_419_21.n4 a_419_21.n3 7.30353
R150 A.n0 A.t1 229.754
R151 A A.n0 159.315
R152 A.n0 A.t0 157.453
C0 SLEEP VPWR 0.07913f
C1 A VPWR 0.055498f
C2 SLEEP X 0.176949f
C3 SLEEP VGND 0.067619f
C4 VPWR X 0.020844f
C5 A VGND 0.051879f
C6 SLEEP VPB 0.119415f
C7 VPWR VGND 0.102679f
C8 A VPB 0.04669f
C9 X VGND 0.544571f
C10 VPWR VPB 0.116357f
C11 X VPB 0.009206f
C12 VGND VPB 0.009839f
C13 VGND VNB 0.651371f
C14 X VNB 0.025042f
C15 VPWR VNB 0.516619f
C16 A VNB 0.150465f
C17 SLEEP VNB 0.389045f
C18 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_2 VPB VNB VGND VPWR X SLEEP A
X0 X.t5 a_251_21.t2 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t3 a_251_21.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t2 SLEEP.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 SLEEP.t1 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X.t0 SLEEP.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X5 VGND.t3 a_251_21.t4 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 SLEEP.t3 a_27_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR.t2 A.t0 a_251_21.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND.t1 A.t1 a_251_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_27_297.t0 a_251_21.t5 X.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 a_251_21.n2 a_251_21.t1 725.646
R1 a_251_21.t0 a_251_21.n2 248.954
R2 a_251_21.n1 a_251_21.t5 212.081
R3 a_251_21.n0 a_251_21.t2 212.081
R4 a_251_21.n2 a_251_21.n1 207.535
R5 a_251_21.n1 a_251_21.t4 139.78
R6 a_251_21.n0 a_251_21.t3 139.78
R7 a_251_21.n1 a_251_21.n0 61.346
R8 a_27_297.t0 a_27_297.n1 298.416
R9 a_27_297.n1 a_27_297.t3 288.245
R10 a_27_297.n1 a_27_297.n0 187.506
R11 a_27_297.n0 a_27_297.t1 26.5955
R12 a_27_297.n0 a_27_297.t2 26.5955
R13 X.n2 X.n1 337.207
R14 X X.n4 186.358
R15 X.n4 X.n3 185
R16 X.n2 X.n0 137.189
R17 X.n1 X.t4 26.5955
R18 X.n1 X.t5 26.5955
R19 X.n4 X.t2 24.9236
R20 X.n4 X.t3 24.9236
R21 X.n0 X.t1 24.9236
R22 X.n0 X.t0 24.9236
R23 X X.n3 11.8308
R24 X.n3 X.n2 3.10353
R25 VPB.t0 VPB.t2 556.386
R26 VPB.t1 VPB.t0 248.599
R27 VPB.t3 VPB.t1 248.599
R28 VPB.t4 VPB.t3 248.599
R29 VPB VPB.t4 201.246
R30 VGND.n4 VGND.t1 264.288
R31 VGND.n8 VGND.n1 207.965
R32 VGND.n3 VGND.t3 160.8
R33 VGND.n10 VGND.t0 151.194
R34 VGND.n7 VGND.n2 34.6358
R35 VGND.n9 VGND.n8 32.377
R36 VGND.n3 VGND.n2 26.3534
R37 VGND.n1 VGND.t4 24.9236
R38 VGND.n1 VGND.t2 24.9236
R39 VGND.n10 VGND.n9 24.4711
R40 VGND.n4 VGND.n3 15.4369
R41 VGND.n11 VGND.n10 9.3005
R42 VGND.n5 VGND.n2 9.3005
R43 VGND.n7 VGND.n6 9.3005
R44 VGND.n9 VGND.n0 9.3005
R45 VGND.n8 VGND.n7 2.25932
R46 VGND.n5 VGND.n4 0.572285
R47 VGND.n6 VGND.n5 0.120292
R48 VGND.n6 VGND.n0 0.120292
R49 VGND.n11 VGND.n0 0.120292
R50 VGND VGND.n11 0.0213333
R51 VNB.t3 VNB.t1 2677.02
R52 VNB.t4 VNB.t3 1196.12
R53 VNB.t2 VNB.t4 1196.12
R54 VNB.t0 VNB.t2 1196.12
R55 VNB VNB.t0 968.285
R56 SLEEP.n0 SLEEP.t0 212.081
R57 SLEEP.n1 SLEEP.t3 212.081
R58 SLEEP SLEEP.n2 153.601
R59 SLEEP.n0 SLEEP.t1 139.78
R60 SLEEP.n1 SLEEP.t2 139.78
R61 SLEEP.n2 SLEEP.n0 38.7066
R62 SLEEP.n2 SLEEP.n1 22.6399
R63 VPWR.n1 VPWR.t2 676.692
R64 VPWR.n1 VPWR.n0 322.19
R65 VPWR.n0 VPWR.t1 26.5955
R66 VPWR.n0 VPWR.t0 26.5955
R67 VPWR VPWR.n1 0.151166
R68 A.n0 A.t0 333.173
R69 A A.n0 164.708
R70 A.n0 A.t1 130.732
C0 VPB A 0.10759f
C1 VPB VPWR 0.080685f
C2 SLEEP VPWR 0.04237f
C3 VPB X 0.005224f
C4 SLEEP X 0.069669f
C5 VPB VGND 0.009577f
C6 A VPWR 0.043028f
C7 SLEEP VGND 0.033005f
C8 A X 0.00143f
C9 VPWR X 0.009649f
C10 A VGND 0.053975f
C11 VPWR VGND 0.064184f
C12 X VGND 0.281397f
C13 VPB SLEEP 0.055356f
C14 VGND VNB 0.466325f
C15 X VNB 0.016372f
C16 VPWR VNB 0.34094f
C17 A VNB 0.206554f
C18 SLEEP VNB 0.203992f
C19 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_1 VPB VNB VGND VPWR A SLEEP X
X0 X.t0 a_74_47.t2 a_265_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR.t1 A.t0 a_74_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1573 pd=1.39 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_265_297.t1 SLEEP.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.1573 ps=1.39 w=1 l=0.15
X3 X.t2 SLEEP.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VGND.t2 A.t1 a_74_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t1 a_74_47.t3 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_74_47.t0 a_74_47.n1 654.968
R1 a_74_47.n1 a_74_47.t1 302.779
R2 a_74_47.n1 a_74_47.n0 246.404
R3 a_74_47.n0 a_74_47.t2 236.18
R4 a_74_47.n0 a_74_47.t3 163.881
R5 a_265_297.t0 a_265_297.t1 41.3705
R6 X X.n0 589.914
R7 X.n2 X.n0 585
R8 X.n2 X.n1 211.56
R9 X.n0 X.t0 26.5955
R10 X.n1 X.t1 24.9236
R11 X.n1 X.t2 24.9236
R12 X X.n2 2.85764
R13 VPB VPB.t0 334.425
R14 VPB.t0 VPB.t2 319.627
R15 VPB.t2 VPB.t1 213.084
R16 A A.n0 221.946
R17 A.n0 A.t1 176.733
R18 A.n0 A.t0 119.624
R19 VPWR VPWR.n0 317.954
R20 VPWR.n0 VPWR.t1 121.953
R21 VPWR.n0 VPWR.t0 25.6105
R22 SLEEP.n0 SLEEP.t0 236.18
R23 SLEEP.n0 SLEEP.t1 163.881
R24 SLEEP SLEEP.n0 156.678
R25 VGND.n1 VGND.t1 282.298
R26 VGND.n1 VGND.n0 129.262
R27 VGND.n0 VGND.t2 57.8133
R28 VGND.n0 VGND.t0 24.7549
R29 VGND VGND.n1 0.55669
R30 VNB VNB.t2 1594.82
R31 VNB.t2 VNB.t0 1381.23
R32 VNB.t0 VNB.t1 1196.12
C0 A VGND 0.027194f
C1 X VGND 0.175424f
C2 VPB SLEEP 0.031643f
C3 VPB VPWR 0.075008f
C4 VPB A 0.061515f
C5 SLEEP VPWR 0.020882f
C6 VPB X 0.02233f
C7 SLEEP A 0.044907f
C8 VPB VGND 0.010151f
C9 VPWR A 0.012306f
C10 SLEEP X 0.019983f
C11 SLEEP VGND 0.027938f
C12 VPWR X 0.102774f
C13 VPWR VGND 0.046161f
C14 A X 0.002335f
C15 VGND VNB 0.329149f
C16 X VNB 0.085029f
C17 A VNB 0.21207f
C18 VPWR VNB 0.268516f
C19 SLEEP VNB 0.09622f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_8 VPB VNB VGND VPWR SLEEP X A
X0 X.t9 a_123_297.t4 VGND.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X.t8 a_123_297.t5 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_321_297.t8 a_123_297.t6 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X.t7 a_123_297.t7 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t6 a_123_297.t8 a_321_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_123_297.t3 A.t0 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_321_297.t6 a_123_297.t9 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t8 a_123_297.t10 X.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR.t4 a_123_297.t11 a_321_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND.t7 a_123_297.t12 X.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_123_297.t0 A.t1 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND.t6 a_123_297.t13 X.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_321_297.t4 a_123_297.t14 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t9 A.t2 a_123_297.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 X.t0 SLEEP.t0 a_321_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X.t1 SLEEP.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t2 a_123_297.t15 a_321_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_321_297.t2 a_123_297.t16 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VGND.t5 a_123_297.t17 X.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t9 A.t3 a_123_297.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR.t0 a_123_297.t18 a_321_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X.t2 a_123_297.t19 VGND.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
R0 a_123_297.n27 a_123_297.n26 230.686
R1 a_123_297.n6 a_123_297.t14 212.081
R2 a_123_297.n8 a_123_297.t15 212.081
R3 a_123_297.n4 a_123_297.t16 212.081
R4 a_123_297.n14 a_123_297.t18 212.081
R5 a_123_297.n16 a_123_297.t6 212.081
R6 a_123_297.n2 a_123_297.t8 212.081
R7 a_123_297.n22 a_123_297.t9 212.081
R8 a_123_297.n23 a_123_297.t11 212.081
R9 a_123_297.n7 a_123_297.n5 172.725
R10 a_123_297.n25 a_123_297.n24 152
R11 a_123_297.n21 a_123_297.n1 152
R12 a_123_297.n20 a_123_297.n19 152
R13 a_123_297.n18 a_123_297.n17 152
R14 a_123_297.n15 a_123_297.n3 152
R15 a_123_297.n13 a_123_297.n12 152
R16 a_123_297.n11 a_123_297.n10 152
R17 a_123_297.n9 a_123_297.n5 152
R18 a_123_297.n6 a_123_297.t13 139.78
R19 a_123_297.n8 a_123_297.t7 139.78
R20 a_123_297.n4 a_123_297.t12 139.78
R21 a_123_297.n14 a_123_297.t5 139.78
R22 a_123_297.n16 a_123_297.t10 139.78
R23 a_123_297.n2 a_123_297.t4 139.78
R24 a_123_297.n22 a_123_297.t17 139.78
R25 a_123_297.n23 a_123_297.t19 139.78
R26 a_123_297.n26 a_123_297.n0 108.678
R27 a_123_297.n26 a_123_297.n25 65.3719
R28 a_123_297.n10 a_123_297.n9 49.6611
R29 a_123_297.n21 a_123_297.n20 49.6611
R30 a_123_297.n8 a_123_297.n7 45.2793
R31 a_123_297.n24 a_123_297.n22 45.2793
R32 a_123_297.n13 a_123_297.n4 42.3581
R33 a_123_297.n17 a_123_297.n2 42.3581
R34 a_123_297.n15 a_123_297.n14 30.6732
R35 a_123_297.n16 a_123_297.n15 30.6732
R36 a_123_297.n27 a_123_297.t2 26.5955
R37 a_123_297.t0 a_123_297.n27 26.5955
R38 a_123_297.n0 a_123_297.t1 24.9236
R39 a_123_297.n0 a_123_297.t3 24.9236
R40 a_123_297.n11 a_123_297.n5 20.7243
R41 a_123_297.n12 a_123_297.n11 20.7243
R42 a_123_297.n12 a_123_297.n3 20.7243
R43 a_123_297.n18 a_123_297.n3 20.7243
R44 a_123_297.n19 a_123_297.n18 20.7243
R45 a_123_297.n19 a_123_297.n1 20.7243
R46 a_123_297.n25 a_123_297.n1 20.7243
R47 a_123_297.n14 a_123_297.n13 18.9884
R48 a_123_297.n17 a_123_297.n16 18.9884
R49 a_123_297.n7 a_123_297.n6 16.0672
R50 a_123_297.n24 a_123_297.n23 16.0672
R51 a_123_297.n10 a_123_297.n4 7.30353
R52 a_123_297.n20 a_123_297.n2 7.30353
R53 a_123_297.n9 a_123_297.n8 4.38232
R54 a_123_297.n22 a_123_297.n21 4.38232
R55 VGND.n10 VGND.n9 219.595
R56 VGND.n11 VGND.n8 207.965
R57 VGND.n6 VGND.n5 207.965
R58 VGND.n17 VGND.n4 207.965
R59 VGND.n25 VGND.t10 159.19
R60 VGND.n2 VGND.n1 60.3054
R61 VGND.n1 VGND.t4 56.3082
R62 VGND.n1 VGND.t9 56.3082
R63 VGND.n13 VGND.n12 34.6358
R64 VGND.n19 VGND.n18 34.6358
R65 VGND.n24 VGND.n23 34.6358
R66 VGND.n16 VGND.n6 33.1299
R67 VGND.n17 VGND.n16 30.1181
R68 VGND.n12 VGND.n11 27.1064
R69 VGND.n9 VGND.t0 24.9236
R70 VGND.n9 VGND.t6 24.9236
R71 VGND.n8 VGND.t1 24.9236
R72 VGND.n8 VGND.t7 24.9236
R73 VGND.n5 VGND.t2 24.9236
R74 VGND.n5 VGND.t8 24.9236
R75 VGND.n4 VGND.t3 24.9236
R76 VGND.n4 VGND.t5 24.9236
R77 VGND.n26 VGND.n25 24.7358
R78 VGND.n19 VGND.n2 17.6946
R79 VGND.n11 VGND.n10 14.4456
R80 VGND.n23 VGND.n2 13.177
R81 VGND.n12 VGND.n7 9.3005
R82 VGND.n14 VGND.n13 9.3005
R83 VGND.n16 VGND.n15 9.3005
R84 VGND.n18 VGND.n3 9.3005
R85 VGND.n20 VGND.n19 9.3005
R86 VGND.n21 VGND.n2 9.3005
R87 VGND.n23 VGND.n22 9.3005
R88 VGND.n24 VGND.n0 9.3005
R89 VGND.n18 VGND.n17 4.51815
R90 VGND.n25 VGND.n24 2.63579
R91 VGND.n13 VGND.n6 1.50638
R92 VGND.n10 VGND.n7 0.832121
R93 VGND.n14 VGND.n7 0.120292
R94 VGND.n15 VGND.n14 0.120292
R95 VGND.n15 VGND.n3 0.120292
R96 VGND.n20 VGND.n3 0.120292
R97 VGND.n21 VGND.n20 0.120292
R98 VGND.n22 VGND.n21 0.120292
R99 VGND.n22 VGND.n0 0.120292
R100 VGND.n26 VGND.n0 0.120292
R101 VGND VGND.n26 0.0226354
R102 X X.t0 463.93
R103 X X.n7 161.041
R104 X.n7 X.t1 136.792
R105 X.n2 X.n0 135.249
R106 X.n2 X.n1 98.982
R107 X.n4 X.n3 98.982
R108 X.n6 X.n5 98.982
R109 X.n4 X.n2 36.2672
R110 X.n6 X.n4 36.2672
R111 X.n7 X.n6 36.2672
R112 X.n0 X.t3 24.9236
R113 X.n0 X.t2 24.9236
R114 X.n1 X.t6 24.9236
R115 X.n1 X.t9 24.9236
R116 X.n3 X.t5 24.9236
R117 X.n3 X.t8 24.9236
R118 X.n5 X.t4 24.9236
R119 X.n5 X.t7 24.9236
R120 VNB.t9 VNB.t1 2164.4
R121 VNB VNB.t10 1808.41
R122 VNB.t3 VNB.t0 1196.12
R123 VNB.t6 VNB.t3 1196.12
R124 VNB.t4 VNB.t6 1196.12
R125 VNB.t7 VNB.t4 1196.12
R126 VNB.t5 VNB.t7 1196.12
R127 VNB.t8 VNB.t5 1196.12
R128 VNB.t2 VNB.t8 1196.12
R129 VNB.t1 VNB.t2 1196.12
R130 VNB.t10 VNB.t9 1196.12
R131 VPWR.n9 VPWR.n8 322.159
R132 VPWR.n3 VPWR.n2 316.245
R133 VPWR.n12 VPWR.n5 316.245
R134 VPWR.n7 VPWR.n6 316.245
R135 VPWR.n20 VPWR.t8 254.663
R136 VPWR.n18 VPWR.t9 251.321
R137 VPWR.n17 VPWR.n3 32.7534
R138 VPWR.n19 VPWR.n18 29.7417
R139 VPWR.n13 VPWR.n12 26.7299
R140 VPWR.n2 VPWR.t5 26.5955
R141 VPWR.n2 VPWR.t4 26.5955
R142 VPWR.n5 VPWR.t7 26.5955
R143 VPWR.n5 VPWR.t6 26.5955
R144 VPWR.n6 VPWR.t1 26.5955
R145 VPWR.n6 VPWR.t0 26.5955
R146 VPWR.n8 VPWR.t3 26.5955
R147 VPWR.n8 VPWR.t2 26.5955
R148 VPWR.n12 VPWR.n11 23.7181
R149 VPWR.n18 VPWR.n17 21.0829
R150 VPWR.n20 VPWR.n19 20.7064
R151 VPWR.n11 VPWR.n7 20.7064
R152 VPWR.n13 VPWR.n3 17.6946
R153 VPWR.n11 VPWR.n10 9.3005
R154 VPWR.n12 VPWR.n4 9.3005
R155 VPWR.n14 VPWR.n13 9.3005
R156 VPWR.n15 VPWR.n3 9.3005
R157 VPWR.n17 VPWR.n16 9.3005
R158 VPWR.n18 VPWR.n1 9.3005
R159 VPWR.n19 VPWR.n0 9.3005
R160 VPWR.n21 VPWR.n20 9.3005
R161 VPWR.n9 VPWR.n7 6.87961
R162 VPWR.n10 VPWR.n9 0.654977
R163 VPWR.n10 VPWR.n4 0.120292
R164 VPWR.n14 VPWR.n4 0.120292
R165 VPWR.n15 VPWR.n14 0.120292
R166 VPWR.n16 VPWR.n15 0.120292
R167 VPWR.n16 VPWR.n1 0.120292
R168 VPWR.n1 VPWR.n0 0.120292
R169 VPWR.n21 VPWR.n0 0.120292
R170 VPWR VPWR.n21 0.0226354
R171 a_321_297.n1 a_321_297.t5 267.354
R172 a_321_297.n4 a_321_297.n2 243.446
R173 a_321_297.n4 a_321_297.n3 207.483
R174 a_321_297.n1 a_321_297.n0 207.483
R175 a_321_297.n6 a_321_297.n5 207.482
R176 a_321_297.n5 a_321_297.n1 35.9624
R177 a_321_297.n5 a_321_297.n4 35.9624
R178 a_321_297.n2 a_321_297.t0 26.5955
R179 a_321_297.n2 a_321_297.t4 26.5955
R180 a_321_297.n3 a_321_297.t3 26.5955
R181 a_321_297.n3 a_321_297.t2 26.5955
R182 a_321_297.n0 a_321_297.t7 26.5955
R183 a_321_297.n0 a_321_297.t6 26.5955
R184 a_321_297.n6 a_321_297.t1 26.5955
R185 a_321_297.t8 a_321_297.n6 26.5955
R186 VPB.t10 VPB.t5 591.9
R187 VPB.t4 VPB.t0 248.599
R188 VPB.t3 VPB.t4 248.599
R189 VPB.t2 VPB.t3 248.599
R190 VPB.t1 VPB.t2 248.599
R191 VPB.t8 VPB.t1 248.599
R192 VPB.t7 VPB.t8 248.599
R193 VPB.t6 VPB.t7 248.599
R194 VPB.t5 VPB.t6 248.599
R195 VPB.t9 VPB.t10 248.599
R196 VPB VPB.t9 233.802
R197 SLEEP.n18 SLEEP.n16 212.081
R198 SLEEP.n19 SLEEP.n14 212.081
R199 SLEEP.n13 SLEEP.n11 212.081
R200 SLEEP.n23 SLEEP.n9 212.081
R201 SLEEP.n25 SLEEP.n7 212.081
R202 SLEEP.n5 SLEEP.n3 212.081
R203 SLEEP.n31 SLEEP.n1 212.081
R204 SLEEP.n32 SLEEP.t0 212.081
R205 SLEEP SLEEP.n33 166.081
R206 SLEEP.n22 SLEEP.n21 152
R207 SLEEP.n24 SLEEP.n6 152
R208 SLEEP.n27 SLEEP.n26 152
R209 SLEEP.n29 SLEEP.n28 152
R210 SLEEP.n30 SLEEP.n0 152
R211 SLEEP.n18 SLEEP.n17 139.78
R212 SLEEP.n19 SLEEP.n15 139.78
R213 SLEEP.n13 SLEEP.n12 139.78
R214 SLEEP.n23 SLEEP.n10 139.78
R215 SLEEP.n25 SLEEP.n8 139.78
R216 SLEEP.n5 SLEEP.n4 139.78
R217 SLEEP.n31 SLEEP.n2 139.78
R218 SLEEP.n32 SLEEP.t1 139.78
R219 SLEEP.n21 SLEEP.n20 92.1128
R220 SLEEP.n19 SLEEP.n18 61.346
R221 SLEEP.n30 SLEEP.n29 49.6611
R222 SLEEP.n26 SLEEP.n5 44.549
R223 SLEEP.n33 SLEEP.n31 43.0884
R224 SLEEP.n22 SLEEP.n13 40.1672
R225 SLEEP.n25 SLEEP.n24 32.8641
R226 SLEEP.n20 SLEEP.n13 29.6015
R227 SLEEP.n24 SLEEP.n23 28.4823
R228 SLEEP.n20 SLEEP.n19 25.1769
R229 SLEEP.n21 SLEEP.n6 21.7605
R230 SLEEP.n27 SLEEP.n6 21.7605
R231 SLEEP.n28 SLEEP.n27 21.7605
R232 SLEEP.n28 SLEEP.n0 21.7605
R233 SLEEP.n23 SLEEP.n22 21.1793
R234 SLEEP.n33 SLEEP.n32 18.2581
R235 SLEEP.n26 SLEEP.n25 16.7975
R236 SLEEP SLEEP.n0 7.6805
R237 SLEEP.n31 SLEEP.n30 6.57323
R238 SLEEP.n29 SLEEP.n5 5.11262
R239 A.n0 A.t3 212.081
R240 A.n2 A.t1 212.081
R241 A A.n2 188.474
R242 A.n0 A.t2 174.835
R243 A.n1 A.t0 139.78
R244 A.n2 A.n1 35.055
R245 A.n1 A.n0 26.2914
C0 A VPWR 0.070552f
C1 VPB X 0.016952f
C2 VPB VGND 0.01305f
C3 A X 1.82e-20
C4 SLEEP VPWR 0.065416f
C5 SLEEP X 0.74429f
C6 A VGND 0.127449f
C7 VPWR X 0.045024f
C8 SLEEP VGND 0.109725f
C9 VPWR VGND 0.17328f
C10 X VGND 1.07228f
C11 VPB A 0.088792f
C12 VPB SLEEP 0.246125f
C13 VPB VPWR 0.181362f
C14 VGND VNB 0.965865f
C15 X VNB 0.073273f
C16 VPWR VNB 0.806797f
C17 SLEEP VNB 0.74645f
C18 A VNB 0.307748f
C19 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_16 VPB VNB VGND VPWR SLEEP X A
X0 X.t20 SLEEP.t0 a_505_297# VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t6 a_143_297.t8 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X.t5 a_143_297.t9 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_505_297# SLEEP.t1 X.t19 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_143_297.t4 A.t0 VGND.t23 VNB.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND.t20 SLEEP.t2 X.t34 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X.t18 SLEEP.t3 a_505_297# VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_143_297.t5 A.t1 VGND.t24 VNB.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_505_297# a_143_297.t10 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t5 a_143_297.t11 a_505_297# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 X.t17 SLEEP.t4 a_505_297# VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t19 SLEEP.t5 X.t33 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t18 SLEEP.t6 X.t32 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t9 A.t2 a_143_297.t6 VPB.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t17 SLEEP.t7 X.t31 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_143_297.t7 A.t3 VPWR.t10 VPB.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_505_297# SLEEP.t8 X.t16 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND.t16 SLEEP.t9 X.t30 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR.t4 a_143_297.t12 a_505_297# VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_505_297# SLEEP.t10 X.t15 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 X.t14 SLEEP.t11 a_505_297# VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 X.t13 SLEEP.t12 a_505_297# VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t7 A.t4 a_143_297.t0 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_505_297# SLEEP.t13 X.t12 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND.t21 A.t5 a_143_297.t1 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_505_297# SLEEP.t14 X.t11 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 X.t29 SLEEP.t15 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 X.t10 SLEEP.t16 a_505_297# VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 X.t4 a_143_297.t13 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X30 X.t28 SLEEP.t17 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 X.t27 SLEEP.t18 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 X.t9 SLEEP.t19 a_505_297# VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 X.t26 SLEEP.t20 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_505_297# a_143_297.t14 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_505_297# SLEEP.t21 X.t8 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_143_297.t2 A.t6 VPWR.t8 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR.t2 a_143_297.t15 a_505_297# VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X40 VGND.t3 a_143_297.t16 X.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 VGND.t2 a_143_297.t17 X.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X42 VGND.t11 SLEEP.t22 X.t25 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 a_505_297# a_143_297.t18 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 a_505_297# SLEEP.t23 X.t7 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X45 VGND.t1 a_143_297.t19 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 VGND.t10 SLEEP.t24 X.t24 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 X.t23 SLEEP.t25 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X48 VPWR.t0 a_143_297.t20 a_505_297# VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X49 VGND.t22 A.t7 a_143_297.t3 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X50 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X51 X.t22 SLEEP.t26 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 X.t0 a_143_297.t21 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X53 X.t21 SLEEP.t27 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_143_297.n77 a_143_297.n76 231.56
R1 a_143_297.n75 a_143_297.n1 215.172
R2 a_143_297.n30 a_143_297.n28 212.081
R3 a_143_297.n32 a_143_297.n26 212.081
R4 a_143_297.n24 a_143_297.n22 212.081
R5 a_143_297.n38 a_143_297.n20 212.081
R6 a_143_297.n40 a_143_297.n18 212.081
R7 a_143_297.n43 a_143_297.n41 212.081
R8 a_143_297.n49 a_143_297.n14 212.081
R9 a_143_297.n51 a_143_297.n12 212.081
R10 a_143_297.n10 a_143_297.n8 212.081
R11 a_143_297.n56 a_143_297.t11 212.081
R12 a_143_297.n6 a_143_297.t10 212.081
R13 a_143_297.n62 a_143_297.t12 212.081
R14 a_143_297.n64 a_143_297.t14 212.081
R15 a_143_297.n4 a_143_297.t15 212.081
R16 a_143_297.n70 a_143_297.t18 212.081
R17 a_143_297.n71 a_143_297.t20 212.081
R18 a_143_297.n31 a_143_297.n25 172.725
R19 a_143_297.n73 a_143_297.n72 152
R20 a_143_297.n69 a_143_297.n3 152
R21 a_143_297.n68 a_143_297.n67 152
R22 a_143_297.n66 a_143_297.n65 152
R23 a_143_297.n63 a_143_297.n5 152
R24 a_143_297.n61 a_143_297.n60 152
R25 a_143_297.n59 a_143_297.n58 152
R26 a_143_297.n57 a_143_297.n7 152
R27 a_143_297.n55 a_143_297.n54 152
R28 a_143_297.n53 a_143_297.n52 152
R29 a_143_297.n50 a_143_297.n11 152
R30 a_143_297.n48 a_143_297.n47 152
R31 a_143_297.n46 a_143_297.n16 152
R32 a_143_297.n45 a_143_297.n44 152
R33 a_143_297.n39 a_143_297.n17 152
R34 a_143_297.n37 a_143_297.n36 152
R35 a_143_297.n35 a_143_297.n34 152
R36 a_143_297.n33 a_143_297.n25 152
R37 a_143_297.n30 a_143_297.n29 139.78
R38 a_143_297.n32 a_143_297.n27 139.78
R39 a_143_297.n24 a_143_297.n23 139.78
R40 a_143_297.n38 a_143_297.n21 139.78
R41 a_143_297.n40 a_143_297.n19 139.78
R42 a_143_297.n43 a_143_297.n42 139.78
R43 a_143_297.n49 a_143_297.n15 139.78
R44 a_143_297.n51 a_143_297.n13 139.78
R45 a_143_297.n10 a_143_297.n9 139.78
R46 a_143_297.n56 a_143_297.t21 139.78
R47 a_143_297.n6 a_143_297.t19 139.78
R48 a_143_297.n62 a_143_297.t9 139.78
R49 a_143_297.n64 a_143_297.t17 139.78
R50 a_143_297.n4 a_143_297.t8 139.78
R51 a_143_297.n70 a_143_297.t16 139.78
R52 a_143_297.n71 a_143_297.t13 139.78
R53 a_143_297.n76 a_143_297.n0 115.999
R54 a_143_297.n74 a_143_297.n2 112.273
R55 a_143_297.n74 a_143_297.n73 64.2637
R56 a_143_297.n34 a_143_297.n33 49.6611
R57 a_143_297.n48 a_143_297.n16 49.6611
R58 a_143_297.n58 a_143_297.n57 49.6611
R59 a_143_297.n69 a_143_297.n68 49.6611
R60 a_143_297.n32 a_143_297.n31 48.2005
R61 a_143_297.n72 a_143_297.n70 48.2005
R62 a_143_297.n44 a_143_297.n43 45.2793
R63 a_143_297.n61 a_143_297.n6 45.2793
R64 a_143_297.n50 a_143_297.n49 42.3581
R65 a_143_297.n56 a_143_297.n55 42.3581
R66 a_143_297.n37 a_143_297.n24 39.4369
R67 a_143_297.n65 a_143_297.n4 39.4369
R68 a_143_297.n76 a_143_297.n75 34.9096
R69 a_143_297.n40 a_143_297.n39 33.5944
R70 a_143_297.n63 a_143_297.n62 33.5944
R71 a_143_297.n52 a_143_297.n51 30.6732
R72 a_143_297.n52 a_143_297.n10 30.6732
R73 a_143_297.n39 a_143_297.n38 27.752
R74 a_143_297.n64 a_143_297.n63 27.752
R75 a_143_297.n1 a_143_297.t6 26.5955
R76 a_143_297.n1 a_143_297.t7 26.5955
R77 a_143_297.t0 a_143_297.n77 26.5955
R78 a_143_297.n77 a_143_297.t2 26.5955
R79 a_143_297.n2 a_143_297.t1 24.9236
R80 a_143_297.n2 a_143_297.t5 24.9236
R81 a_143_297.n0 a_143_297.t3 24.9236
R82 a_143_297.n0 a_143_297.t4 24.9236
R83 a_143_297.n38 a_143_297.n37 21.9096
R84 a_143_297.n65 a_143_297.n64 21.9096
R85 a_143_297.n35 a_143_297.n25 20.7243
R86 a_143_297.n36 a_143_297.n35 20.7243
R87 a_143_297.n36 a_143_297.n17 20.7243
R88 a_143_297.n45 a_143_297.n17 20.7243
R89 a_143_297.n46 a_143_297.n45 20.7243
R90 a_143_297.n47 a_143_297.n46 20.7243
R91 a_143_297.n47 a_143_297.n11 20.7243
R92 a_143_297.n53 a_143_297.n11 20.7243
R93 a_143_297.n54 a_143_297.n53 20.7243
R94 a_143_297.n54 a_143_297.n7 20.7243
R95 a_143_297.n59 a_143_297.n7 20.7243
R96 a_143_297.n60 a_143_297.n59 20.7243
R97 a_143_297.n60 a_143_297.n5 20.7243
R98 a_143_297.n66 a_143_297.n5 20.7243
R99 a_143_297.n67 a_143_297.n66 20.7243
R100 a_143_297.n67 a_143_297.n3 20.7243
R101 a_143_297.n73 a_143_297.n3 20.7243
R102 a_143_297.n51 a_143_297.n50 18.9884
R103 a_143_297.n55 a_143_297.n10 18.9884
R104 a_143_297.n44 a_143_297.n40 16.0672
R105 a_143_297.n62 a_143_297.n61 16.0672
R106 a_143_297.n31 a_143_297.n30 13.146
R107 a_143_297.n72 a_143_297.n71 13.146
R108 a_143_297.n75 a_143_297.n74 12.8005
R109 a_143_297.n34 a_143_297.n24 10.2247
R110 a_143_297.n68 a_143_297.n4 10.2247
R111 a_143_297.n49 a_143_297.n48 7.30353
R112 a_143_297.n57 a_143_297.n56 7.30353
R113 a_143_297.n43 a_143_297.n16 4.38232
R114 a_143_297.n58 a_143_297.n6 4.38232
R115 a_143_297.n33 a_143_297.n32 1.46111
R116 a_143_297.n70 a_143_297.n69 1.46111
R117 VPWR.n10 VPWR.t5 348.74
R118 VPWR.n5 VPWR.n4 316.245
R119 VPWR.n13 VPWR.n7 316.245
R120 VPWR.n9 VPWR.n8 316.245
R121 VPWR.n25 VPWR.t8 255.113
R122 VPWR.n19 VPWR.t9 251.321
R123 VPWR.n2 VPWR.n1 231.264
R124 VPWR.n24 VPWR.n23 34.6358
R125 VPWR.n18 VPWR.n5 32.7534
R126 VPWR.n20 VPWR.n19 31.2476
R127 VPWR.n14 VPWR.n13 26.7299
R128 VPWR.n1 VPWR.t10 26.5955
R129 VPWR.n1 VPWR.t7 26.5955
R130 VPWR.n4 VPWR.t1 26.5955
R131 VPWR.n4 VPWR.t0 26.5955
R132 VPWR.n7 VPWR.t3 26.5955
R133 VPWR.n7 VPWR.t2 26.5955
R134 VPWR.n8 VPWR.t6 26.5955
R135 VPWR.n8 VPWR.t4 26.5955
R136 VPWR.n20 VPWR.n2 25.6005
R137 VPWR.n13 VPWR.n12 23.7181
R138 VPWR.n12 VPWR.n9 20.7064
R139 VPWR.n19 VPWR.n18 19.577
R140 VPWR.n14 VPWR.n5 17.6946
R141 VPWR.n26 VPWR.n25 14.5711
R142 VPWR.n25 VPWR.n24 13.177
R143 VPWR.n12 VPWR.n11 9.3005
R144 VPWR.n13 VPWR.n6 9.3005
R145 VPWR.n15 VPWR.n14 9.3005
R146 VPWR.n16 VPWR.n5 9.3005
R147 VPWR.n18 VPWR.n17 9.3005
R148 VPWR.n19 VPWR.n3 9.3005
R149 VPWR.n21 VPWR.n20 9.3005
R150 VPWR.n23 VPWR.n22 9.3005
R151 VPWR.n24 VPWR.n0 9.3005
R152 VPWR.n23 VPWR.n2 9.03579
R153 VPWR.n10 VPWR.n9 6.88081
R154 VPWR.n11 VPWR.n10 0.653676
R155 VPWR.n11 VPWR.n6 0.120292
R156 VPWR.n15 VPWR.n6 0.120292
R157 VPWR.n16 VPWR.n15 0.120292
R158 VPWR.n17 VPWR.n16 0.120292
R159 VPWR.n17 VPWR.n3 0.120292
R160 VPWR.n21 VPWR.n3 0.120292
R161 VPWR.n22 VPWR.n21 0.120292
R162 VPWR.n22 VPWR.n0 0.120292
R163 VPWR.n26 VPWR.n0 0.120292
R164 VPWR VPWR.n26 0.0226354
R165 VPB.t5 VPB.t11 2983.18
R166 VPB.t23 VPB.t0 580.062
R167 VPB VPB.t20 292.991
R168 VPB.t15 VPB.t13 248.599
R169 VPB.t18 VPB.t15 248.599
R170 VPB.t8 VPB.t18 248.599
R171 VPB.t10 VPB.t8 248.599
R172 VPB.t12 VPB.t10 248.599
R173 VPB.t14 VPB.t12 248.599
R174 VPB.t16 VPB.t14 248.599
R175 VPB.t17 VPB.t16 248.599
R176 VPB.t22 VPB.t17 248.599
R177 VPB.t21 VPB.t22 248.599
R178 VPB.t7 VPB.t21 248.599
R179 VPB.t9 VPB.t7 248.599
R180 VPB.t11 VPB.t9 248.599
R181 VPB.t6 VPB.t5 248.599
R182 VPB.t4 VPB.t6 248.599
R183 VPB.t3 VPB.t4 248.599
R184 VPB.t2 VPB.t3 248.599
R185 VPB.t1 VPB.t2 248.599
R186 VPB.t0 VPB.t1 248.599
R187 VPB.t24 VPB.t23 248.599
R188 VPB.t19 VPB.t24 248.599
R189 VPB.t20 VPB.t19 248.599
R190 SLEEP.n6 SLEEP.t13 212.081
R191 SLEEP.n7 SLEEP.t16 212.081
R192 SLEEP.n9 SLEEP.t23 212.081
R193 SLEEP.n11 SLEEP.t4 212.081
R194 SLEEP.n4 SLEEP.t10 212.081
R195 SLEEP.n16 SLEEP.t12 212.081
R196 SLEEP.n2 SLEEP.t14 212.081
R197 SLEEP.n22 SLEEP.t19 212.081
R198 SLEEP.n24 SLEEP.t21 212.081
R199 SLEEP.n49 SLEEP.t0 212.081
R200 SLEEP.n25 SLEEP.t1 212.081
R201 SLEEP.n43 SLEEP.t3 212.081
R202 SLEEP.n41 SLEEP.t8 212.081
R203 SLEEP.n27 SLEEP.t11 212.081
R204 SLEEP.n35 SLEEP.n29 212.081
R205 SLEEP.n33 SLEEP.n31 212.081
R206 SLEEP.n34 SLEEP.n28 172.725
R207 SLEEP.n10 SLEEP.n5 152
R208 SLEEP.n13 SLEEP.n12 152
R209 SLEEP.n15 SLEEP.n14 152
R210 SLEEP.n17 SLEEP.n3 152
R211 SLEEP.n19 SLEEP.n18 152
R212 SLEEP.n21 SLEEP.n20 152
R213 SLEEP.n23 SLEEP.n0 152
R214 SLEEP.n51 SLEEP.n50 152
R215 SLEEP.n48 SLEEP.n1 152
R216 SLEEP.n47 SLEEP.n46 152
R217 SLEEP.n45 SLEEP.n44 152
R218 SLEEP.n42 SLEEP.n26 152
R219 SLEEP.n40 SLEEP.n39 152
R220 SLEEP.n38 SLEEP.n37 152
R221 SLEEP.n36 SLEEP.n28 152
R222 SLEEP.n6 SLEEP.t2 139.78
R223 SLEEP.n7 SLEEP.t25 139.78
R224 SLEEP.n9 SLEEP.t24 139.78
R225 SLEEP.n11 SLEEP.t20 139.78
R226 SLEEP.n4 SLEEP.t22 139.78
R227 SLEEP.n16 SLEEP.t18 139.78
R228 SLEEP.n2 SLEEP.t9 139.78
R229 SLEEP.n22 SLEEP.t17 139.78
R230 SLEEP.n24 SLEEP.t7 139.78
R231 SLEEP.n49 SLEEP.t15 139.78
R232 SLEEP.n25 SLEEP.t6 139.78
R233 SLEEP.n43 SLEEP.t27 139.78
R234 SLEEP.n41 SLEEP.t5 139.78
R235 SLEEP.n27 SLEEP.t26 139.78
R236 SLEEP.n35 SLEEP.n30 139.78
R237 SLEEP.n33 SLEEP.n32 139.78
R238 SLEEP.n8 SLEEP.n5 90.8506
R239 SLEEP.n7 SLEEP.n6 61.346
R240 SLEEP.n18 SLEEP.n17 49.6611
R241 SLEEP.n48 SLEEP.n47 49.6611
R242 SLEEP.n37 SLEEP.n36 49.6611
R243 SLEEP.n35 SLEEP.n34 48.2005
R244 SLEEP.n16 SLEEP.n15 45.2793
R245 SLEEP.n44 SLEEP.n25 45.2793
R246 SLEEP.n21 SLEEP.n2 42.3581
R247 SLEEP.n50 SLEEP.n49 42.3581
R248 SLEEP.n10 SLEEP.n9 39.4369
R249 SLEEP.n40 SLEEP.n27 39.4369
R250 SLEEP.n12 SLEEP.n4 33.5944
R251 SLEEP.n43 SLEEP.n42 33.5944
R252 SLEEP.n23 SLEEP.n22 30.6732
R253 SLEEP.n24 SLEEP.n23 30.6732
R254 SLEEP.n9 SLEEP.n8 30.3874
R255 SLEEP.n12 SLEEP.n11 27.752
R256 SLEEP.n42 SLEEP.n41 27.752
R257 SLEEP.n8 SLEEP.n7 24.3727
R258 SLEEP.n11 SLEEP.n10 21.9096
R259 SLEEP.n41 SLEEP.n40 21.9096
R260 SLEEP.n13 SLEEP.n5 20.7243
R261 SLEEP.n14 SLEEP.n13 20.7243
R262 SLEEP.n14 SLEEP.n3 20.7243
R263 SLEEP.n19 SLEEP.n3 20.7243
R264 SLEEP.n20 SLEEP.n19 20.7243
R265 SLEEP.n20 SLEEP.n0 20.7243
R266 SLEEP.n51 SLEEP.n1 20.7243
R267 SLEEP.n46 SLEEP.n1 20.7243
R268 SLEEP.n46 SLEEP.n45 20.7243
R269 SLEEP.n45 SLEEP.n26 20.7243
R270 SLEEP.n39 SLEEP.n26 20.7243
R271 SLEEP.n39 SLEEP.n38 20.7243
R272 SLEEP.n38 SLEEP.n28 20.7243
R273 SLEEP.n22 SLEEP.n21 18.9884
R274 SLEEP.n50 SLEEP.n24 18.9884
R275 SLEEP.n15 SLEEP.n4 16.0672
R276 SLEEP.n44 SLEEP.n43 16.0672
R277 SLEEP SLEEP.n0 15.5434
R278 SLEEP.n34 SLEEP.n33 13.146
R279 SLEEP.n37 SLEEP.n27 10.2247
R280 SLEEP.n18 SLEEP.n2 7.30353
R281 SLEEP.n49 SLEEP.n48 7.30353
R282 SLEEP SLEEP.n51 5.18145
R283 SLEEP.n17 SLEEP.n16 4.38232
R284 SLEEP.n47 SLEEP.n25 4.38232
R285 SLEEP.n36 SLEEP.n35 1.46111
R286 X.n2 X.n0 345.308
R287 X.n2 X.n1 300.885
R288 X.n4 X.n3 300.885
R289 X.n6 X.n5 300.885
R290 X.n8 X.n7 300.885
R291 X.n10 X.n9 300.885
R292 X.n12 X.n11 300.885
R293 X.n20 X.n18 217.601
R294 X.n18 X.t0 136.792
R295 X.n15 X.n13 135.249
R296 X.n32 X.n31 98.9924
R297 X.n15 X.n14 98.982
R298 X.n17 X.n16 98.982
R299 X.n20 X.n19 98.982
R300 X.n22 X.n21 98.982
R301 X.n24 X.n23 98.982
R302 X.n26 X.n25 98.982
R303 X.n28 X.n27 98.982
R304 X.n30 X.n29 98.982
R305 X.n4 X.n2 44.424
R306 X.n6 X.n4 44.424
R307 X.n8 X.n6 44.424
R308 X.n10 X.n8 44.424
R309 X.n12 X.n10 44.424
R310 X.n17 X.n15 36.2672
R311 X.n18 X.n17 36.2672
R312 X.n22 X.n20 36.2672
R313 X.n24 X.n22 36.2672
R314 X.n26 X.n24 36.2672
R315 X.n28 X.n26 36.2672
R316 X.n30 X.n28 36.2672
R317 X.n32 X.n30 36.2672
R318 X.n0 X.t16 26.5955
R319 X.n0 X.t14 26.5955
R320 X.n1 X.t19 26.5955
R321 X.n1 X.t18 26.5955
R322 X.n3 X.t8 26.5955
R323 X.n3 X.t20 26.5955
R324 X.n5 X.t11 26.5955
R325 X.n5 X.t9 26.5955
R326 X.n7 X.t15 26.5955
R327 X.n7 X.t13 26.5955
R328 X.n9 X.t7 26.5955
R329 X.n9 X.t17 26.5955
R330 X.n11 X.t12 26.5955
R331 X.n11 X.t10 26.5955
R332 X.n13 X.t3 24.9236
R333 X.n13 X.t4 24.9236
R334 X.n14 X.t2 24.9236
R335 X.n14 X.t6 24.9236
R336 X.n16 X.t1 24.9236
R337 X.n16 X.t5 24.9236
R338 X.n19 X.t33 24.9236
R339 X.n19 X.t22 24.9236
R340 X.n21 X.t32 24.9236
R341 X.n21 X.t21 24.9236
R342 X.n23 X.t31 24.9236
R343 X.n23 X.t29 24.9236
R344 X.n25 X.t30 24.9236
R345 X.n25 X.t28 24.9236
R346 X.n27 X.t25 24.9236
R347 X.n27 X.t27 24.9236
R348 X.n29 X.t24 24.9236
R349 X.n29 X.t26 24.9236
R350 X.n31 X.t34 24.9236
R351 X.n31 X.t23 24.9236
R352 X X.n32 12.312
R353 X X.n12 2.23346
R354 VGND.n26 VGND.t20 288.839
R355 VGND.n15 VGND.t8 283.521
R356 VGND.n25 VGND.n24 207.965
R357 VGND.n30 VGND.n23 207.965
R358 VGND.n32 VGND.n31 207.965
R359 VGND.n38 VGND.n20 207.965
R360 VGND.n41 VGND.n40 207.965
R361 VGND.n47 VGND.n17 207.965
R362 VGND.n9 VGND.n8 207.965
R363 VGND.n71 VGND.n7 207.965
R364 VGND.n5 VGND.n4 207.965
R365 VGND.n84 VGND.t23 150.077
R366 VGND.n82 VGND.n2 116.624
R367 VGND.n78 VGND.n77 59.2832
R368 VGND.n77 VGND.t4 56.3082
R369 VGND.n77 VGND.t21 56.3082
R370 VGND.n65 VGND.n64 34.6358
R371 VGND.n29 VGND.n28 34.6358
R372 VGND.n37 VGND.n21 34.6358
R373 VGND.n42 VGND.n39 34.6358
R374 VGND.n46 VGND.n18 34.6358
R375 VGND.n49 VGND.n48 34.6358
R376 VGND.n53 VGND.n52 34.6358
R377 VGND.n54 VGND.n53 34.6358
R378 VGND.n54 VGND.n13 34.6358
R379 VGND.n58 VGND.n13 34.6358
R380 VGND.n59 VGND.n58 34.6358
R381 VGND.n60 VGND.n59 34.6358
R382 VGND.n60 VGND.n11 34.6358
R383 VGND.n64 VGND.n11 34.6358
R384 VGND.n66 VGND.n65 34.6358
R385 VGND.n70 VGND.n69 34.6358
R386 VGND.n76 VGND.n75 34.6358
R387 VGND.n82 VGND.n1 34.2593
R388 VGND.n33 VGND.n32 33.1299
R389 VGND.n72 VGND.n71 33.1299
R390 VGND.n33 VGND.n30 30.1181
R391 VGND.n72 VGND.n5 30.1181
R392 VGND.n38 VGND.n37 27.1064
R393 VGND.n69 VGND.n9 27.1064
R394 VGND.n52 VGND.n15 25.6005
R395 VGND.n84 VGND.n83 25.224
R396 VGND.n24 VGND.t9 24.9236
R397 VGND.n24 VGND.t10 24.9236
R398 VGND.n23 VGND.t12 24.9236
R399 VGND.n23 VGND.t11 24.9236
R400 VGND.n31 VGND.t13 24.9236
R401 VGND.n31 VGND.t16 24.9236
R402 VGND.n20 VGND.t14 24.9236
R403 VGND.n20 VGND.t17 24.9236
R404 VGND.n40 VGND.t15 24.9236
R405 VGND.n40 VGND.t18 24.9236
R406 VGND.n17 VGND.t7 24.9236
R407 VGND.n17 VGND.t19 24.9236
R408 VGND.n8 VGND.t0 24.9236
R409 VGND.n8 VGND.t1 24.9236
R410 VGND.n7 VGND.t5 24.9236
R411 VGND.n7 VGND.t2 24.9236
R412 VGND.n4 VGND.t6 24.9236
R413 VGND.n4 VGND.t3 24.9236
R414 VGND.n2 VGND.t24 24.9236
R415 VGND.n2 VGND.t22 24.9236
R416 VGND.n28 VGND.n25 24.0946
R417 VGND.n42 VGND.n41 21.0829
R418 VGND.n48 VGND.n47 19.577
R419 VGND.n78 VGND.n76 17.6946
R420 VGND.n26 VGND.n25 17.4932
R421 VGND.n83 VGND.n82 16.1887
R422 VGND.n47 VGND.n46 15.0593
R423 VGND.n41 VGND.n18 13.5534
R424 VGND.n78 VGND.n1 10.1652
R425 VGND.n28 VGND.n27 9.3005
R426 VGND.n29 VGND.n22 9.3005
R427 VGND.n34 VGND.n33 9.3005
R428 VGND.n35 VGND.n21 9.3005
R429 VGND.n37 VGND.n36 9.3005
R430 VGND.n39 VGND.n19 9.3005
R431 VGND.n43 VGND.n42 9.3005
R432 VGND.n44 VGND.n18 9.3005
R433 VGND.n46 VGND.n45 9.3005
R434 VGND.n48 VGND.n16 9.3005
R435 VGND.n50 VGND.n49 9.3005
R436 VGND.n52 VGND.n51 9.3005
R437 VGND.n53 VGND.n14 9.3005
R438 VGND.n55 VGND.n54 9.3005
R439 VGND.n56 VGND.n13 9.3005
R440 VGND.n58 VGND.n57 9.3005
R441 VGND.n59 VGND.n12 9.3005
R442 VGND.n61 VGND.n60 9.3005
R443 VGND.n62 VGND.n11 9.3005
R444 VGND.n64 VGND.n63 9.3005
R445 VGND.n65 VGND.n10 9.3005
R446 VGND.n67 VGND.n66 9.3005
R447 VGND.n69 VGND.n68 9.3005
R448 VGND.n70 VGND.n6 9.3005
R449 VGND.n73 VGND.n72 9.3005
R450 VGND.n75 VGND.n74 9.3005
R451 VGND.n76 VGND.n3 9.3005
R452 VGND.n79 VGND.n78 9.3005
R453 VGND.n80 VGND.n1 9.3005
R454 VGND.n82 VGND.n81 9.3005
R455 VGND.n83 VGND.n0 9.3005
R456 VGND.n49 VGND.n15 9.03579
R457 VGND.n39 VGND.n38 7.52991
R458 VGND.n66 VGND.n9 7.52991
R459 VGND.n85 VGND.n84 6.99075
R460 VGND.n30 VGND.n29 4.51815
R461 VGND.n75 VGND.n5 4.51815
R462 VGND.n32 VGND.n21 1.50638
R463 VGND.n71 VGND.n70 1.50638
R464 VGND.n27 VGND.n26 0.765081
R465 VGND.n85 VGND.n0 0.150171
R466 VGND.n27 VGND.n22 0.120292
R467 VGND.n34 VGND.n22 0.120292
R468 VGND.n35 VGND.n34 0.120292
R469 VGND.n36 VGND.n35 0.120292
R470 VGND.n36 VGND.n19 0.120292
R471 VGND.n43 VGND.n19 0.120292
R472 VGND.n44 VGND.n43 0.120292
R473 VGND.n45 VGND.n44 0.120292
R474 VGND.n45 VGND.n16 0.120292
R475 VGND.n50 VGND.n16 0.120292
R476 VGND.n51 VGND.n50 0.120292
R477 VGND.n51 VGND.n14 0.120292
R478 VGND.n55 VGND.n14 0.120292
R479 VGND.n56 VGND.n55 0.120292
R480 VGND.n57 VGND.n56 0.120292
R481 VGND.n57 VGND.n12 0.120292
R482 VGND.n61 VGND.n12 0.120292
R483 VGND.n62 VGND.n61 0.120292
R484 VGND.n63 VGND.n62 0.120292
R485 VGND.n63 VGND.n10 0.120292
R486 VGND.n67 VGND.n10 0.120292
R487 VGND.n68 VGND.n67 0.120292
R488 VGND.n68 VGND.n6 0.120292
R489 VGND.n73 VGND.n6 0.120292
R490 VGND.n74 VGND.n73 0.120292
R491 VGND.n74 VGND.n3 0.120292
R492 VGND.n79 VGND.n3 0.120292
R493 VGND.n80 VGND.n79 0.120292
R494 VGND.n81 VGND.n80 0.120292
R495 VGND.n81 VGND.n0 0.120292
R496 VGND VGND.n85 0.113169
R497 VNB.t0 VNB.t8 14353.4
R498 VNB.t21 VNB.t4 2164.4
R499 VNB VNB.t23 2036.25
R500 VNB.t9 VNB.t20 1196.12
R501 VNB.t10 VNB.t9 1196.12
R502 VNB.t12 VNB.t10 1196.12
R503 VNB.t11 VNB.t12 1196.12
R504 VNB.t13 VNB.t11 1196.12
R505 VNB.t16 VNB.t13 1196.12
R506 VNB.t14 VNB.t16 1196.12
R507 VNB.t17 VNB.t14 1196.12
R508 VNB.t15 VNB.t17 1196.12
R509 VNB.t18 VNB.t15 1196.12
R510 VNB.t7 VNB.t18 1196.12
R511 VNB.t19 VNB.t7 1196.12
R512 VNB.t8 VNB.t19 1196.12
R513 VNB.t1 VNB.t0 1196.12
R514 VNB.t5 VNB.t1 1196.12
R515 VNB.t2 VNB.t5 1196.12
R516 VNB.t6 VNB.t2 1196.12
R517 VNB.t3 VNB.t6 1196.12
R518 VNB.t4 VNB.t3 1196.12
R519 VNB.t24 VNB.t21 1196.12
R520 VNB.t22 VNB.t24 1196.12
R521 VNB.t23 VNB.t22 1196.12
R522 A.n0 A.t2 212.081
R523 A.n2 A.t3 212.081
R524 A.n4 A.t4 212.081
R525 A.n6 A.t6 212.081
R526 A.n0 A.t5 171.913
R527 A.n5 A.t0 139.78
R528 A.n3 A.t7 139.78
R529 A.n1 A.t1 139.78
R530 A A.n6 99.3452
R531 A.n2 A.n1 32.1338
R532 A.n4 A.n3 32.1338
R533 A.n6 A.n5 32.1338
R534 A.n1 A.n0 29.2126
R535 A.n3 A.n2 29.2126
R536 A.n5 A.n4 29.2126
C0 a_505_297# VPB 0.050054f
C1 VGND VPB 0.021259f
C2 a_505_297# A 1.18e-19
C3 VGND A 0.189894f
C4 a_505_297# SLEEP 0.244631f
C5 VGND SLEEP 0.225121f
C6 VPB A 0.161223f
C7 a_505_297# VPWR 2.27951f
C8 VGND VPWR 0.324815f
C9 VPB SLEEP 0.503433f
C10 a_505_297# X 0.986312f
C11 VGND X 2.12056f
C12 VPB VPWR 0.313074f
C13 A VPWR 0.104224f
C14 VPB X 0.029846f
C15 SLEEP VPWR 0.131568f
C16 SLEEP X 1.57762f
C17 VPWR X 0.092292f
C18 VGND a_505_297# 0.03618f
C19 VGND VNB 1.777767f
C20 X VNB 0.142439f
C21 VPWR VNB 1.463692f
C22 SLEEP VNB 1.48019f
C23 A VNB 0.506977f
C24 VPB VNB 3.26264f
C25 a_505_297# VNB 0.022326f
C26 VGND.n0 VNB 0.037649f
C27 VGND.n1 VNB 0.007128f
C28 VGND.t24 VNB 0.006236f
C29 VGND.t22 VNB 0.006236f
C30 VGND.n2 VNB 0.01758f
C31 VGND.n3 VNB 0.031384f
C32 VGND.t6 VNB 0.006236f
C33 VGND.t3 VNB 0.006236f
C34 VGND.n4 VNB 0.01332f
C35 VGND.n5 VNB 0.016067f
C36 VGND.n6 VNB 0.031384f
C37 VGND.t5 VNB 0.006236f
C38 VGND.t2 VNB 0.006236f
C39 VGND.n7 VNB 0.01332f
C40 VGND.t0 VNB 0.006236f
C41 VGND.t1 VNB 0.006236f
C42 VGND.n8 VNB 0.01332f
C43 VGND.n9 VNB 0.016067f
C44 VGND.n10 VNB 0.031384f
C45 VGND.n11 VNB 0.003435f
C46 VGND.n12 VNB 0.031384f
C47 VGND.n13 VNB -0.001292f
C48 VGND.n14 VNB 0.031384f
C49 VGND.t8 VNB 0.023112f
C50 VGND.n15 VNB 0.018747f
C51 VGND.n16 VNB 0.031384f
C52 VGND.t7 VNB 0.006236f
C53 VGND.t19 VNB 0.006236f
C54 VGND.n17 VNB 0.01332f
C55 VGND.n18 VNB 0.007732f
C56 VGND.n19 VNB 0.031384f
C57 VGND.t14 VNB 0.006236f
C58 VGND.t17 VNB 0.006236f
C59 VGND.n20 VNB 0.01332f
C60 VGND.n21 VNB 0.005799f
C61 VGND.n22 VNB 0.031384f
C62 VGND.t12 VNB 0.006236f
C63 VGND.t11 VNB 0.006236f
C64 VGND.n23 VNB 0.01332f
C65 VGND.t9 VNB 0.006236f
C66 VGND.t10 VNB 0.006236f
C67 VGND.n24 VNB 0.01332f
C68 VGND.n25 VNB 0.019204f
C69 VGND.t20 VNB 0.023337f
C70 VGND.n26 VNB 0.060808f
C71 VGND.n27 VNB 0.10979f
C72 VGND.n28 VNB 0.009424f
C73 VGND.n29 VNB 0.006282f
C74 VGND.n30 VNB 0.016067f
C75 VGND.t13 VNB 0.006236f
C76 VGND.t16 VNB 0.006236f
C77 VGND.n31 VNB 0.01332f
C78 VGND.n32 VNB 0.016067f
C79 VGND.n33 VNB 0.010149f
C80 VGND.n34 VNB 0.031384f
C81 VGND.n35 VNB 0.031384f
C82 VGND.n36 VNB 0.031384f
C83 VGND.n37 VNB 0.009907f
C84 VGND.n38 VNB 0.016067f
C85 VGND.n39 VNB 0.006766f
C86 VGND.t15 VNB 0.006236f
C87 VGND.t18 VNB 0.006236f
C88 VGND.n40 VNB 0.01332f
C89 VGND.n41 VNB 0.016067f
C90 VGND.n42 VNB 0.00894f
C91 VGND.n43 VNB 0.031384f
C92 VGND.n44 VNB 0.031384f
C93 VGND.n45 VNB 0.031384f
C94 VGND.n46 VNB 0.007974f
C95 VGND.n47 VNB 0.016067f
C96 VGND.n48 VNB 0.008699f
C97 VGND.n49 VNB 0.007007f
C98 VGND.n50 VNB 0.031384f
C99 VGND.n51 VNB 0.031384f
C100 VGND.n52 VNB 0.009665f
C101 VGND.n53 VNB -0.001292f
C102 VGND.n54 VNB 0.008752f
C103 VGND.n55 VNB 0.031384f
C104 VGND.n56 VNB 0.031384f
C105 VGND.n57 VNB 0.031384f
C106 VGND.n58 VNB 0.00757f
C107 VGND.n59 VNB 0.001072f
C108 VGND.n60 VNB 0.005207f
C109 VGND.n61 VNB 0.031384f
C110 VGND.n62 VNB 0.031384f
C111 VGND.n63 VNB 0.031384f
C112 VGND.n64 VNB 0.002844f
C113 VGND.n65 VNB 0.005798f
C114 VGND.n66 VNB 0.006766f
C115 VGND.n67 VNB 0.031384f
C116 VGND.n68 VNB 0.031384f
C117 VGND.n69 VNB 0.009907f
C118 VGND.n70 VNB 0.005799f
C119 VGND.n71 VNB 0.016067f
C120 VGND.n72 VNB 0.010149f
C121 VGND.n73 VNB 0.031384f
C122 VGND.n74 VNB 0.031384f
C123 VGND.n75 VNB 0.006282f
C124 VGND.n76 VNB 0.008397f
C125 VGND.t4 VNB 0.014089f
C126 VGND.t21 VNB 0.014089f
C127 VGND.n77 VNB 0.03892f
C128 VGND.n78 VNB 0.071122f
C129 VGND.n79 VNB 0.031384f
C130 VGND.n80 VNB 0.031384f
C131 VGND.n81 VNB 0.031384f
C132 VGND.n82 VNB 0.037811f
C133 VGND.n83 VNB 0.006645f
C134 VGND.t23 VNB 0.022895f
C135 VGND.n84 VNB 0.053756f
C136 VGND.n85 VNB 0.029914f
C137 X.t16 VNB 0.011429f
C138 X.t14 VNB 0.011429f
C139 X.n0 VNB 0.039938f
C140 X.t19 VNB 0.011429f
C141 X.t18 VNB 0.011429f
C142 X.n1 VNB 0.023576f
C143 X.n2 VNB 0.15545f
C144 X.t8 VNB 0.011429f
C145 X.t20 VNB 0.011429f
C146 X.n3 VNB 0.023576f
C147 X.n4 VNB 0.044624f
C148 X.t11 VNB 0.011429f
C149 X.t9 VNB 0.011429f
C150 X.n5 VNB 0.023576f
C151 X.n6 VNB 0.044624f
C152 X.t15 VNB 0.011429f
C153 X.t13 VNB 0.011429f
C154 X.n7 VNB 0.023576f
C155 X.n8 VNB 0.044624f
C156 X.t7 VNB 0.011429f
C157 X.t17 VNB 0.011429f
C158 X.n9 VNB 0.023576f
C159 X.n10 VNB 0.044624f
C160 X.t12 VNB 0.011429f
C161 X.t10 VNB 0.011429f
C162 X.n11 VNB 0.023576f
C163 X.n12 VNB 0.04848f
C164 X.t3 VNB 0.007429f
C165 X.t4 VNB 0.007429f
C166 X.n13 VNB 0.028187f
C167 X.t2 VNB 0.007429f
C168 X.t6 VNB 0.007429f
C169 X.n14 VNB 0.016917f
C170 X.n15 VNB 0.080561f
C171 X.t1 VNB 0.007429f
C172 X.t5 VNB 0.007429f
C173 X.n16 VNB 0.016917f
C174 X.n17 VNB 0.049801f
C175 X.t0 VNB 0.025152f
C176 X.n18 VNB 0.26036f
C177 X.t33 VNB 0.007429f
C178 X.t22 VNB 0.007429f
C179 X.n19 VNB 0.016917f
C180 X.n20 VNB 0.253738f
C181 X.t32 VNB 0.007429f
C182 X.t21 VNB 0.007429f
C183 X.n21 VNB 0.016917f
C184 X.n22 VNB 0.049801f
C185 X.t31 VNB 0.007429f
C186 X.t29 VNB 0.007429f
C187 X.n23 VNB 0.016917f
C188 X.n24 VNB 0.049801f
C189 X.t30 VNB 0.007429f
C190 X.t28 VNB 0.007429f
C191 X.n25 VNB 0.016917f
C192 X.n26 VNB 0.049801f
C193 X.t25 VNB 0.007429f
C194 X.t27 VNB 0.007429f
C195 X.n27 VNB 0.016917f
C196 X.n28 VNB 0.049801f
C197 X.t24 VNB 0.007429f
C198 X.t26 VNB 0.007429f
C199 X.n29 VNB 0.016917f
C200 X.n30 VNB 0.049801f
C201 X.t34 VNB 0.007429f
C202 X.t23 VNB 0.007429f
C203 X.n31 VNB 0.016842f
C204 X.n32 VNB 0.085943f
C205 VPWR.n0 VNB 0.031604f
C206 VPWR.t8 VNB 0.038496f
C207 VPWR.t10 VNB 0.009662f
C208 VPWR.t7 VNB 0.009662f
C209 VPWR.n1 VNB 0.023315f
C210 VPWR.n2 VNB 0.030318f
C211 VPWR.n3 VNB 0.031604f
C212 VPWR.t9 VNB 0.041308f
C213 VPWR.t1 VNB 0.009662f
C214 VPWR.t0 VNB 0.009662f
C215 VPWR.n4 VNB 0.021178f
C216 VPWR.n5 VNB 0.041006f
C217 VPWR.n6 VNB 0.031604f
C218 VPWR.t3 VNB 0.009662f
C219 VPWR.t2 VNB 0.009662f
C220 VPWR.n7 VNB 0.021178f
C221 VPWR.t6 VNB 0.009662f
C222 VPWR.t4 VNB 0.009662f
C223 VPWR.n8 VNB 0.021178f
C224 VPWR.n9 VNB 0.041887f
C225 VPWR.t5 VNB 0.039703f
C226 VPWR.n10 VNB 0.367392f
C227 VPWR.n11 VNB 1.06074f
C228 VPWR.n12 VNB 0.007178f
C229 VPWR.n13 VNB 0.041006f
C230 VPWR.n14 VNB 0.007178f
C231 VPWR.n15 VNB 0.031604f
C232 VPWR.n16 VNB 0.031604f
C233 VPWR.n17 VNB 0.031604f
C234 VPWR.n18 VNB 0.008456f
C235 VPWR.n19 VNB 0.054324f
C236 VPWR.n20 VNB 0.009186f
C237 VPWR.n21 VNB 0.031604f
C238 VPWR.n22 VNB 0.031604f
C239 VPWR.n23 VNB 0.007057f
C240 VPWR.n24 VNB 0.007726f
C241 VPWR.n25 VNB 0.046129f
C242 VPWR.n26 VNB 0.021055f
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 VNB VPB VGND VPWR KAPWR X A SLEEP
X0 VPWR.t3 SLEEP.t0 a_255_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 KAPWR.t15 a_1122_47.t8 X.t10 VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VGND.t4 SLEEP.t1 a_341_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t20 a_1122_47.t9 X.t3 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VGND.t19 a_1122_47.t10 X.t2 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 a_255_297.t2 SLEEP.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t18 a_1122_47.t11 X.t1 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 X.t9 a_1122_47.t12 KAPWR.t14 VPB.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_341_47.t0 a_147_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR.t1 SLEEP.t3 a_255_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 KAPWR.t19 a_341_47.t12 a_1122_47.t6 VPB.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 KAPWR.t13 a_1122_47.t13 X.t8 VPB.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND.t17 a_1122_47.t14 X.t0 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 X.t7 a_1122_47.t15 KAPWR.t12 VPB.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 VGND.t26 a_341_47.t13 a_1122_47.t7 VNB.t26 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 a_255_297.t7 a_147_47.t3 a_341_47.t10 VPB.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 KAPWR.t11 a_1122_47.t16 X.t6 VPB.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X17 X.t22 a_1122_47.t17 VGND.t16 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VGND.t15 a_1122_47.t18 X.t21 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X.t5 a_1122_47.t19 KAPWR.t10 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X20 a_341_47.t9 a_147_47.t4 a_255_297.t6 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 KAPWR.t9 a_1122_47.t20 X.t4 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 X.t20 a_1122_47.t21 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_147_47.t1 A.t0 VGND.t27 VNB.t27 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1755 ps=1.84 w=0.65 l=0.15
X24 VGND.t22 a_147_47.t5 a_341_47.t8 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VGND.t13 a_1122_47.t22 X.t19 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 a_147_47.t0 A.t1 VPWR.t4 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.28 ps=2.56 w=1 l=0.15
X27 a_255_297.t5 a_147_47.t6 a_341_47.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1122_47.t3 a_341_47.t14 KAPWR.t18 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VGND.t28 a_147_47.t7 a_341_47.t11 VNB.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 X.t31 a_1122_47.t23 KAPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 KAPWR.t7 a_1122_47.t24 X.t30 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 VGND.t3 SLEEP.t4 a_341_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 X.t18 a_1122_47.t25 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 a_1122_47.t4 a_341_47.t15 VGND.t25 VNB.t25 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 KAPWR.t6 a_1122_47.t26 X.t29 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 X.t28 a_1122_47.t27 KAPWR.t5 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X37 X.t17 a_1122_47.t28 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X.t16 a_1122_47.t29 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 a_1122_47.t5 a_341_47.t16 VGND.t24 VNB.t24 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X40 a_255_297.t0 SLEEP.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X41 KAPWR.t16 a_341_47.t17 a_1122_47.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X42 X.t27 a_1122_47.t30 KAPWR.t4 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X43 a_341_47.t6 a_147_47.t8 VGND.t21 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X44 X.t26 a_1122_47.t31 KAPWR.t3 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X45 a_341_47.t2 SLEEP.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 a_341_47.t1 SLEEP.t7 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 X.t15 a_1122_47.t32 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X48 X.t14 a_1122_47.t33 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X49 a_341_47.t5 a_147_47.t9 a_255_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X50 VGND.t23 a_341_47.t18 a_1122_47.t1 VNB.t23 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X51 X.t13 a_1122_47.t34 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X52 KAPWR.t2 a_1122_47.t35 X.t25 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X53 KAPWR.t1 a_1122_47.t36 X.t24 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X54 a_1122_47.t2 a_341_47.t19 KAPWR.t17 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X55 VGND.t6 a_1122_47.t37 X.t12 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X56 X.t23 a_1122_47.t38 KAPWR.t0 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X57 VGND.t5 a_1122_47.t39 X.t11 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 SLEEP.n0 SLEEP.t5 212.081
R1 SLEEP.n3 SLEEP.t0 212.081
R2 SLEEP.n6 SLEEP.t2 212.081
R3 SLEEP.n4 SLEEP.t3 212.081
R4 SLEEP.n5 SLEEP.n2 173.761
R5 SLEEP SLEEP.n1 163.52
R6 SLEEP.n9 SLEEP.n8 152
R7 SLEEP.n7 SLEEP.n2 152
R8 SLEEP.n0 SLEEP.t1 139.78
R9 SLEEP.n3 SLEEP.t7 139.78
R10 SLEEP.n6 SLEEP.t4 139.78
R11 SLEEP.n4 SLEEP.t6 139.78
R12 SLEEP.n8 SLEEP.n7 49.6611
R13 SLEEP.n3 SLEEP.n1 45.2793
R14 SLEEP.n6 SLEEP.n5 42.3581
R15 SLEEP.n9 SLEEP.n2 21.7605
R16 SLEEP.n5 SLEEP.n4 18.9884
R17 SLEEP.n1 SLEEP.n0 16.0672
R18 SLEEP SLEEP.n9 10.2405
R19 SLEEP.n7 SLEEP.n6 7.30353
R20 SLEEP.n8 SLEEP.n3 4.38232
R21 a_255_297.n3 a_255_297.n2 296.538
R22 a_255_297.t0 a_255_297.n5 278.784
R23 a_255_297.n3 a_255_297.t4 267.592
R24 a_255_297.n5 a_255_297.n0 207.26
R25 a_255_297.n4 a_255_297.n1 188.952
R26 a_255_297.n5 a_255_297.n4 57.3601
R27 a_255_297.n4 a_255_297.n3 53.34
R28 a_255_297.n0 a_255_297.t3 26.5955
R29 a_255_297.n0 a_255_297.t2 26.5955
R30 a_255_297.n1 a_255_297.t1 26.5955
R31 a_255_297.n1 a_255_297.t7 26.5955
R32 a_255_297.n2 a_255_297.t6 26.5955
R33 a_255_297.n2 a_255_297.t5 26.5955
R34 VPWR.n4 VPWR.n3 316.245
R35 VPWR.n6 VPWR.n5 315.86
R36 VPWR.n16 VPWR.t4 239.476
R37 VPWR.n9 VPWR.n8 34.6358
R38 VPWR.n10 VPWR.n9 34.6358
R39 VPWR.n10 VPWR.n1 34.6358
R40 VPWR.n14 VPWR.n1 34.6358
R41 VPWR.n15 VPWR.n14 34.6358
R42 VPWR.n8 VPWR.n4 33.5064
R43 VPWR.n3 VPWR.t2 26.5955
R44 VPWR.n3 VPWR.t1 26.5955
R45 VPWR.n5 VPWR.t0 26.5955
R46 VPWR.n5 VPWR.t3 26.5955
R47 VPWR.n16 VPWR.n15 11.6711
R48 VPWR.n8 VPWR.n7 9.3005
R49 VPWR.n9 VPWR.n2 9.3005
R50 VPWR.n11 VPWR.n10 9.3005
R51 VPWR.n12 VPWR.n1 9.3005
R52 VPWR.n14 VPWR.n13 9.3005
R53 VPWR.n15 VPWR.n0 9.3005
R54 VPWR.n17 VPWR.n16 9.3005
R55 VPWR.n6 VPWR.n4 6.18238
R56 VPWR.n7 VPWR.n6 0.64888
R57 VPWR.n7 VPWR.n2 0.120292
R58 VPWR.n11 VPWR.n2 0.120292
R59 VPWR.n12 VPWR.n11 0.120292
R60 VPWR.n13 VPWR.n12 0.120292
R61 VPWR.n13 VPWR.n0 0.120292
R62 VPWR.n17 VPWR.n0 0.120292
R63 VPWR VPWR.n17 0.0213333
R64 VPB.t20 VPB.t4 574.144
R65 VPB.t0 VPB 375.858
R66 VPB VPB.t20 301.87
R67 VPB.t15 VPB.t18 254.518
R68 VPB.t10 VPB.t15 254.518
R69 VPB.t23 VPB.t10 254.518
R70 VPB.t17 VPB.t23 254.518
R71 VPB.t14 VPB.t17 254.518
R72 VPB.t13 VPB.t14 254.518
R73 VPB.t9 VPB.t13 254.518
R74 VPB.t25 VPB.t26 254.518
R75 VPB.t22 VPB.t25 254.518
R76 VPB.t16 VPB.t22 254.518
R77 VPB.t12 VPB.t16 254.518
R78 VPB.t11 VPB.t12 254.518
R79 VPB.t24 VPB.t11 254.518
R80 VPB.t19 VPB.t24 254.518
R81 VPB.t5 VPB.t19 254.518
R82 VPB.t7 VPB.t5 254.518
R83 VPB.t27 VPB.t7 254.518
R84 VPB.t6 VPB.t27 254.518
R85 VPB.t26 VPB.t9 251.559
R86 VPB.t3 VPB.t0 248.599
R87 VPB.t2 VPB.t3 248.599
R88 VPB.t1 VPB.t2 248.599
R89 VPB.t28 VPB.t1 248.599
R90 VPB.t21 VPB.t28 248.599
R91 VPB.t8 VPB.t21 248.599
R92 VPB.t4 VPB.t8 248.599
R93 VPB VPB.t6 145.017
R94 a_1122_47.n49 a_1122_47.n48 227.921
R95 a_1122_47.n50 a_1122_47.n2 226.815
R96 a_1122_47.n49 a_1122_47.n47 220.84
R97 a_1122_47.n2 a_1122_47.n3 217.256
R98 a_1122_47.n11 a_1122_47.t36 212.081
R99 a_1122_47.n12 a_1122_47.t30 212.081
R100 a_1122_47.n13 a_1122_47.t20 212.081
R101 a_1122_47.n15 a_1122_47.t12 212.081
R102 a_1122_47.n17 a_1122_47.t35 212.081
R103 a_1122_47.n1 a_1122_47.t27 212.081
R104 a_1122_47.n22 a_1122_47.t26 212.081
R105 a_1122_47.n8 a_1122_47.t19 212.081
R106 a_1122_47.n27 a_1122_47.t16 212.081
R107 a_1122_47.n0 a_1122_47.t15 212.081
R108 a_1122_47.n32 a_1122_47.t8 212.081
R109 a_1122_47.n34 a_1122_47.t31 212.081
R110 a_1122_47.n35 a_1122_47.t24 212.081
R111 a_1122_47.n41 a_1122_47.t23 212.081
R112 a_1122_47.n43 a_1122_47.t13 212.081
R113 a_1122_47.n44 a_1122_47.t38 212.081
R114 a_1122_47.n14 a_1122_47.n10 169.409
R115 a_1122_47.n11 a_1122_47.t14 162.274
R116 a_1122_47.n12 a_1122_47.t25 162.274
R117 a_1122_47.n13 a_1122_47.t18 162.274
R118 a_1122_47.n15 a_1122_47.t29 162.274
R119 a_1122_47.n17 a_1122_47.t22 162.274
R120 a_1122_47.n1 a_1122_47.t33 162.274
R121 a_1122_47.n22 a_1122_47.t39 162.274
R122 a_1122_47.n8 a_1122_47.t34 162.274
R123 a_1122_47.n27 a_1122_47.t10 162.274
R124 a_1122_47.n0 a_1122_47.t28 162.274
R125 a_1122_47.n32 a_1122_47.t37 162.274
R126 a_1122_47.n34 a_1122_47.t32 162.274
R127 a_1122_47.n35 a_1122_47.t9 162.274
R128 a_1122_47.n41 a_1122_47.t17 162.274
R129 a_1122_47.n43 a_1122_47.t11 162.274
R130 a_1122_47.n44 a_1122_47.t21 162.274
R131 a_1122_47.n46 a_1122_47.n45 152
R132 a_1122_47.n42 a_1122_47.n4 152
R133 a_1122_47.n40 a_1122_47.n39 152
R134 a_1122_47.n38 a_1122_47.n5 152
R135 a_1122_47.n37 a_1122_47.n36 152
R136 a_1122_47.n33 a_1122_47.n6 152
R137 a_1122_47.n31 a_1122_47.n30 152
R138 a_1122_47.n29 a_1122_47.n0 152
R139 a_1122_47.n28 a_1122_47.n7 152
R140 a_1122_47.n26 a_1122_47.n25 152
R141 a_1122_47.n24 a_1122_47.n23 152
R142 a_1122_47.n21 a_1122_47.n9 152
R143 a_1122_47.n1 a_1122_47.n20 152
R144 a_1122_47.n19 a_1122_47.n18 152
R145 a_1122_47.n16 a_1122_47.n10 152
R146 a_1122_47.n12 a_1122_47.n11 55.2698
R147 a_1122_47.n13 a_1122_47.n12 55.2698
R148 a_1122_47.n18 a_1122_47.n1 43.7018
R149 a_1122_47.n21 a_1122_47.n1 43.7018
R150 a_1122_47.n0 a_1122_47.n28 43.7018
R151 a_1122_47.n40 a_1122_47.n5 43.7018
R152 a_1122_47.n31 a_1122_47.n0 43.7018
R153 a_1122_47.n2 a_1122_47.n46 43.5205
R154 a_1122_47.n2 a_1122_47.n49 43.5205
R155 a_1122_47.n47 a_1122_47.t1 40.0005
R156 a_1122_47.n47 a_1122_47.t5 40.0005
R157 a_1122_47.n3 a_1122_47.t7 40.0005
R158 a_1122_47.n3 a_1122_47.t4 40.0005
R159 a_1122_47.n42 a_1122_47.n41 39.8458
R160 a_1122_47.n36 a_1122_47.n35 35.9898
R161 a_1122_47.n14 a_1122_47.n13 35.3472
R162 a_1122_47.n27 a_1122_47.n26 33.4192
R163 a_1122_47.n23 a_1122_47.n22 32.7765
R164 a_1122_47.n17 a_1122_47.n16 31.4912
R165 a_1122_47.n33 a_1122_47.n32 30.8485
R166 a_1122_47.n45 a_1122_47.n43 28.2778
R167 a_1122_47.n48 a_1122_47.t6 27.5805
R168 a_1122_47.n48 a_1122_47.t2 27.5805
R169 a_1122_47.t0 a_1122_47.n50 27.5805
R170 a_1122_47.n50 a_1122_47.t3 27.5805
R171 a_1122_47.n45 a_1122_47.n44 26.9925
R172 a_1122_47.n34 a_1122_47.n33 24.4218
R173 a_1122_47.n16 a_1122_47.n15 23.7792
R174 a_1122_47.n23 a_1122_47.n8 22.4938
R175 a_1122_47.n26 a_1122_47.n8 21.2085
R176 a_1122_47.n15 a_1122_47.n14 19.9232
R177 a_1122_47.n36 a_1122_47.n34 19.2805
R178 a_1122_47.n19 a_1122_47.n10 17.4085
R179 a_1122_47.n20 a_1122_47.n19 17.4085
R180 a_1122_47.n20 a_1122_47.n9 17.4085
R181 a_1122_47.n24 a_1122_47.n9 17.4085
R182 a_1122_47.n25 a_1122_47.n24 17.4085
R183 a_1122_47.n25 a_1122_47.n7 17.4085
R184 a_1122_47.n29 a_1122_47.n7 17.4085
R185 a_1122_47.n30 a_1122_47.n29 17.4085
R186 a_1122_47.n30 a_1122_47.n6 17.4085
R187 a_1122_47.n37 a_1122_47.n6 17.4085
R188 a_1122_47.n38 a_1122_47.n37 17.4085
R189 a_1122_47.n39 a_1122_47.n38 17.4085
R190 a_1122_47.n39 a_1122_47.n4 17.4085
R191 a_1122_47.n46 a_1122_47.n4 17.4085
R192 a_1122_47.n43 a_1122_47.n42 15.4245
R193 a_1122_47.n32 a_1122_47.n31 12.8538
R194 a_1122_47.n18 a_1122_47.n17 12.2112
R195 a_1122_47.n22 a_1122_47.n21 10.9258
R196 a_1122_47.n28 a_1122_47.n27 10.2832
R197 a_1122_47.n35 a_1122_47.n5 7.7125
R198 a_1122_47.n41 a_1122_47.n40 3.8565
R199 X.n15 X.n13 338.599
R200 X.n15 X.n14 303.454
R201 X.n17 X.n16 303.454
R202 X.n19 X.n18 303.454
R203 X.n21 X.n20 303.454
R204 X.n23 X.n22 303.454
R205 X.n25 X.n24 303.454
R206 X.n27 X.n26 299.724
R207 X.n2 X.n0 248.638
R208 X.n2 X.n1 203.463
R209 X.n4 X.n3 203.463
R210 X.n8 X.n7 203.463
R211 X.n10 X.n9 203.463
R212 X.n12 X.n11 203.463
R213 X.n6 X.n5 202.456
R214 X X.n29 199.607
R215 X.n4 X.n2 45.177
R216 X.n10 X.n8 45.177
R217 X.n12 X.n10 45.177
R218 X.n6 X.n4 44.0476
R219 X.n8 X.n6 44.0476
R220 X.n0 X.t1 40.0005
R221 X.n0 X.t20 40.0005
R222 X.n1 X.t3 40.0005
R223 X.n1 X.t22 40.0005
R224 X.n3 X.t12 40.0005
R225 X.n3 X.t15 40.0005
R226 X.n5 X.t2 40.0005
R227 X.n5 X.t17 40.0005
R228 X.n7 X.t11 40.0005
R229 X.n7 X.t13 40.0005
R230 X.n9 X.t19 40.0005
R231 X.n9 X.t14 40.0005
R232 X.n11 X.t21 40.0005
R233 X.n11 X.t16 40.0005
R234 X.n29 X.t0 40.0005
R235 X.n29 X.t18 40.0005
R236 X.n17 X.n15 32.0005
R237 X.n19 X.n17 32.0005
R238 X.n23 X.n21 32.0005
R239 X.n25 X.n23 32.0005
R240 X.n21 X.n19 31.2005
R241 X.n24 X.t4 27.5805
R242 X.n24 X.t9 27.5805
R243 X.n13 X.t8 27.5805
R244 X.n13 X.t23 27.5805
R245 X.n14 X.t30 27.5805
R246 X.n14 X.t31 27.5805
R247 X.n16 X.t10 27.5805
R248 X.n16 X.t26 27.5805
R249 X.n18 X.t6 27.5805
R250 X.n18 X.t7 27.5805
R251 X.n20 X.t29 27.5805
R252 X.n20 X.t5 27.5805
R253 X.n22 X.t25 27.5805
R254 X.n22 X.t28 27.5805
R255 X.n26 X.t24 27.5805
R256 X.n26 X.t27 27.5805
R257 X.n28 X.n12 13.177
R258 X.n27 X.n25 10.4484
R259 X.n28 X 3.13183
R260 X X.n27 1.75844
R261 X X.n28 0.604792
R262 KAPWR.n1 KAPWR.t1 769.73
R263 KAPWR.n7 KAPWR.n6 594.822
R264 KAPWR.n5 KAPWR.n4 594.822
R265 KAPWR.n3 KAPWR.n2 594.822
R266 KAPWR.n11 KAPWR.n10 594.793
R267 KAPWR.n9 KAPWR.n8 594.793
R268 KAPWR.n13 KAPWR.n12 594.644
R269 KAPWR.n1 KAPWR.n0 594.529
R270 KAPWR.n18 KAPWR.t17 237.472
R271 KAPWR.n17 KAPWR.n16 209.893
R272 KAPWR.n15 KAPWR.n14 209.893
R273 KAPWR.n16 KAPWR.t18 27.5805
R274 KAPWR.n16 KAPWR.t19 27.5805
R275 KAPWR.n14 KAPWR.t0 27.5805
R276 KAPWR.n14 KAPWR.t16 27.5805
R277 KAPWR.n12 KAPWR.t8 27.5805
R278 KAPWR.n12 KAPWR.t13 27.5805
R279 KAPWR.n10 KAPWR.t3 27.5805
R280 KAPWR.n10 KAPWR.t7 27.5805
R281 KAPWR.n8 KAPWR.t12 27.5805
R282 KAPWR.n8 KAPWR.t15 27.5805
R283 KAPWR.n6 KAPWR.t11 27.5805
R284 KAPWR.n4 KAPWR.t5 27.5805
R285 KAPWR.n4 KAPWR.t6 27.5805
R286 KAPWR.n2 KAPWR.t14 27.5805
R287 KAPWR.n2 KAPWR.t2 27.5805
R288 KAPWR.n0 KAPWR.t4 27.5805
R289 KAPWR.n0 KAPWR.t9 27.5805
R290 KAPWR.n6 KAPWR.t10 26.5955
R291 KAPWR KAPWR.n18 3.22334
R292 KAPWR.n13 KAPWR.n11 0.508673
R293 KAPWR.n7 KAPWR.n5 0.496173
R294 KAPWR.n11 KAPWR.n9 0.496173
R295 KAPWR.n18 KAPWR.n17 0.496173
R296 KAPWR.n5 KAPWR.n3 0.493048
R297 KAPWR.n9 KAPWR.n7 0.493048
R298 KAPWR.n17 KAPWR.n15 0.493048
R299 KAPWR.n3 KAPWR.n1 0.489923
R300 KAPWR.n15 KAPWR.n13 0.489923
R301 a_341_47.n15 a_341_47.n14 321.88
R302 a_341_47.n14 a_341_47.n1 298.637
R303 a_341_47.n12 a_341_47.n7 195.246
R304 a_341_47.n4 a_341_47.t17 184.768
R305 a_341_47.n5 a_341_47.t14 184.768
R306 a_341_47.n6 a_341_47.t12 184.768
R307 a_341_47.n7 a_341_47.t19 184.768
R308 a_341_47.n4 a_341_47.t13 146.208
R309 a_341_47.n5 a_341_47.t15 146.208
R310 a_341_47.n6 a_341_47.t18 146.208
R311 a_341_47.n7 a_341_47.t16 146.208
R312 a_341_47.n0 a_341_47.n13 138.359
R313 a_341_47.n10 a_341_47.n8 135.249
R314 a_341_47.n10 a_341_47.n9 98.982
R315 a_341_47.n3 a_341_47.n2 95.6388
R316 a_341_47.n5 a_341_47.n4 40.6397
R317 a_341_47.n6 a_341_47.n5 40.6397
R318 a_341_47.n7 a_341_47.n6 40.6397
R319 a_341_47.n1 a_341_47.t10 26.5955
R320 a_341_47.n1 a_341_47.t9 26.5955
R321 a_341_47.n15 a_341_47.t7 26.5955
R322 a_341_47.t5 a_341_47.n15 26.5955
R323 a_341_47.n11 a_341_47.n10 25.1561
R324 a_341_47.n2 a_341_47.t11 24.9236
R325 a_341_47.n2 a_341_47.t6 24.9236
R326 a_341_47.n13 a_341_47.t8 24.9236
R327 a_341_47.n13 a_341_47.t0 24.9236
R328 a_341_47.n8 a_341_47.t4 24.9236
R329 a_341_47.n8 a_341_47.t1 24.9236
R330 a_341_47.n9 a_341_47.t3 24.9236
R331 a_341_47.n9 a_341_47.t2 24.9236
R332 a_341_47.n14 a_341_47.n0 24.4369
R333 a_341_47.n11 a_341_47.n3 15.4672
R334 a_341_47.n0 a_341_47.n12 9.49615
R335 a_341_47.n12 a_341_47.n11 9.3005
R336 a_341_47.n0 a_341_47.n3 4.26717
R337 VGND.n57 VGND.t4 265.401
R338 VGND.t4 VGND.n7 257.858
R339 VGND.n22 VGND.t17 248.373
R340 VGND.n55 VGND.t24 225
R341 VGND.n62 VGND.n6 207.965
R342 VGND.n65 VGND.n64 207.965
R343 VGND.n71 VGND.n3 207.965
R344 VGND.n49 VGND.n48 206.909
R345 VGND.n10 VGND.n9 206.909
R346 VGND.n33 VGND.n32 205.899
R347 VGND.n35 VGND.n34 205.899
R348 VGND.n26 VGND.n25 205.481
R349 VGND.n18 VGND.n17 205.481
R350 VGND.n21 VGND.n20 204.692
R351 VGND.n42 VGND.n41 204.692
R352 VGND.n13 VGND.n12 204.692
R353 VGND.n1 VGND.t0 152.594
R354 VGND.n78 VGND.t27 151.139
R355 VGND.n20 VGND.t12 40.0005
R356 VGND.n20 VGND.t15 40.0005
R357 VGND.n25 VGND.t10 40.0005
R358 VGND.n25 VGND.t13 40.0005
R359 VGND.n17 VGND.t8 40.0005
R360 VGND.n17 VGND.t5 40.0005
R361 VGND.n32 VGND.t19 40.0005
R362 VGND.n34 VGND.t11 40.0005
R363 VGND.n34 VGND.t6 40.0005
R364 VGND.n41 VGND.t9 40.0005
R365 VGND.n41 VGND.t20 40.0005
R366 VGND.n12 VGND.t16 40.0005
R367 VGND.n12 VGND.t18 40.0005
R368 VGND.n48 VGND.t14 40.0005
R369 VGND.n48 VGND.t26 40.0005
R370 VGND.n9 VGND.t25 40.0005
R371 VGND.n9 VGND.t23 40.0005
R372 VGND.n32 VGND.t7 38.5719
R373 VGND.n36 VGND.n33 34.6358
R374 VGND.n40 VGND.n15 34.6358
R375 VGND.n44 VGND.n43 34.6358
R376 VGND.n66 VGND.n63 34.6358
R377 VGND.n70 VGND.n4 34.6358
R378 VGND.n73 VGND.n72 34.6358
R379 VGND.n77 VGND.n76 34.6358
R380 VGND.n62 VGND.n61 32.377
R381 VGND.n49 VGND.n47 31.624
R382 VGND.n31 VGND.n18 29.7417
R383 VGND.n50 VGND.n10 27.1064
R384 VGND.n66 VGND.n65 26.3534
R385 VGND.n61 VGND.n7 26.1449
R386 VGND.n26 VGND.n24 25.224
R387 VGND.n27 VGND.n26 25.224
R388 VGND.n55 VGND.n54 25.1487
R389 VGND.n6 VGND.t1 24.9236
R390 VGND.n6 VGND.t3 24.9236
R391 VGND.n64 VGND.t2 24.9236
R392 VGND.n64 VGND.t28 24.9236
R393 VGND.n3 VGND.t21 24.9236
R394 VGND.n3 VGND.t22 24.9236
R395 VGND.n54 VGND.n10 22.5887
R396 VGND.n24 VGND.n21 20.7064
R397 VGND.n27 VGND.n18 20.7064
R398 VGND.n71 VGND.n70 20.3299
R399 VGND.n50 VGND.n49 18.0711
R400 VGND.n33 VGND.n31 16.1887
R401 VGND.n72 VGND.n71 14.3064
R402 VGND.n47 VGND.n13 13.5534
R403 VGND.n36 VGND.n35 11.6711
R404 VGND.n78 VGND.n77 11.6711
R405 VGND.n79 VGND.n78 10.4299
R406 VGND.n24 VGND.n23 9.3005
R407 VGND.n26 VGND.n19 9.3005
R408 VGND.n28 VGND.n27 9.3005
R409 VGND.n29 VGND.n18 9.3005
R410 VGND.n31 VGND.n30 9.3005
R411 VGND.n33 VGND.n16 9.3005
R412 VGND.n37 VGND.n36 9.3005
R413 VGND.n38 VGND.n15 9.3005
R414 VGND.n40 VGND.n39 9.3005
R415 VGND.n43 VGND.n14 9.3005
R416 VGND.n45 VGND.n44 9.3005
R417 VGND.n47 VGND.n46 9.3005
R418 VGND.n49 VGND.n11 9.3005
R419 VGND.n51 VGND.n50 9.3005
R420 VGND.n52 VGND.n10 9.3005
R421 VGND.n54 VGND.n53 9.3005
R422 VGND.n56 VGND.n8 9.3005
R423 VGND.n59 VGND.n58 9.3005
R424 VGND.n61 VGND.n60 9.3005
R425 VGND.n63 VGND.n5 9.3005
R426 VGND.n67 VGND.n66 9.3005
R427 VGND.n68 VGND.n4 9.3005
R428 VGND.n70 VGND.n69 9.3005
R429 VGND.n72 VGND.n2 9.3005
R430 VGND.n74 VGND.n73 9.3005
R431 VGND.n76 VGND.n75 9.3005
R432 VGND.n77 VGND.n0 9.3005
R433 VGND.n43 VGND.n42 9.03579
R434 VGND.n57 VGND.n56 8.9605
R435 VGND.n65 VGND.n4 8.28285
R436 VGND.n73 VGND.n1 7.90638
R437 VGND.n22 VGND.n21 6.84811
R438 VGND.n42 VGND.n40 6.02403
R439 VGND.n76 VGND.n1 4.89462
R440 VGND.n35 VGND.n15 4.51815
R441 VGND.n63 VGND.n62 2.25932
R442 VGND.n44 VGND.n13 1.50638
R443 VGND.n58 VGND.n7 0.985115
R444 VGND.n23 VGND.n22 0.661516
R445 VGND.n56 VGND.n55 0.591269
R446 VGND.n23 VGND.n19 0.120292
R447 VGND.n28 VGND.n19 0.120292
R448 VGND.n29 VGND.n28 0.120292
R449 VGND.n30 VGND.n29 0.120292
R450 VGND.n30 VGND.n16 0.120292
R451 VGND.n37 VGND.n16 0.120292
R452 VGND.n38 VGND.n37 0.120292
R453 VGND.n39 VGND.n38 0.120292
R454 VGND.n39 VGND.n14 0.120292
R455 VGND.n45 VGND.n14 0.120292
R456 VGND.n46 VGND.n45 0.120292
R457 VGND.n46 VGND.n11 0.120292
R458 VGND.n51 VGND.n11 0.120292
R459 VGND.n52 VGND.n51 0.120292
R460 VGND.n53 VGND.n52 0.120292
R461 VGND.n53 VGND.n8 0.120292
R462 VGND.n59 VGND.n8 0.120292
R463 VGND.n60 VGND.n59 0.120292
R464 VGND.n60 VGND.n5 0.120292
R465 VGND.n67 VGND.n5 0.120292
R466 VGND.n68 VGND.n67 0.120292
R467 VGND.n69 VGND.n68 0.120292
R468 VGND.n69 VGND.n2 0.120292
R469 VGND.n74 VGND.n2 0.120292
R470 VGND.n75 VGND.n74 0.120292
R471 VGND.n75 VGND.n0 0.120292
R472 VGND.n79 VGND.n0 0.120292
R473 VGND.n58 VGND.n57 0.0989615
R474 VGND VGND.n79 0.0213333
R475 VNB.t27 VNB.t0 2762.46
R476 VNB.t4 VNB 1808.41
R477 VNB VNB.t27 1452.43
R478 VNB.t12 VNB.t17 1224.6
R479 VNB.t15 VNB.t12 1224.6
R480 VNB.t10 VNB.t15 1224.6
R481 VNB.t13 VNB.t10 1224.6
R482 VNB.t8 VNB.t13 1224.6
R483 VNB.t5 VNB.t8 1224.6
R484 VNB.t7 VNB.t5 1224.6
R485 VNB.t11 VNB.t19 1224.6
R486 VNB.t6 VNB.t11 1224.6
R487 VNB.t9 VNB.t6 1224.6
R488 VNB.t20 VNB.t9 1224.6
R489 VNB.t16 VNB.t20 1224.6
R490 VNB.t18 VNB.t16 1224.6
R491 VNB.t14 VNB.t18 1224.6
R492 VNB.t26 VNB.t14 1224.6
R493 VNB.t25 VNB.t26 1224.6
R494 VNB.t23 VNB.t25 1224.6
R495 VNB.t24 VNB.t23 1224.6
R496 VNB.t19 VNB.t7 1210.36
R497 VNB.t1 VNB.t4 1196.12
R498 VNB.t3 VNB.t1 1196.12
R499 VNB.t2 VNB.t3 1196.12
R500 VNB.t28 VNB.t2 1196.12
R501 VNB.t21 VNB.t28 1196.12
R502 VNB.t22 VNB.t21 1196.12
R503 VNB.t0 VNB.t22 1196.12
R504 VNB VNB.t24 697.736
R505 a_147_47.t0 a_147_47.n8 252.549
R506 a_147_47.n1 a_147_47.t3 212.081
R507 a_147_47.n2 a_147_47.t4 212.081
R508 a_147_47.n4 a_147_47.t6 212.081
R509 a_147_47.n0 a_147_47.t9 212.081
R510 a_147_47.n6 a_147_47.n3 173.761
R511 a_147_47.n8 a_147_47.t1 153.874
R512 a_147_47.n6 a_147_47.n5 152
R513 a_147_47.n1 a_147_47.t7 139.78
R514 a_147_47.n2 a_147_47.t8 139.78
R515 a_147_47.n4 a_147_47.t5 139.78
R516 a_147_47.n0 a_147_47.t2 139.78
R517 a_147_47.n7 a_147_47.n0 112.322
R518 a_147_47.n2 a_147_47.n1 61.346
R519 a_147_47.n3 a_147_47.n2 54.0429
R520 a_147_47.n5 a_147_47.n4 42.3581
R521 a_147_47.n7 a_147_47.n6 30.5712
R522 a_147_47.n5 a_147_47.n0 18.9884
R523 a_147_47.n8 a_147_47.n7 14.5696
R524 a_147_47.n4 a_147_47.n3 7.30353
R525 A.n0 A.t1 229.754
R526 A A.n0 162.45
R527 A.n0 A.t0 157.453
C0 KAPWR SLEEP 0.021826f
C1 VGND VPB 0.01726f
C2 VGND A 0.05163f
C3 VGND SLEEP 0.055482f
C4 VPB A 0.04669f
C5 VPWR KAPWR 1.99558f
C6 VPB SLEEP 0.120132f
C7 VPWR X 0.277351f
C8 VPWR VGND 0.011604f
C9 KAPWR X 1.27396f
C10 KAPWR VGND 0.250559f
C11 X VGND 0.973835f
C12 VPWR VPB 0.247844f
C13 VPWR A 0.050363f
C14 KAPWR VPB 0.043789f
C15 KAPWR A 0.008158f
C16 VPWR SLEEP 0.064161f
C17 X VPB 0.031597f
C18 VGND VNB 1.55771f
C19 X VNB 0.110579f
C20 KAPWR VNB 0.028251f
C21 VPWR VNB 1.28044f
C22 SLEEP VNB 0.362171f
C23 A VNB 0.150465f
C24 VPB VNB 2.81966f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47.t1 a_27_47.t2 a_1108_47.t2 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 VGND.t3 a_1283_21.t3 Q.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_1283_21.t1 a_1108_47.t4 a_1462_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 a_651_413.t2 a_27_47.t3 a_543_47.t2 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 VPWR.t4 a_1283_21.t4 Q.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_1108_47.t0 a_193_47.t2 a_761_289.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND.t5 RESET_B.t0 a_805_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q.t0 a_1283_21.t5 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X9 VPWR.t2 CLK.t0 a_27_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 a_448_47.t0 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_761_289.t1 a_543_47.t4 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 a_193_47.t1 a_27_47.t4 VGND.t8 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47.t1 a_27_47.t5 a_761_289.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X14 a_1462_47.t1 RESET_B.t1 VGND.t6 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X15 a_543_47.t1 a_27_47.t6 a_448_47.t3 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_543_47.t0 a_193_47.t3 a_448_47.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47.t1 D.t1 VGND.t7 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X18 VPWR.t5 a_1283_21.t6 a_1270_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR.t8 a_1108_47.t5 a_1283_21.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413.t1 a_193_47.t4 a_1108_47.t3 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47.t0 a_27_47.t7 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21.t0 RESET_B.t2 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR.t1 a_761_289.t5 a_651_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X24 Q.t1 a_1283_21.t7 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X25 a_639_47.t1 a_193_47.t5 a_543_47.t3 VNB.t14 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND.t4 a_1283_21.t8 a_1217_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413.t1 RESET_B.t3 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_761_289.t0 a_543_47.t5 VPWR.t9 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
R0 a_761_289.n3 a_761_289.n2 647.119
R1 a_761_289.n1 a_761_289.t4 350.253
R2 a_761_289.n2 a_761_289.n0 260.339
R3 a_761_289.n2 a_761_289.n1 246.119
R4 a_761_289.n1 a_761_289.t5 189.588
R5 a_761_289.n3 a_761_289.t2 89.1195
R6 a_761_289.n0 a_761_289.t3 63.3338
R7 a_761_289.t0 a_761_289.n3 41.0422
R8 a_761_289.n0 a_761_289.t1 31.9797
R9 a_639_47.t0 a_639_47.t1 198.571
R10 a_805_47.t0 a_805_47.t1 60.0005
R11 VNB.t7 VNB.t13 3631.07
R12 VNB.t2 VNB.t4 2961.81
R13 VNB.t14 VNB.t1 2363.75
R14 VNB.t5 VNB.t12 2121.68
R15 VNB.t9 VNB.t3 1879.61
R16 VNB.t11 VNB.t6 1552.1
R17 VNB.t3 VNB.t11 1409.71
R18 VNB.t6 VNB.t5 1366.99
R19 VNB.t8 VNB.t14 1366.99
R20 VNB.t13 VNB.t8 1352.75
R21 VNB.t12 VNB.t2 1295.79
R22 VNB.t4 VNB.t10 1196.12
R23 VNB.t0 VNB.t7 1196.12
R24 VNB.t1 VNB.t9 1025.24
R25 VNB VNB.t0 925.567
R26 a_27_47.n1 a_27_47.t3 530.01
R27 a_27_47.t1 a_27_47.n5 421.021
R28 a_27_47.n0 a_27_47.t5 337.142
R29 a_27_47.n3 a_27_47.t0 280.223
R30 a_27_47.n4 a_27_47.t7 263.173
R31 a_27_47.n4 a_27_47.t4 227.826
R32 a_27_47.n0 a_27_47.t2 199.762
R33 a_27_47.n2 a_27_47.n1 170.81
R34 a_27_47.n2 a_27_47.n0 167.321
R35 a_27_47.n5 a_27_47.n4 152
R36 a_27_47.n1 a_27_47.t6 141.923
R37 a_27_47.n3 a_27_47.n2 10.8376
R38 a_27_47.n5 a_27_47.n3 2.50485
R39 a_1108_47.n3 a_1108_47.n2 636.953
R40 a_1108_47.n1 a_1108_47.t4 366.856
R41 a_1108_47.n2 a_1108_47.n0 300.2
R42 a_1108_47.n2 a_1108_47.n1 225.036
R43 a_1108_47.n1 a_1108_47.t5 174.056
R44 a_1108_47.n0 a_1108_47.t0 70.0005
R45 a_1108_47.t1 a_1108_47.n3 68.0124
R46 a_1108_47.n3 a_1108_47.t3 63.3219
R47 a_1108_47.n0 a_1108_47.t2 61.6672
R48 a_1217_47.t0 a_1217_47.t1 94.7268
R49 a_1283_21.n5 a_1283_21.n4 807.871
R50 a_1283_21.n2 a_1283_21.t6 389.183
R51 a_1283_21.n3 a_1283_21.n2 251.167
R52 a_1283_21.n3 a_1283_21.t1 223.571
R53 a_1283_21.n0 a_1283_21.t4 212.081
R54 a_1283_21.n1 a_1283_21.t5 212.081
R55 a_1283_21.n4 a_1283_21.n1 176.576
R56 a_1283_21.n2 a_1283_21.t8 174.891
R57 a_1283_21.n0 a_1283_21.t3 139.78
R58 a_1283_21.n1 a_1283_21.t7 139.78
R59 a_1283_21.n5 a_1283_21.t2 63.3219
R60 a_1283_21.t0 a_1283_21.n5 63.3219
R61 a_1283_21.n1 a_1283_21.n0 61.346
R62 a_1283_21.n4 a_1283_21.n3 37.7195
R63 Q Q.n0 586.793
R64 Q.n3 Q.n0 585
R65 Q.n2 Q.n1 185
R66 Q Q.n2 49.0339
R67 Q.n0 Q.t3 26.5955
R68 Q.n0 Q.t0 26.5955
R69 Q.n1 Q.t2 24.9236
R70 Q.n1 Q.t1 24.9236
R71 Q Q.n3 15.6165
R72 Q.n2 Q 10.4965
R73 Q.n3 Q 1.7925
R74 VGND.n36 VGND.t7 307.536
R75 VGND.n8 VGND.t3 244.825
R76 VGND.n9 VGND.t2 226.882
R77 VGND.n16 VGND.n15 209.254
R78 VGND.n25 VGND.n24 199.739
R79 VGND.n39 VGND.n38 199.739
R80 VGND.n15 VGND.t6 100.001
R81 VGND.n24 VGND.t5 72.8576
R82 VGND.n15 VGND.t4 70.0005
R83 VGND.n24 VGND.t1 60.5809
R84 VGND.n38 VGND.t8 38.5719
R85 VGND.n38 VGND.t0 38.5719
R86 VGND.n10 VGND.n7 34.6358
R87 VGND.n14 VGND.n7 34.6358
R88 VGND.n18 VGND.n17 34.6358
R89 VGND.n18 VGND.n5 34.6358
R90 VGND.n22 VGND.n5 34.6358
R91 VGND.n23 VGND.n22 34.6358
R92 VGND.n26 VGND.n3 34.6358
R93 VGND.n30 VGND.n3 34.6358
R94 VGND.n31 VGND.n30 34.6358
R95 VGND.n32 VGND.n31 34.6358
R96 VGND.n32 VGND.n1 34.6358
R97 VGND.n37 VGND.n36 29.7417
R98 VGND.n10 VGND.n9 24.8476
R99 VGND.n39 VGND.n37 22.9652
R100 VGND.n16 VGND.n14 17.6946
R101 VGND.n36 VGND.n1 14.6829
R102 VGND.n37 VGND.n0 9.3005
R103 VGND.n36 VGND.n35 9.3005
R104 VGND.n34 VGND.n1 9.3005
R105 VGND.n33 VGND.n32 9.3005
R106 VGND.n31 VGND.n2 9.3005
R107 VGND.n30 VGND.n29 9.3005
R108 VGND.n28 VGND.n3 9.3005
R109 VGND.n27 VGND.n26 9.3005
R110 VGND.n23 VGND.n4 9.3005
R111 VGND.n22 VGND.n21 9.3005
R112 VGND.n20 VGND.n5 9.3005
R113 VGND.n19 VGND.n18 9.3005
R114 VGND.n17 VGND.n6 9.3005
R115 VGND.n14 VGND.n13 9.3005
R116 VGND.n12 VGND.n7 9.3005
R117 VGND.n11 VGND.n10 9.3005
R118 VGND.n26 VGND.n25 7.90638
R119 VGND.n40 VGND.n39 7.12063
R120 VGND.n9 VGND.n8 6.48892
R121 VGND.n17 VGND.n16 2.63579
R122 VGND.n25 VGND.n23 1.88285
R123 VGND.n11 VGND.n8 0.663075
R124 VGND.n40 VGND.n0 0.148519
R125 VGND.n12 VGND.n11 0.120292
R126 VGND.n13 VGND.n12 0.120292
R127 VGND.n13 VGND.n6 0.120292
R128 VGND.n19 VGND.n6 0.120292
R129 VGND.n20 VGND.n19 0.120292
R130 VGND.n21 VGND.n20 0.120292
R131 VGND.n21 VGND.n4 0.120292
R132 VGND.n27 VGND.n4 0.120292
R133 VGND.n28 VGND.n27 0.120292
R134 VGND.n29 VGND.n28 0.120292
R135 VGND.n29 VGND.n2 0.120292
R136 VGND.n33 VGND.n2 0.120292
R137 VGND.n34 VGND.n33 0.120292
R138 VGND.n35 VGND.n34 0.120292
R139 VGND.n35 VGND.n0 0.120292
R140 VGND VGND.n40 0.114842
R141 a_1462_47.t0 a_1462_47.t1 87.1434
R142 a_543_47.n3 a_543_47.n2 674.338
R143 a_543_47.n1 a_543_47.t5 332.58
R144 a_543_47.n2 a_543_47.n0 284.012
R145 a_543_47.n2 a_543_47.n1 253.648
R146 a_543_47.n1 a_543_47.t4 168.701
R147 a_543_47.n3 a_543_47.t2 96.1553
R148 a_543_47.t0 a_543_47.n3 65.6672
R149 a_543_47.n0 a_543_47.t1 65.0005
R150 a_543_47.n0 a_543_47.t3 45.0005
R151 a_651_413.n0 a_651_413.t1 1327.82
R152 a_651_413.n0 a_651_413.t2 194.655
R153 a_651_413.t0 a_651_413.n0 63.3219
R154 VPB.t11 VPB.t0 790.188
R155 VPB.t9 VPB.t5 636.293
R156 VPB.t7 VPB.t10 583.023
R157 VPB.t13 VPB.t2 414.33
R158 VPB.t4 VPB.t8 319.627
R159 VPB.t10 VPB.t12 292.991
R160 VPB.t1 VPB.t13 292.991
R161 VPB.t2 VPB.t7 287.072
R162 VPB.t0 VPB.t1 272.274
R163 VPB.t12 VPB.t14 254.518
R164 VPB.t5 VPB.t6 248.599
R165 VPB.t8 VPB.t9 248.599
R166 VPB.t14 VPB.t4 248.599
R167 VPB.t3 VPB.t11 248.599
R168 VPB VPB.t3 192.369
R169 VPWR.n23 VPWR.t9 806.511
R170 VPWR.n2 VPWR.t0 667.778
R171 VPWR.n10 VPWR.t8 667.751
R172 VPWR.n17 VPWR.n9 604.457
R173 VPWR.n39 VPWR.n1 604.394
R174 VPWR.n26 VPWR.n25 601.679
R175 VPWR.n12 VPWR.t3 343.579
R176 VPWR.n11 VPWR.t4 257.204
R177 VPWR.n9 VPWR.t5 119.608
R178 VPWR.n25 VPWR.t1 93.81
R179 VPWR.n25 VPWR.t6 63.3219
R180 VPWR.n9 VPWR.t7 63.3219
R181 VPWR.n1 VPWR.t10 41.5552
R182 VPWR.n1 VPWR.t2 41.5552
R183 VPWR.n38 VPWR.n37 34.6358
R184 VPWR.n31 VPWR.n4 34.6358
R185 VPWR.n32 VPWR.n31 34.6358
R186 VPWR.n33 VPWR.n32 34.6358
R187 VPWR.n27 VPWR.n24 34.6358
R188 VPWR.n18 VPWR.n7 34.6358
R189 VPWR.n22 VPWR.n7 34.6358
R190 VPWR.n33 VPWR.n2 32.377
R191 VPWR.n23 VPWR.n22 32.0005
R192 VPWR.n17 VPWR.n16 30.1181
R193 VPWR.n13 VPWR.n12 24.8476
R194 VPWR.n39 VPWR.n38 22.9652
R195 VPWR.n18 VPWR.n17 20.3299
R196 VPWR.n37 VPWR.n2 18.0711
R197 VPWR.n24 VPWR.n23 9.41227
R198 VPWR.n14 VPWR.n13 9.3005
R199 VPWR.n16 VPWR.n15 9.3005
R200 VPWR.n17 VPWR.n8 9.3005
R201 VPWR.n19 VPWR.n18 9.3005
R202 VPWR.n20 VPWR.n7 9.3005
R203 VPWR.n22 VPWR.n21 9.3005
R204 VPWR.n23 VPWR.n6 9.3005
R205 VPWR.n24 VPWR.n5 9.3005
R206 VPWR.n28 VPWR.n27 9.3005
R207 VPWR.n29 VPWR.n4 9.3005
R208 VPWR.n31 VPWR.n30 9.3005
R209 VPWR.n32 VPWR.n3 9.3005
R210 VPWR.n34 VPWR.n33 9.3005
R211 VPWR.n35 VPWR.n2 9.3005
R212 VPWR.n37 VPWR.n36 9.3005
R213 VPWR.n38 VPWR.n0 9.3005
R214 VPWR.n16 VPWR.n10 9.03579
R215 VPWR.n40 VPWR.n39 7.12063
R216 VPWR.n12 VPWR.n11 6.48892
R217 VPWR.n26 VPWR.n4 6.02403
R218 VPWR.n27 VPWR.n26 3.76521
R219 VPWR.n13 VPWR.n10 0.753441
R220 VPWR.n14 VPWR.n11 0.663075
R221 VPWR.n40 VPWR.n0 0.148519
R222 VPWR.n15 VPWR.n14 0.120292
R223 VPWR.n15 VPWR.n8 0.120292
R224 VPWR.n19 VPWR.n8 0.120292
R225 VPWR.n20 VPWR.n19 0.120292
R226 VPWR.n21 VPWR.n20 0.120292
R227 VPWR.n21 VPWR.n6 0.120292
R228 VPWR.n6 VPWR.n5 0.120292
R229 VPWR.n28 VPWR.n5 0.120292
R230 VPWR.n29 VPWR.n28 0.120292
R231 VPWR.n30 VPWR.n29 0.120292
R232 VPWR.n30 VPWR.n3 0.120292
R233 VPWR.n34 VPWR.n3 0.120292
R234 VPWR.n35 VPWR.n34 0.120292
R235 VPWR.n36 VPWR.n35 0.120292
R236 VPWR.n36 VPWR.n0 0.120292
R237 VPWR VPWR.n40 0.114842
R238 a_193_47.t0 a_193_47.n3 370.026
R239 a_193_47.n0 a_193_47.t2 351.356
R240 a_193_47.n1 a_193_47.t5 334.717
R241 a_193_47.n3 a_193_47.t1 325.971
R242 a_193_47.n1 a_193_47.t3 309.935
R243 a_193_47.n0 a_193_47.t4 305.683
R244 a_193_47.n2 a_193_47.n0 16.879
R245 a_193_47.n3 a_193_47.n2 10.8867
R246 a_193_47.n2 a_193_47.n1 9.3005
R247 RESET_B.n1 RESET_B.t3 408.63
R248 RESET_B.n3 RESET_B.t2 347.577
R249 RESET_B.n3 RESET_B.t1 193.337
R250 RESET_B.n2 RESET_B.n1 167.575
R251 RESET_B.n4 RESET_B.n3 152
R252 RESET_B.n1 RESET_B.t0 132.282
R253 RESET_B RESET_B.n0 14.0185
R254 RESET_B.n4 RESET_B.n2 12.1952
R255 RESET_B.n2 RESET_B.n0 9.38606
R256 RESET_B RESET_B.n4 4.67077
R257 RESET_B.n0 RESET_B 4.53383
R258 CLK.n0 CLK.t0 294.557
R259 CLK.n0 CLK.t1 211.01
R260 CLK.n1 CLK.n0 152
R261 CLK.n1 CLK 10.4234
R262 CLK CLK.n1 2.01193
R263 D.n0 D.t1 333.651
R264 D.n0 D.t0 297.233
R265 D D.n0 196.737
R266 a_448_47.n1 a_448_47.n0 926.024
R267 a_448_47.n1 a_448_47.t2 82.0838
R268 a_448_47.n0 a_448_47.t3 63.3338
R269 a_448_47.t0 a_448_47.n1 63.3219
R270 a_448_47.n0 a_448_47.t1 29.7268
R271 a_1270_413.t0 a_1270_413.t1 126.644
C0 RESET_B VGND 0.288034f
C1 VPWR VGND 0.071912f
C2 RESET_B Q 8.96e-19
C3 VPWR Q 0.169355f
C4 VGND Q 0.109665f
C5 VPB CLK 0.069345f
C6 VPB D 0.137565f
C7 VPB RESET_B 0.138482f
C8 VPB VPWR 0.233696f
C9 CLK RESET_B 1.09e-19
C10 CLK VPWR 0.017406f
C11 VPB VGND 0.012153f
C12 D RESET_B 4.72e-19
C13 D VPWR 0.081188f
C14 VPB Q 0.005549f
C15 CLK VGND 0.017208f
C16 D VGND 0.051614f
C17 RESET_B VPWR 0.065186f
C18 Q VNB 0.029557f
C19 VGND VNB 1.09584f
C20 VPWR VNB 0.902284f
C21 RESET_B VNB 0.262848f
C22 D VNB 0.159894f
C23 CLK VNB 0.195254f
C24 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47.t0 a_27_47.t2 a_1108_47.t1 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21.t2 a_1108_47.t4 a_1462_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413.t0 a_27_47.t3 a_543_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47.t2 a_193_47.t2 a_761_289.t1 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND.t4 RESET_B.t0 a_805_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR.t11 a_1283_21.t3 Q.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47.t3 D.t0 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 Q.t6 a_1283_21.t4 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t9 a_1283_21.t5 Q.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289.t2 a_543_47.t4 VGND.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 Q.t3 a_1283_21.t6 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47.t0 a_27_47.t4 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47.t0 a_27_47.t5 a_761_289.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 a_1462_47.t0 RESET_B.t1 VGND.t5 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47.t0 a_27_47.t6 a_448_47.t0 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_543_47.t2 a_193_47.t3 a_448_47.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47.t2 D.t1 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X19 VPWR.t7 a_1283_21.t7 a_1270_413.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR.t12 a_1108_47.t5 a_1283_21.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q.t4 a_1283_21.t8 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413.t0 a_193_47.t4 a_1108_47.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47.t1 a_27_47.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21.t0 RESET_B.t2 VPWR.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND.t6 a_1283_21.t9 Q.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VGND.t8 a_1283_21.t10 Q.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR.t1 a_761_289.t5 a_651_413.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 a_639_47.t1 a_193_47.t5 a_543_47.t3 VNB.t16 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND.t10 a_1283_21.t11 a_1217_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413.t2 RESET_B.t3 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X31 VGND.t3 CLK.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_761_289.t3 a_543_47.t5 VPWR.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X33 Q.t0 a_1283_21.t12 VGND.t9 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_761_289.n3 a_761_289.n2 647.119
R1 a_761_289.n1 a_761_289.t4 350.253
R2 a_761_289.n2 a_761_289.n0 260.339
R3 a_761_289.n2 a_761_289.n1 246.119
R4 a_761_289.n1 a_761_289.t5 189.588
R5 a_761_289.n3 a_761_289.t0 89.1195
R6 a_761_289.n0 a_761_289.t1 63.3338
R7 a_761_289.t3 a_761_289.n3 41.0422
R8 a_761_289.n0 a_761_289.t2 31.9797
R9 a_639_47.t0 a_639_47.t1 198.571
R10 a_805_47.t0 a_805_47.t1 60.0005
R11 VNB.t3 VNB.t6 3631.07
R12 VNB.t9 VNB.t10 2677.02
R13 VNB.t16 VNB.t0 2363.75
R14 VNB.t13 VNB.t15 2121.68
R15 VNB.t1 VNB.t8 1879.61
R16 VNB.t5 VNB.t2 1552.1
R17 VNB.t8 VNB.t5 1409.71
R18 VNB.t2 VNB.t13 1366.99
R19 VNB.t4 VNB.t16 1366.99
R20 VNB.t6 VNB.t4 1352.75
R21 VNB.t15 VNB.t9 1295.79
R22 VNB.t14 VNB.t12 1196.12
R23 VNB.t11 VNB.t14 1196.12
R24 VNB.t10 VNB.t11 1196.12
R25 VNB.t7 VNB.t3 1196.12
R26 VNB.t0 VNB.t1 1025.24
R27 VNB VNB.t7 925.567
R28 a_27_47.n1 a_27_47.t3 530.01
R29 a_27_47.t0 a_27_47.n5 421.021
R30 a_27_47.n0 a_27_47.t5 337.142
R31 a_27_47.n3 a_27_47.t1 280.223
R32 a_27_47.n4 a_27_47.t7 263.173
R33 a_27_47.n4 a_27_47.t4 227.826
R34 a_27_47.n0 a_27_47.t2 199.762
R35 a_27_47.n2 a_27_47.n1 170.81
R36 a_27_47.n2 a_27_47.n0 167.321
R37 a_27_47.n5 a_27_47.n4 152
R38 a_27_47.n1 a_27_47.t6 141.923
R39 a_27_47.n3 a_27_47.n2 10.8376
R40 a_27_47.n5 a_27_47.n3 2.50485
R41 a_1108_47.n3 a_1108_47.n2 636.953
R42 a_1108_47.n1 a_1108_47.t4 366.856
R43 a_1108_47.n2 a_1108_47.n0 300.2
R44 a_1108_47.n2 a_1108_47.n1 225.036
R45 a_1108_47.n1 a_1108_47.t5 174.056
R46 a_1108_47.n0 a_1108_47.t2 70.0005
R47 a_1108_47.t0 a_1108_47.n3 68.0124
R48 a_1108_47.n3 a_1108_47.t3 63.3219
R49 a_1108_47.n0 a_1108_47.t1 61.6672
R50 a_1217_47.t1 a_1217_47.t0 94.7268
R51 a_1462_47.t0 a_1462_47.t1 87.1434
R52 a_1283_21.n14 a_1283_21.n13 692.797
R53 a_1283_21.n11 a_1283_21.t7 389.183
R54 a_1283_21.n12 a_1283_21.n11 251.167
R55 a_1283_21.n12 a_1283_21.t2 223.571
R56 a_1283_21.n2 a_1283_21.t3 212.081
R57 a_1283_21.n1 a_1283_21.t4 212.081
R58 a_1283_21.n6 a_1283_21.t5 212.081
R59 a_1283_21.n8 a_1283_21.t8 212.081
R60 a_1283_21.n11 a_1283_21.t11 174.891
R61 a_1283_21.n4 a_1283_21.n3 172.725
R62 a_1283_21.n10 a_1283_21.n9 152
R63 a_1283_21.n7 a_1283_21.n0 152
R64 a_1283_21.n5 a_1283_21.n4 152
R65 a_1283_21.n2 a_1283_21.t10 139.78
R66 a_1283_21.n1 a_1283_21.t12 139.78
R67 a_1283_21.n6 a_1283_21.t9 139.78
R68 a_1283_21.n8 a_1283_21.t6 139.78
R69 a_1283_21.n14 a_1283_21.t1 63.3219
R70 a_1283_21.t0 a_1283_21.n14 63.3219
R71 a_1283_21.n9 a_1283_21.n7 49.6611
R72 a_1283_21.n6 a_1283_21.n5 42.3581
R73 a_1283_21.n3 a_1283_21.n2 30.6732
R74 a_1283_21.n3 a_1283_21.n1 30.6732
R75 a_1283_21.n13 a_1283_21.n10 30.4767
R76 a_1283_21.n13 a_1283_21.n12 28.3392
R77 a_1283_21.n4 a_1283_21.n0 20.7243
R78 a_1283_21.n10 a_1283_21.n0 20.7243
R79 a_1283_21.n5 a_1283_21.n1 18.9884
R80 a_1283_21.n7 a_1283_21.n6 7.30353
R81 a_1283_21.n9 a_1283_21.n8 4.38232
R82 a_543_47.n3 a_543_47.n2 674.338
R83 a_543_47.n1 a_543_47.t5 332.58
R84 a_543_47.n2 a_543_47.n0 284.012
R85 a_543_47.n2 a_543_47.n1 253.648
R86 a_543_47.n1 a_543_47.t4 168.701
R87 a_543_47.t1 a_543_47.n3 96.1553
R88 a_543_47.n3 a_543_47.t2 65.6672
R89 a_543_47.n0 a_543_47.t0 65.0005
R90 a_543_47.n0 a_543_47.t3 45.0005
R91 a_651_413.n0 a_651_413.t2 1327.82
R92 a_651_413.t0 a_651_413.n0 194.655
R93 a_651_413.n0 a_651_413.t1 63.3219
R94 VPB.t0 VPB.t10 790.188
R95 VPB.t5 VPB.t7 583.023
R96 VPB.t16 VPB.t11 577.104
R97 VPB.t2 VPB.t3 414.33
R98 VPB.t12 VPB.t4 319.627
R99 VPB.t7 VPB.t1 292.991
R100 VPB.t6 VPB.t2 292.991
R101 VPB.t3 VPB.t5 287.072
R102 VPB.t10 VPB.t6 272.274
R103 VPB.t1 VPB.t9 254.518
R104 VPB.t14 VPB.t15 248.599
R105 VPB.t13 VPB.t14 248.599
R106 VPB.t11 VPB.t13 248.599
R107 VPB.t4 VPB.t16 248.599
R108 VPB.t9 VPB.t12 248.599
R109 VPB.t8 VPB.t0 248.599
R110 VPB VPB.t8 192.369
R111 a_193_47.t1 a_193_47.n3 370.026
R112 a_193_47.n0 a_193_47.t2 351.356
R113 a_193_47.n1 a_193_47.t5 334.717
R114 a_193_47.n3 a_193_47.t0 325.971
R115 a_193_47.n1 a_193_47.t3 309.935
R116 a_193_47.n0 a_193_47.t4 305.683
R117 a_193_47.n2 a_193_47.n0 16.879
R118 a_193_47.n3 a_193_47.n2 10.8867
R119 a_193_47.n2 a_193_47.n1 9.3005
R120 RESET_B.n1 RESET_B.t3 408.63
R121 RESET_B.n3 RESET_B.t2 347.577
R122 RESET_B.n3 RESET_B.t1 193.337
R123 RESET_B.n2 RESET_B.n1 167.575
R124 RESET_B.n4 RESET_B.n3 152
R125 RESET_B.n1 RESET_B.t0 132.282
R126 RESET_B RESET_B.n0 14.0185
R127 RESET_B.n4 RESET_B.n2 12.1952
R128 RESET_B.n2 RESET_B.n0 9.38606
R129 RESET_B RESET_B.n4 4.67077
R130 RESET_B.n0 RESET_B 4.53383
R131 VGND.n42 VGND.t2 307.536
R132 VGND.n11 VGND.t8 292.839
R133 VGND.n22 VGND.n21 209.254
R134 VGND.n10 VGND.n9 207.965
R135 VGND.n31 VGND.n30 199.739
R136 VGND.n45 VGND.n44 199.739
R137 VGND.n15 VGND.t7 160.8
R138 VGND.n21 VGND.t5 100.001
R139 VGND.n30 VGND.t4 72.8576
R140 VGND.n21 VGND.t10 70.0005
R141 VGND.n30 VGND.t1 60.5809
R142 VGND.n44 VGND.t0 38.5719
R143 VGND.n44 VGND.t3 38.5719
R144 VGND.n14 VGND.n13 34.6358
R145 VGND.n16 VGND.n7 34.6358
R146 VGND.n20 VGND.n7 34.6358
R147 VGND.n24 VGND.n23 34.6358
R148 VGND.n24 VGND.n5 34.6358
R149 VGND.n28 VGND.n5 34.6358
R150 VGND.n29 VGND.n28 34.6358
R151 VGND.n32 VGND.n3 34.6358
R152 VGND.n36 VGND.n3 34.6358
R153 VGND.n37 VGND.n36 34.6358
R154 VGND.n38 VGND.n37 34.6358
R155 VGND.n38 VGND.n1 34.6358
R156 VGND.n43 VGND.n42 29.7417
R157 VGND.n16 VGND.n15 27.8593
R158 VGND.n9 VGND.t9 24.9236
R159 VGND.n9 VGND.t6 24.9236
R160 VGND.n45 VGND.n43 22.9652
R161 VGND.n13 VGND.n10 21.8358
R162 VGND.n11 VGND.n10 19.5226
R163 VGND.n22 VGND.n20 17.6946
R164 VGND.n42 VGND.n1 14.6829
R165 VGND.n43 VGND.n0 9.3005
R166 VGND.n42 VGND.n41 9.3005
R167 VGND.n40 VGND.n1 9.3005
R168 VGND.n39 VGND.n38 9.3005
R169 VGND.n37 VGND.n2 9.3005
R170 VGND.n36 VGND.n35 9.3005
R171 VGND.n34 VGND.n3 9.3005
R172 VGND.n33 VGND.n32 9.3005
R173 VGND.n13 VGND.n12 9.3005
R174 VGND.n14 VGND.n8 9.3005
R175 VGND.n17 VGND.n16 9.3005
R176 VGND.n18 VGND.n7 9.3005
R177 VGND.n20 VGND.n19 9.3005
R178 VGND.n23 VGND.n6 9.3005
R179 VGND.n25 VGND.n24 9.3005
R180 VGND.n26 VGND.n5 9.3005
R181 VGND.n28 VGND.n27 9.3005
R182 VGND.n29 VGND.n4 9.3005
R183 VGND.n32 VGND.n31 7.90638
R184 VGND.n46 VGND.n45 7.12063
R185 VGND.n15 VGND.n14 6.77697
R186 VGND.n23 VGND.n22 2.63579
R187 VGND.n31 VGND.n29 1.88285
R188 VGND.n12 VGND.n11 1.02737
R189 VGND.n46 VGND.n0 0.148519
R190 VGND.n12 VGND.n8 0.120292
R191 VGND.n17 VGND.n8 0.120292
R192 VGND.n18 VGND.n17 0.120292
R193 VGND.n19 VGND.n18 0.120292
R194 VGND.n19 VGND.n6 0.120292
R195 VGND.n25 VGND.n6 0.120292
R196 VGND.n26 VGND.n25 0.120292
R197 VGND.n27 VGND.n26 0.120292
R198 VGND.n27 VGND.n4 0.120292
R199 VGND.n33 VGND.n4 0.120292
R200 VGND.n34 VGND.n33 0.120292
R201 VGND.n35 VGND.n34 0.120292
R202 VGND.n35 VGND.n2 0.120292
R203 VGND.n39 VGND.n2 0.120292
R204 VGND.n40 VGND.n39 0.120292
R205 VGND.n41 VGND.n40 0.120292
R206 VGND.n41 VGND.n0 0.120292
R207 VGND VGND.n46 0.114842
R208 Q.n2 Q.n0 248.088
R209 Q.n2 Q.n1 208.507
R210 Q.n5 Q.n3 137.576
R211 Q.n5 Q.n4 99.1759
R212 Q.n0 Q.t5 26.5955
R213 Q.n0 Q.t4 26.5955
R214 Q.n1 Q.t7 26.5955
R215 Q.n1 Q.t6 26.5955
R216 Q.n3 Q.t2 24.9236
R217 Q.n3 Q.t3 24.9236
R218 Q.n4 Q.t1 24.9236
R219 Q.n4 Q.t0 24.9236
R220 Q Q.n5 22.8275
R221 Q Q.n2 19.9075
R222 VPWR.n29 VPWR.t2 806.511
R223 VPWR.n2 VPWR.t6 667.778
R224 VPWR.n10 VPWR.t12 667.751
R225 VPWR.n23 VPWR.n9 604.457
R226 VPWR.n45 VPWR.n1 604.394
R227 VPWR.n32 VPWR.n31 601.679
R228 VPWR.n14 VPWR.t11 362.599
R229 VPWR.n18 VPWR.t8 347.572
R230 VPWR.n13 VPWR.n12 323.988
R231 VPWR.n9 VPWR.t7 119.608
R232 VPWR.n31 VPWR.t1 93.81
R233 VPWR.n31 VPWR.t4 63.3219
R234 VPWR.n9 VPWR.t5 63.3219
R235 VPWR.n1 VPWR.t0 41.5552
R236 VPWR.n1 VPWR.t3 41.5552
R237 VPWR.n44 VPWR.n43 34.6358
R238 VPWR.n37 VPWR.n4 34.6358
R239 VPWR.n38 VPWR.n37 34.6358
R240 VPWR.n39 VPWR.n38 34.6358
R241 VPWR.n33 VPWR.n30 34.6358
R242 VPWR.n24 VPWR.n7 34.6358
R243 VPWR.n28 VPWR.n7 34.6358
R244 VPWR.n17 VPWR.n16 34.6358
R245 VPWR.n39 VPWR.n2 32.377
R246 VPWR.n29 VPWR.n28 32.0005
R247 VPWR.n23 VPWR.n22 30.1181
R248 VPWR.n19 VPWR.n18 27.8593
R249 VPWR.n12 VPWR.t10 26.5955
R250 VPWR.n12 VPWR.t9 26.5955
R251 VPWR.n45 VPWR.n44 22.9652
R252 VPWR.n16 VPWR.n13 21.8358
R253 VPWR.n24 VPWR.n23 20.3299
R254 VPWR.n14 VPWR.n13 19.5226
R255 VPWR.n43 VPWR.n2 18.0711
R256 VPWR.n30 VPWR.n29 9.41227
R257 VPWR.n16 VPWR.n15 9.3005
R258 VPWR.n17 VPWR.n11 9.3005
R259 VPWR.n20 VPWR.n19 9.3005
R260 VPWR.n22 VPWR.n21 9.3005
R261 VPWR.n23 VPWR.n8 9.3005
R262 VPWR.n25 VPWR.n24 9.3005
R263 VPWR.n26 VPWR.n7 9.3005
R264 VPWR.n28 VPWR.n27 9.3005
R265 VPWR.n29 VPWR.n6 9.3005
R266 VPWR.n30 VPWR.n5 9.3005
R267 VPWR.n34 VPWR.n33 9.3005
R268 VPWR.n35 VPWR.n4 9.3005
R269 VPWR.n37 VPWR.n36 9.3005
R270 VPWR.n38 VPWR.n3 9.3005
R271 VPWR.n40 VPWR.n39 9.3005
R272 VPWR.n41 VPWR.n2 9.3005
R273 VPWR.n43 VPWR.n42 9.3005
R274 VPWR.n44 VPWR.n0 9.3005
R275 VPWR.n22 VPWR.n10 9.03579
R276 VPWR.n46 VPWR.n45 7.12063
R277 VPWR.n18 VPWR.n17 6.77697
R278 VPWR.n32 VPWR.n4 6.02403
R279 VPWR.n33 VPWR.n32 3.76521
R280 VPWR.n15 VPWR.n14 1.02737
R281 VPWR.n19 VPWR.n10 0.753441
R282 VPWR.n46 VPWR.n0 0.148519
R283 VPWR.n15 VPWR.n11 0.120292
R284 VPWR.n20 VPWR.n11 0.120292
R285 VPWR.n21 VPWR.n20 0.120292
R286 VPWR.n21 VPWR.n8 0.120292
R287 VPWR.n25 VPWR.n8 0.120292
R288 VPWR.n26 VPWR.n25 0.120292
R289 VPWR.n27 VPWR.n26 0.120292
R290 VPWR.n27 VPWR.n6 0.120292
R291 VPWR.n6 VPWR.n5 0.120292
R292 VPWR.n34 VPWR.n5 0.120292
R293 VPWR.n35 VPWR.n34 0.120292
R294 VPWR.n36 VPWR.n35 0.120292
R295 VPWR.n36 VPWR.n3 0.120292
R296 VPWR.n40 VPWR.n3 0.120292
R297 VPWR.n41 VPWR.n40 0.120292
R298 VPWR.n42 VPWR.n41 0.120292
R299 VPWR.n42 VPWR.n0 0.120292
R300 VPWR VPWR.n46 0.114842
R301 CLK.n0 CLK.t0 294.557
R302 CLK.n0 CLK.t1 211.01
R303 CLK.n1 CLK.n0 152
R304 CLK.n1 CLK 10.4234
R305 CLK CLK.n1 2.01193
R306 D.n0 D.t1 333.651
R307 D.n0 D.t0 297.233
R308 D D.n0 196.737
R309 a_448_47.n1 a_448_47.n0 926.024
R310 a_448_47.t1 a_448_47.n1 82.0838
R311 a_448_47.n0 a_448_47.t0 63.3338
R312 a_448_47.n1 a_448_47.t3 63.3219
R313 a_448_47.n0 a_448_47.t2 29.7268
R314 a_1270_413.t0 a_1270_413.t1 126.644
C0 VGND CLK 0.017208f
C1 Q VPB 0.017629f
C2 RESET_B VPWR 0.065186f
C3 VGND D 0.051614f
C4 VGND RESET_B 0.288033f
C5 Q RESET_B 0.001878f
C6 VGND VPWR 0.077885f
C7 Q VPWR 0.3679f
C8 VPB CLK 0.069345f
C9 VGND Q 0.295568f
C10 VPB D 0.137565f
C11 VPB RESET_B 0.138482f
C12 VPB VPWR 0.242331f
C13 CLK RESET_B 1.09e-19
C14 D RESET_B 4.72e-19
C15 CLK VPWR 0.017406f
C16 VGND VPB 0.012277f
C17 D VPWR 0.081188f
C18 Q VNB 0.061504f
C19 VGND VNB 1.18004f
C20 VPWR VNB 0.977124f
C21 RESET_B VNB 0.260102f
C22 D VNB 0.159894f
C23 CLK VNB 0.195254f
C24 VPB VNB 2.1109f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfsbp_1 VPB VNB VGND VPWR Q Q_N SET_B D CLK
X0 a_1178_261.t0 a_1028_413.t5 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X1 VGND.t8 a_652_21.t3 a_586_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X2 a_1178_261.t1 a_1028_413.t6 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X3 a_956_413.t1 a_476_47.t4 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1136_413.t1 a_193_47.t2 a_1028_413.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X5 VPWR.t4 a_476_47.t5 a_652_21.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR.t10 CLK.t0 a_27_47.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_586_47.t0 a_193_47.t3 a_476_47.t3 VNB.t13 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X8 a_1056_47.t0 a_476_47.t6 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_476_47.t0 a_27_47.t2 a_381_47.t3 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X10 a_381_47.t2 D.t0 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X11 a_652_21.t2 SET_B.t0 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X12 a_1224_47.t1 a_27_47.t3 a_1028_413.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 VGND.t3 a_1028_413.t7 a_1786_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_562_413.t0 a_27_47.t4 a_476_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VPWR.t2 a_1028_413.t8 a_1786_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 a_1028_413.t2 a_193_47.t4 a_1056_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47.t2 a_193_47.t5 a_381_47.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X18 a_1296_47.t1 a_1178_261.t2 a_1224_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 Q_N.t1 a_1028_413.t9 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X20 a_193_47.t0 a_27_47.t5 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR.t6 a_652_21.t4 a_562_413.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X22 VGND.t9 SET_B.t1 a_1296_47.t0 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 a_1028_413.t1 a_27_47.t6 a_956_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 VPWR.t5 a_1178_261.t3 a_1136_413.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 a_193_47.t1 a_27_47.t7 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 Q_N.t0 a_1028_413.t10 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X27 a_796_47.t0 SET_B.t2 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X28 a_381_47.t0 D.t1 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 a_652_21.t1 a_476_47.t7 a_796_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VPWR.t11 SET_B.t3 a_1028_413.t4 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND.t4 CLK.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1028_413.n5 a_1028_413.t4 724.652
R1 a_1028_413.n5 a_1028_413.n4 611.504
R2 a_1028_413.n7 a_1028_413.n6 287.401
R3 a_1028_413.n3 a_1028_413.t5 258.673
R4 a_1028_413.n0 a_1028_413.t8 257.182
R5 a_1028_413.n1 a_1028_413.t10 221.72
R6 a_1028_413.n6 a_1028_413.n3 217.255
R7 a_1028_413.n2 a_1028_413.t6 210.474
R8 a_1028_413.n0 a_1028_413.t7 163.995
R9 a_1028_413.n2 a_1028_413.n1 154.419
R10 a_1028_413.n1 a_1028_413.t9 149.421
R11 a_1028_413.n1 a_1028_413.n0 144.601
R12 a_1028_413.n4 a_1028_413.t3 119.608
R13 a_1028_413.n6 a_1028_413.n5 93.3652
R14 a_1028_413.n4 a_1028_413.t1 63.3219
R15 a_1028_413.t0 a_1028_413.n7 47.1434
R16 a_1028_413.n7 a_1028_413.t2 47.1434
R17 a_1028_413.n3 a_1028_413.n2 32.1338
R18 VPWR.n36 VPWR.t7 721.837
R19 VPWR.n8 VPWR.t5 648.322
R20 VPWR.n16 VPWR.n11 604.783
R21 VPWR.n38 VPWR.n1 604.394
R22 VPWR.n6 VPWR.n5 599.74
R23 VPWR.n29 VPWR.n28 585
R24 VPWR.n13 VPWR.t2 390.272
R25 VPWR.n12 VPWR.t0 261.553
R26 VPWR.n28 VPWR.t8 91.4648
R27 VPWR.n11 VPWR.t11 91.4648
R28 VPWR.n28 VPWR.t6 86.7743
R29 VPWR.n5 VPWR.t3 63.3219
R30 VPWR.n5 VPWR.t4 63.3219
R31 VPWR.n1 VPWR.t9 41.5552
R32 VPWR.n1 VPWR.t10 41.5552
R33 VPWR.n31 VPWR.n3 34.6358
R34 VPWR.n35 VPWR.n3 34.6358
R35 VPWR.n22 VPWR.n21 34.6358
R36 VPWR.n23 VPWR.n22 34.6358
R37 VPWR.n31 VPWR.n30 33.5954
R38 VPWR.n11 VPWR.t1 32.8338
R39 VPWR.n15 VPWR.n12 32.377
R40 VPWR.n27 VPWR.n6 31.624
R41 VPWR.n18 VPWR.n17 27.873
R42 VPWR.n17 VPWR.n16 25.6005
R43 VPWR.n37 VPWR.n36 22.9652
R44 VPWR.n38 VPWR.n37 22.9652
R45 VPWR.n36 VPWR.n35 21.4593
R46 VPWR.n21 VPWR.n8 19.2553
R47 VPWR.n16 VPWR.n15 18.824
R48 VPWR.n23 VPWR.n6 12.8005
R49 VPWR.n29 VPWR.n27 12.5335
R50 VPWR.n15 VPWR.n14 9.3005
R51 VPWR.n16 VPWR.n10 9.3005
R52 VPWR.n17 VPWR.n9 9.3005
R53 VPWR.n19 VPWR.n18 9.3005
R54 VPWR.n21 VPWR.n20 9.3005
R55 VPWR.n22 VPWR.n7 9.3005
R56 VPWR.n24 VPWR.n23 9.3005
R57 VPWR.n25 VPWR.n6 9.3005
R58 VPWR.n27 VPWR.n26 9.3005
R59 VPWR.n30 VPWR.n4 9.3005
R60 VPWR.n32 VPWR.n31 9.3005
R61 VPWR.n33 VPWR.n3 9.3005
R62 VPWR.n35 VPWR.n34 9.3005
R63 VPWR.n36 VPWR.n2 9.3005
R64 VPWR.n37 VPWR.n0 9.3005
R65 VPWR.n39 VPWR.n38 7.12063
R66 VPWR.n13 VPWR.n12 7.07919
R67 VPWR.n30 VPWR.n29 3.37505
R68 VPWR.n18 VPWR.n8 0.815045
R69 VPWR.n14 VPWR.n13 0.201153
R70 VPWR.n39 VPWR.n0 0.148519
R71 VPWR.n14 VPWR.n10 0.120292
R72 VPWR.n10 VPWR.n9 0.120292
R73 VPWR.n19 VPWR.n9 0.120292
R74 VPWR.n20 VPWR.n19 0.120292
R75 VPWR.n20 VPWR.n7 0.120292
R76 VPWR.n24 VPWR.n7 0.120292
R77 VPWR.n25 VPWR.n24 0.120292
R78 VPWR.n26 VPWR.n25 0.120292
R79 VPWR.n26 VPWR.n4 0.120292
R80 VPWR.n32 VPWR.n4 0.120292
R81 VPWR.n33 VPWR.n32 0.120292
R82 VPWR.n34 VPWR.n33 0.120292
R83 VPWR.n34 VPWR.n2 0.120292
R84 VPWR.n2 VPWR.n0 0.120292
R85 VPWR VPWR.n39 0.0927068
R86 a_1178_261.n0 a_1178_261.t2 372.274
R87 a_1178_261.t0 a_1178_261.n1 371.185
R88 a_1178_261.n1 a_1178_261.t1 291.327
R89 a_1178_261.n1 a_1178_261.n0 264.267
R90 a_1178_261.n0 a_1178_261.t3 167.992
R91 VPB.t2 VPB.t3 556.386
R92 VPB.t4 VPB.t2 556.386
R93 VPB.t5 VPB.t15 556.386
R94 VPB.t13 VPB.t10 556.386
R95 VPB.t0 VPB.t9 355.14
R96 VPB.t1 VPB.t12 319.627
R97 VPB.t9 VPB.t11 313.707
R98 VPB.t10 VPB.t8 287.072
R99 VPB.t15 VPB.t4 284.113
R100 VPB.t7 VPB.t6 248.599
R101 VPB.t11 VPB.t7 248.599
R102 VPB.t8 VPB.t0 248.599
R103 VPB.t14 VPB.t13 248.599
R104 VPB.t12 VPB.t5 213.084
R105 VPB.t6 VPB.t1 213.084
R106 VPB VPB.t14 142.056
R107 a_652_21.n2 a_652_21.n1 594.413
R108 a_652_21.n0 a_652_21.t3 387.961
R109 a_652_21.n1 a_652_21.t1 334.156
R110 a_652_21.n1 a_652_21.n0 187.072
R111 a_652_21.n0 a_652_21.t4 143.746
R112 a_652_21.t0 a_652_21.n2 63.3219
R113 a_652_21.n2 a_652_21.t2 63.3219
R114 a_586_47.t1 a_586_47.t0 93.5174
R115 VGND.n34 VGND.t7 280.51
R116 VGND.n11 VGND.t3 272.31
R117 VGND.n23 VGND.t5 237.877
R118 VGND.n37 VGND.n36 199.739
R119 VGND.n9 VGND.n8 185
R120 VGND.n4 VGND.n3 185
R121 VGND.n12 VGND.t2 165.714
R122 VGND.n3 VGND.t8 81.4291
R123 VGND.n8 VGND.t9 67.1434
R124 VGND.n8 VGND.t1 55.3018
R125 VGND.n3 VGND.t6 38.5719
R126 VGND.n36 VGND.t0 38.5719
R127 VGND.n36 VGND.t4 38.5719
R128 VGND.n18 VGND.n17 34.6358
R129 VGND.n19 VGND.n18 34.6358
R130 VGND.n19 VGND.n6 34.6358
R131 VGND.n29 VGND.n28 34.6358
R132 VGND.n30 VGND.n29 34.6358
R133 VGND.n30 VGND.n1 34.6358
R134 VGND.n13 VGND.n12 32.377
R135 VGND.n25 VGND.n24 28.6616
R136 VGND.n24 VGND.n23 27.8593
R137 VGND.n14 VGND.n13 23.5154
R138 VGND.n35 VGND.n34 22.9652
R139 VGND.n37 VGND.n35 22.9652
R140 VGND.n34 VGND.n1 21.4593
R141 VGND.n23 VGND.n6 15.8123
R142 VGND.n28 VGND.n4 13.8312
R143 VGND.n35 VGND.n0 9.3005
R144 VGND.n34 VGND.n33 9.3005
R145 VGND.n32 VGND.n1 9.3005
R146 VGND.n31 VGND.n30 9.3005
R147 VGND.n29 VGND.n2 9.3005
R148 VGND.n28 VGND.n27 9.3005
R149 VGND.n26 VGND.n25 9.3005
R150 VGND.n24 VGND.n5 9.3005
R151 VGND.n23 VGND.n22 9.3005
R152 VGND.n21 VGND.n6 9.3005
R153 VGND.n20 VGND.n19 9.3005
R154 VGND.n18 VGND.n7 9.3005
R155 VGND.n17 VGND.n16 9.3005
R156 VGND.n15 VGND.n14 9.3005
R157 VGND.n13 VGND.n10 9.3005
R158 VGND.n17 VGND.n9 7.97588
R159 VGND.n38 VGND.n37 7.12063
R160 VGND.n12 VGND.n11 7.07919
R161 VGND.n25 VGND.n4 4.51198
R162 VGND.n14 VGND.n9 1.08358
R163 VGND.n11 VGND.n10 0.201153
R164 VGND.n38 VGND.n0 0.148519
R165 VGND.n15 VGND.n10 0.120292
R166 VGND.n16 VGND.n15 0.120292
R167 VGND.n16 VGND.n7 0.120292
R168 VGND.n20 VGND.n7 0.120292
R169 VGND.n21 VGND.n20 0.120292
R170 VGND.n22 VGND.n21 0.120292
R171 VGND.n22 VGND.n5 0.120292
R172 VGND.n26 VGND.n5 0.120292
R173 VGND.n27 VGND.n26 0.120292
R174 VGND.n27 VGND.n2 0.120292
R175 VGND.n31 VGND.n2 0.120292
R176 VGND.n32 VGND.n31 0.120292
R177 VGND.n33 VGND.n32 0.120292
R178 VGND.n33 VGND.n0 0.120292
R179 VGND VGND.n38 0.0927068
R180 VNB.t3 VNB.t4 2677.02
R181 VNB.t5 VNB.t3 2677.02
R182 VNB.t9 VNB.t8 2677.02
R183 VNB.t2 VNB.t12 2677.02
R184 VNB.t15 VNB.t5 1765.7
R185 VNB.t14 VNB.t11 1623.3
R186 VNB.t0 VNB.t13 1566.34
R187 VNB.t10 VNB.t1 1366.99
R188 VNB.t13 VNB.t14 1366.99
R189 VNB.t12 VNB.t0 1352.75
R190 VNB.t6 VNB.t2 1196.12
R191 VNB.t7 VNB.t15 1025.24
R192 VNB.t1 VNB.t7 1025.24
R193 VNB.t8 VNB.t10 1025.24
R194 VNB.t11 VNB.t9 1025.24
R195 VNB VNB.t6 683.495
R196 a_476_47.n4 a_476_47.n3 707.533
R197 a_476_47.n1 a_476_47.t6 344.899
R198 a_476_47.n2 a_476_47.t4 289.493
R199 a_476_47.n3 a_476_47.n0 288.925
R200 a_476_47.n2 a_476_47.t5 228.148
R201 a_476_47.n3 a_476_47.n2 214.781
R202 a_476_47.n2 a_476_47.n1 105.749
R203 a_476_47.n1 a_476_47.t7 93.1872
R204 a_476_47.n0 a_476_47.t0 70.0005
R205 a_476_47.n0 a_476_47.t3 63.3338
R206 a_476_47.t1 a_476_47.n4 63.3219
R207 a_476_47.n4 a_476_47.t2 63.3219
R208 a_956_413.t0 a_956_413.t1 98.5005
R209 a_193_47.n1 a_193_47.t5 533.949
R210 a_193_47.t1 a_193_47.n3 424.863
R211 a_193_47.n0 a_193_47.t2 368.31
R212 a_193_47.n0 a_193_47.t4 261.351
R213 a_193_47.n3 a_193_47.t0 242.915
R214 a_193_47.n2 a_193_47.n0 187.082
R215 a_193_47.n2 a_193_47.n1 164.226
R216 a_193_47.n1 a_193_47.t3 141.923
R217 a_193_47.n3 a_193_47.n2 10.842
R218 a_1136_413.t0 a_1136_413.t1 98.5005
R219 CLK.n0 CLK.t0 270.457
R220 CLK.n0 CLK.t1 235.109
R221 CLK.n1 CLK.n0 152
R222 CLK.n1 CLK 7.6805
R223 CLK CLK.n1 4.75479
R224 a_27_47.n2 a_27_47.t3 418.678
R225 a_27_47.t0 a_27_47.n5 390.067
R226 a_27_47.n3 a_27_47.t2 311.954
R227 a_27_47.n3 a_27_47.t4 308.168
R228 a_27_47.n2 a_27_47.t6 300.252
R229 a_27_47.n1 a_27_47.t1 287.998
R230 a_27_47.n0 a_27_47.t7 263.173
R231 a_27_47.n0 a_27_47.t5 227.826
R232 a_27_47.n1 a_27_47.n0 152
R233 a_27_47.n5 a_27_47.n1 35.3396
R234 a_27_47.n4 a_27_47.n2 17.2377
R235 a_27_47.n5 a_27_47.n4 10.8063
R236 a_27_47.n4 a_27_47.n3 9.3005
R237 a_1056_47.t0 a_1056_47.t1 60.0005
R238 a_1786_47.t0 a_1786_47.n3 386.31
R239 a_1786_47.n3 a_1786_47.t1 242.385
R240 a_1786_47.n2 a_1786_47.n0 239.04
R241 a_1786_47.n3 a_1786_47.n2 175.274
R242 a_1786_47.n2 a_1786_47.n1 166.739
R243 a_381_47.n1 a_381_47.n0 644.056
R244 a_381_47.n1 a_381_47.t1 95.0032
R245 a_381_47.n0 a_381_47.t3 63.3338
R246 a_381_47.t2 a_381_47.n1 31.6371
R247 a_381_47.n0 a_381_47.t0 26.7713
R248 D.n0 D.t0 264.029
R249 D.n0 D.t1 174.056
R250 D.n1 D.n0 152
R251 D.n1 D 8.58587
R252 D D.n1 2.02977
R253 SET_B.n0 SET_B.t0 389.618
R254 SET_B.n1 SET_B.t3 386.892
R255 SET_B.n2 SET_B.n1 186.411
R256 SET_B.n2 SET_B.n0 156.06
R257 SET_B.n1 SET_B.t1 148.35
R258 SET_B.n0 SET_B.t2 142.569
R259 SET_B SET_B.n2 2.65416
R260 a_1224_47.t0 a_1224_47.t1 60.0005
R261 a_562_413.t0 a_562_413.t1 211.071
R262 a_1296_47.t0 a_1296_47.t1 60.0005
R263 Q_N Q_N.n0 593.34
R264 Q_N.n3 Q_N.n0 585
R265 Q_N.n2 Q_N.n0 585
R266 Q_N.n1 Q_N.t1 128.958
R267 Q_N.n0 Q_N.t0 26.5955
R268 Q_N.n3 Q_N 8.33989
R269 Q_N.n2 Q_N 8.33989
R270 Q_N Q_N.n1 7.03503
R271 Q_N.n1 Q_N 5.87845
R272 Q_N Q_N.n3 4.84898
R273 Q_N Q_N.n2 4.84898
R274 a_796_47.t0 a_796_47.t1 60.0005
C0 SET_B Q 2.15e-19
C1 VPWR Q_N 0.129301f
C2 VGND Q_N 0.101213f
C3 VPWR Q 0.082253f
C4 VPB CLK 0.070197f
C5 VGND Q 0.061147f
C6 VPB D 0.048468f
C7 VPB SET_B 0.143314f
C8 VPB VPWR 0.246766f
C9 VPB VGND 0.022829f
C10 CLK VPWR 0.019428f
C11 VPB Q_N 0.009855f
C12 D VPWR 0.015788f
C13 CLK VGND 0.019435f
C14 SET_B VPWR 0.079222f
C15 VPB Q 0.019769f
C16 D VGND 0.013952f
C17 SET_B VGND 0.336296f
C18 SET_B Q_N 0.001264f
C19 VPWR VGND 0.101436f
C20 Q VNB 0.087852f
C21 Q_N VNB 0.007304f
C22 VGND VNB 1.17804f
C23 VPWR VNB 0.954075f
C24 SET_B VNB 0.244635f
C25 D VNB 0.107124f
C26 CLK VNB 0.195843f
C27 VPB VNB 2.1109f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfsbp_2 VPB VNB VGND VPWR Q Q_N SET_B D CLK
X0 a_1178_261.t1 a_1028_413.t5 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X1 VPWR.t5 a_1028_413.t6 a_1870_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VGND.t2 a_652_21.t3 a_586_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X3 a_1178_261.t0 a_1028_413.t7 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X4 VGND.t5 a_1028_413.t8 a_1870_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_956_413.t0 a_476_47.t4 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_1136_413.t0 a_193_47.t2 a_1028_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR.t11 a_476_47.t5 a_652_21.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR.t1 CLK.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_586_47.t1 a_193_47.t3 a_476_47.t2 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X10 a_1056_47.t0 a_476_47.t6 VGND.t12 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_476_47.t0 a_27_47.t2 a_381_47.t3 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X12 a_381_47.t0 D.t0 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X13 a_652_21.t0 SET_B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X14 a_1224_47.t1 a_27_47.t3 a_1028_413.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_562_413.t1 a_27_47.t4 a_476_47.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 VPWR.t14 a_1870_47.t2 Q.t1 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_1028_413.t2 a_193_47.t4 a_1056_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 VGND.t7 a_1870_47.t3 Q.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_476_47.t3 a_193_47.t5 a_381_47.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X20 a_1296_47.t1 a_1178_261.t2 a_1224_47.t0 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 Q_N.t3 a_1028_413.t9 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_193_47.t0 a_27_47.t5 VGND.t11 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 VPWR.t12 a_652_21.t4 a_562_413.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X24 VGND.t0 SET_B.t1 a_1296_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 Q.t2 a_1870_47.t4 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_1028_413.t4 a_27_47.t6 a_956_413.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X27 VPWR.t8 a_1178_261.t3 a_1136_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 Q.t0 a_1870_47.t5 VPWR.t13 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR.t2 a_1028_413.t10 Q_N.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND.t4 a_1028_413.t11 Q_N.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_193_47.t1 a_27_47.t7 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 Q_N.t0 a_1028_413.t12 VPWR.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_796_47.t0 SET_B.t2 VGND.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X34 a_381_47.t1 D.t1 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X35 a_652_21.t2 a_476_47.t7 a_796_47.t1 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 VPWR.t7 SET_B.t3 a_1028_413.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 VGND.t1 CLK.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1028_413.n6 a_1028_413.t3 724.652
R1 a_1028_413.n6 a_1028_413.n5 611.504
R2 a_1028_413.n8 a_1028_413.n7 287.401
R3 a_1028_413.n4 a_1028_413.t5 258.673
R4 a_1028_413.n0 a_1028_413.t6 221.72
R5 a_1028_413.n1 a_1028_413.t10 221.72
R6 a_1028_413.n2 a_1028_413.t12 221.72
R7 a_1028_413.n7 a_1028_413.n4 217.255
R8 a_1028_413.n3 a_1028_413.t7 210.474
R9 a_1028_413.n1 a_1028_413.n0 167.808
R10 a_1028_413.n3 a_1028_413.n2 154.419
R11 a_1028_413.n0 a_1028_413.t8 149.421
R12 a_1028_413.n1 a_1028_413.t11 149.421
R13 a_1028_413.n2 a_1028_413.t9 149.421
R14 a_1028_413.n5 a_1028_413.t1 119.608
R15 a_1028_413.n7 a_1028_413.n6 93.3652
R16 a_1028_413.n2 a_1028_413.n1 74.9783
R17 a_1028_413.n5 a_1028_413.t4 63.3219
R18 a_1028_413.t0 a_1028_413.n8 47.1434
R19 a_1028_413.n8 a_1028_413.t2 47.1434
R20 a_1028_413.n4 a_1028_413.n3 32.1338
R21 VPWR.n47 VPWR.t6 721.837
R22 VPWR.n8 VPWR.t8 648.322
R23 VPWR.n27 VPWR.n11 604.783
R24 VPWR.n49 VPWR.n1 604.394
R25 VPWR.n6 VPWR.n5 599.74
R26 VPWR.n40 VPWR.n39 585
R27 VPWR.n17 VPWR.t14 346.651
R28 VPWR.n12 VPWR.t4 261.553
R29 VPWR.n21 VPWR.t2 250.464
R30 VPWR.n16 VPWR.n15 230.879
R31 VPWR.n39 VPWR.t0 91.4648
R32 VPWR.n11 VPWR.t7 91.4648
R33 VPWR.n39 VPWR.t12 86.7743
R34 VPWR.n5 VPWR.t10 63.3219
R35 VPWR.n5 VPWR.t11 63.3219
R36 VPWR.n1 VPWR.t9 41.5552
R37 VPWR.n1 VPWR.t1 41.5552
R38 VPWR.n17 VPWR.n16 39.3453
R39 VPWR.n42 VPWR.n3 34.6358
R40 VPWR.n46 VPWR.n3 34.6358
R41 VPWR.n33 VPWR.n32 34.6358
R42 VPWR.n34 VPWR.n33 34.6358
R43 VPWR.n20 VPWR.n14 34.6358
R44 VPWR.n42 VPWR.n41 33.5954
R45 VPWR.n11 VPWR.t3 32.8338
R46 VPWR.n26 VPWR.n12 32.377
R47 VPWR.n38 VPWR.n6 31.624
R48 VPWR.n29 VPWR.n28 27.873
R49 VPWR.n22 VPWR.n21 27.1064
R50 VPWR.n15 VPWR.t13 26.5955
R51 VPWR.n15 VPWR.t5 26.5955
R52 VPWR.n28 VPWR.n27 25.6005
R53 VPWR.n22 VPWR.n12 23.3417
R54 VPWR.n21 VPWR.n20 23.3417
R55 VPWR.n48 VPWR.n47 22.9652
R56 VPWR.n49 VPWR.n48 22.9652
R57 VPWR.n47 VPWR.n46 21.4593
R58 VPWR.n32 VPWR.n8 19.2553
R59 VPWR.n27 VPWR.n26 18.824
R60 VPWR.n34 VPWR.n6 12.8005
R61 VPWR.n40 VPWR.n38 12.5335
R62 VPWR.n18 VPWR.n14 9.3005
R63 VPWR.n20 VPWR.n19 9.3005
R64 VPWR.n21 VPWR.n13 9.3005
R65 VPWR.n23 VPWR.n22 9.3005
R66 VPWR.n24 VPWR.n12 9.3005
R67 VPWR.n26 VPWR.n25 9.3005
R68 VPWR.n27 VPWR.n10 9.3005
R69 VPWR.n28 VPWR.n9 9.3005
R70 VPWR.n30 VPWR.n29 9.3005
R71 VPWR.n32 VPWR.n31 9.3005
R72 VPWR.n33 VPWR.n7 9.3005
R73 VPWR.n35 VPWR.n34 9.3005
R74 VPWR.n36 VPWR.n6 9.3005
R75 VPWR.n38 VPWR.n37 9.3005
R76 VPWR.n41 VPWR.n4 9.3005
R77 VPWR.n43 VPWR.n42 9.3005
R78 VPWR.n44 VPWR.n3 9.3005
R79 VPWR.n46 VPWR.n45 9.3005
R80 VPWR.n47 VPWR.n2 9.3005
R81 VPWR.n48 VPWR.n0 9.3005
R82 VPWR.n50 VPWR.n49 7.12063
R83 VPWR.n41 VPWR.n40 3.37505
R84 VPWR.n18 VPWR.n17 2.24154
R85 VPWR.n29 VPWR.n8 0.815045
R86 VPWR.n16 VPWR.n14 0.376971
R87 VPWR.n50 VPWR.n0 0.148519
R88 VPWR.n19 VPWR.n18 0.120292
R89 VPWR.n19 VPWR.n13 0.120292
R90 VPWR.n23 VPWR.n13 0.120292
R91 VPWR.n24 VPWR.n23 0.120292
R92 VPWR.n25 VPWR.n24 0.120292
R93 VPWR.n25 VPWR.n10 0.120292
R94 VPWR.n10 VPWR.n9 0.120292
R95 VPWR.n30 VPWR.n9 0.120292
R96 VPWR.n31 VPWR.n30 0.120292
R97 VPWR.n31 VPWR.n7 0.120292
R98 VPWR.n35 VPWR.n7 0.120292
R99 VPWR.n36 VPWR.n35 0.120292
R100 VPWR.n37 VPWR.n36 0.120292
R101 VPWR.n37 VPWR.n4 0.120292
R102 VPWR.n43 VPWR.n4 0.120292
R103 VPWR.n44 VPWR.n43 0.120292
R104 VPWR.n45 VPWR.n44 0.120292
R105 VPWR.n45 VPWR.n2 0.120292
R106 VPWR.n2 VPWR.n0 0.120292
R107 VPWR VPWR.n50 0.0927068
R108 a_1178_261.n0 a_1178_261.t2 372.274
R109 a_1178_261.t1 a_1178_261.n1 371.185
R110 a_1178_261.n1 a_1178_261.t0 291.327
R111 a_1178_261.n1 a_1178_261.n0 264.267
R112 a_1178_261.n0 a_1178_261.t3 167.992
R113 VPB.t3 VPB.t4 556.386
R114 VPB.t5 VPB.t2 556.386
R115 VPB.t11 VPB.t10 556.386
R116 VPB.t13 VPB.t9 556.386
R117 VPB.t6 VPB.t16 355.14
R118 VPB.t12 VPB.t7 319.627
R119 VPB.t16 VPB.t0 313.707
R120 VPB.t9 VPB.t8 287.072
R121 VPB.t10 VPB.t5 284.113
R122 VPB.t17 VPB.t18 248.599
R123 VPB.t4 VPB.t17 248.599
R124 VPB.t2 VPB.t3 248.599
R125 VPB.t15 VPB.t14 248.599
R126 VPB.t0 VPB.t15 248.599
R127 VPB.t8 VPB.t6 248.599
R128 VPB.t1 VPB.t13 248.599
R129 VPB.t7 VPB.t11 213.084
R130 VPB.t14 VPB.t12 213.084
R131 VPB VPB.t1 142.056
R132 a_1870_47.t1 a_1870_47.n2 241.767
R133 a_1870_47.n2 a_1870_47.t0 236.308
R134 a_1870_47.n1 a_1870_47.t5 212.081
R135 a_1870_47.n0 a_1870_47.t2 212.081
R136 a_1870_47.n2 a_1870_47.n1 176.436
R137 a_1870_47.n1 a_1870_47.t4 139.78
R138 a_1870_47.n0 a_1870_47.t3 139.78
R139 a_1870_47.n1 a_1870_47.n0 61.346
R140 a_652_21.n2 a_652_21.n1 594.413
R141 a_652_21.n0 a_652_21.t3 387.961
R142 a_652_21.n1 a_652_21.t2 334.156
R143 a_652_21.n1 a_652_21.n0 187.072
R144 a_652_21.n0 a_652_21.t4 143.746
R145 a_652_21.n2 a_652_21.t1 63.3219
R146 a_652_21.t0 a_652_21.n2 63.3219
R147 a_586_47.t0 a_586_47.t1 93.5174
R148 VGND.n13 VGND.t7 291.087
R149 VGND.n43 VGND.t9 280.51
R150 VGND.n32 VGND.t12 237.877
R151 VGND.n46 VGND.n45 199.739
R152 VGND.n9 VGND.n8 185
R153 VGND.n4 VGND.n3 185
R154 VGND.n21 VGND.t3 165.714
R155 VGND.n17 VGND.t4 156.238
R156 VGND.n15 VGND.n14 110.424
R157 VGND.n3 VGND.t2 81.4291
R158 VGND.n8 VGND.t0 67.1434
R159 VGND.n8 VGND.t6 55.3018
R160 VGND.n3 VGND.t10 38.5719
R161 VGND.n45 VGND.t11 38.5719
R162 VGND.n45 VGND.t1 38.5719
R163 VGND.n27 VGND.n26 34.6358
R164 VGND.n28 VGND.n27 34.6358
R165 VGND.n28 VGND.n6 34.6358
R166 VGND.n38 VGND.n37 34.6358
R167 VGND.n39 VGND.n38 34.6358
R168 VGND.n39 VGND.n1 34.6358
R169 VGND.n22 VGND.n21 32.377
R170 VGND.n34 VGND.n33 28.6616
R171 VGND.n33 VGND.n32 27.8593
R172 VGND.n17 VGND.n11 27.1064
R173 VGND.n14 VGND.t8 24.9236
R174 VGND.n14 VGND.t5 24.9236
R175 VGND.n23 VGND.n22 23.5154
R176 VGND.n17 VGND.n16 23.3417
R177 VGND.n21 VGND.n11 23.3417
R178 VGND.n44 VGND.n43 22.9652
R179 VGND.n46 VGND.n44 22.9652
R180 VGND.n16 VGND.n15 22.5887
R181 VGND.n43 VGND.n1 21.4593
R182 VGND.n32 VGND.n6 15.8123
R183 VGND.n37 VGND.n4 13.8312
R184 VGND.n44 VGND.n0 9.3005
R185 VGND.n43 VGND.n42 9.3005
R186 VGND.n41 VGND.n1 9.3005
R187 VGND.n40 VGND.n39 9.3005
R188 VGND.n38 VGND.n2 9.3005
R189 VGND.n37 VGND.n36 9.3005
R190 VGND.n35 VGND.n34 9.3005
R191 VGND.n33 VGND.n5 9.3005
R192 VGND.n32 VGND.n31 9.3005
R193 VGND.n30 VGND.n6 9.3005
R194 VGND.n29 VGND.n28 9.3005
R195 VGND.n27 VGND.n7 9.3005
R196 VGND.n26 VGND.n25 9.3005
R197 VGND.n24 VGND.n23 9.3005
R198 VGND.n22 VGND.n10 9.3005
R199 VGND.n21 VGND.n20 9.3005
R200 VGND.n16 VGND.n12 9.3005
R201 VGND.n18 VGND.n17 9.3005
R202 VGND.n19 VGND.n11 9.3005
R203 VGND.n26 VGND.n9 7.97588
R204 VGND.n47 VGND.n46 7.12063
R205 VGND.n15 VGND.n13 6.51043
R206 VGND.n34 VGND.n4 4.51198
R207 VGND.n23 VGND.n9 1.08358
R208 VGND.n13 VGND.n12 0.662665
R209 VGND.n47 VGND.n0 0.148519
R210 VGND.n18 VGND.n12 0.120292
R211 VGND.n19 VGND.n18 0.120292
R212 VGND.n20 VGND.n19 0.120292
R213 VGND.n20 VGND.n10 0.120292
R214 VGND.n24 VGND.n10 0.120292
R215 VGND.n25 VGND.n24 0.120292
R216 VGND.n25 VGND.n7 0.120292
R217 VGND.n29 VGND.n7 0.120292
R218 VGND.n30 VGND.n29 0.120292
R219 VGND.n31 VGND.n30 0.120292
R220 VGND.n31 VGND.n5 0.120292
R221 VGND.n35 VGND.n5 0.120292
R222 VGND.n36 VGND.n35 0.120292
R223 VGND.n36 VGND.n2 0.120292
R224 VGND.n40 VGND.n2 0.120292
R225 VGND.n41 VGND.n40 0.120292
R226 VGND.n42 VGND.n41 0.120292
R227 VGND.n42 VGND.n0 0.120292
R228 VGND VGND.n47 0.0927068
R229 VNB.t3 VNB.t5 2677.02
R230 VNB.t6 VNB.t4 2677.02
R231 VNB.t18 VNB.t17 2677.02
R232 VNB.t16 VNB.t13 2677.02
R233 VNB.t0 VNB.t6 1765.7
R234 VNB.t2 VNB.t14 1623.3
R235 VNB.t7 VNB.t9 1566.34
R236 VNB.t10 VNB.t8 1366.99
R237 VNB.t9 VNB.t2 1366.99
R238 VNB.t13 VNB.t7 1352.75
R239 VNB.t11 VNB.t12 1196.12
R240 VNB.t5 VNB.t11 1196.12
R241 VNB.t4 VNB.t3 1196.12
R242 VNB.t1 VNB.t16 1196.12
R243 VNB.t15 VNB.t0 1025.24
R244 VNB.t8 VNB.t15 1025.24
R245 VNB.t17 VNB.t10 1025.24
R246 VNB.t14 VNB.t18 1025.24
R247 VNB VNB.t1 683.495
R248 a_476_47.n4 a_476_47.n3 707.533
R249 a_476_47.n1 a_476_47.t6 344.899
R250 a_476_47.n2 a_476_47.t4 289.493
R251 a_476_47.n3 a_476_47.n0 288.925
R252 a_476_47.n2 a_476_47.t5 228.148
R253 a_476_47.n3 a_476_47.n2 214.781
R254 a_476_47.n2 a_476_47.n1 105.749
R255 a_476_47.n1 a_476_47.t7 93.1872
R256 a_476_47.n0 a_476_47.t0 70.0005
R257 a_476_47.n0 a_476_47.t2 63.3338
R258 a_476_47.t1 a_476_47.n4 63.3219
R259 a_476_47.n4 a_476_47.t3 63.3219
R260 a_956_413.t0 a_956_413.t1 98.5005
R261 a_193_47.n1 a_193_47.t5 533.949
R262 a_193_47.t1 a_193_47.n3 424.863
R263 a_193_47.n0 a_193_47.t2 368.31
R264 a_193_47.n0 a_193_47.t4 261.351
R265 a_193_47.n3 a_193_47.t0 242.915
R266 a_193_47.n2 a_193_47.n0 187.082
R267 a_193_47.n2 a_193_47.n1 164.226
R268 a_193_47.n1 a_193_47.t3 141.923
R269 a_193_47.n3 a_193_47.n2 10.842
R270 a_1136_413.t0 a_1136_413.t1 98.5005
R271 CLK.n0 CLK.t0 270.457
R272 CLK.n0 CLK.t1 235.109
R273 CLK.n1 CLK.n0 152
R274 CLK.n1 CLK 7.6805
R275 CLK CLK.n1 4.75479
R276 a_27_47.n2 a_27_47.t3 418.678
R277 a_27_47.t0 a_27_47.n5 390.067
R278 a_27_47.n3 a_27_47.t2 311.954
R279 a_27_47.n3 a_27_47.t4 308.168
R280 a_27_47.n2 a_27_47.t6 300.252
R281 a_27_47.n1 a_27_47.t1 287.998
R282 a_27_47.n0 a_27_47.t7 263.173
R283 a_27_47.n0 a_27_47.t5 227.826
R284 a_27_47.n1 a_27_47.n0 152
R285 a_27_47.n5 a_27_47.n1 35.3396
R286 a_27_47.n4 a_27_47.n2 17.2377
R287 a_27_47.n5 a_27_47.n4 10.8063
R288 a_27_47.n4 a_27_47.n3 9.3005
R289 a_1056_47.t0 a_1056_47.t1 60.0005
R290 a_381_47.n1 a_381_47.n0 644.056
R291 a_381_47.n1 a_381_47.t2 95.0032
R292 a_381_47.n0 a_381_47.t3 63.3338
R293 a_381_47.t0 a_381_47.n1 31.6371
R294 a_381_47.n0 a_381_47.t1 26.7713
R295 D.n0 D.t0 264.029
R296 D.n0 D.t1 174.056
R297 D.n1 D.n0 152
R298 D.n1 D 8.58587
R299 D D.n1 2.02977
R300 SET_B.n0 SET_B.t0 389.618
R301 SET_B.n1 SET_B.t3 386.892
R302 SET_B.n2 SET_B.n1 186.411
R303 SET_B.n2 SET_B.n0 156.06
R304 SET_B.n1 SET_B.t1 148.35
R305 SET_B.n0 SET_B.t2 142.569
R306 SET_B SET_B.n2 2.65416
R307 a_1224_47.t0 a_1224_47.t1 60.0005
R308 a_562_413.t0 a_562_413.t1 211.071
R309 Q Q.n0 593.34
R310 Q.n3 Q.n0 585
R311 Q.n4 Q.n0 585
R312 Q.n2 Q.n1 185
R313 Q Q.n2 48.1618
R314 Q.n3 Q 33.0892
R315 Q.n0 Q.t1 26.5955
R316 Q.n0 Q.t0 26.5955
R317 Q.n1 Q.t3 24.9236
R318 Q.n1 Q.t2 24.9236
R319 Q.n4 Q 8.33989
R320 Q.n2 Q 6.9125
R321 Q Q.n4 4.84898
R322 Q Q.n3 4.65505
R323 a_1296_47.t0 a_1296_47.t1 60.0005
R324 Q_N Q_N.n0 593.34
R325 Q_N.n4 Q_N.n0 585
R326 Q_N.n3 Q_N.n0 585
R327 Q_N.n1 Q_N 185.97
R328 Q_N.n2 Q_N.n1 185
R329 Q_N.n0 Q_N.t1 26.5955
R330 Q_N.n0 Q_N.t0 26.5955
R331 Q_N.n1 Q_N.t2 24.9236
R332 Q_N.n1 Q_N.t3 24.9236
R333 Q_N.n2 Q_N 12.2187
R334 Q_N.n4 Q_N 8.33989
R335 Q_N.n3 Q_N 8.33989
R336 Q_N Q_N.n4 4.84898
R337 Q_N Q_N.n3 4.84898
R338 Q_N Q_N.n2 0.970197
R339 a_796_47.t0 a_796_47.t1 60.0005
C0 SET_B Q_N 0.001264f
C1 VPWR VGND 0.120553f
C2 SET_B Q 4.05e-19
C3 VPWR Q_N 0.211897f
C4 VGND Q_N 0.155721f
C5 VPWR Q 0.215894f
C6 VPB CLK 0.070197f
C7 VGND Q 0.150182f
C8 VPB D 0.048468f
C9 VPB SET_B 0.144174f
C10 VPB VPWR 0.257687f
C11 VPB VGND 0.019396f
C12 CLK VPWR 0.019428f
C13 CLK VGND 0.019435f
C14 D VPWR 0.015788f
C15 VPB Q_N 0.005444f
C16 VPB Q 0.009433f
C17 D VGND 0.013952f
C18 SET_B VPWR 0.079485f
C19 SET_B VGND 0.336607f
C20 Q VNB 0.055453f
C21 Q_N VNB 0.004442f
C22 VGND VNB 1.22369f
C23 VPWR VNB 1.00278f
C24 SET_B VNB 0.245456f
C25 D VNB 0.107124f
C26 CLK VNB 0.195843f
C27 VPB VNB 2.19949f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_1 VPB VNB VPWR VGND Q SET_B D CLK
X0 VGND.t3 a_652_21.t3 a_586_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413.t1 a_476_47.t4 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR.t8 a_476_47.t5 a_652_21.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR.t3 CLK.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_586_47.t0 a_193_47.t2 a_476_47.t2 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1056_47.t1 a_476_47.t6 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 a_476_47.t0 a_27_47.t2 a_381_47.t3 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X7 a_381_47.t0 D.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X8 a_652_21.t2 SET_B.t0 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47.t1 a_27_47.t3 a_1032_413.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413.t1 a_27_47.t4 a_476_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND.t4 a_1032_413.t5 a_1602_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 VPWR.t1 a_1182_261.t2 a_1140_413.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 a_1032_413.t1 a_193_47.t3 a_1056_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 a_476_47.t3 a_193_47.t4 a_381_47.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X15 a_1296_47.t1 a_1182_261.t3 a_1224_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_193_47.t0 a_27_47.t5 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR.t5 a_652_21.t4 a_562_413.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X18 VPWR.t2 SET_B.t1 a_1032_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 a_1032_413.t3 a_27_47.t6 a_956_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X20 a_1182_261.t1 a_1032_413.t6 VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X21 a_193_47.t1 a_27_47.t7 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1140_413.t1 a_193_47.t5 a_1032_413.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR.t10 a_1032_413.t7 a_1602_47.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X24 a_796_47.t0 SET_B.t2 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X25 a_381_47.t2 D.t1 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 a_1182_261.t0 a_1032_413.t8 VGND.t8 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X27 a_652_21.t1 a_476_47.t7 a_796_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 VGND.t1 CLK.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VGND.t6 SET_B.t3 a_1296_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
R0 a_652_21.n2 a_652_21.n1 594.413
R1 a_652_21.n0 a_652_21.t3 387.961
R2 a_652_21.n1 a_652_21.t1 328.048
R3 a_652_21.n1 a_652_21.n0 187.072
R4 a_652_21.n0 a_652_21.t4 143.746
R5 a_652_21.t0 a_652_21.n2 63.3219
R6 a_652_21.n2 a_652_21.t2 63.3219
R7 a_586_47.t1 a_586_47.t0 93.5174
R8 VGND.n29 VGND.t5 280.51
R9 VGND.n10 VGND.t4 262.281
R10 VGND.n18 VGND.t7 238.772
R11 VGND.n32 VGND.n31 199.739
R12 VGND.n9 VGND.n8 185
R13 VGND.n4 VGND.n3 185
R14 VGND.n3 VGND.t3 81.4291
R15 VGND.n8 VGND.t6 67.1434
R16 VGND.n8 VGND.t8 55.3018
R17 VGND.n3 VGND.t2 38.5719
R18 VGND.n31 VGND.t0 38.5719
R19 VGND.n31 VGND.t1 38.5719
R20 VGND.n13 VGND.n12 34.6358
R21 VGND.n14 VGND.n13 34.6358
R22 VGND.n14 VGND.n6 34.6358
R23 VGND.n24 VGND.n23 34.6358
R24 VGND.n25 VGND.n24 34.6358
R25 VGND.n25 VGND.n1 34.6358
R26 VGND.n19 VGND.n18 29.3652
R27 VGND.n20 VGND.n19 28.6616
R28 VGND.n30 VGND.n29 22.9652
R29 VGND.n32 VGND.n30 22.9652
R30 VGND.n29 VGND.n1 21.4593
R31 VGND.n18 VGND.n6 15.8123
R32 VGND.n23 VGND.n4 13.8312
R33 VGND.n12 VGND.n9 9.48177
R34 VGND.n12 VGND.n11 9.3005
R35 VGND.n13 VGND.n7 9.3005
R36 VGND.n15 VGND.n14 9.3005
R37 VGND.n16 VGND.n6 9.3005
R38 VGND.n18 VGND.n17 9.3005
R39 VGND.n19 VGND.n5 9.3005
R40 VGND.n21 VGND.n20 9.3005
R41 VGND.n23 VGND.n22 9.3005
R42 VGND.n24 VGND.n2 9.3005
R43 VGND.n26 VGND.n25 9.3005
R44 VGND.n27 VGND.n1 9.3005
R45 VGND.n29 VGND.n28 9.3005
R46 VGND.n30 VGND.n0 9.3005
R47 VGND.n10 VGND.n9 7.70898
R48 VGND.n33 VGND.n32 7.12063
R49 VGND.n20 VGND.n4 4.51198
R50 VGND.n11 VGND.n10 0.20946
R51 VGND.n33 VGND.n0 0.148519
R52 VGND.n11 VGND.n7 0.120292
R53 VGND.n15 VGND.n7 0.120292
R54 VGND.n16 VGND.n15 0.120292
R55 VGND.n17 VGND.n16 0.120292
R56 VGND.n17 VGND.n5 0.120292
R57 VGND.n21 VGND.n5 0.120292
R58 VGND.n22 VGND.n21 0.120292
R59 VGND.n22 VGND.n2 0.120292
R60 VGND.n26 VGND.n2 0.120292
R61 VGND.n27 VGND.n26 0.120292
R62 VGND.n28 VGND.n27 0.120292
R63 VGND.n28 VGND.n0 0.120292
R64 VGND VGND.n33 0.114842
R65 VNB.t14 VNB.t8 2677.02
R66 VNB.t13 VNB.t12 2677.02
R67 VNB.t2 VNB.t10 2677.02
R68 VNB.t11 VNB.t14 1765.7
R69 VNB.t7 VNB.t5 1623.3
R70 VNB.t0 VNB.t6 1566.34
R71 VNB.t9 VNB.t1 1366.99
R72 VNB.t6 VNB.t7 1366.99
R73 VNB.t10 VNB.t0 1352.75
R74 VNB.t4 VNB.t2 1196.12
R75 VNB.t3 VNB.t11 1082.2
R76 VNB.t1 VNB.t3 1025.24
R77 VNB.t12 VNB.t9 1025.24
R78 VNB.t5 VNB.t13 1025.24
R79 VNB VNB.t4 683.495
R80 a_476_47.n4 a_476_47.n3 707.533
R81 a_476_47.n1 a_476_47.t6 344.899
R82 a_476_47.n2 a_476_47.t4 289.493
R83 a_476_47.n3 a_476_47.n0 288.925
R84 a_476_47.n2 a_476_47.t5 228.148
R85 a_476_47.n3 a_476_47.n2 214.781
R86 a_476_47.n2 a_476_47.n1 105.749
R87 a_476_47.n1 a_476_47.t7 93.1872
R88 a_476_47.n0 a_476_47.t0 70.0005
R89 a_476_47.n0 a_476_47.t2 63.3338
R90 a_476_47.t1 a_476_47.n4 63.3219
R91 a_476_47.n4 a_476_47.t3 63.3219
R92 VPWR.n32 VPWR.t4 721.837
R93 VPWR.n8 VPWR.t1 648.322
R94 VPWR.n12 VPWR.n11 604.783
R95 VPWR.n34 VPWR.n1 604.394
R96 VPWR.n6 VPWR.n5 599.74
R97 VPWR.n25 VPWR.n24 585
R98 VPWR.n10 VPWR.t10 377.736
R99 VPWR.n24 VPWR.t6 91.4648
R100 VPWR.n11 VPWR.t2 91.4648
R101 VPWR.n24 VPWR.t5 86.7743
R102 VPWR.n5 VPWR.t7 63.3219
R103 VPWR.n5 VPWR.t8 63.3219
R104 VPWR.n1 VPWR.t0 41.5552
R105 VPWR.n1 VPWR.t3 41.5552
R106 VPWR.n27 VPWR.n3 34.6358
R107 VPWR.n31 VPWR.n3 34.6358
R108 VPWR.n18 VPWR.n17 34.6358
R109 VPWR.n19 VPWR.n18 34.6358
R110 VPWR.n27 VPWR.n26 33.5954
R111 VPWR.n11 VPWR.t9 32.8338
R112 VPWR.n23 VPWR.n6 31.624
R113 VPWR.n13 VPWR.n12 27.1064
R114 VPWR.n14 VPWR.n13 26.8326
R115 VPWR.n33 VPWR.n32 22.9652
R116 VPWR.n34 VPWR.n33 22.9652
R117 VPWR.n32 VPWR.n31 21.4593
R118 VPWR.n17 VPWR.n8 20.2409
R119 VPWR.n19 VPWR.n6 12.8005
R120 VPWR.n25 VPWR.n23 12.5335
R121 VPWR.n13 VPWR.n9 9.3005
R122 VPWR.n15 VPWR.n14 9.3005
R123 VPWR.n17 VPWR.n16 9.3005
R124 VPWR.n18 VPWR.n7 9.3005
R125 VPWR.n20 VPWR.n19 9.3005
R126 VPWR.n21 VPWR.n6 9.3005
R127 VPWR.n23 VPWR.n22 9.3005
R128 VPWR.n26 VPWR.n4 9.3005
R129 VPWR.n28 VPWR.n27 9.3005
R130 VPWR.n29 VPWR.n3 9.3005
R131 VPWR.n31 VPWR.n30 9.3005
R132 VPWR.n32 VPWR.n2 9.3005
R133 VPWR.n33 VPWR.n0 9.3005
R134 VPWR.n35 VPWR.n34 7.12063
R135 VPWR.n12 VPWR.n10 6.68214
R136 VPWR.n26 VPWR.n25 3.37505
R137 VPWR.n14 VPWR.n8 0.349591
R138 VPWR.n10 VPWR.n9 0.222582
R139 VPWR.n35 VPWR.n0 0.148519
R140 VPWR.n15 VPWR.n9 0.120292
R141 VPWR.n16 VPWR.n15 0.120292
R142 VPWR.n16 VPWR.n7 0.120292
R143 VPWR.n20 VPWR.n7 0.120292
R144 VPWR.n21 VPWR.n20 0.120292
R145 VPWR.n22 VPWR.n21 0.120292
R146 VPWR.n22 VPWR.n4 0.120292
R147 VPWR.n28 VPWR.n4 0.120292
R148 VPWR.n29 VPWR.n28 0.120292
R149 VPWR.n30 VPWR.n29 0.120292
R150 VPWR.n30 VPWR.n2 0.120292
R151 VPWR.n2 VPWR.n0 0.120292
R152 VPWR VPWR.n35 0.114842
R153 a_956_413.t0 a_956_413.t1 107.882
R154 VPB.t13 VPB.t14 556.386
R155 VPB.t3 VPB.t4 556.386
R156 VPB.t2 VPB.t6 556.386
R157 VPB.t0 VPB.t7 355.14
R158 VPB.t1 VPB.t9 319.627
R159 VPB.t7 VPB.t10 313.707
R160 VPB.t6 VPB.t8 287.072
R161 VPB.t4 VPB.t13 284.113
R162 VPB.t11 VPB.t12 248.599
R163 VPB.t10 VPB.t11 248.599
R164 VPB.t8 VPB.t0 248.599
R165 VPB.t5 VPB.t2 248.599
R166 VPB.t12 VPB.t1 224.923
R167 VPB.t9 VPB.t3 213.084
R168 VPB VPB.t5 142.056
R169 CLK.n0 CLK.t0 270.457
R170 CLK.n0 CLK.t1 235.109
R171 CLK.n1 CLK.n0 152
R172 CLK.n1 CLK 7.6805
R173 CLK CLK.n1 4.75479
R174 a_27_47.n2 a_27_47.t3 419.505
R175 a_27_47.t1 a_27_47.n5 390.067
R176 a_27_47.n3 a_27_47.t2 312.796
R177 a_27_47.n3 a_27_47.t4 307.325
R178 a_27_47.n2 a_27_47.t6 300.252
R179 a_27_47.n1 a_27_47.t0 287.998
R180 a_27_47.n0 a_27_47.t7 263.173
R181 a_27_47.n0 a_27_47.t5 227.826
R182 a_27_47.n1 a_27_47.n0 152
R183 a_27_47.n5 a_27_47.n1 35.3396
R184 a_27_47.n4 a_27_47.n2 18.2878
R185 a_27_47.n5 a_27_47.n4 10.8599
R186 a_27_47.n4 a_27_47.n3 9.3005
R187 a_193_47.n1 a_193_47.t4 533.949
R188 a_193_47.t1 a_193_47.n3 424.863
R189 a_193_47.n0 a_193_47.t5 379.021
R190 a_193_47.n0 a_193_47.t3 261.351
R191 a_193_47.n3 a_193_47.t0 242.915
R192 a_193_47.n2 a_193_47.n0 187.064
R193 a_193_47.n2 a_193_47.n1 164.76
R194 a_193_47.n1 a_193_47.t2 141.923
R195 a_193_47.n3 a_193_47.n2 10.8599
R196 a_1056_47.t0 a_1056_47.t1 60.0005
R197 a_381_47.n1 a_381_47.n0 644.056
R198 a_381_47.n1 a_381_47.t1 95.0032
R199 a_381_47.n0 a_381_47.t3 63.3338
R200 a_381_47.t0 a_381_47.n1 31.6371
R201 a_381_47.n0 a_381_47.t2 26.7713
R202 D.n0 D.t0 264.029
R203 D.n0 D.t1 174.056
R204 D.n1 D.n0 152
R205 D.n1 D 8.58587
R206 D D.n1 2.02977
R207 SET_B.n0 SET_B.t0 389.618
R208 SET_B.n1 SET_B.t1 386.892
R209 SET_B.n2 SET_B.n1 188.581
R210 SET_B.n2 SET_B.n0 156.06
R211 SET_B.n1 SET_B.t3 148.35
R212 SET_B.n0 SET_B.t2 142.569
R213 SET_B SET_B.n2 2.65416
R214 a_1032_413.t0 a_1032_413.n5 726.158
R215 a_1032_413.n5 a_1032_413.n0 610.48
R216 a_1032_413.n4 a_1032_413.n1 287.401
R217 a_1032_413.n2 a_1032_413.t7 237.787
R218 a_1032_413.n4 a_1032_413.n3 229.714
R219 a_1032_413.n2 a_1032_413.t5 208.868
R220 a_1032_413.n3 a_1032_413.t6 205.654
R221 a_1032_413.n3 a_1032_413.t8 189.588
R222 a_1032_413.n3 a_1032_413.n2 137.298
R223 a_1032_413.n0 a_1032_413.t2 119.608
R224 a_1032_413.n5 a_1032_413.n4 93.3652
R225 a_1032_413.n0 a_1032_413.t3 63.3219
R226 a_1032_413.n1 a_1032_413.t4 47.1434
R227 a_1032_413.n1 a_1032_413.t1 47.1434
R228 a_1224_47.t0 a_1224_47.t1 60.0005
R229 a_562_413.t0 a_562_413.t1 211.071
R230 a_1602_47.t1 a_1602_47.n3 393.632
R231 a_1602_47.n3 a_1602_47.t0 248.404
R232 a_1602_47.n2 a_1602_47.n0 241.536
R233 a_1602_47.n3 a_1602_47.n2 174.886
R234 a_1602_47.n2 a_1602_47.n1 169.237
R235 a_1182_261.n0 a_1182_261.t3 374.755
R236 a_1182_261.t1 a_1182_261.n1 371.185
R237 a_1182_261.n1 a_1182_261.t0 291.327
R238 a_1182_261.n1 a_1182_261.n0 265.774
R239 a_1182_261.n0 a_1182_261.t2 169.453
R240 a_1140_413.t0 a_1140_413.t1 98.5005
R241 a_1296_47.t0 a_1296_47.t1 65.7148
R242 a_796_47.t0 a_796_47.t1 60.0005
C0 VPWR Q 0.070378f
C1 VGND Q 0.059486f
C2 VPB CLK 0.070197f
C3 VPB D 0.048468f
C4 VPB SET_B 0.142745f
C5 VPB VPWR 0.218217f
C6 VPB VGND 0.017329f
C7 CLK VPWR 0.019428f
C8 VPB Q 0.017394f
C9 D VPWR 0.015788f
C10 CLK VGND 0.019435f
C11 SET_B VPWR 0.080687f
C12 D VGND 0.013952f
C13 SET_B VGND 0.337887f
C14 VPWR VGND 0.068713f
C15 SET_B Q 4.58e-19
C16 Q VNB 0.083407f
C17 VGND VNB 1.07774f
C18 VPWR VNB 0.874725f
C19 SET_B VNB 0.246768f
C20 D VNB 0.107124f
C21 CLK VNB 0.195843f
C22 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_2 VPB VNB VPWR VGND Q SET_B D CLK
X0 VGND.t7 a_652_21.t3 a_586_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413.t0 a_476_47.t4 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413.t1 a_193_47.t2 a_1028_413.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR.t4 a_476_47.t5 a_652_21.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1228_47.t1 a_27_47.t2 a_1028_413.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X5 VPWR.t6 CLK.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_586_47.t1 a_193_47.t3 a_476_47.t1 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X7 a_1056_47.t1 a_476_47.t6 VGND.t9 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_476_47.t2 a_27_47.t3 a_381_47.t0 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X9 a_381_47.t1 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X10 a_652_21.t0 SET_B.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR.t7 a_1602_47.t2 Q.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413.t0 a_27_47.t4 a_476_47.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND.t5 a_1028_413.t5 a_1602_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND.t4 a_1602_47.t3 Q.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Q.t2 a_1602_47.t4 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413.t0 a_193_47.t4 a_1056_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47.t0 a_193_47.t5 a_381_47.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X18 a_193_47.t0 a_27_47.t5 VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR.t9 a_1028_413.t6 a_1602_47.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR.t10 a_652_21.t4 a_562_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q.t0 a_1602_47.t5 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_1028_413.t4 a_27_47.t6 a_956_413.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR.t0 a_1178_261# a_1136_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47.t1 a_27_47.t7 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_796_47.t0 SET_B.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X26 a_1300_47.t0 a_1178_261# a_1228_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X27 a_381_47.t3 D.t1 VGND.t10 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 a_1178_261# a_1028_413.t7 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X29 a_652_21.t2 a_476_47.t7 a_796_47.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VPWR.t3 SET_B.t2 a_1028_413.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND.t3 CLK.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 VGND.t2 SET_B.t3 a_1300_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
R0 a_652_21.n2 a_652_21.n1 594.413
R1 a_652_21.n0 a_652_21.t3 387.961
R2 a_652_21.n1 a_652_21.t2 334.156
R3 a_652_21.n1 a_652_21.n0 187.072
R4 a_652_21.n0 a_652_21.t4 143.746
R5 a_652_21.n2 a_652_21.t1 63.3219
R6 a_652_21.t0 a_652_21.n2 63.3219
R7 a_586_47.t0 a_586_47.t1 93.5174
R8 VGND.n13 VGND.t4 292.935
R9 VGND.n37 VGND.t10 280.51
R10 VGND.n26 VGND.t9 238.772
R11 VGND.n40 VGND.n39 199.739
R12 VGND.n9 VGND.n8 185
R13 VGND.n4 VGND.n3 185
R14 VGND.n12 VGND.n11 110.424
R15 VGND.n3 VGND.t7 81.4291
R16 VGND.n8 VGND.t2 67.1434
R17 VGND.n8 VGND.t6 55.3018
R18 VGND.n3 VGND.t1 38.5719
R19 VGND.n39 VGND.t8 38.5719
R20 VGND.n39 VGND.t3 38.5719
R21 VGND.n16 VGND.n15 34.6358
R22 VGND.n21 VGND.n20 34.6358
R23 VGND.n22 VGND.n21 34.6358
R24 VGND.n22 VGND.n6 34.6358
R25 VGND.n32 VGND.n31 34.6358
R26 VGND.n33 VGND.n32 34.6358
R27 VGND.n33 VGND.n1 34.6358
R28 VGND.n27 VGND.n26 29.3652
R29 VGND.n28 VGND.n27 28.6616
R30 VGND.n15 VGND.n12 25.6005
R31 VGND.n11 VGND.t0 24.9236
R32 VGND.n11 VGND.t5 24.9236
R33 VGND.n17 VGND.n16 23.5154
R34 VGND.n38 VGND.n37 22.9652
R35 VGND.n40 VGND.n38 22.9652
R36 VGND.n37 VGND.n1 21.4593
R37 VGND.n26 VGND.n6 15.8123
R38 VGND.n31 VGND.n4 13.8312
R39 VGND.n20 VGND.n9 9.48177
R40 VGND.n38 VGND.n0 9.3005
R41 VGND.n37 VGND.n36 9.3005
R42 VGND.n35 VGND.n1 9.3005
R43 VGND.n34 VGND.n33 9.3005
R44 VGND.n32 VGND.n2 9.3005
R45 VGND.n31 VGND.n30 9.3005
R46 VGND.n29 VGND.n28 9.3005
R47 VGND.n27 VGND.n5 9.3005
R48 VGND.n26 VGND.n25 9.3005
R49 VGND.n24 VGND.n6 9.3005
R50 VGND.n23 VGND.n22 9.3005
R51 VGND.n21 VGND.n7 9.3005
R52 VGND.n20 VGND.n19 9.3005
R53 VGND.n18 VGND.n17 9.3005
R54 VGND.n16 VGND.n10 9.3005
R55 VGND.n15 VGND.n14 9.3005
R56 VGND.n41 VGND.n40 7.12063
R57 VGND.n13 VGND.n12 6.31729
R58 VGND.n28 VGND.n4 4.51198
R59 VGND.n17 VGND.n9 0.689731
R60 VGND.n14 VGND.n13 0.673379
R61 VGND.n41 VGND.n0 0.148519
R62 VGND.n14 VGND.n10 0.120292
R63 VGND.n18 VGND.n10 0.120292
R64 VGND.n19 VGND.n18 0.120292
R65 VGND.n19 VGND.n7 0.120292
R66 VGND.n23 VGND.n7 0.120292
R67 VGND.n24 VGND.n23 0.120292
R68 VGND.n25 VGND.n24 0.120292
R69 VGND.n25 VGND.n5 0.120292
R70 VGND.n29 VGND.n5 0.120292
R71 VGND.n30 VGND.n29 0.120292
R72 VGND.n30 VGND.n2 0.120292
R73 VGND.n34 VGND.n2 0.120292
R74 VGND.n35 VGND.n34 0.120292
R75 VGND.n36 VGND.n35 0.120292
R76 VGND.n36 VGND.n0 0.120292
R77 VGND VGND.n41 0.114842
R78 VNB.t8 VNB.t7 2677.02
R79 VNB.t15 VNB.t14 2677.02
R80 VNB.t13 VNB.t16 2677.02
R81 VNB.t3 VNB.t8 1765.7
R82 VNB.t9 VNB.t2 1623.3
R83 VNB.t12 VNB.t10 1566.34
R84 VNB.t5 VNB.t11 1423.95
R85 VNB.t10 VNB.t9 1366.99
R86 VNB.t16 VNB.t12 1352.75
R87 VNB.t1 VNB.t6 1196.12
R88 VNB.t7 VNB.t1 1196.12
R89 VNB.t4 VNB.t13 1196.12
R90 VNB.t0 VNB.t3 1025.24
R91 VNB.t11 VNB.t0 1025.24
R92 VNB.t14 VNB.t5 1025.24
R93 VNB.t2 VNB.t15 1025.24
R94 VNB VNB.t4 683.495
R95 a_476_47.n4 a_476_47.n3 707.533
R96 a_476_47.n1 a_476_47.t6 344.899
R97 a_476_47.n2 a_476_47.t4 289.493
R98 a_476_47.n3 a_476_47.n0 288.925
R99 a_476_47.n2 a_476_47.t5 228.148
R100 a_476_47.n3 a_476_47.n2 214.781
R101 a_476_47.n2 a_476_47.n1 105.749
R102 a_476_47.n1 a_476_47.t7 93.1872
R103 a_476_47.n0 a_476_47.t2 70.0005
R104 a_476_47.n0 a_476_47.t1 63.3338
R105 a_476_47.n4 a_476_47.t3 63.3219
R106 a_476_47.t0 a_476_47.n4 63.3219
R107 VPWR.n40 VPWR.t1 721.837
R108 VPWR.n20 VPWR.t3 693.902
R109 VPWR.n8 VPWR.t0 648.322
R110 VPWR.n42 VPWR.n1 604.394
R111 VPWR.n6 VPWR.n5 599.74
R112 VPWR.n33 VPWR.n32 585
R113 VPWR.n12 VPWR.t7 347.469
R114 VPWR.n14 VPWR.n13 230.879
R115 VPWR.n32 VPWR.t2 91.4648
R116 VPWR.n32 VPWR.t10 86.7743
R117 VPWR.n5 VPWR.t5 63.3219
R118 VPWR.n5 VPWR.t4 63.3219
R119 VPWR.n1 VPWR.t11 41.5552
R120 VPWR.n1 VPWR.t6 41.5552
R121 VPWR.n14 VPWR.n12 36.6199
R122 VPWR.n35 VPWR.n3 34.6358
R123 VPWR.n39 VPWR.n3 34.6358
R124 VPWR.n26 VPWR.n25 34.6358
R125 VPWR.n27 VPWR.n26 34.6358
R126 VPWR.n15 VPWR.n11 34.6358
R127 VPWR.n19 VPWR.n11 34.6358
R128 VPWR.n35 VPWR.n34 33.5954
R129 VPWR.n31 VPWR.n6 31.624
R130 VPWR.n22 VPWR.n21 27.873
R131 VPWR.n13 VPWR.t8 26.5955
R132 VPWR.n13 VPWR.t9 26.5955
R133 VPWR.n21 VPWR.n20 25.6005
R134 VPWR.n41 VPWR.n40 22.9652
R135 VPWR.n42 VPWR.n41 22.9652
R136 VPWR.n40 VPWR.n39 21.4593
R137 VPWR.n20 VPWR.n19 18.824
R138 VPWR.n25 VPWR.n8 18.735
R139 VPWR.n27 VPWR.n6 12.8005
R140 VPWR.n33 VPWR.n31 12.5335
R141 VPWR.n16 VPWR.n15 9.3005
R142 VPWR.n17 VPWR.n11 9.3005
R143 VPWR.n19 VPWR.n18 9.3005
R144 VPWR.n20 VPWR.n10 9.3005
R145 VPWR.n21 VPWR.n9 9.3005
R146 VPWR.n23 VPWR.n22 9.3005
R147 VPWR.n25 VPWR.n24 9.3005
R148 VPWR.n26 VPWR.n7 9.3005
R149 VPWR.n28 VPWR.n27 9.3005
R150 VPWR.n29 VPWR.n6 9.3005
R151 VPWR.n31 VPWR.n30 9.3005
R152 VPWR.n34 VPWR.n4 9.3005
R153 VPWR.n36 VPWR.n35 9.3005
R154 VPWR.n37 VPWR.n3 9.3005
R155 VPWR.n39 VPWR.n38 9.3005
R156 VPWR.n40 VPWR.n2 9.3005
R157 VPWR.n41 VPWR.n0 9.3005
R158 VPWR.n43 VPWR.n42 7.12063
R159 VPWR.n15 VPWR.n14 3.38874
R160 VPWR.n34 VPWR.n33 3.37505
R161 VPWR.n16 VPWR.n12 2.09743
R162 VPWR.n22 VPWR.n8 0.815045
R163 VPWR.n43 VPWR.n0 0.148519
R164 VPWR.n17 VPWR.n16 0.120292
R165 VPWR.n18 VPWR.n17 0.120292
R166 VPWR.n18 VPWR.n10 0.120292
R167 VPWR.n10 VPWR.n9 0.120292
R168 VPWR.n23 VPWR.n9 0.120292
R169 VPWR.n24 VPWR.n23 0.120292
R170 VPWR.n24 VPWR.n7 0.120292
R171 VPWR.n28 VPWR.n7 0.120292
R172 VPWR.n29 VPWR.n28 0.120292
R173 VPWR.n30 VPWR.n29 0.120292
R174 VPWR.n30 VPWR.n4 0.120292
R175 VPWR.n36 VPWR.n4 0.120292
R176 VPWR.n37 VPWR.n36 0.120292
R177 VPWR.n38 VPWR.n37 0.120292
R178 VPWR.n38 VPWR.n2 0.120292
R179 VPWR.n2 VPWR.n0 0.120292
R180 VPWR VPWR.n43 0.114842
R181 a_956_413.t0 a_956_413.t1 98.5005
R182 VPB.t3 VPB.t10 852.337
R183 VPB.t0 VPB.t3 556.386
R184 VPB.t15 VPB.t1 556.386
R185 VPB.t13 VPB.t11 355.14
R186 VPB.t14 VPB.t12 319.627
R187 VPB.t11 VPB.t2 313.707
R188 VPB.t1 VPB.t8 287.072
R189 VPB.t9 VPB.t7 248.599
R190 VPB.t10 VPB.t9 248.599
R191 VPB.t4 VPB.t5 248.599
R192 VPB.t2 VPB.t4 248.599
R193 VPB.t8 VPB.t13 248.599
R194 VPB.t6 VPB.t15 248.599
R195 VPB.t12 VPB.t0 213.084
R196 VPB.t5 VPB.t14 213.084
R197 VPB VPB.t6 142.056
R198 a_193_47.n1 a_193_47.t5 533.949
R199 a_193_47.t1 a_193_47.n3 423.546
R200 a_193_47.n0 a_193_47.t2 373.666
R201 a_193_47.n0 a_193_47.t4 264.029
R202 a_193_47.n3 a_193_47.t0 242.632
R203 a_193_47.n2 a_193_47.n0 189.742
R204 a_193_47.n2 a_193_47.n1 164.226
R205 a_193_47.n1 a_193_47.t3 141.923
R206 a_193_47.n3 a_193_47.n2 10.842
R207 a_1028_413.n5 a_1028_413.t2 726.158
R208 a_1028_413.n5 a_1028_413.n4 610.48
R209 a_1028_413.n3 a_1028_413.n2 399.219
R210 a_1028_413.n7 a_1028_413.n6 287.401
R211 a_1028_413.n6 a_1028_413.n3 217.637
R212 a_1028_413.n1 a_1028_413.t7 189.588
R213 a_1028_413.n0 a_1028_413.t6 184.768
R214 a_1028_413.n0 a_1028_413.t5 171.913
R215 a_1028_413.n1 a_1028_413.n0 143.835
R216 a_1028_413.n4 a_1028_413.t1 119.608
R217 a_1028_413.n6 a_1028_413.n5 94.8711
R218 a_1028_413.n4 a_1028_413.t4 63.3219
R219 a_1028_413.n7 a_1028_413.t3 52.8576
R220 a_1028_413.t0 a_1028_413.n7 47.1434
R221 a_1028_413.n3 a_1028_413.n1 12.2418
R222 a_1136_413.t0 a_1136_413.t1 98.5005
R223 a_27_47.n2 a_27_47.t2 418.356
R224 a_27_47.t0 a_27_47.n5 385.147
R225 a_27_47.n3 a_27_47.t3 311.954
R226 a_27_47.n3 a_27_47.t4 308.168
R227 a_27_47.n2 a_27_47.t6 300.252
R228 a_27_47.n1 a_27_47.t1 282.147
R229 a_27_47.n0 a_27_47.t7 262.945
R230 a_27_47.n0 a_27_47.t5 227.597
R231 a_27_47.n1 a_27_47.n0 152
R232 a_27_47.n5 a_27_47.n1 35.3396
R233 a_27_47.n4 a_27_47.n2 17.2377
R234 a_27_47.n5 a_27_47.n4 10.842
R235 a_27_47.n4 a_27_47.n3 9.3005
R236 a_1228_47.t0 a_1228_47.t1 60.0005
R237 CLK.n0 CLK.t0 272.062
R238 CLK.n0 CLK.t1 236.716
R239 CLK.n1 CLK.n0 152
R240 CLK.n1 CLK 7.6805
R241 CLK CLK.n1 4.75479
R242 a_1056_47.t0 a_1056_47.t1 60.0005
R243 a_381_47.n1 a_381_47.n0 644.056
R244 a_381_47.n1 a_381_47.t2 95.0032
R245 a_381_47.n0 a_381_47.t0 63.3338
R246 a_381_47.t1 a_381_47.n1 31.6371
R247 a_381_47.n0 a_381_47.t3 26.7713
R248 D.n0 D.t0 264.029
R249 D.n0 D.t1 174.056
R250 D.n1 D.n0 152
R251 D.n1 D 8.58587
R252 D D.n1 2.02977
R253 SET_B.n0 SET_B.t0 389.618
R254 SET_B.n1 SET_B.t2 372.149
R255 SET_B.n2 SET_B.n1 185.464
R256 SET_B.n2 SET_B.n0 156.06
R257 SET_B.n1 SET_B.t3 148.35
R258 SET_B.n0 SET_B.t1 142.569
R259 SET_B SET_B.n2 2.65416
R260 a_1602_47.n2 a_1602_47.t0 247.993
R261 a_1602_47.t1 a_1602_47.n2 247.275
R262 a_1602_47.n1 a_1602_47.t4 212.081
R263 a_1602_47.n0 a_1602_47.t2 212.081
R264 a_1602_47.n2 a_1602_47.n1 174.886
R265 a_1602_47.n1 a_1602_47.t5 139.78
R266 a_1602_47.n0 a_1602_47.t3 139.78
R267 a_1602_47.n1 a_1602_47.n0 61.346
R268 Q.n5 Q 593.34
R269 Q.n5 Q.n4 585
R270 Q.n6 Q.n5 585
R271 Q.n2 Q.n0 186.352
R272 Q.n3 Q.n2 39.8639
R273 Q.n7 Q.n6 33.746
R274 Q.n5 Q.t3 26.5955
R275 Q.n5 Q.t2 26.5955
R276 Q.n0 Q.t1 24.9236
R277 Q.n0 Q.t0 24.9236
R278 Q.n1 Q 13.5534
R279 Q.n8 Q 12.8005
R280 Q.n3 Q 9.24494
R281 Q.n4 Q 8.33989
R282 Q Q.n8 7.84194
R283 Q.n7 Q 7.46717
R284 Q.n1 Q 7.2005
R285 Q.n2 Q.n1 6.69904
R286 Q.n8 Q.n7 5.1205
R287 Q.n4 Q 4.84898
R288 Q.n6 Q 4.84898
R289 Q.n9 Q 4.84374
R290 Q Q.n9 2.9987
R291 Q.n3 Q 1.96973
R292 Q.n9 Q.n3 0.875714
R293 a_562_413.t0 a_562_413.t1 211.071
R294 a_796_47.t0 a_796_47.t1 60.0005
R295 a_1300_47.t0 a_1300_47.t1 60.0005
C0 SET_B VGND 0.335297f
C1 VPWR VGND 0.066998f
C2 SET_B Q 9.77e-19
C3 VPWR Q 0.217422f
C4 VGND Q 0.14947f
C5 a_1178_261# VPB 0.11585f
C6 VPB CLK 0.069834f
C7 VPB D 0.048468f
C8 VPB SET_B 0.143014f
C9 a_1178_261# SET_B 0.124895f
C10 VPB VPWR 0.21143f
C11 a_1178_261# VPWR 0.125191f
C12 VPB VGND 0.011162f
C13 CLK VPWR 0.017454f
C14 a_1178_261# VGND 0.065287f
C15 CLK VGND 0.017215f
C16 VPB Q 0.008678f
C17 D VPWR 0.015788f
C18 D VGND 0.013952f
C19 SET_B VPWR 0.079638f
C20 Q VNB 0.052086f
C21 VGND VNB 1.07496f
C22 VPWR VNB 0.888166f
C23 SET_B VNB 0.246461f
C24 D VNB 0.107124f
C25 CLK VNB 0.195914f
C26 VPB VNB 1.9337f
C27 a_1178_261# VNB 0.129158f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_4 VPB VNB VPWR VGND Q CLK D SET_B
X0 a_1178_261.t1 a_1028_413.t5 VPWR.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X1 VGND.t1 a_652_21.t3 a_586_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X2 VPWR.t5 a_1028_413.t6 a_1598_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_1178_261.t0 a_1028_413.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X4 a_956_413.t0 a_476_47.t4 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_1136_413.t0 a_193_47.t2 a_1028_413.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X6 VPWR.t8 a_476_47.t5 a_652_21.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR.t2 CLK.t0 a_27_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_586_47.t1 a_193_47.t3 a_476_47.t0 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X9 Q.t0 a_1598_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_1056_47.t1 a_476_47.t6 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_476_47.t1 a_27_47.t2 a_381_47.t1 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X12 a_381_47.t3 D.t0 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X13 a_652_21.t0 SET_B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X14 a_1224_47.t0 a_27_47.t3 a_1028_413.t3 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_562_413.t1 a_27_47.t4 a_476_47.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_1028_413.t1 a_193_47.t4 a_1056_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47.t2 a_193_47.t5 a_381_47.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X18 a_1296_47.t1 a_1178_261.t2 a_1224_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 VGND.t2 a_1028_413.t8 a_1598_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 a_193_47.t0 a_27_47.t5 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR.t4 a_652_21.t4 a_562_413.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X22 VGND.t5 SET_B.t1 a_1296_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 a_1028_413.t4 a_27_47.t6 a_956_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 VPWR.t3 a_1178_261.t3 a_1136_413.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 a_193_47.t1 a_27_47.t7 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 Q.t1 a_1598_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X27 a_796_47.t0 SET_B.t2 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X28 a_381_47.t2 D.t1 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 a_652_21.t2 a_476_47.t7 a_796_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VPWR.t9 SET_B.t3 a_1028_413.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND.t8 CLK.t1 a_27_47.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1028_413.n4 a_1028_413.t2 726.158
R1 a_1028_413.n5 a_1028_413.n4 610.48
R2 a_1028_413.n3 a_1028_413.n0 287.401
R3 a_1028_413.n1 a_1028_413.t6 237.787
R4 a_1028_413.n3 a_1028_413.n2 228.209
R5 a_1028_413.n1 a_1028_413.t8 208.868
R6 a_1028_413.n2 a_1028_413.t5 205.654
R7 a_1028_413.n2 a_1028_413.t7 189.588
R8 a_1028_413.n2 a_1028_413.n1 137.298
R9 a_1028_413.t0 a_1028_413.n5 119.608
R10 a_1028_413.n4 a_1028_413.n3 94.8711
R11 a_1028_413.n5 a_1028_413.t4 63.3219
R12 a_1028_413.n0 a_1028_413.t3 47.1434
R13 a_1028_413.n0 a_1028_413.t1 47.1434
R14 VPWR.n38 VPWR.t10 721.837
R15 VPWR.n8 VPWR.t3 648.322
R16 VPWR.n18 VPWR.n11 604.783
R17 VPWR.n40 VPWR.n1 604.394
R18 VPWR.n6 VPWR.n5 599.74
R19 VPWR.n31 VPWR.n30 585
R20 VPWR.n13 VPWR.t5 371.82
R21 VPWR.n14 VPWR.t1 342.308
R22 VPWR.n30 VPWR.t0 91.4648
R23 VPWR.n11 VPWR.t9 91.4648
R24 VPWR.n30 VPWR.t4 86.7743
R25 VPWR.n5 VPWR.t7 63.3219
R26 VPWR.n5 VPWR.t8 63.3219
R27 VPWR.n1 VPWR.t11 41.5552
R28 VPWR.n1 VPWR.t2 41.5552
R29 VPWR.n33 VPWR.n3 34.6358
R30 VPWR.n37 VPWR.n3 34.6358
R31 VPWR.n24 VPWR.n23 34.6358
R32 VPWR.n25 VPWR.n24 34.6358
R33 VPWR.n17 VPWR.n12 34.6358
R34 VPWR.n33 VPWR.n32 33.5954
R35 VPWR.n11 VPWR.t6 32.8338
R36 VPWR.n29 VPWR.n6 31.624
R37 VPWR.n13 VPWR.n12 30.8711
R38 VPWR.n20 VPWR.n19 27.873
R39 VPWR.n19 VPWR.n18 25.6005
R40 VPWR.n39 VPWR.n38 22.9652
R41 VPWR.n40 VPWR.n39 22.9652
R42 VPWR.n38 VPWR.n37 21.4593
R43 VPWR.n18 VPWR.n17 18.824
R44 VPWR.n23 VPWR.n8 18.735
R45 VPWR.n25 VPWR.n6 12.8005
R46 VPWR.n31 VPWR.n29 12.5335
R47 VPWR.n15 VPWR.n12 9.3005
R48 VPWR.n17 VPWR.n16 9.3005
R49 VPWR.n18 VPWR.n10 9.3005
R50 VPWR.n19 VPWR.n9 9.3005
R51 VPWR.n21 VPWR.n20 9.3005
R52 VPWR.n23 VPWR.n22 9.3005
R53 VPWR.n24 VPWR.n7 9.3005
R54 VPWR.n26 VPWR.n25 9.3005
R55 VPWR.n27 VPWR.n6 9.3005
R56 VPWR.n29 VPWR.n28 9.3005
R57 VPWR.n32 VPWR.n4 9.3005
R58 VPWR.n34 VPWR.n33 9.3005
R59 VPWR.n35 VPWR.n3 9.3005
R60 VPWR.n37 VPWR.n36 9.3005
R61 VPWR.n38 VPWR.n2 9.3005
R62 VPWR.n39 VPWR.n0 9.3005
R63 VPWR.n41 VPWR.n40 7.12063
R64 VPWR.n14 VPWR.n13 6.66355
R65 VPWR.n32 VPWR.n31 3.37505
R66 VPWR.n20 VPWR.n8 0.815045
R67 VPWR.n15 VPWR.n14 0.192575
R68 VPWR.n41 VPWR.n0 0.148519
R69 VPWR.n16 VPWR.n15 0.120292
R70 VPWR.n16 VPWR.n10 0.120292
R71 VPWR.n10 VPWR.n9 0.120292
R72 VPWR.n21 VPWR.n9 0.120292
R73 VPWR.n22 VPWR.n21 0.120292
R74 VPWR.n22 VPWR.n7 0.120292
R75 VPWR.n26 VPWR.n7 0.120292
R76 VPWR.n27 VPWR.n26 0.120292
R77 VPWR.n28 VPWR.n27 0.120292
R78 VPWR.n28 VPWR.n4 0.120292
R79 VPWR.n34 VPWR.n4 0.120292
R80 VPWR.n35 VPWR.n34 0.120292
R81 VPWR.n36 VPWR.n35 0.120292
R82 VPWR.n36 VPWR.n2 0.120292
R83 VPWR.n2 VPWR.n0 0.120292
R84 VPWR VPWR.n41 0.114842
R85 a_1178_261.n0 a_1178_261.t2 381.183
R86 a_1178_261.t1 a_1178_261.n1 371.185
R87 a_1178_261.n1 a_1178_261.t0 285.87
R88 a_1178_261.n1 a_1178_261.n0 265.774
R89 a_1178_261.n0 a_1178_261.t3 169.453
R90 VPB.t4 VPB.t1 1275.55
R91 VPB.t5 VPB.t4 556.386
R92 VPB.t9 VPB.t10 556.386
R93 VPB.t15 VPB.t14 556.386
R94 VPB.t12 VPB.t3 355.14
R95 VPB.t13 VPB.t6 319.627
R96 VPB.t3 VPB.t0 313.707
R97 VPB.t14 VPB.t11 287.072
R98 VPB.t10 VPB.t5 284.113
R99 VPB.t8 VPB.t7 248.599
R100 VPB.t0 VPB.t8 248.599
R101 VPB.t11 VPB.t12 248.599
R102 VPB.t2 VPB.t15 248.599
R103 VPB.t6 VPB.t9 213.084
R104 VPB.t7 VPB.t13 213.084
R105 VPB VPB.t2 142.056
R106 a_652_21.n2 a_652_21.n1 594.413
R107 a_652_21.n0 a_652_21.t3 387.961
R108 a_652_21.n1 a_652_21.t2 334.156
R109 a_652_21.n1 a_652_21.n0 187.072
R110 a_652_21.n0 a_652_21.t4 143.746
R111 a_652_21.n2 a_652_21.t1 63.3219
R112 a_652_21.t0 a_652_21.n2 63.3219
R113 a_586_47.t0 a_586_47.t1 93.5174
R114 VGND.n12 VGND.t0 285.728
R115 VGND.n36 VGND.t7 280.51
R116 VGND.n11 VGND.t2 256.353
R117 VGND.n25 VGND.t4 237.877
R118 VGND.n39 VGND.n38 199.739
R119 VGND.n9 VGND.n8 185
R120 VGND.n4 VGND.n3 185
R121 VGND.n3 VGND.t1 81.4291
R122 VGND.n8 VGND.t5 67.1434
R123 VGND.n8 VGND.t3 55.3018
R124 VGND.n3 VGND.t6 38.5719
R125 VGND.n38 VGND.t9 38.5719
R126 VGND.n38 VGND.t8 38.5719
R127 VGND.n15 VGND.n14 34.6358
R128 VGND.n20 VGND.n19 34.6358
R129 VGND.n21 VGND.n20 34.6358
R130 VGND.n21 VGND.n6 34.6358
R131 VGND.n31 VGND.n30 34.6358
R132 VGND.n32 VGND.n31 34.6358
R133 VGND.n32 VGND.n1 34.6358
R134 VGND.n14 VGND.n11 30.8711
R135 VGND.n27 VGND.n26 28.6616
R136 VGND.n26 VGND.n25 27.8593
R137 VGND.n16 VGND.n15 23.5154
R138 VGND.n37 VGND.n36 22.9652
R139 VGND.n39 VGND.n37 22.9652
R140 VGND.n36 VGND.n1 21.4593
R141 VGND.n25 VGND.n6 15.8123
R142 VGND.n30 VGND.n4 13.8312
R143 VGND.n14 VGND.n13 9.3005
R144 VGND.n15 VGND.n10 9.3005
R145 VGND.n17 VGND.n16 9.3005
R146 VGND.n19 VGND.n18 9.3005
R147 VGND.n20 VGND.n7 9.3005
R148 VGND.n22 VGND.n21 9.3005
R149 VGND.n23 VGND.n6 9.3005
R150 VGND.n25 VGND.n24 9.3005
R151 VGND.n26 VGND.n5 9.3005
R152 VGND.n28 VGND.n27 9.3005
R153 VGND.n30 VGND.n29 9.3005
R154 VGND.n31 VGND.n2 9.3005
R155 VGND.n33 VGND.n32 9.3005
R156 VGND.n34 VGND.n1 9.3005
R157 VGND.n36 VGND.n35 9.3005
R158 VGND.n37 VGND.n0 9.3005
R159 VGND.n19 VGND.n9 7.97588
R160 VGND.n40 VGND.n39 7.12063
R161 VGND.n12 VGND.n11 6.66355
R162 VGND.n27 VGND.n4 4.51198
R163 VGND.n16 VGND.n9 1.08358
R164 VGND.n13 VGND.n12 0.192575
R165 VGND.n40 VGND.n0 0.148519
R166 VGND.n13 VGND.n10 0.120292
R167 VGND.n17 VGND.n10 0.120292
R168 VGND.n18 VGND.n17 0.120292
R169 VGND.n18 VGND.n7 0.120292
R170 VGND.n22 VGND.n7 0.120292
R171 VGND.n23 VGND.n22 0.120292
R172 VGND.n24 VGND.n23 0.120292
R173 VGND.n24 VGND.n5 0.120292
R174 VGND.n28 VGND.n5 0.120292
R175 VGND.n29 VGND.n28 0.120292
R176 VGND.n29 VGND.n2 0.120292
R177 VGND.n33 VGND.n2 0.120292
R178 VGND.n34 VGND.n33 0.120292
R179 VGND.n35 VGND.n34 0.120292
R180 VGND.n35 VGND.n0 0.120292
R181 VGND VGND.n40 0.114842
R182 VNB.t2 VNB.t0 6137.22
R183 VNB.t3 VNB.t2 2677.02
R184 VNB.t7 VNB.t6 2677.02
R185 VNB.t15 VNB.t12 2677.02
R186 VNB.t10 VNB.t3 1765.7
R187 VNB.t1 VNB.t11 1623.3
R188 VNB.t9 VNB.t4 1566.34
R189 VNB.t5 VNB.t14 1366.99
R190 VNB.t4 VNB.t1 1366.99
R191 VNB.t12 VNB.t9 1352.75
R192 VNB.t13 VNB.t15 1196.12
R193 VNB.t8 VNB.t10 1025.24
R194 VNB.t14 VNB.t8 1025.24
R195 VNB.t6 VNB.t5 1025.24
R196 VNB.t11 VNB.t7 1025.24
R197 VNB VNB.t13 683.495
R198 a_1598_47.t1 a_1598_47.n21 401.825
R199 a_1598_47.n21 a_1598_47.t0 257.108
R200 a_1598_47.n7 a_1598_47.t3 221.72
R201 a_1598_47.n11 a_1598_47.n9 221.72
R202 a_1598_47.n6 a_1598_47.n4 221.72
R203 a_1598_47.n1 a_1598_47.n2 221.72
R204 a_1598_47.n18 a_1598_47.n16 221.72
R205 a_1598_47.n13 a_1598_47.n8 171.782
R206 a_1598_47.n20 a_1598_47.n19 152
R207 a_1598_47.n1 a_1598_47.n0 152
R208 a_1598_47.n15 a_1598_47.n14 152
R209 a_1598_47.n13 a_1598_47.n12 152
R210 a_1598_47.n7 a_1598_47.t2 149.421
R211 a_1598_47.n11 a_1598_47.n10 149.421
R212 a_1598_47.n6 a_1598_47.n5 149.421
R213 a_1598_47.n1 a_1598_47.n3 149.421
R214 a_1598_47.n18 a_1598_47.n17 149.421
R215 a_1598_47.n1 a_1598_47.n15 60.6968
R216 a_1598_47.n19 a_1598_47.n1 60.6968
R217 a_1598_47.n12 a_1598_47.n6 48.2005
R218 a_1598_47.n8 a_1598_47.n7 41.0598
R219 a_1598_47.n21 a_1598_47.n20 35.4914
R220 a_1598_47.n11 a_1598_47.n8 33.919
R221 a_1598_47.n12 a_1598_47.n11 26.7783
R222 a_1598_47.n14 a_1598_47.n13 19.7823
R223 a_1598_47.n14 a_1598_47.n0 19.7823
R224 a_1598_47.n20 a_1598_47.n0 19.7823
R225 a_1598_47.n19 a_1598_47.n18 16.0672
R226 a_1598_47.n15 a_1598_47.n6 12.4968
R227 Q.n2 Q.t1 354.445
R228 Q.n0 Q.t0 209.923
R229 Q.n1 Q 127.639
R230 Q.n3 Q 120.064
R231 Q.n5 Q 12.244
R232 Q.n3 Q 8.41193
R233 Q.n0 Q 7.49764
R234 Q Q.n2 6.78064
R235 Q Q.n5 6.67876
R236 Q.n2 Q 5.56925
R237 Q Q.n0 4.93764
R238 Q.n4 Q.n3 3.10907
R239 Q.n5 Q.n1 3.10907
R240 Q Q.n4 1.3918
R241 Q.n1 Q 1.2805
R242 Q.n4 Q 0.914786
R243 a_476_47.n4 a_476_47.n3 707.533
R244 a_476_47.n1 a_476_47.t6 344.899
R245 a_476_47.n2 a_476_47.t4 289.493
R246 a_476_47.n3 a_476_47.n0 288.925
R247 a_476_47.n2 a_476_47.t5 228.148
R248 a_476_47.n3 a_476_47.n2 214.781
R249 a_476_47.n2 a_476_47.n1 105.749
R250 a_476_47.n1 a_476_47.t7 93.1872
R251 a_476_47.n0 a_476_47.t1 70.0005
R252 a_476_47.n0 a_476_47.t0 63.3338
R253 a_476_47.n4 a_476_47.t3 63.3219
R254 a_476_47.t2 a_476_47.n4 63.3219
R255 a_956_413.t0 a_956_413.t1 98.5005
R256 a_193_47.n1 a_193_47.t5 533.949
R257 a_193_47.t1 a_193_47.n3 424.863
R258 a_193_47.n0 a_193_47.t2 373.666
R259 a_193_47.n0 a_193_47.t4 264.029
R260 a_193_47.n3 a_193_47.t0 242.915
R261 a_193_47.n2 a_193_47.n0 189.742
R262 a_193_47.n2 a_193_47.n1 164.226
R263 a_193_47.n1 a_193_47.t3 141.923
R264 a_193_47.n3 a_193_47.n2 10.842
R265 a_1136_413.t0 a_1136_413.t1 98.5005
R266 CLK.n0 CLK.t0 270.457
R267 CLK.n0 CLK.t1 235.109
R268 CLK.n1 CLK.n0 152
R269 CLK.n1 CLK 7.6805
R270 CLK CLK.n1 4.75479
R271 a_27_47.n2 a_27_47.t3 421.01
R272 a_27_47.t1 a_27_47.n5 390.067
R273 a_27_47.n3 a_27_47.t2 311.954
R274 a_27_47.n3 a_27_47.t4 308.168
R275 a_27_47.n2 a_27_47.t6 300.252
R276 a_27_47.n1 a_27_47.t0 287.998
R277 a_27_47.n0 a_27_47.t7 263.173
R278 a_27_47.n0 a_27_47.t5 227.826
R279 a_27_47.n1 a_27_47.n0 152
R280 a_27_47.n5 a_27_47.n1 35.3396
R281 a_27_47.n4 a_27_47.n2 17.2377
R282 a_27_47.n5 a_27_47.n4 10.8331
R283 a_27_47.n4 a_27_47.n3 9.3005
R284 a_1056_47.t0 a_1056_47.t1 60.0005
R285 a_381_47.n1 a_381_47.n0 644.056
R286 a_381_47.n1 a_381_47.t0 95.0032
R287 a_381_47.n0 a_381_47.t1 63.3338
R288 a_381_47.t3 a_381_47.n1 31.6371
R289 a_381_47.n0 a_381_47.t2 26.7713
R290 D.n0 D.t0 264.029
R291 D.n0 D.t1 174.056
R292 D.n1 D.n0 152
R293 D.n1 D 8.58587
R294 D D.n1 2.02977
R295 SET_B.n0 SET_B.t0 389.618
R296 SET_B.n1 SET_B.t3 386.892
R297 SET_B.n2 SET_B.n1 186.411
R298 SET_B.n2 SET_B.n0 156.06
R299 SET_B.n1 SET_B.t1 148.35
R300 SET_B.n0 SET_B.t2 142.569
R301 SET_B SET_B.n2 2.65416
R302 a_1224_47.t0 a_1224_47.t1 60.0005
R303 a_562_413.t0 a_562_413.t1 211.071
R304 a_1296_47.t0 a_1296_47.t1 60.0005
R305 a_796_47.t0 a_796_47.t1 60.0005
C0 VPB SET_B 0.142976f
C1 VPB VPWR 0.231731f
C2 VPB VGND 0.013642f
C3 CLK VPWR 0.019428f
C4 VPB Q 0.023621f
C5 CLK VGND 0.019435f
C6 D VPWR 0.015788f
C7 SET_B VPWR 0.079577f
C8 D VGND 0.013952f
C9 SET_B VGND 0.335541f
C10 VPWR VGND 0.09407f
C11 SET_B Q 0.00107f
C12 VPWR Q 0.464678f
C13 VGND Q 0.315177f
C14 VPB CLK 0.070197f
C15 VPB D 0.048468f
C16 Q VNB 0.117532f
C17 VGND VNB 1.19869f
C18 VPWR VNB 0.971775f
C19 SET_B VNB 0.243523f
C20 D VNB 0.107124f
C21 CLK VNB 0.195843f
C22 VPB VNB 2.19949f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxbp_1 VGND VPWR VNB VPB Q_N Q D CLK
X0 Q.t1 a_1059_315.t2 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413.t1 a_193_47.t2 a_634_159.t1 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413.t0 a_27_47.t2 a_466_413.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR.t1 CLK.t0 a_27_47.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_381_47.t2 D.t0 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t1 a_634_159.t4 a_592_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6 a_466_413.t1 a_193_47.t3 a_381_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7 VPWR.t9 a_634_159.t5 a_561_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8 a_634_159.t3 a_466_413.t4 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9 Q.t0 a_1059_315.t3 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t5 a_1059_315.t4 a_1490_369.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_634_159.t0 a_466_413.t5 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413.t0 a_193_47.t4 a_891_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND.t6 a_1059_315.t5 a_1017_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47.t0 a_27_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413.t2 a_27_47.t4 a_634_159.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 VPWR.t0 a_891_413.t4 a_1059_315.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X17 a_592_47.t0 a_193_47.t5 a_466_413.t0 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X18 VPWR.t7 a_1059_315.t6 a_975_413.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_1017_47.t0 a_27_47.t5 a_891_413.t3 VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 a_193_47.t1 a_27_47.t6 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 a_466_413.t3 a_27_47.t7 a_381_47.t1 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 VGND.t0 a_891_413.t5 a_1059_315.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 Q_N.t1 a_1490_369.t2 VGND.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X24 a_381_47.t3 D.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 Q_N.t0 a_1490_369.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X26 VGND.t8 CLK.t1 a_27_47.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR.t6 a_1059_315.t7 a_1490_369.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
R0 a_1059_315.n3 a_1059_315.t5 382.745
R1 a_1059_315.n0 a_1059_315.t7 258.798
R2 a_1059_315.t0 a_1059_315.n4 226.315
R3 a_1059_315.n1 a_1059_315.t3 213.542
R4 a_1059_315.n4 a_1059_315.n3 173.959
R5 a_1059_315.n2 a_1059_315.n1 173.916
R6 a_1059_315.n0 a_1059_315.t4 166.388
R7 a_1059_315.n2 a_1059_315.t1 149.642
R8 a_1059_315.n1 a_1059_315.t2 139.78
R9 a_1059_315.n3 a_1059_315.t6 138.53
R10 a_1059_315.n1 a_1059_315.n0 129.264
R11 a_1059_315.n4 a_1059_315.n2 16.6232
R12 VGND.n6 VGND.t6 251
R13 VGND.n27 VGND.t3 243.028
R14 VGND.n10 VGND.n9 218.506
R15 VGND.n8 VGND.n7 206.251
R16 VGND.n30 VGND.n29 199.739
R17 VGND.n21 VGND.n4 199.53
R18 VGND.n4 VGND.t9 74.8666
R19 VGND.n7 VGND.t5 54.2862
R20 VGND.n4 VGND.t1 40.0005
R21 VGND.n29 VGND.t2 38.5719
R22 VGND.n29 VGND.t8 38.5719
R23 VGND.n16 VGND.n15 34.6358
R24 VGND.n17 VGND.n16 34.6358
R25 VGND.n17 VGND.n3 34.6358
R26 VGND.n23 VGND.n22 34.6358
R27 VGND.n23 VGND.n1 34.6358
R28 VGND.n11 VGND.n10 32.7534
R29 VGND.n11 VGND.n6 31.2476
R30 VGND.n22 VGND.n21 30.8711
R31 VGND.n27 VGND.n1 27.4829
R32 VGND.n7 VGND.t4 25.9346
R33 VGND.n9 VGND.t7 24.9236
R34 VGND.n9 VGND.t0 24.9236
R35 VGND.n28 VGND.n27 22.9652
R36 VGND.n30 VGND.n28 22.9652
R37 VGND.n15 VGND.n6 22.2123
R38 VGND.n21 VGND.n3 10.5417
R39 VGND.n10 VGND.n8 9.42894
R40 VGND.n28 VGND.n0 9.3005
R41 VGND.n27 VGND.n26 9.3005
R42 VGND.n12 VGND.n11 9.3005
R43 VGND.n13 VGND.n6 9.3005
R44 VGND.n15 VGND.n14 9.3005
R45 VGND.n16 VGND.n5 9.3005
R46 VGND.n18 VGND.n17 9.3005
R47 VGND.n19 VGND.n3 9.3005
R48 VGND.n21 VGND.n20 9.3005
R49 VGND.n22 VGND.n2 9.3005
R50 VGND.n24 VGND.n23 9.3005
R51 VGND.n25 VGND.n1 9.3005
R52 VGND.n31 VGND.n30 7.12063
R53 VGND.n12 VGND.n8 0.201218
R54 VGND.n31 VGND.n0 0.148519
R55 VGND.n13 VGND.n12 0.120292
R56 VGND.n14 VGND.n13 0.120292
R57 VGND.n14 VGND.n5 0.120292
R58 VGND.n18 VGND.n5 0.120292
R59 VGND.n19 VGND.n18 0.120292
R60 VGND.n20 VGND.n19 0.120292
R61 VGND.n20 VGND.n2 0.120292
R62 VGND.n24 VGND.n2 0.120292
R63 VGND.n25 VGND.n24 0.120292
R64 VGND.n26 VGND.n25 0.120292
R65 VGND.n26 VGND.n0 0.120292
R66 VGND VGND.n31 0.114842
R67 Q.n0 Q.t0 317.469
R68 Q.n0 Q.t1 129.078
R69 Q Q.n0 5.84085
R70 VNB.t9 VNB.t0 2705.5
R71 VNB.t11 VNB.t10 2677.02
R72 VNB.t2 VNB.t5 2677.02
R73 VNB.t1 VNB.t13 1694.5
R74 VNB.t5 VNB.t4 1594.82
R75 VNB.t6 VNB.t3 1509.39
R76 VNB.t13 VNB.t6 1438.19
R77 VNB.t7 VNB.t1 1409.71
R78 VNB.t4 VNB.t7 1409.71
R79 VNB.t10 VNB.t8 1352.75
R80 VNB.t3 VNB.t9 1352.75
R81 VNB.t0 VNB.t11 1196.12
R82 VNB.t12 VNB.t2 1196.12
R83 VNB VNB.t12 683.495
R84 a_193_47.n1 a_193_47.t5 407.217
R85 a_193_47.t1 a_193_47.n3 392.493
R86 a_193_47.n0 a_193_47.t4 308.651
R87 a_193_47.n0 a_193_47.t2 298.373
R88 a_193_47.n3 a_193_47.t0 294.144
R89 a_193_47.n1 a_193_47.t3 273.572
R90 a_193_47.n2 a_193_47.n1 170.9
R91 a_193_47.n2 a_193_47.n0 11.4492
R92 a_193_47.n3 a_193_47.n2 10.2617
R93 a_634_159.n3 a_634_159.n2 674.014
R94 a_634_159.n1 a_634_159.t5 406.401
R95 a_634_159.n2 a_634_159.n0 213.988
R96 a_634_159.n2 a_634_159.n1 180.161
R97 a_634_159.n1 a_634_159.t4 130.054
R98 a_634_159.n3 a_634_159.t2 89.1195
R99 a_634_159.n0 a_634_159.t1 71.6672
R100 a_634_159.t0 a_634_159.n3 37.5243
R101 a_634_159.n0 a_634_159.t3 28.438
R102 a_891_413.n3 a_891_413.n2 696.059
R103 a_891_413.n2 a_891_413.n0 258.788
R104 a_891_413.n2 a_891_413.n1 251.109
R105 a_891_413.n1 a_891_413.t4 212.081
R106 a_891_413.n1 a_891_413.t5 141.242
R107 a_891_413.n0 a_891_413.t3 76.6672
R108 a_891_413.t0 a_891_413.n3 63.3219
R109 a_891_413.n3 a_891_413.t2 63.3219
R110 a_891_413.n0 a_891_413.t1 50.0005
R111 a_27_47.n2 a_27_47.t5 443.44
R112 a_27_47.t1 a_27_47.n5 390.067
R113 a_27_47.n3 a_27_47.t7 345.305
R114 a_27_47.n3 a_27_47.t2 296.969
R115 a_27_47.n1 a_27_47.t0 287.998
R116 a_27_47.n0 a_27_47.t6 263.173
R117 a_27_47.n2 a_27_47.t4 254.389
R118 a_27_47.n0 a_27_47.t3 227.826
R119 a_27_47.n4 a_27_47.n2 193.59
R120 a_27_47.n1 a_27_47.n0 152
R121 a_27_47.n5 a_27_47.n1 35.3396
R122 a_27_47.n4 a_27_47.n3 12.4401
R123 a_27_47.n5 a_27_47.n4 11.0742
R124 a_466_413.n3 a_466_413.n2 695.683
R125 a_466_413.n2 a_466_413.n1 298.361
R126 a_466_413.n0 a_466_413.t4 230.484
R127 a_466_413.n0 a_466_413.t5 196.013
R128 a_466_413.n2 a_466_413.n0 168.738
R129 a_466_413.t1 a_466_413.n3 79.7386
R130 a_466_413.n3 a_466_413.t2 72.7029
R131 a_466_413.n1 a_466_413.t0 70.0005
R132 a_466_413.n1 a_466_413.t3 45.0005
R133 a_561_413.t0 a_561_413.t1 171.202
R134 VPB.t10 VPB.t0 624.456
R135 VPB.t11 VPB.t9 556.386
R136 VPB.t5 VPB.t8 556.386
R137 VPB.t13 VPB.t4 390.654
R138 VPB.t1 VPB.t10 337.384
R139 VPB.t7 VPB.t13 304.829
R140 VPB.t9 VPB.t3 287.072
R141 VPB.t4 VPB.t6 281.154
R142 VPB.t2 VPB.t7 281.154
R143 VPB.t8 VPB.t2 251.559
R144 VPB.t0 VPB.t11 248.599
R145 VPB.t6 VPB.t1 248.599
R146 VPB.t12 VPB.t5 248.599
R147 VPB VPB.t12 142.056
R148 CLK.n0 CLK.t0 294.557
R149 CLK.n0 CLK.t1 211.01
R150 CLK CLK.n0 153.97
R151 VPWR.n15 VPWR.t7 667.734
R152 VPWR.n29 VPWR.t5 666.677
R153 VPWR.n31 VPWR.n1 604.394
R154 VPWR.n10 VPWR.n9 333.348
R155 VPWR.n22 VPWR.n5 320.976
R156 VPWR.n12 VPWR.n11 246.825
R157 VPWR.n5 VPWR.t9 113.98
R158 VPWR.n11 VPWR.t6 61.9872
R159 VPWR.n1 VPWR.t4 41.5552
R160 VPWR.n1 VPWR.t1 41.5552
R161 VPWR.n5 VPWR.t3 35.4605
R162 VPWR.n17 VPWR.n16 34.6358
R163 VPWR.n17 VPWR.n6 34.6358
R164 VPWR.n21 VPWR.n6 34.6358
R165 VPWR.n24 VPWR.n23 34.6358
R166 VPWR.n24 VPWR.n3 34.6358
R167 VPWR.n28 VPWR.n3 34.6358
R168 VPWR.n14 VPWR.n10 32.0005
R169 VPWR.n15 VPWR.n14 30.4946
R170 VPWR.n11 VPWR.t2 30.1692
R171 VPWR.n29 VPWR.n28 27.4829
R172 VPWR.n9 VPWR.t8 26.5955
R173 VPWR.n9 VPWR.t0 26.5955
R174 VPWR.n31 VPWR.n30 22.9652
R175 VPWR.n30 VPWR.n29 21.8358
R176 VPWR.n23 VPWR.n22 18.4476
R177 VPWR.n22 VPWR.n21 16.1887
R178 VPWR.n16 VPWR.n15 15.0593
R179 VPWR.n12 VPWR.n10 10.1829
R180 VPWR.n14 VPWR.n13 9.3005
R181 VPWR.n15 VPWR.n8 9.3005
R182 VPWR.n16 VPWR.n7 9.3005
R183 VPWR.n18 VPWR.n17 9.3005
R184 VPWR.n19 VPWR.n6 9.3005
R185 VPWR.n21 VPWR.n20 9.3005
R186 VPWR.n23 VPWR.n4 9.3005
R187 VPWR.n25 VPWR.n24 9.3005
R188 VPWR.n26 VPWR.n3 9.3005
R189 VPWR.n28 VPWR.n27 9.3005
R190 VPWR.n29 VPWR.n2 9.3005
R191 VPWR.n30 VPWR.n0 9.3005
R192 VPWR.n32 VPWR.n31 7.12063
R193 VPWR.n13 VPWR.n12 0.200304
R194 VPWR.n32 VPWR.n0 0.148519
R195 VPWR.n13 VPWR.n8 0.120292
R196 VPWR.n8 VPWR.n7 0.120292
R197 VPWR.n18 VPWR.n7 0.120292
R198 VPWR.n19 VPWR.n18 0.120292
R199 VPWR.n20 VPWR.n19 0.120292
R200 VPWR.n20 VPWR.n4 0.120292
R201 VPWR.n25 VPWR.n4 0.120292
R202 VPWR.n26 VPWR.n25 0.120292
R203 VPWR.n27 VPWR.n26 0.120292
R204 VPWR.n27 VPWR.n2 0.120292
R205 VPWR.n2 VPWR.n0 0.120292
R206 VPWR VPWR.n32 0.114842
R207 D.n0 D.t1 302.731
R208 D.n0 D.t0 212.757
R209 D D.n0 170.058
R210 a_381_47.n1 a_381_47.n0 896.306
R211 a_381_47.n0 a_381_47.t1 90.0005
R212 a_381_47.t0 a_381_47.n1 65.6672
R213 a_381_47.n1 a_381_47.t2 63.3219
R214 a_381_47.n0 a_381_47.t3 31.3935
R215 a_592_47.t1 a_592_47.t0 99.7268
R216 a_1490_369.t0 a_1490_369.n1 389.671
R217 a_1490_369.n1 a_1490_369.t1 254.625
R218 a_1490_369.n0 a_1490_369.t3 236.934
R219 a_1490_369.n1 a_1490_369.n0 173.528
R220 a_1490_369.n0 a_1490_369.t2 164.633
R221 a_975_413.t0 a_975_413.t1 197
R222 a_1017_47.t1 a_1017_47.t0 93.0601
R223 Q_N Q_N.t1 259.565
R224 Q_N Q_N.t0 233.177
C0 VGND VPB 0.015716f
C1 VPB CLK 0.070057f
C2 VGND CLK 0.019463f
C3 Q VPB 0.011402f
C4 VGND Q 0.079189f
C5 VPB D 0.096334f
C6 Q_N VPB 0.011861f
C7 VGND D 0.038993f
C8 VGND Q_N 0.065009f
C9 VPB VPWR 0.200637f
C10 VGND VPWR 0.093137f
C11 CLK VPWR 0.019411f
C12 Q VPWR 0.111692f
C13 D VPWR 0.025067f
C14 Q_N VPWR 0.128202f
C15 Q_N VNB 0.093273f
C16 Q VNB 0.007853f
C17 VGND VNB 0.985366f
C18 VPWR VNB 0.794315f
C19 D VNB 0.142509f
C20 CLK VNB 0.195983f
C21 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxbp_2 VGND VPWR VNB VPB Q_N Q D CLK
X0 Q.t2 a_1059_315.t2 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413.t1 a_193_47.t2 a_634_159.t0 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413.t0 a_27_47.t2 a_466_413.t3 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_381_47.t1 D.t0 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t2 a_634_159.t4 a_592_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6 VPWR.t10 a_1589_47# Q_N.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t6 a_1059_315.t3 Q.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t10 a_1589_47# Q_N.t3 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_466_413.t0 a_193_47.t3 a_381_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10 VPWR.t8 a_634_159.t5 a_561_413.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11 a_634_159.t1 a_466_413.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12 Q.t0 a_1059_315.t4 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_634_159.t2 a_466_413.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14 a_975_413.t0 a_193_47.t4 a_891_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 Q_N.t0 a_1589_47# VPWR.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X16 VGND.t5 a_1059_315.t5 a_1017_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X17 a_193_47.t0 a_27_47.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_891_413.t2 a_27_47.t4 a_634_159.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X19 VPWR.t2 a_891_413.t4 a_1059_315.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X20 a_592_47.t0 a_193_47.t5 a_466_413.t1 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X21 Q_N.t2 a_1589_47# VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X22 VPWR.t4 a_1059_315.t6 a_975_413.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X23 a_1017_47.t1 a_27_47.t5 a_891_413.t3 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X24 a_193_47.t1 a_27_47.t6 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_466_413.t2 a_27_47.t7 a_381_47.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X26 VGND.t1 a_891_413.t5 a_1059_315.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 VGND.t6 a_1059_315.t7 Q.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_381_47.t2 D.t1 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VGND.t0 CLK.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_1059_315.n7 a_1059_315.t5 382.745
R1 a_1059_315.n2 a_1059_315.n0 258.798
R2 a_1059_315.t1 a_1059_315.n8 226.315
R3 a_1059_315.n5 a_1059_315.t4 213.542
R4 a_1059_315.n4 a_1059_315.t3 212.081
R5 a_1059_315.n8 a_1059_315.n7 173.959
R6 a_1059_315.n6 a_1059_315.n5 173.916
R7 a_1059_315.n2 a_1059_315.n1 167.835
R8 a_1059_315.n6 a_1059_315.t0 149.642
R9 a_1059_315.n3 a_1059_315.n2 140.219
R10 a_1059_315.n5 a_1059_315.t2 139.78
R11 a_1059_315.n3 a_1059_315.t7 139.78
R12 a_1059_315.n7 a_1059_315.t6 138.53
R13 a_1059_315.n5 a_1059_315.n4 59.8853
R14 a_1059_315.n8 a_1059_315.n6 16.6232
R15 a_1059_315.n4 a_1059_315.n3 1.46111
R16 VGND.n6 VGND.t5 251
R17 VGND.n36 VGND.t8 243.028
R18 VGND.n9 VGND.t6 236.276
R19 VGND.n19 VGND.n8 218.506
R20 VGND.n39 VGND.n38 199.739
R21 VGND.n30 VGND.n4 199.53
R22 VGND.n11 VGND.t10 164.058
R23 VGND.n12 VGND.t9 135.594
R24 VGND.n4 VGND.t3 74.8666
R25 VGND.n4 VGND.t2 40.0005
R26 VGND.n38 VGND.t4 38.5719
R27 VGND.n38 VGND.t0 38.5719
R28 VGND.n14 VGND.n13 34.6358
R29 VGND.n18 VGND.n17 34.6358
R30 VGND.n25 VGND.n24 34.6358
R31 VGND.n26 VGND.n25 34.6358
R32 VGND.n26 VGND.n3 34.6358
R33 VGND.n32 VGND.n31 34.6358
R34 VGND.n32 VGND.n1 34.6358
R35 VGND.n20 VGND.n19 32.7534
R36 VGND.n20 VGND.n6 31.2476
R37 VGND.n31 VGND.n30 30.8711
R38 VGND.n36 VGND.n1 27.4829
R39 VGND.n17 VGND.n9 26.7299
R40 VGND.n13 VGND.n12 25.6005
R41 VGND.n8 VGND.t7 24.9236
R42 VGND.n8 VGND.t1 24.9236
R43 VGND.n37 VGND.n36 22.9652
R44 VGND.n39 VGND.n37 22.9652
R45 VGND.n24 VGND.n6 22.2123
R46 VGND.n30 VGND.n3 10.5417
R47 VGND.n37 VGND.n0 9.3005
R48 VGND.n36 VGND.n35 9.3005
R49 VGND.n34 VGND.n1 9.3005
R50 VGND.n33 VGND.n32 9.3005
R51 VGND.n31 VGND.n2 9.3005
R52 VGND.n30 VGND.n29 9.3005
R53 VGND.n28 VGND.n3 9.3005
R54 VGND.n27 VGND.n26 9.3005
R55 VGND.n25 VGND.n5 9.3005
R56 VGND.n24 VGND.n23 9.3005
R57 VGND.n22 VGND.n6 9.3005
R58 VGND.n21 VGND.n20 9.3005
R59 VGND.n18 VGND.n7 9.3005
R60 VGND.n17 VGND.n16 9.3005
R61 VGND.n15 VGND.n14 9.3005
R62 VGND.n13 VGND.n10 9.3005
R63 VGND.n14 VGND.n9 7.90638
R64 VGND.n40 VGND.n39 7.12063
R65 VGND.n12 VGND.n11 6.32884
R66 VGND.n19 VGND.n18 1.88285
R67 VGND.n11 VGND.n10 0.664094
R68 VGND.n40 VGND.n0 0.148519
R69 VGND.n15 VGND.n10 0.120292
R70 VGND.n16 VGND.n15 0.120292
R71 VGND.n16 VGND.n7 0.120292
R72 VGND.n21 VGND.n7 0.120292
R73 VGND.n22 VGND.n21 0.120292
R74 VGND.n23 VGND.n22 0.120292
R75 VGND.n23 VGND.n5 0.120292
R76 VGND.n27 VGND.n5 0.120292
R77 VGND.n28 VGND.n27 0.120292
R78 VGND.n29 VGND.n28 0.120292
R79 VGND.n29 VGND.n2 0.120292
R80 VGND.n33 VGND.n2 0.120292
R81 VGND.n34 VGND.n33 0.120292
R82 VGND.n35 VGND.n34 0.120292
R83 VGND.n35 VGND.n0 0.120292
R84 VGND VGND.n40 0.114842
R85 Q.n1 Q.n0 284.957
R86 Q Q.n2 186.165
R87 Q.n2 Q.n1 185
R88 Q.n0 Q.t3 26.5955
R89 Q.n0 Q.t0 26.5955
R90 Q.n2 Q.t1 24.9236
R91 Q.n2 Q.t2 24.9236
R92 Q Q.n1 12.0247
R93 VNB.t7 VNB.t13 4243.37
R94 VNB.t8 VNB.t1 2705.5
R95 VNB.t6 VNB.t12 2677.02
R96 VNB.t2 VNB.t3 1694.5
R97 VNB.t12 VNB.t11 1594.82
R98 VNB.t4 VNB.t10 1509.39
R99 VNB.t3 VNB.t4 1438.19
R100 VNB.t5 VNB.t2 1409.71
R101 VNB.t11 VNB.t5 1409.71
R102 VNB.t10 VNB.t8 1352.75
R103 VNB.t13 VNB.t14 1196.12
R104 VNB.t9 VNB.t7 1196.12
R105 VNB.t1 VNB.t9 1196.12
R106 VNB.t0 VNB.t6 1196.12
R107 VNB VNB.t0 683.495
R108 a_193_47.n1 a_193_47.t5 407.217
R109 a_193_47.t1 a_193_47.n3 392.493
R110 a_193_47.n0 a_193_47.t4 308.651
R111 a_193_47.n0 a_193_47.t2 298.373
R112 a_193_47.n3 a_193_47.t0 294.144
R113 a_193_47.n1 a_193_47.t3 273.572
R114 a_193_47.n2 a_193_47.n1 170.9
R115 a_193_47.n2 a_193_47.n0 11.4492
R116 a_193_47.n3 a_193_47.n2 10.2617
R117 a_634_159.n3 a_634_159.n2 674.014
R118 a_634_159.n1 a_634_159.t5 406.401
R119 a_634_159.n2 a_634_159.n0 213.988
R120 a_634_159.n2 a_634_159.n1 180.161
R121 a_634_159.n1 a_634_159.t4 130.054
R122 a_634_159.n3 a_634_159.t3 89.1195
R123 a_634_159.n0 a_634_159.t0 71.6672
R124 a_634_159.t2 a_634_159.n3 37.5243
R125 a_634_159.n0 a_634_159.t1 28.438
R126 a_891_413.n3 a_891_413.n2 696.059
R127 a_891_413.n2 a_891_413.n0 258.788
R128 a_891_413.n2 a_891_413.n1 251.109
R129 a_891_413.n1 a_891_413.t4 212.081
R130 a_891_413.n1 a_891_413.t5 141.242
R131 a_891_413.n0 a_891_413.t3 76.6672
R132 a_891_413.t0 a_891_413.n3 63.3219
R133 a_891_413.n3 a_891_413.t2 63.3219
R134 a_891_413.n0 a_891_413.t1 50.0005
R135 a_27_47.n2 a_27_47.t5 443.44
R136 a_27_47.t0 a_27_47.n5 390.067
R137 a_27_47.n3 a_27_47.t7 345.305
R138 a_27_47.n3 a_27_47.t2 296.969
R139 a_27_47.n1 a_27_47.t1 287.998
R140 a_27_47.n0 a_27_47.t6 263.173
R141 a_27_47.n2 a_27_47.t4 254.389
R142 a_27_47.n0 a_27_47.t3 227.826
R143 a_27_47.n4 a_27_47.n2 193.59
R144 a_27_47.n1 a_27_47.n0 152
R145 a_27_47.n5 a_27_47.n1 35.3396
R146 a_27_47.n4 a_27_47.n3 12.4401
R147 a_27_47.n5 a_27_47.n4 11.0742
R148 a_466_413.n3 a_466_413.n2 695.683
R149 a_466_413.n2 a_466_413.n1 298.361
R150 a_466_413.n0 a_466_413.t4 230.484
R151 a_466_413.n0 a_466_413.t5 196.013
R152 a_466_413.n2 a_466_413.n0 168.738
R153 a_466_413.t0 a_466_413.n3 79.7386
R154 a_466_413.n3 a_466_413.t3 72.7029
R155 a_466_413.n1 a_466_413.t1 70.0005
R156 a_466_413.n1 a_466_413.t2 45.0005
R157 a_561_413.t0 a_561_413.t1 171.202
R158 VPB.t8 VPB.t13 887.851
R159 VPB.t6 VPB.t4 624.456
R160 VPB.t9 VPB.t5 556.386
R161 VPB.t12 VPB.t1 390.654
R162 VPB.t2 VPB.t6 337.384
R163 VPB.t11 VPB.t12 304.829
R164 VPB.t1 VPB.t10 281.154
R165 VPB.t3 VPB.t11 281.154
R166 VPB.t5 VPB.t3 251.559
R167 VPB.t13 VPB.t14 248.599
R168 VPB.t7 VPB.t8 248.599
R169 VPB.t4 VPB.t7 248.599
R170 VPB.t10 VPB.t2 248.599
R171 VPB.t0 VPB.t9 248.599
R172 VPB VPB.t0 142.056
R173 CLK.n0 CLK.t0 294.557
R174 CLK.n0 CLK.t1 211.01
R175 CLK CLK.n0 153.97
R176 VPWR.n24 VPWR.t4 667.734
R177 VPWR.n38 VPWR.t3 666.677
R178 VPWR.n40 VPWR.n1 604.394
R179 VPWR.n18 VPWR.t6 361.389
R180 VPWR.n10 VPWR.n9 333.348
R181 VPWR.n31 VPWR.n5 320.976
R182 VPWR.n13 VPWR.t9 270.69
R183 VPWR.n14 VPWR.t10 258.435
R184 VPWR.n5 VPWR.t8 113.98
R185 VPWR.n1 VPWR.t7 41.5552
R186 VPWR.n1 VPWR.t0 41.5552
R187 VPWR.n5 VPWR.t1 35.4605
R188 VPWR.n26 VPWR.n25 34.6358
R189 VPWR.n26 VPWR.n6 34.6358
R190 VPWR.n30 VPWR.n6 34.6358
R191 VPWR.n33 VPWR.n32 34.6358
R192 VPWR.n33 VPWR.n3 34.6358
R193 VPWR.n37 VPWR.n3 34.6358
R194 VPWR.n20 VPWR.n19 34.6358
R195 VPWR.n17 VPWR.n12 34.6358
R196 VPWR.n23 VPWR.n10 32.0005
R197 VPWR.n24 VPWR.n23 30.4946
R198 VPWR.n13 VPWR.n12 28.2358
R199 VPWR.n38 VPWR.n37 27.4829
R200 VPWR.n9 VPWR.t5 26.5955
R201 VPWR.n9 VPWR.t2 26.5955
R202 VPWR.n40 VPWR.n39 22.9652
R203 VPWR.n39 VPWR.n38 21.8358
R204 VPWR.n19 VPWR.n18 19.577
R205 VPWR.n32 VPWR.n31 18.4476
R206 VPWR.n31 VPWR.n30 16.1887
R207 VPWR.n25 VPWR.n24 15.0593
R208 VPWR.n15 VPWR.n12 9.3005
R209 VPWR.n17 VPWR.n16 9.3005
R210 VPWR.n19 VPWR.n11 9.3005
R211 VPWR.n21 VPWR.n20 9.3005
R212 VPWR.n23 VPWR.n22 9.3005
R213 VPWR.n24 VPWR.n8 9.3005
R214 VPWR.n25 VPWR.n7 9.3005
R215 VPWR.n27 VPWR.n26 9.3005
R216 VPWR.n28 VPWR.n6 9.3005
R217 VPWR.n30 VPWR.n29 9.3005
R218 VPWR.n32 VPWR.n4 9.3005
R219 VPWR.n34 VPWR.n33 9.3005
R220 VPWR.n35 VPWR.n3 9.3005
R221 VPWR.n37 VPWR.n36 9.3005
R222 VPWR.n38 VPWR.n2 9.3005
R223 VPWR.n39 VPWR.n0 9.3005
R224 VPWR.n41 VPWR.n40 7.12063
R225 VPWR.n14 VPWR.n13 6.75886
R226 VPWR.n20 VPWR.n10 2.63579
R227 VPWR.n18 VPWR.n17 1.88285
R228 VPWR.n15 VPWR.n14 0.585488
R229 VPWR.n41 VPWR.n0 0.148519
R230 VPWR.n16 VPWR.n15 0.120292
R231 VPWR.n16 VPWR.n11 0.120292
R232 VPWR.n21 VPWR.n11 0.120292
R233 VPWR.n22 VPWR.n21 0.120292
R234 VPWR.n22 VPWR.n8 0.120292
R235 VPWR.n8 VPWR.n7 0.120292
R236 VPWR.n27 VPWR.n7 0.120292
R237 VPWR.n28 VPWR.n27 0.120292
R238 VPWR.n29 VPWR.n28 0.120292
R239 VPWR.n29 VPWR.n4 0.120292
R240 VPWR.n34 VPWR.n4 0.120292
R241 VPWR.n35 VPWR.n34 0.120292
R242 VPWR.n36 VPWR.n35 0.120292
R243 VPWR.n36 VPWR.n2 0.120292
R244 VPWR.n2 VPWR.n0 0.120292
R245 VPWR VPWR.n41 0.114842
R246 D.n0 D.t1 302.731
R247 D.n0 D.t0 212.757
R248 D D.n0 170.058
R249 a_381_47.n1 a_381_47.n0 896.306
R250 a_381_47.n0 a_381_47.t3 90.0005
R251 a_381_47.t0 a_381_47.n1 65.6672
R252 a_381_47.n1 a_381_47.t1 63.3219
R253 a_381_47.n0 a_381_47.t2 31.3935
R254 a_592_47.t1 a_592_47.t0 99.7268
R255 Q_N Q_N.n1 238.083
R256 Q_N Q_N.n0 206.582
R257 Q_N.n0 Q_N.t1 26.5955
R258 Q_N.n0 Q_N.t0 26.5955
R259 Q_N.n1 Q_N.t3 24.9236
R260 Q_N.n1 Q_N.t2 24.9236
R261 a_975_413.t0 a_975_413.t1 197
R262 a_1017_47.t0 a_1017_47.t1 93.0601
C0 CLK VPWR 0.019411f
C1 VPB VGND 0.020423f
C2 CLK VGND 0.019463f
C3 D VPWR 0.025067f
C4 VPB Q 0.006781f
C5 VPB a_1589_47# 0.082201f
C6 VPB Q_N 0.005492f
C7 D VGND 0.038993f
C8 VPWR VGND 0.134094f
C9 VPWR Q 0.172468f
C10 VPWR a_1589_47# 0.224154f
C11 VGND Q 0.105043f
C12 VPWR Q_N 0.209726f
C13 VGND a_1589_47# 0.160615f
C14 VGND Q_N 0.139334f
C15 Q a_1589_47# 0.034766f
C16 Q_N a_1589_47# 0.098975f
C17 VPB CLK 0.070057f
C18 VPB D 0.096334f
C19 VPB VPWR 0.23281f
C20 Q_N VNB 0.024053f
C21 Q VNB 0.005604f
C22 VGND VNB 1.1138f
C23 VPWR VNB 0.910748f
C24 D VNB 0.142509f
C25 CLK VNB 0.195983f
C26 VPB VNB 1.9337f
C27 a_1589_47# VNB 0.22524f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q.t0 a_1059_315# VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413.t2 a_193_47.t2 a_634_159.t3 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413.t1 a_27_47.t2 a_466_413.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR.t3 CLK.t0 a_27_47.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47.t2 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND.t2 a_634_159.t4 a_592_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 a_466_413.t2 a_193_47.t3 a_381_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8 VPWR.t0 a_634_159.t5 a_561_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9 a_634_159.t0 a_466_413.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10 a_634_159.t1 a_466_413.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11 a_975_413.t1 a_193_47.t4 a_891_413.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VGND.t5 a_1059_315# a_1017_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13 a_193_47.t0 a_27_47.t3 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_891_413.t0 a_27_47.t4 a_634_159.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15 a_592_47.t1 a_193_47.t5 a_466_413.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X16 VPWR.t4 a_1059_315# a_975_413.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X17 a_1017_47.t1 a_27_47.t5 a_891_413.t1 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 a_193_47.t1 a_27_47.t6 VPWR.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 a_466_413.t1 a_27_47.t7 a_381_47.t0 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 VGND.t6 a_891_413.t4 a_1059_315# VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_381_47.t3 D.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X22 VGND.t3 CLK.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 VGND.n6 VGND.t5 251
R1 VGND.n22 VGND.t1 243.028
R2 VGND.n8 VGND.n7 226.281
R3 VGND.n25 VGND.n24 199.739
R4 VGND.n16 VGND.n4 199.53
R5 VGND.n4 VGND.t0 74.8666
R6 VGND.n4 VGND.t2 40.0005
R7 VGND.n24 VGND.t7 38.5719
R8 VGND.n24 VGND.t3 38.5719
R9 VGND.n11 VGND.n10 34.6358
R10 VGND.n12 VGND.n11 34.6358
R11 VGND.n12 VGND.n3 34.6358
R12 VGND.n18 VGND.n17 34.6358
R13 VGND.n18 VGND.n1 34.6358
R14 VGND.n17 VGND.n16 30.8711
R15 VGND.n22 VGND.n1 27.4829
R16 VGND.n7 VGND.t4 24.9236
R17 VGND.n7 VGND.t6 24.9236
R18 VGND.n23 VGND.n22 22.9652
R19 VGND.n25 VGND.n23 22.9652
R20 VGND.n10 VGND.n6 22.2123
R21 VGND.n16 VGND.n3 10.5417
R22 VGND.n23 VGND.n0 9.3005
R23 VGND.n22 VGND.n21 9.3005
R24 VGND.n10 VGND.n9 9.3005
R25 VGND.n11 VGND.n5 9.3005
R26 VGND.n13 VGND.n12 9.3005
R27 VGND.n14 VGND.n3 9.3005
R28 VGND.n16 VGND.n15 9.3005
R29 VGND.n17 VGND.n2 9.3005
R30 VGND.n19 VGND.n18 9.3005
R31 VGND.n20 VGND.n1 9.3005
R32 VGND.n8 VGND.n6 7.13885
R33 VGND.n26 VGND.n25 7.12063
R34 VGND.n9 VGND.n8 0.49211
R35 VGND.n26 VGND.n0 0.148519
R36 VGND.n9 VGND.n5 0.120292
R37 VGND.n13 VGND.n5 0.120292
R38 VGND.n14 VGND.n13 0.120292
R39 VGND.n15 VGND.n14 0.120292
R40 VGND.n15 VGND.n2 0.120292
R41 VGND.n19 VGND.n2 0.120292
R42 VGND.n20 VGND.n19 0.120292
R43 VGND.n21 VGND.n20 0.120292
R44 VGND.n21 VGND.n0 0.120292
R45 VGND VGND.n26 0.114842
R46 Q Q.t0 134.917
R47 VNB.t4 VNB.t6 2691.26
R48 VNB.t7 VNB.t1 2677.02
R49 VNB.t2 VNB.t0 1694.5
R50 VNB.t1 VNB.t9 1594.82
R51 VNB.t10 VNB.t8 1509.39
R52 VNB.t0 VNB.t10 1438.19
R53 VNB.t11 VNB.t2 1409.71
R54 VNB.t9 VNB.t11 1409.71
R55 VNB.t8 VNB.t4 1352.75
R56 VNB.t6 VNB.t5 1196.12
R57 VNB.t3 VNB.t7 1196.12
R58 VNB VNB.t3 683.495
R59 a_193_47.n1 a_193_47.t5 407.217
R60 a_193_47.t1 a_193_47.n3 392.493
R61 a_193_47.n0 a_193_47.t4 308.651
R62 a_193_47.n0 a_193_47.t2 298.373
R63 a_193_47.n3 a_193_47.t0 294.144
R64 a_193_47.n1 a_193_47.t3 273.572
R65 a_193_47.n2 a_193_47.n1 170.9
R66 a_193_47.n2 a_193_47.n0 11.4492
R67 a_193_47.n3 a_193_47.n2 10.2617
R68 a_634_159.n3 a_634_159.n2 674.014
R69 a_634_159.n1 a_634_159.t5 406.401
R70 a_634_159.n2 a_634_159.n0 213.988
R71 a_634_159.n2 a_634_159.n1 180.161
R72 a_634_159.n1 a_634_159.t4 130.054
R73 a_634_159.n3 a_634_159.t2 89.1195
R74 a_634_159.n0 a_634_159.t3 71.6672
R75 a_634_159.t1 a_634_159.n3 37.5243
R76 a_634_159.n0 a_634_159.t0 28.438
R77 a_891_413.n4 a_891_413.n3 696.059
R78 a_891_413.n3 a_891_413.n0 258.788
R79 a_891_413.n3 a_891_413.n2 250.916
R80 a_891_413.n2 a_891_413.n1 212.081
R81 a_891_413.n2 a_891_413.t4 141.242
R82 a_891_413.n0 a_891_413.t1 76.6672
R83 a_891_413.n4 a_891_413.t3 63.3219
R84 a_891_413.t0 a_891_413.n4 63.3219
R85 a_891_413.n0 a_891_413.t2 50.0005
R86 a_27_47.n2 a_27_47.t5 443.44
R87 a_27_47.t1 a_27_47.n5 390.067
R88 a_27_47.n3 a_27_47.t7 345.305
R89 a_27_47.n3 a_27_47.t2 296.969
R90 a_27_47.n1 a_27_47.t0 287.998
R91 a_27_47.n0 a_27_47.t6 263.173
R92 a_27_47.n2 a_27_47.t4 254.389
R93 a_27_47.n0 a_27_47.t3 227.826
R94 a_27_47.n4 a_27_47.n2 193.59
R95 a_27_47.n1 a_27_47.n0 152
R96 a_27_47.n5 a_27_47.n1 35.3396
R97 a_27_47.n4 a_27_47.n3 12.4401
R98 a_27_47.n5 a_27_47.n4 11.0742
R99 a_466_413.n3 a_466_413.n2 695.683
R100 a_466_413.n2 a_466_413.n1 298.361
R101 a_466_413.n0 a_466_413.t4 230.484
R102 a_466_413.n0 a_466_413.t5 196.013
R103 a_466_413.n2 a_466_413.n0 168.738
R104 a_466_413.n3 a_466_413.t2 79.7386
R105 a_466_413.t0 a_466_413.n3 72.7029
R106 a_466_413.n1 a_466_413.t3 70.0005
R107 a_466_413.n1 a_466_413.t1 45.0005
R108 a_561_413.t0 a_561_413.t1 171.202
R109 VPB.t4 VPB.t1 556.386
R110 VPB.t0 VPB.t2 390.654
R111 VPB.t8 VPB.t3 337.384
R112 VPB.t6 VPB.t0 304.829
R113 VPB.t2 VPB.t5 281.154
R114 VPB.t9 VPB.t6 281.154
R115 VPB.t1 VPB.t9 251.559
R116 VPB.t5 VPB.t8 248.599
R117 VPB.t7 VPB.t4 248.599
R118 VPB VPB.t7 142.056
R119 CLK.n0 CLK.t0 294.557
R120 CLK.n0 CLK.t1 211.01
R121 CLK CLK.n0 153.97
R122 VPWR.n6 VPWR.t4 673.736
R123 VPWR.n14 VPWR.t1 666.677
R124 VPWR.n16 VPWR.n1 604.394
R125 VPWR.n7 VPWR.n5 320.976
R126 VPWR.n5 VPWR.t0 113.98
R127 VPWR.n1 VPWR.t5 41.5552
R128 VPWR.n1 VPWR.t3 41.5552
R129 VPWR.n5 VPWR.t2 35.4605
R130 VPWR.n9 VPWR.n8 34.6358
R131 VPWR.n9 VPWR.n3 34.6358
R132 VPWR.n13 VPWR.n3 34.6358
R133 VPWR.n14 VPWR.n13 27.4829
R134 VPWR.n7 VPWR.n6 23.7763
R135 VPWR.n16 VPWR.n15 22.9652
R136 VPWR.n15 VPWR.n14 21.8358
R137 VPWR.n8 VPWR.n7 18.4476
R138 VPWR.n8 VPWR.n4 9.3005
R139 VPWR.n10 VPWR.n9 9.3005
R140 VPWR.n11 VPWR.n3 9.3005
R141 VPWR.n13 VPWR.n12 9.3005
R142 VPWR.n14 VPWR.n2 9.3005
R143 VPWR.n15 VPWR.n0 9.3005
R144 VPWR.n17 VPWR.n16 7.12063
R145 VPWR.n6 VPWR.n4 0.16021
R146 VPWR.n17 VPWR.n0 0.148519
R147 VPWR.n10 VPWR.n4 0.120292
R148 VPWR.n11 VPWR.n10 0.120292
R149 VPWR.n12 VPWR.n11 0.120292
R150 VPWR.n12 VPWR.n2 0.120292
R151 VPWR.n2 VPWR.n0 0.120292
R152 VPWR VPWR.n17 0.114842
R153 D.n0 D.t1 302.731
R154 D.n0 D.t0 212.757
R155 D D.n0 170.058
R156 a_381_47.n1 a_381_47.n0 896.306
R157 a_381_47.n0 a_381_47.t0 90.0005
R158 a_381_47.t1 a_381_47.n1 65.6672
R159 a_381_47.n1 a_381_47.t2 63.3219
R160 a_381_47.n0 a_381_47.t3 31.3935
R161 a_592_47.t0 a_592_47.t1 99.7268
R162 a_975_413.t0 a_975_413.t1 197
R163 a_1017_47.t0 a_1017_47.t1 93.0601
C0 CLK VGND 0.019463f
C1 D VPWR 0.025067f
C2 VPB Q 0.013828f
C3 D VGND 0.038993f
C4 a_1059_315# VPB 0.154738f
C5 VPWR VGND 0.063886f
C6 VPWR Q 0.110929f
C7 VGND Q 0.076612f
C8 a_1059_315# VPWR 0.232446f
C9 a_1059_315# VGND 0.155119f
C10 a_1059_315# Q 0.081249f
C11 VPB CLK 0.070057f
C12 VPB D 0.096334f
C13 VPB VPWR 0.168181f
C14 VPB VGND 0.012227f
C15 CLK VPWR 0.019411f
C16 Q VNB 0.088256f
C17 VGND VNB 0.84362f
C18 VPWR VNB 0.681368f
C19 D VNB 0.142509f
C20 CLK VNB 0.195983f
C21 VPB VNB 1.49072f
C22 a_1059_315# VNB 0.248849f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q.t1 a_1059_315# VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_891_413.t0 a_193_47.t2 a_634_159.t2 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3 a_561_413.t1 a_27_47.t2 a_466_413.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4 VPWR.t4 CLK.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47.t3 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND.t1 a_634_159.t4 a_592_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND.t5 a_1059_315# Q.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_466_413.t2 a_193_47.t3 a_381_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10 VPWR.t2 a_634_159.t5 a_561_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11 a_634_159.t0 a_466_413.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12 a_634_159.t1 a_466_413.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13 a_975_413.t0 a_193_47.t4 a_891_413.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VGND.t4 a_1059_315# a_1017_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15 a_193_47.t1 a_27_47.t3 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_891_413.t2 a_27_47.t4 a_634_159.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X17 a_592_47.t1 a_193_47.t5 a_466_413.t3 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X18 VPWR.t5 a_1059_315# a_975_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_1017_47.t0 a_27_47.t5 a_891_413.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 a_193_47.t0 a_27_47.t6 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 a_466_413.t1 a_27_47.t7 a_381_47.t0 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 VGND.t3 a_891_413.t4 a_1059_315# VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_381_47.t2 D.t1 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VGND.t2 CLK.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 VGND.n6 VGND.t4 251
R1 VGND.n7 VGND.t5 247.452
R2 VGND.n26 VGND.t8 243.028
R3 VGND.n9 VGND.n8 218.506
R4 VGND.n29 VGND.n28 199.739
R5 VGND.n20 VGND.n4 199.53
R6 VGND.n4 VGND.t0 74.8666
R7 VGND.n4 VGND.t1 40.0005
R8 VGND.n28 VGND.t7 38.5719
R9 VGND.n28 VGND.t2 38.5719
R10 VGND.n15 VGND.n14 34.6358
R11 VGND.n16 VGND.n15 34.6358
R12 VGND.n16 VGND.n3 34.6358
R13 VGND.n22 VGND.n21 34.6358
R14 VGND.n22 VGND.n1 34.6358
R15 VGND.n10 VGND.n9 32.377
R16 VGND.n10 VGND.n6 31.2476
R17 VGND.n21 VGND.n20 30.8711
R18 VGND.n26 VGND.n1 27.4829
R19 VGND.n8 VGND.t6 24.9236
R20 VGND.n8 VGND.t3 24.9236
R21 VGND.n27 VGND.n26 22.9652
R22 VGND.n29 VGND.n27 22.9652
R23 VGND.n14 VGND.n6 22.2123
R24 VGND.n20 VGND.n3 10.5417
R25 VGND.n9 VGND.n7 9.31175
R26 VGND.n27 VGND.n0 9.3005
R27 VGND.n26 VGND.n25 9.3005
R28 VGND.n11 VGND.n10 9.3005
R29 VGND.n12 VGND.n6 9.3005
R30 VGND.n14 VGND.n13 9.3005
R31 VGND.n15 VGND.n5 9.3005
R32 VGND.n17 VGND.n16 9.3005
R33 VGND.n18 VGND.n3 9.3005
R34 VGND.n20 VGND.n19 9.3005
R35 VGND.n21 VGND.n2 9.3005
R36 VGND.n23 VGND.n22 9.3005
R37 VGND.n24 VGND.n1 9.3005
R38 VGND.n30 VGND.n29 7.12063
R39 VGND.n11 VGND.n7 0.697081
R40 VGND.n30 VGND.n0 0.148519
R41 VGND.n12 VGND.n11 0.120292
R42 VGND.n13 VGND.n12 0.120292
R43 VGND.n13 VGND.n5 0.120292
R44 VGND.n17 VGND.n5 0.120292
R45 VGND.n18 VGND.n17 0.120292
R46 VGND.n19 VGND.n18 0.120292
R47 VGND.n19 VGND.n2 0.120292
R48 VGND.n23 VGND.n2 0.120292
R49 VGND.n24 VGND.n23 0.120292
R50 VGND.n25 VGND.n24 0.120292
R51 VGND.n25 VGND.n0 0.120292
R52 VGND VGND.n30 0.114842
R53 Q Q.n0 95.7215
R54 Q.n0 Q.t0 24.9236
R55 Q.n0 Q.t1 24.9236
R56 VNB.t7 VNB.t4 2691.26
R57 VNB.t10 VNB.t12 2677.02
R58 VNB.t1 VNB.t0 1694.5
R59 VNB.t12 VNB.t2 1594.82
R60 VNB.t5 VNB.t11 1509.39
R61 VNB.t0 VNB.t5 1438.19
R62 VNB.t6 VNB.t1 1409.71
R63 VNB.t2 VNB.t6 1409.71
R64 VNB.t11 VNB.t7 1352.75
R65 VNB.t9 VNB.t8 1196.12
R66 VNB.t4 VNB.t9 1196.12
R67 VNB.t3 VNB.t10 1196.12
R68 VNB VNB.t3 683.495
R69 VPWR.n6 VPWR.t5 673.736
R70 VPWR.n14 VPWR.t0 666.677
R71 VPWR.n16 VPWR.n1 604.394
R72 VPWR.n7 VPWR.n5 320.976
R73 VPWR.n5 VPWR.t2 113.98
R74 VPWR.n1 VPWR.t3 41.5552
R75 VPWR.n1 VPWR.t4 41.5552
R76 VPWR.n5 VPWR.t1 35.4605
R77 VPWR.n9 VPWR.n8 34.6358
R78 VPWR.n9 VPWR.n3 34.6358
R79 VPWR.n13 VPWR.n3 34.6358
R80 VPWR.n14 VPWR.n13 27.4829
R81 VPWR.n7 VPWR.n6 23.7763
R82 VPWR.n16 VPWR.n15 22.9652
R83 VPWR.n15 VPWR.n14 21.8358
R84 VPWR.n8 VPWR.n7 18.4476
R85 VPWR.n8 VPWR.n4 9.3005
R86 VPWR.n10 VPWR.n9 9.3005
R87 VPWR.n11 VPWR.n3 9.3005
R88 VPWR.n13 VPWR.n12 9.3005
R89 VPWR.n14 VPWR.n2 9.3005
R90 VPWR.n15 VPWR.n0 9.3005
R91 VPWR.n17 VPWR.n16 7.12063
R92 VPWR.n6 VPWR.n4 0.16021
R93 VPWR.n17 VPWR.n0 0.148519
R94 VPWR.n10 VPWR.n4 0.120292
R95 VPWR.n11 VPWR.n10 0.120292
R96 VPWR.n12 VPWR.n11 0.120292
R97 VPWR.n12 VPWR.n2 0.120292
R98 VPWR.n2 VPWR.n0 0.120292
R99 VPWR VPWR.n17 0.114842
R100 VPB.t3 VPB.t0 556.386
R101 VPB.t2 VPB.t1 390.654
R102 VPB.t6 VPB.t7 337.384
R103 VPB.t8 VPB.t2 304.829
R104 VPB.t1 VPB.t9 281.154
R105 VPB.t5 VPB.t8 281.154
R106 VPB.t0 VPB.t5 251.559
R107 VPB.t9 VPB.t6 248.599
R108 VPB.t4 VPB.t3 248.599
R109 VPB VPB.t4 142.056
R110 a_193_47.n1 a_193_47.t5 407.217
R111 a_193_47.t0 a_193_47.n3 392.493
R112 a_193_47.n0 a_193_47.t4 308.651
R113 a_193_47.n0 a_193_47.t2 298.373
R114 a_193_47.n3 a_193_47.t1 294.144
R115 a_193_47.n1 a_193_47.t3 273.572
R116 a_193_47.n2 a_193_47.n1 170.9
R117 a_193_47.n2 a_193_47.n0 11.4492
R118 a_193_47.n3 a_193_47.n2 10.2617
R119 a_634_159.n3 a_634_159.n2 674.014
R120 a_634_159.n1 a_634_159.t5 406.401
R121 a_634_159.n2 a_634_159.n0 213.988
R122 a_634_159.n2 a_634_159.n1 180.161
R123 a_634_159.n1 a_634_159.t4 130.054
R124 a_634_159.n3 a_634_159.t3 89.1195
R125 a_634_159.n0 a_634_159.t2 71.6672
R126 a_634_159.t1 a_634_159.n3 37.5243
R127 a_634_159.n0 a_634_159.t0 28.438
R128 a_891_413.n4 a_891_413.n3 696.059
R129 a_891_413.n3 a_891_413.n0 258.788
R130 a_891_413.n3 a_891_413.n2 250.916
R131 a_891_413.n2 a_891_413.n1 212.081
R132 a_891_413.n2 a_891_413.t4 141.242
R133 a_891_413.n0 a_891_413.t3 76.6672
R134 a_891_413.t1 a_891_413.n4 63.3219
R135 a_891_413.n4 a_891_413.t2 63.3219
R136 a_891_413.n0 a_891_413.t0 50.0005
R137 a_27_47.n2 a_27_47.t5 443.44
R138 a_27_47.t1 a_27_47.n5 390.067
R139 a_27_47.n3 a_27_47.t7 345.305
R140 a_27_47.n3 a_27_47.t2 296.969
R141 a_27_47.n1 a_27_47.t0 287.998
R142 a_27_47.n0 a_27_47.t6 263.173
R143 a_27_47.n2 a_27_47.t4 254.389
R144 a_27_47.n0 a_27_47.t3 227.826
R145 a_27_47.n4 a_27_47.n2 193.59
R146 a_27_47.n1 a_27_47.n0 152
R147 a_27_47.n5 a_27_47.n1 35.3396
R148 a_27_47.n4 a_27_47.n3 12.4401
R149 a_27_47.n5 a_27_47.n4 11.0742
R150 a_466_413.n3 a_466_413.n2 695.683
R151 a_466_413.n2 a_466_413.n1 298.361
R152 a_466_413.n0 a_466_413.t4 230.484
R153 a_466_413.n0 a_466_413.t5 196.013
R154 a_466_413.n2 a_466_413.n0 168.738
R155 a_466_413.n3 a_466_413.t2 79.7386
R156 a_466_413.t0 a_466_413.n3 72.7029
R157 a_466_413.n1 a_466_413.t3 70.0005
R158 a_466_413.n1 a_466_413.t1 45.0005
R159 a_561_413.t0 a_561_413.t1 171.202
R160 CLK.n0 CLK.t0 294.557
R161 CLK.n0 CLK.t1 211.01
R162 CLK CLK.n0 153.97
R163 D.n0 D.t1 302.731
R164 D.n0 D.t0 212.757
R165 D D.n0 170.058
R166 a_381_47.n1 a_381_47.n0 896.306
R167 a_381_47.n0 a_381_47.t0 90.0005
R168 a_381_47.t1 a_381_47.n1 65.6672
R169 a_381_47.n1 a_381_47.t3 63.3219
R170 a_381_47.n0 a_381_47.t2 31.3935
R171 a_592_47.t0 a_592_47.t1 99.7268
R172 a_975_413.t0 a_975_413.t1 197
R173 a_1017_47.t1 a_1017_47.t0 93.0601
C0 CLK VPWR 0.019411f
C1 VPB VGND 0.014667f
C2 VPB Q 0.007287f
C3 CLK VGND 0.019463f
C4 D VPWR 0.025067f
C5 a_1059_315# VPWR 0.250757f
C6 D VGND 0.038993f
C7 a_1059_315# VGND 0.171637f
C8 VPWR VGND 0.082807f
C9 a_1059_315# Q 0.121751f
C10 VPWR Q 0.171866f
C11 VGND Q 0.10404f
C12 VPB CLK 0.070057f
C13 VPB D 0.096334f
C14 a_1059_315# VPB 0.184378f
C15 VPB VPWR 0.181734f
C16 Q VNB 0.040388f
C17 VGND VNB 0.908998f
C18 VPWR VNB 0.751085f
C19 D VNB 0.142509f
C20 CLK VNB 0.195983f
C21 VPB VNB 1.57932f
C22 a_1059_315# VNB 0.332253f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR VNB VPB Q D CLK
X0 Q.t1 a_1062_300.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_1020_47# a_27_47.t2 a_891_413.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47.t1 a_193_47.t2 a_475_413.t1 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR.t2 a_1062_300.t3 a_975_413.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X4 a_634_183.t0 a_475_413.t4 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X5 VPWR.t8 CLK.t0 a_27_47.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_381_47.t1 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_475_413.t3 a_27_47.t3 a_381_47.t3 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VPWR.t1 a_634_183.t4 a_568_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 Q.t3 a_1062_300.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X10 a_568_413.t1 a_27_47.t4 a_475_413.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X11 a_634_183.t1 a_475_413.t5 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413.t1 a_193_47.t3 a_891_413.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_193_47.t1 a_27_47.t5 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_891_413.t2 a_27_47.t6 a_634_183.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15 VGND.t6 a_891_413.t4 a_1062_300.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VGND.t2 a_1062_300.t5 Q.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_193_47.t0 a_27_47.t7 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X18 a_381_47.t0 D.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 VPWR.t7 a_891_413.t5 a_1062_300.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X20 a_475_413.t0 a_193_47.t4 a_381_47.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X21 a_891_413.t1 a_193_47.t5 a_634_183.t2 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X22 VGND.t1 a_634_183.t5 a_572_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X23 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VPWR.t3 a_1062_300.t6 Q.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
R0 a_1062_300.n17 a_1062_300.n16 359.399
R1 a_1062_300.t1 a_1062_300.n18 228.28
R2 a_1062_300.n4 a_1062_300.t6 212.081
R3 a_1062_300.n3 a_1062_300.t2 212.081
R4 a_1062_300.n9 a_1062_300.n1 212.081
R5 a_1062_300.n12 a_1062_300.n10 212.081
R6 a_1062_300.n18 a_1062_300.n17 178.764
R7 a_1062_300.n6 a_1062_300.n5 177.601
R8 a_1062_300.n15 a_1062_300.t0 165.512
R9 a_1062_300.n17 a_1062_300.t3 163.387
R10 a_1062_300.n14 a_1062_300.n13 152
R11 a_1062_300.n8 a_1062_300.n0 152
R12 a_1062_300.n7 a_1062_300.n6 152
R13 a_1062_300.n4 a_1062_300.t5 139.78
R14 a_1062_300.n3 a_1062_300.t4 139.78
R15 a_1062_300.n9 a_1062_300.n2 139.78
R16 a_1062_300.n12 a_1062_300.n11 139.78
R17 a_1062_300.n8 a_1062_300.n7 49.6611
R18 a_1062_300.n13 a_1062_300.n9 44.549
R19 a_1062_300.n15 a_1062_300.n14 41.4123
R20 a_1062_300.n5 a_1062_300.n3 40.8975
R21 a_1062_300.n18 a_1062_300.n15 34.921
R22 a_1062_300.n6 a_1062_300.n0 25.6005
R23 a_1062_300.n14 a_1062_300.n0 25.6005
R24 a_1062_300.n5 a_1062_300.n4 20.449
R25 a_1062_300.n13 a_1062_300.n12 16.7975
R26 a_1062_300.n7 a_1062_300.n3 8.76414
R27 a_1062_300.n9 a_1062_300.n8 5.11262
R28 VPWR.n18 VPWR.t2 673.327
R29 VPWR.n32 VPWR.t0 666.677
R30 VPWR.n34 VPWR.n1 604.394
R31 VPWR.n10 VPWR.t3 360.404
R32 VPWR.n13 VPWR.t7 357.514
R33 VPWR.n11 VPWR.t4 349.83
R34 VPWR.n25 VPWR.n5 320.976
R35 VPWR.n5 VPWR.t1 113.98
R36 VPWR.n1 VPWR.t5 41.5552
R37 VPWR.n1 VPWR.t8 41.5552
R38 VPWR.n5 VPWR.t6 35.4605
R39 VPWR.n20 VPWR.n19 34.6358
R40 VPWR.n20 VPWR.n6 34.6358
R41 VPWR.n24 VPWR.n6 34.6358
R42 VPWR.n27 VPWR.n26 34.6358
R43 VPWR.n27 VPWR.n3 34.6358
R44 VPWR.n31 VPWR.n3 34.6358
R45 VPWR.n17 VPWR.n8 34.6358
R46 VPWR.n12 VPWR.n11 34.2593
R47 VPWR.n13 VPWR.n8 31.2476
R48 VPWR.n32 VPWR.n31 27.4829
R49 VPWR.n13 VPWR.n12 24.4711
R50 VPWR.n34 VPWR.n33 22.9652
R51 VPWR.n33 VPWR.n32 21.8358
R52 VPWR.n26 VPWR.n25 18.4476
R53 VPWR.n25 VPWR.n24 16.1887
R54 VPWR.n19 VPWR.n18 15.0593
R55 VPWR.n12 VPWR.n9 9.3005
R56 VPWR.n14 VPWR.n13 9.3005
R57 VPWR.n15 VPWR.n8 9.3005
R58 VPWR.n17 VPWR.n16 9.3005
R59 VPWR.n19 VPWR.n7 9.3005
R60 VPWR.n21 VPWR.n20 9.3005
R61 VPWR.n22 VPWR.n6 9.3005
R62 VPWR.n24 VPWR.n23 9.3005
R63 VPWR.n26 VPWR.n4 9.3005
R64 VPWR.n28 VPWR.n27 9.3005
R65 VPWR.n29 VPWR.n3 9.3005
R66 VPWR.n31 VPWR.n30 9.3005
R67 VPWR.n32 VPWR.n2 9.3005
R68 VPWR.n33 VPWR.n0 9.3005
R69 VPWR.n11 VPWR.n10 7.48837
R70 VPWR.n35 VPWR.n34 7.12063
R71 VPWR.n18 VPWR.n17 3.38874
R72 VPWR.n10 VPWR.n9 0.638101
R73 VPWR.n35 VPWR.n0 0.148519
R74 VPWR.n14 VPWR.n9 0.120292
R75 VPWR.n15 VPWR.n14 0.120292
R76 VPWR.n16 VPWR.n15 0.120292
R77 VPWR.n16 VPWR.n7 0.120292
R78 VPWR.n21 VPWR.n7 0.120292
R79 VPWR.n22 VPWR.n21 0.120292
R80 VPWR.n23 VPWR.n22 0.120292
R81 VPWR.n23 VPWR.n4 0.120292
R82 VPWR.n28 VPWR.n4 0.120292
R83 VPWR.n29 VPWR.n28 0.120292
R84 VPWR.n30 VPWR.n29 0.120292
R85 VPWR.n30 VPWR.n2 0.120292
R86 VPWR.n2 VPWR.n0 0.120292
R87 VPWR VPWR.n35 0.114842
R88 Q.n5 Q.n4 1176.51
R89 Q.n3 Q.n2 205.28
R90 Q.n1 Q.n0 98.6958
R91 Q.n3 Q.n1 74.1652
R92 Q.n1 Q 53.7923
R93 Q.n4 Q.n3 42.2102
R94 Q.n2 Q.t0 26.5955
R95 Q.n2 Q.t1 26.5955
R96 Q.n0 Q.t2 24.9236
R97 Q.n0 Q.t3 24.9236
R98 Q.n5 Q 9.49065
R99 Q.n4 Q 5.92289
R100 Q Q.n5 3.47789
R101 VPB.t9 VPB.t4 787.227
R102 VPB.t3 VPB.t9 639.253
R103 VPB.t7 VPB.t0 556.386
R104 VPB.t1 VPB.t8 390.654
R105 VPB.t11 VPB.t3 346.262
R106 VPB.t5 VPB.t1 284.113
R107 VPB.t8 VPB.t6 281.154
R108 VPB.t0 VPB.t12 278.193
R109 VPB.t12 VPB.t5 275.235
R110 VPB.t4 VPB.t2 248.599
R111 VPB.t6 VPB.t11 248.599
R112 VPB.t10 VPB.t7 248.599
R113 VPB VPB.t10 142.056
R114 a_27_47.n3 a_27_47.t3 501.817
R115 a_27_47.n2 a_27_47.t2 448.26
R116 a_27_47.t1 a_27_47.n5 390.067
R117 a_27_47.n1 a_27_47.t0 287.998
R118 a_27_47.n0 a_27_47.t7 263.173
R119 a_27_47.n2 a_27_47.t6 254.389
R120 a_27_47.n0 a_27_47.t5 227.826
R121 a_27_47.n4 a_27_47.n2 193.421
R122 a_27_47.n4 a_27_47.n3 168.151
R123 a_27_47.n1 a_27_47.n0 152
R124 a_27_47.n3 a_27_47.t4 148.35
R125 a_27_47.n5 a_27_47.n1 35.3396
R126 a_27_47.n5 a_27_47.n4 11.2706
R127 a_891_413.n3 a_891_413.n2 702.082
R128 a_891_413.n2 a_891_413.n1 273.671
R129 a_891_413.n2 a_891_413.n0 257.283
R130 a_891_413.n1 a_891_413.t5 212.081
R131 a_891_413.n1 a_891_413.t4 139.78
R132 a_891_413.n0 a_891_413.t1 73.3338
R133 a_891_413.t0 a_891_413.n3 63.3219
R134 a_891_413.n3 a_891_413.t2 63.3219
R135 a_891_413.n0 a_891_413.t3 48.3338
R136 VNB.t11 VNB.t5 4100.97
R137 VNB.t5 VNB.t3 3787.7
R138 VNB.t9 VNB.t4 2677.02
R139 VNB.t1 VNB.t6 2078.96
R140 VNB.t8 VNB.t11 1466.67
R141 VNB.t6 VNB.t8 1438.19
R142 VNB.t7 VNB.t1 1395.47
R143 VNB.t10 VNB.t7 1366.99
R144 VNB.t4 VNB.t10 1352.75
R145 VNB.t3 VNB.t2 1196.12
R146 VNB.t0 VNB.t9 1196.12
R147 VNB VNB.t0 683.495
R148 a_193_47.t0 a_193_47.n3 424.863
R149 a_193_47.n0 a_193_47.t3 348.661
R150 a_193_47.n1 a_193_47.t4 345.803
R151 a_193_47.n1 a_193_47.t2 281.236
R152 a_193_47.n0 a_193_47.t5 271.262
R153 a_193_47.n3 a_193_47.t1 242.915
R154 a_193_47.n2 a_193_47.n0 18.9875
R155 a_193_47.n3 a_193_47.n2 10.4492
R156 a_193_47.n2 a_193_47.n1 9.3005
R157 a_475_413.n3 a_475_413.n2 693.048
R158 a_475_413.n2 a_475_413.n1 300.997
R159 a_475_413.n0 a_475_413.t4 226.541
R160 a_475_413.n0 a_475_413.t5 196.013
R161 a_475_413.n2 a_475_413.n0 168.738
R162 a_475_413.t0 a_475_413.n3 75.0481
R163 a_475_413.n3 a_475_413.t2 72.7029
R164 a_475_413.n1 a_475_413.t3 61.6672
R165 a_475_413.n1 a_475_413.t1 48.3338
R166 a_572_47.t0 a_572_47.t1 98.0601
R167 a_975_413.t0 a_975_413.t1 204.036
R168 VGND.n9 VGND.t2 288.252
R169 VGND.n8 VGND.t3 277.815
R170 VGND.n30 VGND.t4 243.028
R171 VGND.n12 VGND.t6 240.102
R172 VGND.n33 VGND.n32 199.739
R173 VGND.n24 VGND.n4 199.53
R174 VGND.n4 VGND.t1 87.1434
R175 VGND.n4 VGND.t5 66.2951
R176 VGND.n32 VGND.t7 38.5719
R177 VGND.n32 VGND.t0 38.5719
R178 VGND.n14 VGND.n13 34.6358
R179 VGND.n14 VGND.n6 34.6358
R180 VGND.n18 VGND.n6 34.6358
R181 VGND.n19 VGND.n18 34.6358
R182 VGND.n20 VGND.n19 34.6358
R183 VGND.n20 VGND.n3 34.6358
R184 VGND.n26 VGND.n25 34.6358
R185 VGND.n26 VGND.n1 34.6358
R186 VGND.n11 VGND.n8 33.8829
R187 VGND.n12 VGND.n11 31.624
R188 VGND.n25 VGND.n24 30.8711
R189 VGND.n30 VGND.n1 27.4829
R190 VGND.n31 VGND.n30 22.9652
R191 VGND.n33 VGND.n31 22.9652
R192 VGND.n24 VGND.n3 10.5417
R193 VGND.n31 VGND.n0 9.3005
R194 VGND.n30 VGND.n29 9.3005
R195 VGND.n11 VGND.n10 9.3005
R196 VGND.n13 VGND.n7 9.3005
R197 VGND.n15 VGND.n14 9.3005
R198 VGND.n16 VGND.n6 9.3005
R199 VGND.n18 VGND.n17 9.3005
R200 VGND.n19 VGND.n5 9.3005
R201 VGND.n21 VGND.n20 9.3005
R202 VGND.n22 VGND.n3 9.3005
R203 VGND.n24 VGND.n23 9.3005
R204 VGND.n25 VGND.n2 9.3005
R205 VGND.n27 VGND.n26 9.3005
R206 VGND.n28 VGND.n1 9.3005
R207 VGND.n9 VGND.n8 7.87664
R208 VGND.n34 VGND.n33 7.12063
R209 VGND.n13 VGND.n12 3.01226
R210 VGND.n10 VGND.n9 0.626305
R211 VGND.n34 VGND.n0 0.148519
R212 VGND.n10 VGND.n7 0.120292
R213 VGND.n15 VGND.n7 0.120292
R214 VGND.n16 VGND.n15 0.120292
R215 VGND.n17 VGND.n16 0.120292
R216 VGND.n17 VGND.n5 0.120292
R217 VGND.n21 VGND.n5 0.120292
R218 VGND.n22 VGND.n21 0.120292
R219 VGND.n23 VGND.n22 0.120292
R220 VGND.n23 VGND.n2 0.120292
R221 VGND.n27 VGND.n2 0.120292
R222 VGND.n28 VGND.n27 0.120292
R223 VGND.n29 VGND.n28 0.120292
R224 VGND.n29 VGND.n0 0.120292
R225 VGND VGND.n34 0.114842
R226 a_634_183.n3 a_634_183.n2 674.014
R227 a_634_183.n1 a_634_183.t4 433.8
R228 a_634_183.n2 a_634_183.n0 218.13
R229 a_634_183.n2 a_634_183.n1 185.308
R230 a_634_183.n1 a_634_183.t5 128.1
R231 a_634_183.n3 a_634_183.t3 89.1195
R232 a_634_183.n0 a_634_183.t2 63.3338
R233 a_634_183.t1 a_634_183.n3 37.5243
R234 a_634_183.n0 a_634_183.t0 36.7713
R235 CLK.n0 CLK.t0 294.557
R236 CLK.n0 CLK.t1 211.01
R237 CLK.n1 CLK.n0 152
R238 CLK.n1 CLK 10.4234
R239 CLK CLK.n1 2.01193
R240 D.n0 D.t1 305.625
R241 D.n0 D.t0 215.65
R242 D D.n0 154.514
R243 a_381_47.n1 a_381_47.n0 899.936
R244 a_381_47.n0 a_381_47.t2 86.7743
R245 a_381_47.n0 a_381_47.t1 63.3219
R246 a_381_47.n1 a_381_47.t3 58.3338
R247 a_381_47.n2 a_381_47.t0 26.3935
R248 a_381_47.n3 a_381_47.n2 14.4005
R249 a_381_47.n2 a_381_47.n1 8.33383
R250 a_568_413.t0 a_568_413.t1 154.786
C0 D VGND 0.026396f
C1 VPWR VGND 0.100633f
C2 VPWR Q 0.335782f
C3 VGND Q 0.242058f
C4 a_1020_47# VPWR 4.79e-19
C5 VPB CLK 0.070057f
C6 a_1020_47# VGND 0.004151f
C7 VPB D 0.09609f
C8 VPB VPWR 0.198564f
C9 CLK VPWR 0.019411f
C10 VPB VGND 0.014659f
C11 D VPWR 0.027256f
C12 CLK VGND 0.019463f
C13 VPB Q 0.013356f
C14 Q VNB 0.060797f
C15 VGND VNB 0.988933f
C16 VPWR VNB 0.823111f
C17 D VNB 0.129726f
C18 CLK VNB 0.195983f
C19 VPB VNB 1.75651f
.ends

* NGSPICE file created from sky130_fd_sc_hd__diode_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
X0 VNB.t0 DIODE.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
R0 DIODE.n0 DIODE.t0 45.2995
R1 DIODE DIODE.n0 3.29771
R2 DIODE.n0 DIODE 2.38297
R3 VNB VNB.t0 2115.38
C0 VPWR VPB 0.02381f
C1 VGND VPB 0.003161f
C2 VPWR DIODE 0.105447f
C3 VGND DIODE 0.107068f
C4 VPB DIODE 0.046677f
C5 VGND VPWR 0.017949f
C6 VGND VNB 0.147223f
C7 VPWR VNB 0.127718f
C8 DIODE VNB 0.183985f
C9 VPB VNB 0.25038f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlclkp_1 VGND VPWR GCLK GATE CLK VPB VNB
X0 a_381_369.t0 GATE.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_476_413.t3 a_193_47.t2 a_381_369.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.09575 ps=0.965 w=0.42 l=0.15
X2 a_957_369.t1 a_642_307.t2 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2032 pd=1.275 as=0.149 ps=1.325 w=0.64 l=0.15
X3 VPWR.t7 CLK.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_1042_47.t1 a_642_307.t3 a_957_369.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 GCLK.t1 a_957_369.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X6 VGND.t2 CLK.t1 a_1042_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_193_47.t1 a_27_47.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_651_47.t1 a_193_47.t3 a_476_413.t2 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.067125 pd=0.745 as=0.1192 ps=1.09 w=0.39 l=0.15
X9 a_193_47.t0 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 GCLK.t0 a_957_369.t4 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11 VPWR.t5 a_642_307.t4 a_600_413.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 a_476_413.t0 a_27_47.t4 a_396_119.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1192 pd=1.09 as=0.117125 ps=1.085 w=0.42 l=0.15
X13 VPWR.t6 CLK.t2 a_957_369.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.2032 ps=1.275 w=0.64 l=0.15
X14 a_642_307.t0 a_476_413.t4 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.118125 ps=1.04 w=0.65 l=0.15
X15 a_600_413.t0 a_27_47.t5 a_476_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0987 ps=0.89 w=0.42 l=0.15
X16 VPWR.t2 a_476_413.t5 a_642_307.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.27 ps=2.54 w=1 l=0.15
X17 VGND.t3 a_642_307.t5 a_651_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.067125 ps=0.745 w=0.42 l=0.15
X18 VGND.t1 CLK.t3 a_27_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 a_396_119.t1 GATE.t1 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.117125 pd=1.085 as=0.1281 ps=1.45 w=0.42 l=0.15
R0 GATE.n0 GATE.t1 189.588
R1 GATE.n0 GATE.t0 183.161
R2 GATE GATE.n0 164.288
R3 VPWR.n17 VPWR.t3 730.923
R4 VPWR.n11 VPWR.t5 666.241
R5 VPWR.n8 VPWR.n7 606.458
R6 VPWR.n6 VPWR.n5 605.212
R7 VPWR.n19 VPWR.n1 604.394
R8 VPWR.n7 VPWR.t6 58.4849
R9 VPWR.n5 VPWR.t4 53.8677
R10 VPWR.n1 VPWR.t0 41.5552
R11 VPWR.n1 VPWR.t7 41.5552
R12 VPWR.n5 VPWR.t2 36.2229
R13 VPWR.n12 VPWR.n3 34.6358
R14 VPWR.n16 VPWR.n3 34.6358
R15 VPWR.n7 VPWR.t1 31.6057
R16 VPWR.n12 VPWR.n11 30.4946
R17 VPWR.n10 VPWR.n6 30.1181
R18 VPWR.n19 VPWR.n18 22.9652
R19 VPWR.n18 VPWR.n17 22.5887
R20 VPWR.n17 VPWR.n16 19.2005
R21 VPWR.n11 VPWR.n10 16.1887
R22 VPWR.n10 VPWR.n9 9.3005
R23 VPWR.n11 VPWR.n4 9.3005
R24 VPWR.n13 VPWR.n12 9.3005
R25 VPWR.n14 VPWR.n3 9.3005
R26 VPWR.n16 VPWR.n15 9.3005
R27 VPWR.n17 VPWR.n2 9.3005
R28 VPWR.n18 VPWR.n0 9.3005
R29 VPWR.n20 VPWR.n19 7.12063
R30 VPWR.n8 VPWR.n6 6.68414
R31 VPWR.n9 VPWR.n8 0.246649
R32 VPWR.n20 VPWR.n0 0.148519
R33 VPWR.n9 VPWR.n4 0.120292
R34 VPWR.n13 VPWR.n4 0.120292
R35 VPWR.n14 VPWR.n13 0.120292
R36 VPWR.n15 VPWR.n14 0.120292
R37 VPWR.n15 VPWR.n2 0.120292
R38 VPWR.n2 VPWR.n0 0.120292
R39 VPWR VPWR.n20 0.11354
R40 a_381_369.t0 a_381_369.t1 132.286
R41 VPB.t0 VPB.t4 574.277
R42 VPB.t6 VPB.t3 562.306
R43 VPB.t5 VPB.t7 464.642
R44 VPB.t8 VPB.t1 372.974
R45 VPB.t4 VPB.t8 290.193
R46 VPB.t7 VPB.t2 281.154
R47 VPB.t3 VPB.t5 281.154
R48 VPB.t9 VPB.t0 256.592
R49 VPB.t1 VPB.t6 213.084
R50 VPB VPB.t9 198.554
R51 a_193_47.n0 a_193_47.t3 366.247
R52 a_193_47.t0 a_193_47.n1 362.546
R53 a_193_47.n0 a_193_47.t2 310.882
R54 a_193_47.n1 a_193_47.t1 296.75
R55 a_193_47.n1 a_193_47.n0 96.377
R56 a_476_413.n2 a_476_413.n1 727.216
R57 a_476_413.n3 a_476_413.n2 273.046
R58 a_476_413.n0 a_476_413.t5 234.483
R59 a_476_413.n2 a_476_413.n0 169.456
R60 a_476_413.n0 a_476_413.t4 162.184
R61 a_476_413.n1 a_476_413.t3 121.953
R62 a_476_413.n4 a_476_413.n3 117.081
R63 a_476_413.n1 a_476_413.t1 98.5005
R64 a_476_413.n3 a_476_413.t2 46.1549
R65 a_476_413.n5 a_476_413.n4 28.8005
R66 a_476_413.n4 a_476_413.t0 22.637
R67 a_642_307.t1 a_642_307.n0 391.685
R68 a_642_307.n1 a_642_307.t5 370.702
R69 a_642_307.n2 a_642_307.t2 299.377
R70 a_642_307.n2 a_642_307.t3 292.95
R71 a_642_307.n3 a_642_307.t0 244.53
R72 a_642_307.n0 a_642_307.n1 171.589
R73 a_642_307.n1 a_642_307.t4 165.341
R74 a_642_307.n3 a_642_307.n2 152
R75 a_642_307.n0 a_642_307.n3 31.7011
R76 a_957_369.n2 a_957_369.n1 379.344
R77 a_957_369.n1 a_957_369.t0 304.33
R78 a_957_369.n0 a_957_369.t3 241.536
R79 a_957_369.n0 a_957_369.t4 169.237
R80 a_957_369.n1 a_957_369.n0 152
R81 a_957_369.t1 a_957_369.n2 118.508
R82 a_957_369.n2 a_957_369.t2 76.9536
R83 CLK.n1 CLK.t0 269.921
R84 CLK.n0 CLK.t2 255.502
R85 CLK.n1 CLK.t3 234.573
R86 CLK.n0 CLK.t1 233.01
R87 CLK.n2 CLK.n0 180.571
R88 CLK.n2 CLK.n1 152
R89 CLK CLK.n2 10.9719
R90 a_27_47.n0 a_27_47.t4 747.101
R91 a_27_47.t4 a_27_47.t5 660.341
R92 a_27_47.t1 a_27_47.n2 435.587
R93 a_27_47.n2 a_27_47.t0 300.519
R94 a_27_47.n1 a_27_47.t3 266.385
R95 a_27_47.n2 a_27_47.n1 152
R96 a_27_47.n0 a_27_47.t2 91.5805
R97 a_27_47.n1 a_27_47.n0 84.8325
R98 a_1042_47.t0 a_1042_47.t1 60.0005
R99 VNB.t1 VNB.t6 2809.37
R100 VNB.t7 VNB.t5 2677.02
R101 VNB.t0 VNB.t8 2049.99
R102 VNB.t4 VNB.t7 1537.86
R103 VNB.t6 VNB.t0 1517.24
R104 VNB.t3 VNB.t9 1352.75
R105 VNB.t8 VNB.t4 1352.75
R106 VNB.t2 VNB.t1 1196.12
R107 VNB.t5 VNB.t3 1025.24
R108 VNB VNB.t2 911.327
R109 GCLK.n0 GCLK.t1 831.25
R110 GCLK GCLK.t1 824.067
R111 GCLK GCLK.t0 249.829
R112 GCLK.n0 GCLK 77.4939
R113 GCLK GCLK.n0 6.03824
R114 VGND.n14 VGND.t4 265.132
R115 VGND.n6 VGND.n5 214.362
R116 VGND.n4 VGND.n3 209.917
R117 VGND.n17 VGND.n16 198.964
R118 VGND.n3 VGND.t3 70.3307
R119 VGND.n5 VGND.t2 52.8576
R120 VGND.n16 VGND.t0 38.5719
R121 VGND.n16 VGND.t1 38.5719
R122 VGND.n9 VGND.n8 34.6358
R123 VGND.n10 VGND.n9 34.6358
R124 VGND.n10 VGND.n1 34.6358
R125 VGND.n8 VGND.n4 33.5064
R126 VGND.n5 VGND.t6 27.3631
R127 VGND.n3 VGND.t5 24.9241
R128 VGND.n15 VGND.n14 24.8476
R129 VGND.n17 VGND.n15 22.9652
R130 VGND.n14 VGND.n1 19.577
R131 VGND.n15 VGND.n0 9.3005
R132 VGND.n14 VGND.n13 9.3005
R133 VGND.n8 VGND.n7 9.3005
R134 VGND.n9 VGND.n2 9.3005
R135 VGND.n11 VGND.n10 9.3005
R136 VGND.n12 VGND.n1 9.3005
R137 VGND.n18 VGND.n17 7.12063
R138 VGND.n6 VGND.n4 6.70409
R139 VGND.n7 VGND.n6 0.173011
R140 VGND.n18 VGND.n0 0.148519
R141 VGND.n7 VGND.n2 0.120292
R142 VGND.n11 VGND.n2 0.120292
R143 VGND.n12 VGND.n11 0.120292
R144 VGND.n13 VGND.n12 0.120292
R145 VGND.n13 VGND.n0 0.120292
R146 VGND VGND.n18 0.11354
R147 a_651_47.t0 a_651_47.t1 88.1531
R148 a_600_413.t0 a_600_413.t1 98.5005
R149 a_396_119.t0 a_396_119.t1 121.302
R150 a_396_119.n0 a_396_119.t0 29.539
C0 VPB GATE 0.073513f
C1 VPB VPWR 0.14994f
C2 CLK GATE 0.0372f
C3 VPB VGND 0.006063f
C4 CLK VPWR 0.205635f
C5 CLK VGND 0.25787f
C6 GATE VPWR 0.017803f
C7 VPB GCLK 0.01082f
C8 CLK GCLK 0.004248f
C9 GATE VGND 0.089116f
C10 VPWR VGND 0.026372f
C11 GATE GCLK 1.83e-20
C12 VPWR GCLK 0.067933f
C13 VGND GCLK 0.064125f
C14 VPB CLK 0.159354f
C15 GCLK VNB 0.091301f
C16 VGND VNB 0.737323f
C17 VPWR VNB 0.589994f
C18 GATE VNB 0.106385f
C19 CLK VNB 0.360667f
C20 VPB VNB 1.30378f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlclkp_2 VGND VPWR GCLK GATE CLK VPB VNB
X0 a_381_369.t1 GATE.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_957_369.t1 a_643_307.t2 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2016 pd=1.27 as=0.1506 ps=1.33 w=0.64 l=0.15
X2 a_601_413.t0 a_27_47.t2 a_477_413.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0987 ps=0.89 w=0.42 l=0.15
X3 a_397_119.t1 GATE.t1 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.117125 pd=1.085 as=0.1302 ps=1.46 w=0.42 l=0.15
X4 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_1041_47.t0 a_643_307.t3 a_957_369.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 a_477_413.t2 a_193_47.t2 a_381_369.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0968 ps=0.97 w=0.42 l=0.15
X7 VPWR.t3 a_957_369.t3 GCLK.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X8 GCLK.t0 a_957_369.t4 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1506 ps=1.33 w=1 l=0.15
X9 VGND.t2 CLK.t1 a_1041_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.09805 pd=0.98 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_193_47.t1 a_27_47.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_652_47.t0 a_193_47.t3 a_477_413.t3 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.067125 pd=0.745 as=0.1192 ps=1.09 w=0.39 l=0.15
X12 VGND.t0 a_957_369.t5 GCLK.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR.t6 CLK.t2 a_957_369.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1506 pd=1.33 as=0.2016 ps=1.27 w=0.64 l=0.15
X14 a_193_47.t0 a_27_47.t4 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 GCLK.t2 a_957_369.t6 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09805 ps=0.98 w=0.65 l=0.15
X16 a_477_413.t0 a_27_47.t5 a_397_119.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1192 pd=1.09 as=0.117125 ps=1.085 w=0.42 l=0.15
X17 VPWR.t1 a_477_413.t4 a_643_307.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1506 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X18 VGND.t6 a_643_307.t4 a_652_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.114875 pd=1.03 as=0.067125 ps=0.745 w=0.42 l=0.15
X19 VPWR.t2 a_643_307.t5 a_601_413.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X20 a_643_307.t1 a_477_413.t5 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114875 ps=1.03 w=0.65 l=0.15
X21 VGND.t7 CLK.t3 a_27_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 GATE.n0 GATE.t1 189.424
R1 GATE.n0 GATE.t0 183.696
R2 GATE GATE.n0 164.288
R3 VPWR.n23 VPWR.t5 730.923
R4 VPWR.n17 VPWR.t2 666.241
R5 VPWR.n6 VPWR.n5 605.212
R6 VPWR.n25 VPWR.n1 604.394
R7 VPWR.n10 VPWR.n9 600.543
R8 VPWR.n8 VPWR.t3 260.123
R9 VPWR.n5 VPWR.t7 60.0239
R10 VPWR.n9 VPWR.t6 60.0239
R11 VPWR.n1 VPWR.t8 41.5552
R12 VPWR.n1 VPWR.t0 41.5552
R13 VPWR.n18 VPWR.n3 34.6358
R14 VPWR.n22 VPWR.n3 34.6358
R15 VPWR.n12 VPWR.n11 34.6358
R16 VPWR.n5 VPWR.t1 31.6057
R17 VPWR.n9 VPWR.t4 31.6057
R18 VPWR.n18 VPWR.n17 30.8711
R19 VPWR.n16 VPWR.n6 30.4946
R20 VPWR.n24 VPWR.n23 22.9652
R21 VPWR.n25 VPWR.n24 22.9652
R22 VPWR.n11 VPWR.n10 21.4593
R23 VPWR.n23 VPWR.n22 18.824
R24 VPWR.n12 VPWR.n6 17.3181
R25 VPWR.n17 VPWR.n16 15.8123
R26 VPWR.n11 VPWR.n7 9.3005
R27 VPWR.n13 VPWR.n12 9.3005
R28 VPWR.n14 VPWR.n6 9.3005
R29 VPWR.n16 VPWR.n15 9.3005
R30 VPWR.n17 VPWR.n4 9.3005
R31 VPWR.n19 VPWR.n18 9.3005
R32 VPWR.n20 VPWR.n3 9.3005
R33 VPWR.n22 VPWR.n21 9.3005
R34 VPWR.n23 VPWR.n2 9.3005
R35 VPWR.n24 VPWR.n0 9.3005
R36 VPWR.n26 VPWR.n25 7.12063
R37 VPWR.n10 VPWR.n8 6.50647
R38 VPWR.n8 VPWR.n7 0.648786
R39 VPWR.n26 VPWR.n0 0.148519
R40 VPWR.n13 VPWR.n7 0.120292
R41 VPWR.n14 VPWR.n13 0.120292
R42 VPWR.n15 VPWR.n14 0.120292
R43 VPWR.n15 VPWR.n4 0.120292
R44 VPWR.n19 VPWR.n4 0.120292
R45 VPWR.n20 VPWR.n19 0.120292
R46 VPWR.n21 VPWR.n20 0.120292
R47 VPWR.n21 VPWR.n2 0.120292
R48 VPWR.n2 VPWR.n0 0.120292
R49 VPWR VPWR.n26 0.11354
R50 a_381_369.t1 a_381_369.t0 134.631
R51 VPB.t10 VPB.t6 574.277
R52 VPB.t3 VPB.t1 556.386
R53 VPB.t8 VPB.t7 461.683
R54 VPB.t2 VPB.t9 372.974
R55 VPB.t6 VPB.t2 293.248
R56 VPB.t7 VPB.t5 284.113
R57 VPB.t1 VPB.t8 284.113
R58 VPB.t0 VPB.t10 256.592
R59 VPB.t5 VPB.t4 248.599
R60 VPB.t9 VPB.t3 213.084
R61 VPB VPB.t0 195.499
R62 a_643_307.t0 a_643_307.n0 395.272
R63 a_643_307.n3 a_643_307.t4 370.702
R64 a_643_307.n1 a_643_307.t2 299.377
R65 a_643_307.n1 a_643_307.t3 292.95
R66 a_643_307.n2 a_643_307.t1 243.929
R67 a_643_307.n0 a_643_307.n3 171.394
R68 a_643_307.n3 a_643_307.t5 165.341
R69 a_643_307.n2 a_643_307.n1 152
R70 a_643_307.n0 a_643_307.n2 30.9386
R71 a_957_369.n3 a_957_369.n2 379.697
R72 a_957_369.n2 a_957_369.t0 305.745
R73 a_957_369.n0 a_957_369.t3 212.081
R74 a_957_369.n1 a_957_369.t4 212.081
R75 a_957_369.n2 a_957_369.n1 160.764
R76 a_957_369.n0 a_957_369.t5 139.78
R77 a_957_369.n1 a_957_369.t6 139.78
R78 a_957_369.t1 a_957_369.n3 120.047
R79 a_957_369.n3 a_957_369.t2 73.8755
R80 a_957_369.n1 a_957_369.n0 61.346
R81 a_27_47.n0 a_27_47.t5 748.707
R82 a_27_47.t5 a_27_47.t2 660.341
R83 a_27_47.t0 a_27_47.n2 435.587
R84 a_27_47.n2 a_27_47.t1 300.519
R85 a_27_47.n1 a_27_47.t4 266.385
R86 a_27_47.n2 a_27_47.n1 152
R87 a_27_47.n0 a_27_47.t3 91.5805
R88 a_27_47.n1 a_27_47.n0 84.8325
R89 a_477_413.n2 a_477_413.n1 726.838
R90 a_477_413.n3 a_477_413.n2 272.67
R91 a_477_413.n0 a_477_413.t4 235.132
R92 a_477_413.n2 a_477_413.n0 169.649
R93 a_477_413.n0 a_477_413.t5 162.833
R94 a_477_413.n1 a_477_413.t2 121.953
R95 a_477_413.n4 a_477_413.n3 117.081
R96 a_477_413.n1 a_477_413.t1 98.5005
R97 a_477_413.n3 a_477_413.t3 46.1549
R98 a_477_413.n5 a_477_413.n4 28.8005
R99 a_477_413.n4 a_477_413.t0 22.637
R100 a_601_413.t0 a_601_413.t1 98.5005
R101 VGND.n24 VGND.t5 266.56
R102 VGND.n4 VGND.n3 209.547
R103 VGND.n8 VGND.n7 207.213
R104 VGND.n27 VGND.n26 198.964
R105 VGND.n9 VGND.t0 149.364
R106 VGND.n3 VGND.t6 67.979
R107 VGND.n7 VGND.t2 55.7148
R108 VGND.n9 VGND.n8 39.1171
R109 VGND.n26 VGND.t3 38.5719
R110 VGND.n26 VGND.t7 38.5719
R111 VGND.n12 VGND.n6 34.6358
R112 VGND.n13 VGND.n12 34.6358
R113 VGND.n14 VGND.n13 34.6358
R114 VGND.n19 VGND.n18 34.6358
R115 VGND.n20 VGND.n19 34.6358
R116 VGND.n20 VGND.n1 34.6358
R117 VGND.n18 VGND.n4 33.5064
R118 VGND.n7 VGND.t1 25.9346
R119 VGND.n25 VGND.n24 25.224
R120 VGND.n3 VGND.t4 24.9241
R121 VGND.n27 VGND.n25 22.9652
R122 VGND.n24 VGND.n1 19.2005
R123 VGND.n14 VGND.n4 16.9417
R124 VGND.n25 VGND.n0 9.3005
R125 VGND.n24 VGND.n23 9.3005
R126 VGND.n10 VGND.n6 9.3005
R127 VGND.n12 VGND.n11 9.3005
R128 VGND.n13 VGND.n5 9.3005
R129 VGND.n15 VGND.n14 9.3005
R130 VGND.n16 VGND.n4 9.3005
R131 VGND.n18 VGND.n17 9.3005
R132 VGND.n19 VGND.n2 9.3005
R133 VGND.n21 VGND.n20 9.3005
R134 VGND.n22 VGND.n1 9.3005
R135 VGND.n28 VGND.n27 7.12063
R136 VGND.n10 VGND.n9 2.16695
R137 VGND.n8 VGND.n6 0.753441
R138 VGND.n28 VGND.n0 0.148519
R139 VGND.n11 VGND.n10 0.120292
R140 VGND.n11 VGND.n5 0.120292
R141 VGND.n15 VGND.n5 0.120292
R142 VGND.n16 VGND.n15 0.120292
R143 VGND.n17 VGND.n16 0.120292
R144 VGND.n17 VGND.n2 0.120292
R145 VGND.n21 VGND.n2 0.120292
R146 VGND.n22 VGND.n21 0.120292
R147 VGND.n23 VGND.n22 0.120292
R148 VGND.n23 VGND.n0 0.120292
R149 VGND VGND.n28 0.11354
R150 a_397_119.t0 a_397_119.t1 121.302
R151 a_397_119.n0 a_397_119.t0 29.539
R152 VNB.t4 VNB.t7 2823.17
R153 VNB.t6 VNB.t9 2677.02
R154 VNB.t3 VNB.t5 2049.99
R155 VNB.t7 VNB.t3 1517.24
R156 VNB.t8 VNB.t6 1509.39
R157 VNB.t2 VNB.t0 1366.99
R158 VNB.t5 VNB.t8 1352.75
R159 VNB.t0 VNB.t1 1196.12
R160 VNB.t10 VNB.t4 1196.12
R161 VNB.t9 VNB.t2 1025.24
R162 VNB VNB.t10 911.327
R163 CLK.n1 CLK.t0 270.457
R164 CLK.n0 CLK.t2 255.502
R165 CLK.n1 CLK.t3 235.109
R166 CLK.n0 CLK.t1 233.01
R167 CLK.n2 CLK.n0 181.141
R168 CLK.n2 CLK.n1 152
R169 CLK CLK.n2 11.2005
R170 a_1041_47.t0 a_1041_47.t1 60.0005
R171 a_193_47.t0 a_193_47.n1 362.546
R172 a_193_47.n0 a_193_47.t3 351.729
R173 a_193_47.n0 a_193_47.t2 310.882
R174 a_193_47.n1 a_193_47.t1 296.75
R175 a_193_47.n1 a_193_47.n0 94.1934
R176 GCLK GCLK.n0 592.971
R177 GCLK.n2 GCLK.n0 585
R178 GCLK GCLK.n1 185.214
R179 GCLK.n2 GCLK 74.3006
R180 GCLK.n0 GCLK.t1 26.5955
R181 GCLK.n0 GCLK.t0 26.5955
R182 GCLK.n1 GCLK.t3 24.9236
R183 GCLK.n1 GCLK.t2 24.9236
R184 GCLK GCLK.n2 6.03824
R185 a_652_47.t1 a_652_47.t0 88.1531
C0 GATE GCLK 1.83e-20
C1 VPWR VGND 0.049932f
C2 VPWR GCLK 0.150221f
C3 VGND GCLK 0.117708f
C4 VPB CLK 0.160011f
C5 CLK GATE 0.039931f
C6 VPB GATE 0.073792f
C7 CLK VPWR 0.205914f
C8 VPB VPWR 0.166157f
C9 CLK VGND 0.257714f
C10 GATE VPWR 0.017844f
C11 VPB VGND 0.007782f
C12 GATE VGND 0.108425f
C13 CLK GCLK 0.004273f
C14 VPB GCLK 0.004331f
C15 GCLK VNB 0.024772f
C16 VGND VNB 0.812308f
C17 VPWR VNB 0.66373f
C18 GATE VNB 0.107659f
C19 CLK VNB 0.357188f
C20 VPB VNB 1.39235f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlclkp_4 VPWR VGND GCLK CLK GATE VPB VNB
X0 a_381_369.t0 GATE.t0 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_575_47.t0 a_193_47.t2 a_477_413.t2 VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0513 ps=0.645 w=0.36 l=0.15
X2 a_1046_47.t1 a_627_153.t2 a_953_297.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_953_297.t2 a_627_153.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3375 pd=1.675 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR.t4 a_953_297.t3 GCLK.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 GCLK.t7 a_953_297.t4 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t2 a_627_153.t4 a_585_413.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 GCLK.t4 a_953_297.t5 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t9 CLK.t0 a_27_47.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 VPWR.t0 CLK.t1 a_953_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3375 ps=1.675 w=1 l=0.15
X10 GCLK.t3 a_953_297.t6 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.165 ps=1.33 w=1 l=0.15
X11 a_477_413.t3 a_193_47.t3 a_381_369.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0968 ps=0.97 w=0.42 l=0.15
X12 VPWR.t7 a_953_297.t7 GCLK.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X13 a_585_413.t0 a_27_47.t2 a_477_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X14 VPWR.t3 a_477_413.t4 a_627_153.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.26 ps=2.52 w=1 l=0.15
X15 a_477_413.t1 a_27_47.t3 a_381_47.t0 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0513 pd=0.645 as=0.0768 ps=0.805 w=0.36 l=0.15
X16 a_193_47.t0 a_27_47.t4 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 GCLK.t6 a_953_297.t8 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_193_47.t1 a_27_47.t5 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 VGND.t1 a_477_413.t5 a_627_153.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X20 VGND.t3 a_953_297.t9 GCLK.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X21 VGND.t2 a_953_297.t10 GCLK.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_381_47.t1 GATE.t1 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0768 pd=0.805 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND.t0 CLK.t2 a_1046_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VGND.t7 a_627_153.t5 a_575_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X25 VGND.t6 CLK.t3 a_27_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 GATE.n0 GATE.t1 800.12
R1 GATE.n0 GATE.t0 367.928
R2 GATE GATE.n0 165.056
R3 VPWR.n2 VPWR.t10 730.923
R4 VPWR.n4 VPWR.t2 661.833
R5 VPWR.n19 VPWR.n6 605.212
R6 VPWR.n31 VPWR.n1 604.394
R7 VPWR.n12 VPWR.n11 603.708
R8 VPWR.n14 VPWR.n9 314.906
R9 VPWR.n10 VPWR.t4 255.808
R10 VPWR.n1 VPWR.t8 41.5552
R11 VPWR.n1 VPWR.t9 41.5552
R12 VPWR.n6 VPWR.t1 39.4005
R13 VPWR.n25 VPWR.n24 34.6358
R14 VPWR.n26 VPWR.n25 34.6358
R15 VPWR.n18 VPWR.n7 34.6358
R16 VPWR.n9 VPWR.t6 32.5055
R17 VPWR.n9 VPWR.t0 32.5055
R18 VPWR.n32 VPWR.n31 30.7593
R19 VPWR.n6 VPWR.t3 29.5505
R20 VPWR.n20 VPWR.n19 28.9887
R21 VPWR.n14 VPWR.n13 27.8593
R22 VPWR.n11 VPWR.t5 26.5955
R23 VPWR.n11 VPWR.t7 26.5955
R24 VPWR.n24 VPWR.n4 25.977
R25 VPWR.n13 VPWR.n12 24.8476
R26 VPWR.n31 VPWR.n30 22.9652
R27 VPWR.n30 VPWR.n2 22.5887
R28 VPWR.n14 VPWR.n7 21.4593
R29 VPWR.n26 VPWR.n2 19.2005
R30 VPWR.n19 VPWR.n18 18.824
R31 VPWR.n20 VPWR.n4 16.1887
R32 VPWR.n13 VPWR.n8 9.3005
R33 VPWR.n15 VPWR.n14 9.3005
R34 VPWR.n16 VPWR.n7 9.3005
R35 VPWR.n18 VPWR.n17 9.3005
R36 VPWR.n19 VPWR.n5 9.3005
R37 VPWR.n21 VPWR.n20 9.3005
R38 VPWR.n22 VPWR.n4 9.3005
R39 VPWR.n24 VPWR.n23 9.3005
R40 VPWR.n25 VPWR.n3 9.3005
R41 VPWR.n27 VPWR.n26 9.3005
R42 VPWR.n28 VPWR.n2 9.3005
R43 VPWR.n30 VPWR.n29 9.3005
R44 VPWR.n31 VPWR.n0 9.3005
R45 VPWR.n12 VPWR.n10 6.75413
R46 VPWR.n10 VPWR.n8 0.589392
R47 VPWR.n15 VPWR.n8 0.120292
R48 VPWR.n16 VPWR.n15 0.120292
R49 VPWR.n17 VPWR.n16 0.120292
R50 VPWR.n17 VPWR.n5 0.120292
R51 VPWR.n21 VPWR.n5 0.120292
R52 VPWR.n22 VPWR.n21 0.120292
R53 VPWR.n23 VPWR.n22 0.120292
R54 VPWR.n23 VPWR.n3 0.120292
R55 VPWR.n27 VPWR.n3 0.120292
R56 VPWR.n28 VPWR.n27 0.120292
R57 VPWR.n29 VPWR.n28 0.120292
R58 VPWR.n29 VPWR.n0 0.120292
R59 VPWR.n0 VPWR 0.11899
R60 VPWR VPWR.n32 0.0213333
R61 VPWR.n32 VPWR 0.00180208
R62 a_381_369.t0 a_381_369.t1 134.631
R63 VPB.t3 VPB.t4 580.062
R64 VPB.t9 VPB.t11 556.386
R65 VPB.t2 VPB.t0 488.318
R66 VPB.t12 VPB.t1 319.627
R67 VPB.t7 VPB.t8 301.87
R68 VPB.t4 VPB.t2 295.95
R69 VPB.t0 VPB.t7 284.113
R70 VPB.t11 VPB.t12 284.113
R71 VPB.t6 VPB.t5 248.599
R72 VPB.t8 VPB.t6 248.599
R73 VPB.t10 VPB.t9 248.599
R74 VPB.t1 VPB.t3 213.084
R75 VPB VPB.t10 189.409
R76 a_193_47.n0 a_193_47.t2 435.764
R77 a_193_47.t1 a_193_47.n1 388.606
R78 a_193_47.n1 a_193_47.t0 269.942
R79 a_193_47.n0 a_193_47.t3 219.042
R80 a_193_47.n1 a_193_47.n0 202.525
R81 a_477_413.n3 a_477_413.n2 704.822
R82 a_477_413.n2 a_477_413.n1 281
R83 a_477_413.n2 a_477_413.n0 247.243
R84 a_477_413.n0 a_477_413.t4 212.081
R85 a_477_413.n0 a_477_413.t5 143.433
R86 a_477_413.n3 a_477_413.t3 119.608
R87 a_477_413.t0 a_477_413.n3 63.3219
R88 a_477_413.n1 a_477_413.t2 48.3338
R89 a_477_413.n1 a_477_413.t1 46.6672
R90 a_575_47.t1 a_575_47.t0 93.0601
R91 VNB.t2 VNB.t5 2677.02
R92 VNB.t4 VNB.t2 2677.02
R93 VNB.t11 VNB.t12 2677.02
R94 VNB.t12 VNB.t1 1523.62
R95 VNB.t6 VNB.t8 1452.43
R96 VNB.t3 VNB.t4 1352.75
R97 VNB.t1 VNB.t3 1238.83
R98 VNB.t7 VNB.t9 1196.12
R99 VNB.t8 VNB.t7 1196.12
R100 VNB.t0 VNB.t6 1196.12
R101 VNB.t5 VNB.t0 1196.12
R102 VNB.t10 VNB.t11 1196.12
R103 VNB VNB.t10 911.327
R104 a_627_153.t1 a_627_153.n0 395.272
R105 a_627_153.n3 a_627_153.t5 353.757
R106 a_627_153.n1 a_627_153.t2 291.118
R107 a_627_153.n1 a_627_153.t3 263.39
R108 a_627_153.n2 a_627_153.t0 238.347
R109 a_627_153.n2 a_627_153.n1 175.468
R110 a_627_153.n0 a_627_153.n3 172.946
R111 a_627_153.n3 a_627_153.t4 149.822
R112 a_627_153.n0 a_627_153.n2 17.7517
R113 a_953_297.n5 a_953_297.t1 255.042
R114 a_953_297.n6 a_953_297.n5 226.91
R115 a_953_297.n0 a_953_297.t3 212.081
R116 a_953_297.n1 a_953_297.t5 212.081
R117 a_953_297.n2 a_953_297.t7 212.081
R118 a_953_297.n3 a_953_297.t6 212.081
R119 a_953_297.n0 a_953_297.t10 139.78
R120 a_953_297.n1 a_953_297.t8 139.78
R121 a_953_297.n2 a_953_297.t9 139.78
R122 a_953_297.n3 a_953_297.t4 139.78
R123 a_953_297.n5 a_953_297.n4 104.019
R124 a_953_297.t0 a_953_297.n6 96.5305
R125 a_953_297.n1 a_953_297.n0 61.346
R126 a_953_297.n2 a_953_297.n1 61.346
R127 a_953_297.n6 a_953_297.t2 36.4455
R128 a_953_297.n4 a_953_297.n2 35.8991
R129 a_953_297.n4 a_953_297.n3 31.9675
R130 a_1046_47.t0 a_1046_47.t1 49.8467
R131 GCLK GCLK.n1 591.4
R132 GCLK.n5 GCLK.n4 585
R133 GCLK.n4 GCLK.n3 293.384
R134 GCLK.n6 GCLK.n0 233.54
R135 GCLK GCLK.n7 96.7132
R136 GCLK.n1 GCLK.t2 44.3255
R137 GCLK.n0 GCLK.t1 41.539
R138 GCLK.n1 GCLK.t3 26.5955
R139 GCLK.n4 GCLK.t5 26.5955
R140 GCLK.n4 GCLK.t4 26.5955
R141 GCLK.n0 GCLK.t7 24.9236
R142 GCLK.n7 GCLK.t0 24.9236
R143 GCLK.n7 GCLK.t6 24.9236
R144 GCLK.n2 GCLK 9.6005
R145 GCLK.n6 GCLK 7.09868
R146 GCLK GCLK.n5 5.00414
R147 GCLK.n3 GCLK.n2 4.80366
R148 GCLK.n5 GCLK 2.90959
R149 GCLK.n2 GCLK 2.5605
R150 GCLK.n3 GCLK 2.39365
R151 GCLK GCLK.n6 0.815045
R152 VGND.n22 VGND.t7 240.575
R153 VGND.n28 VGND.t9 238.091
R154 VGND.n20 VGND.t1 230.135
R155 VGND.n9 VGND.n8 207.213
R156 VGND.n15 VGND.n14 202.371
R157 VGND.n32 VGND.n1 199.739
R158 VGND.n10 VGND.t2 159.611
R159 VGND.n1 VGND.t8 38.5719
R160 VGND.n1 VGND.t6 38.5719
R161 VGND.n10 VGND.n9 36.6199
R162 VGND.n13 VGND.n7 34.6358
R163 VGND.n16 VGND.n5 34.6358
R164 VGND.n26 VGND.n3 34.6358
R165 VGND.n27 VGND.n26 34.6358
R166 VGND.n33 VGND.n32 30.7593
R167 VGND.n21 VGND.n20 28.9887
R168 VGND.n15 VGND.n13 25.6005
R169 VGND.n8 VGND.t4 24.9236
R170 VGND.n8 VGND.t3 24.9236
R171 VGND.n14 VGND.t5 24.9236
R172 VGND.n14 VGND.t0 24.9236
R173 VGND.n22 VGND.n3 24.4711
R174 VGND.n32 VGND.n0 22.9652
R175 VGND.n16 VGND.n15 22.5887
R176 VGND.n28 VGND.n0 22.5887
R177 VGND.n28 VGND.n27 21.4593
R178 VGND.n22 VGND.n21 19.577
R179 VGND.n20 VGND.n5 18.824
R180 VGND.n32 VGND.n31 9.3005
R181 VGND.n30 VGND.n0 9.3005
R182 VGND.n29 VGND.n28 9.3005
R183 VGND.n27 VGND.n2 9.3005
R184 VGND.n26 VGND.n25 9.3005
R185 VGND.n24 VGND.n3 9.3005
R186 VGND.n23 VGND.n22 9.3005
R187 VGND.n21 VGND.n4 9.3005
R188 VGND.n20 VGND.n19 9.3005
R189 VGND.n18 VGND.n5 9.3005
R190 VGND.n17 VGND.n16 9.3005
R191 VGND.n15 VGND.n6 9.3005
R192 VGND.n13 VGND.n12 9.3005
R193 VGND.n11 VGND.n7 9.3005
R194 VGND.n9 VGND.n7 3.38874
R195 VGND.n11 VGND.n10 2.09743
R196 VGND.n12 VGND.n11 0.120292
R197 VGND.n12 VGND.n6 0.120292
R198 VGND.n17 VGND.n6 0.120292
R199 VGND.n18 VGND.n17 0.120292
R200 VGND.n19 VGND.n18 0.120292
R201 VGND.n19 VGND.n4 0.120292
R202 VGND.n23 VGND.n4 0.120292
R203 VGND.n24 VGND.n23 0.120292
R204 VGND.n25 VGND.n24 0.120292
R205 VGND.n25 VGND.n2 0.120292
R206 VGND.n29 VGND.n2 0.120292
R207 VGND.n30 VGND.n29 0.120292
R208 VGND.n31 VGND.n30 0.120292
R209 VGND.n31 VGND 0.11899
R210 VGND VGND.n33 0.0213333
R211 VGND.n33 VGND 0.00180208
R212 a_585_413.t0 a_585_413.t1 98.5005
R213 CLK.n0 CLK.t0 269.921
R214 CLK.n2 CLK.t1 241.536
R215 CLK.n0 CLK.t3 234.573
R216 CLK.n3 CLK.n2 187.361
R217 CLK.n2 CLK.t2 169.237
R218 CLK.n1 CLK.n0 152
R219 CLK.n1 CLK 11.2005
R220 CLK CLK.n3 4.53383
R221 CLK.n3 CLK.n1 2.4005
R222 a_27_47.t1 a_27_47.n3 391.366
R223 a_27_47.n2 a_27_47.t3 334.421
R224 a_27_47.n2 a_27_47.t2 301.221
R225 a_27_47.n1 a_27_47.t0 289.399
R226 a_27_47.n0 a_27_47.t5 263.173
R227 a_27_47.n0 a_27_47.t4 227.826
R228 a_27_47.n1 a_27_47.n0 152
R229 a_27_47.n3 a_27_47.n2 97.8348
R230 a_27_47.n3 a_27_47.n1 38.9243
R231 a_381_47.n0 a_381_47.t0 86.6672
R232 a_381_47.n0 a_381_47.t1 26.3935
R233 a_381_47.n1 a_381_47.n0 14.4005
C0 GATE VPWR 0.014145f
C1 VGND GCLK 0.266715f
C2 GCLK VPB 0.009094f
C3 GCLK CLK 0.001648f
C4 VGND VPB 0.006419f
C5 GCLK VPWR 0.324772f
C6 VGND CLK 0.252557f
C7 VPB CLK 0.114097f
C8 VGND GATE 0.039776f
C9 VPB GATE 0.056326f
C10 VGND VPWR 0.065494f
C11 VPB VPWR 0.179421f
C12 CLK GATE 0.015777f
C13 CLK VPWR 0.170124f
C14 GCLK VNB 0.027051f
C15 VGND VNB 0.915469f
C16 VPWR VNB 0.739157f
C17 GATE VNB 0.133267f
C18 CLK VNB 0.323619f
C19 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbn_1 VGND VPWR VPB VNB GATE_N D RESET_B Q Q_N
X0 Q.t0 a_724_21.t3 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.22425 ps=1.34 w=0.65 l=0.15
X1 VPWR.t0 D.t0 a_299_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 a_465_47.t1 a_299_47.t2 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_561_413.t2 a_27_47.t2 a_465_47.t0 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X4 Q.t1 a_724_21.t4 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.345 ps=1.69 w=1 l=0.15
X5 a_561_413.t0 a_193_47.t2 a_465_369.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X6 a_724_21.t0 a_561_413.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t3 a_724_21.t5 a_659_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8 VPWR.t7 GATE_N.t0 a_27_47.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 Q_N.t0 a_1308_47.t2 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X10 a_659_47.t0 a_193_47.t3 a_561_413.t1 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X11 VPWR.t5 a_724_21.t6 a_682_413.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 VGND.t1 a_724_21.t7 a_1308_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_193_47.t1 a_27_47.t3 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_682_413.t1 a_27_47.t4 a_561_413.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X15 VPWR.t9 RESET_B.t0 a_724_21.t2 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.155 ps=1.31 w=1 l=0.15
X16 a_942_47.t1 a_561_413.t5 a_724_21.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VPWR.t4 a_724_21.t8 a_1308_47.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X18 a_193_47.t0 a_27_47.t5 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 Q_N.t1 a_1308_47.t3 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X20 VGND.t4 D.t1 a_299_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VGND.t8 RESET_B.t1 a_942_47.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.22425 pd=1.34 as=0.10075 ps=0.96 w=0.65 l=0.15
X22 a_465_369.t1 a_299_47.t3 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND.t5 GATE_N.t1 a_27_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_724_21.n3 a_724_21.t5 368.329
R1 a_724_21.n2 a_724_21.t1 320.801
R2 a_724_21.n5 a_724_21.n4 298.351
R3 a_724_21.n0 a_724_21.t8 247.542
R4 a_724_21.n1 a_724_21.t4 212.081
R5 a_724_21.n4 a_724_21.n3 188.857
R6 a_724_21.n2 a_724_21.n1 173.179
R7 a_724_21.n0 a_724_21.t7 154.356
R8 a_724_21.n3 a_724_21.t6 149.822
R9 a_724_21.n1 a_724_21.t3 139.78
R10 a_724_21.n1 a_724_21.n0 118.309
R11 a_724_21.n4 a_724_21.n2 65.2178
R12 a_724_21.t0 a_724_21.n5 34.4755
R13 a_724_21.n5 a_724_21.t2 26.5955
R14 VGND.n17 VGND.t3 240.833
R15 VGND.n7 VGND.n6 205.75
R16 VGND.n29 VGND.n1 199.739
R17 VGND.n24 VGND.n23 198.964
R18 VGND.n11 VGND.n10 185
R19 VGND.n9 VGND.n8 185
R20 VGND.n10 VGND.n9 64.6159
R21 VGND.n6 VGND.t1 54.2862
R22 VGND.n23 VGND.t7 38.5719
R23 VGND.n23 VGND.t4 38.5719
R24 VGND.n1 VGND.t0 38.5719
R25 VGND.n1 VGND.t5 38.5719
R26 VGND.n10 VGND.t8 35.0774
R27 VGND.n16 VGND.n5 34.6358
R28 VGND.n18 VGND.n3 34.6358
R29 VGND.n22 VGND.n3 34.6358
R30 VGND.n25 VGND.n0 34.6358
R31 VGND.n30 VGND.n29 30.7593
R32 VGND.n9 VGND.t2 27.6928
R33 VGND.n12 VGND.n5 26.4459
R34 VGND.n6 VGND.t6 25.9346
R35 VGND.n24 VGND.n22 24.4711
R36 VGND.n29 VGND.n0 22.9652
R37 VGND.n17 VGND.n16 22.5887
R38 VGND.n18 VGND.n17 21.8358
R39 VGND.n25 VGND.n24 19.9534
R40 VGND.n29 VGND.n28 9.3005
R41 VGND.n13 VGND.n12 9.3005
R42 VGND.n14 VGND.n5 9.3005
R43 VGND.n16 VGND.n15 9.3005
R44 VGND.n17 VGND.n4 9.3005
R45 VGND.n19 VGND.n18 9.3005
R46 VGND.n20 VGND.n3 9.3005
R47 VGND.n22 VGND.n21 9.3005
R48 VGND.n24 VGND.n2 9.3005
R49 VGND.n26 VGND.n25 9.3005
R50 VGND.n27 VGND.n0 9.3005
R51 VGND.n8 VGND.n7 8.18638
R52 VGND.n11 VGND.n8 7.86015
R53 VGND.n12 VGND.n11 1.57243
R54 VGND.n13 VGND.n7 0.214261
R55 VGND.n14 VGND.n13 0.120292
R56 VGND.n15 VGND.n14 0.120292
R57 VGND.n15 VGND.n4 0.120292
R58 VGND.n19 VGND.n4 0.120292
R59 VGND.n20 VGND.n19 0.120292
R60 VGND.n21 VGND.n20 0.120292
R61 VGND.n21 VGND.n2 0.120292
R62 VGND.n26 VGND.n2 0.120292
R63 VGND.n27 VGND.n26 0.120292
R64 VGND.n28 VGND.n27 0.120292
R65 VGND.n28 VGND 0.11899
R66 VGND VGND.n30 0.0213333
R67 VGND.n30 VGND 0.00180208
R68 Q.n0 Q 592
R69 Q.n1 Q.n0 585
R70 Q.n2 Q.t0 209.923
R71 Q.n0 Q.t1 26.5955
R72 Q Q.n2 10.2005
R73 Q Q.n1 7.0005
R74 Q.n1 Q 6.6005
R75 Q.n2 Q 3.4005
R76 VNB.t6 VNB.t4 2677.02
R77 VNB.t5 VNB.t0 2677.02
R78 VNB.t3 VNB.t7 2677.02
R79 VNB.t11 VNB.t6 2392.23
R80 VNB.t10 VNB.t2 1537.86
R81 VNB.t4 VNB.t9 1352.75
R82 VNB.t1 VNB.t5 1352.75
R83 VNB.t0 VNB.t11 1310.03
R84 VNB.t2 VNB.t1 1224.6
R85 VNB.t7 VNB.t10 1196.12
R86 VNB.t8 VNB.t3 1196.12
R87 VNB VNB.t8 669.256
R88 D.n0 D.t0 327.644
R89 D.n0 D.t1 157.338
R90 D D.n0 154.595
R91 a_299_47.t1 a_299_47.n1 438.971
R92 a_299_47.n0 a_299_47.t3 373.283
R93 a_299_47.n1 a_299_47.t0 275.149
R94 a_299_47.n1 a_299_47.n0 156.462
R95 a_299_47.n0 a_299_47.t2 132.282
R96 VPWR.n15 VPWR.t1 868.721
R97 VPWR.n16 VPWR.t5 668.234
R98 VPWR.n27 VPWR.n1 604.394
R99 VPWR.n11 VPWR.n8 318.733
R100 VPWR.n22 VPWR.n4 311.356
R101 VPWR.n10 VPWR.n9 146.25
R102 VPWR.n9 VPWR.t9 75.8455
R103 VPWR.n9 VPWR.t3 60.0855
R104 VPWR.n8 VPWR.t4 58.4849
R105 VPWR.n1 VPWR.t2 41.5552
R106 VPWR.n1 VPWR.t7 41.5552
R107 VPWR.n4 VPWR.t8 41.5552
R108 VPWR.n4 VPWR.t0 41.5552
R109 VPWR.n26 VPWR.n2 34.6358
R110 VPWR.n20 VPWR.n5 34.6358
R111 VPWR.n21 VPWR.n20 34.6358
R112 VPWR.n8 VPWR.t6 31.6057
R113 VPWR.n28 VPWR.n27 30.7593
R114 VPWR.n16 VPWR.n5 27.8593
R115 VPWR.n14 VPWR.n7 26.1544
R116 VPWR.n22 VPWR.n2 25.977
R117 VPWR.n27 VPWR.n26 22.9652
R118 VPWR.n22 VPWR.n21 19.577
R119 VPWR.n15 VPWR.n14 18.0711
R120 VPWR.n16 VPWR.n15 12.8005
R121 VPWR.n11 VPWR.n10 10.0742
R122 VPWR.n12 VPWR.n7 9.3005
R123 VPWR.n14 VPWR.n13 9.3005
R124 VPWR.n15 VPWR.n6 9.3005
R125 VPWR.n17 VPWR.n16 9.3005
R126 VPWR.n18 VPWR.n5 9.3005
R127 VPWR.n20 VPWR.n19 9.3005
R128 VPWR.n21 VPWR.n3 9.3005
R129 VPWR.n23 VPWR.n22 9.3005
R130 VPWR.n24 VPWR.n2 9.3005
R131 VPWR.n26 VPWR.n25 9.3005
R132 VPWR.n27 VPWR.n0 9.3005
R133 VPWR.n10 VPWR.n7 3.89935
R134 VPWR.n12 VPWR.n11 0.213951
R135 VPWR.n13 VPWR.n12 0.120292
R136 VPWR.n13 VPWR.n6 0.120292
R137 VPWR.n17 VPWR.n6 0.120292
R138 VPWR.n18 VPWR.n17 0.120292
R139 VPWR.n19 VPWR.n18 0.120292
R140 VPWR.n19 VPWR.n3 0.120292
R141 VPWR.n23 VPWR.n3 0.120292
R142 VPWR.n24 VPWR.n23 0.120292
R143 VPWR.n25 VPWR.n24 0.120292
R144 VPWR.n25 VPWR.n0 0.120292
R145 VPWR.n0 VPWR 0.11899
R146 VPWR VPWR.n28 0.0213333
R147 VPWR.n28 VPWR 0.00180208
R148 VPB.t7 VPB.t5 556.386
R149 VPB.t6 VPB.t1 556.386
R150 VPB.t4 VPB.t0 556.386
R151 VPB.t11 VPB.t7 497.197
R152 VPB.t2 VPB.t3 358.101
R153 VPB.t10 VPB.t2 284.113
R154 VPB.t5 VPB.t8 281.154
R155 VPB.t1 VPB.t11 272.274
R156 VPB.t0 VPB.t10 248.599
R157 VPB.t9 VPB.t4 248.599
R158 VPB.t3 VPB.t6 213.084
R159 VPB VPB.t9 139.097
R160 a_465_47.n0 a_465_47.t0 88.3338
R161 a_465_47.n0 a_465_47.t1 26.3935
R162 a_465_47.n1 a_465_47.n0 14.4005
R163 a_27_47.t0 a_27_47.n3 411.32
R164 a_27_47.n2 a_27_47.t4 316.111
R165 a_27_47.n2 a_27_47.t2 315.729
R166 a_27_47.n1 a_27_47.t1 289.399
R167 a_27_47.n0 a_27_47.t5 263.173
R168 a_27_47.n0 a_27_47.t3 227.826
R169 a_27_47.n1 a_27_47.n0 152
R170 a_27_47.n3 a_27_47.n2 20.5706
R171 a_27_47.n3 a_27_47.n1 18.9713
R172 a_561_413.n3 a_561_413.n2 692.672
R173 a_561_413.n2 a_561_413.n1 258.964
R174 a_561_413.n2 a_561_413.n0 247.139
R175 a_561_413.n0 a_561_413.t4 212.081
R176 a_561_413.n0 a_561_413.t5 139.78
R177 a_561_413.t0 a_561_413.n3 121.953
R178 a_561_413.n3 a_561_413.t3 91.4648
R179 a_561_413.n1 a_561_413.t1 46.6672
R180 a_561_413.n1 a_561_413.t2 46.6672
R181 a_193_47.n0 a_193_47.t3 464.327
R182 a_193_47.t0 a_193_47.n1 366.837
R183 a_193_47.n1 a_193_47.t1 322.567
R184 a_193_47.n0 a_193_47.t2 242.607
R185 a_193_47.n1 a_193_47.n0 187.469
R186 a_465_369.t1 a_465_369.t0 134.631
R187 a_659_47.t1 a_659_47.t0 93.0601
R188 GATE_N.n0 GATE_N.t0 269.921
R189 GATE_N.n0 GATE_N.t1 234.573
R190 GATE_N.n1 GATE_N.n0 152
R191 GATE_N GATE_N.n1 10.9719
R192 GATE_N.n1 GATE_N 6.79234
R193 a_1308_47.t0 a_1308_47.n1 669.563
R194 a_1308_47.n1 a_1308_47.t1 310.536
R195 a_1308_47.n0 a_1308_47.t2 237.736
R196 a_1308_47.n1 a_1308_47.n0 175.274
R197 a_1308_47.n0 a_1308_47.t3 165.435
R198 Q_N Q_N.n0 593.615
R199 Q_N.n2 Q_N.n0 585
R200 Q_N.n1 Q_N.t1 209.923
R201 Q_N Q_N.n1 95.1636
R202 Q_N.n0 Q_N.t0 26.5955
R203 Q_N.n2 Q_N 8.61589
R204 Q_N Q_N.n2 8.12358
R205 Q_N.n1 Q_N 0.246654
R206 a_682_413.t0 a_682_413.t1 98.5005
R207 RESET_B.n0 RESET_B.t0 241.536
R208 RESET_B.n0 RESET_B.t1 169.237
R209 RESET_B.n1 RESET_B.n0 152
R210 RESET_B.n1 RESET_B 10.2793
R211 RESET_B RESET_B.n1 7.56414
R212 a_942_47.t0 a_942_47.t1 57.2313
C0 VPB D 0.062359f
C1 VPB RESET_B 0.032759f
C2 VPB VPWR 0.178959f
C3 VPB VGND 0.01802f
C4 GATE_N VPWR 0.017119f
C5 GATE_N VGND 0.016722f
C6 D VPWR 0.014067f
C7 VPB Q 0.010863f
C8 RESET_B VPWR 0.022902f
C9 D VGND 0.018848f
C10 VPB Q_N 0.012588f
C11 RESET_B VGND 0.020616f
C12 VPWR VGND 0.113762f
C13 RESET_B Q 3.7e-19
C14 VPWR Q 0.09374f
C15 VGND Q 0.066748f
C16 VPWR Q_N 0.093603f
C17 VPB GATE_N 0.069313f
C18 VGND Q_N 0.057819f
C19 Q_N VNB 0.094005f
C20 Q VNB 0.012022f
C21 VGND VNB 0.883329f
C22 VPWR VNB 0.702992f
C23 RESET_B VNB 0.101428f
C24 D VNB 0.132433f
C25 GATE_N VNB 0.194986f
C26 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbp_1 VGND VPWR VPB VNB Q_N Q RESET_B D GATE
X0 Q.t0 a_711_307.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.23075 ps=1.36 w=0.65 l=0.15
X1 VPWR.t8 D.t0 a_299_47.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 a_560_47.t3 a_193_47.t2 a_465_47.t1 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0612 pd=0.7 as=0.066 ps=0.745 w=0.36 l=0.15
X3 a_645_413.t1 a_193_47.t3 a_560_47.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR.t2 a_711_307.t4 a_645_413.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_465_47.t0 a_299_47.t2 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND.t6 RESET_B.t0 a_941_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.23075 pd=1.36 as=0.095875 ps=0.945 w=0.65 l=0.15
X7 Q.t1 a_711_307.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.355 ps=1.71 w=1 l=0.15
X8 a_560_47.t0 a_27_47.t2 a_465_369.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0968 ps=0.97 w=0.42 l=0.15
X9 VPWR.t5 GATE.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 VGND.t5 a_711_307.t6 a_658_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11 Q_N.t1 a_1308_47.t2 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X12 a_658_47.t1 a_27_47.t3 a_560_47.t1 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0612 ps=0.7 w=0.36 l=0.15
X13 VGND.t4 a_711_307.t7 a_1308_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_193_47.t0 a_27_47.t4 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_711_307.t1 a_560_47.t4 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X16 a_941_47.t0 a_560_47.t5 a_711_307.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VPWR.t3 a_711_307.t8 a_1308_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X18 a_193_47.t1 a_27_47.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 Q_N.t0 a_1308_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X20 VGND.t0 D.t1 a_299_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VPWR.t1 RESET_B.t1 a_711_307.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.355 pd=1.71 as=0.155 ps=1.31 w=1 l=0.15
X22 a_465_369.t0 a_299_47.t3 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND.t8 GATE.t1 a_27_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_711_307.n3 a_711_307.t6 366.002
R1 a_711_307.n2 a_711_307.t2 324.433
R2 a_711_307.n5 a_711_307.n4 299.93
R3 a_711_307.n0 a_711_307.t8 269.921
R4 a_711_307.n1 a_711_307.t5 212.081
R5 a_711_307.n4 a_711_307.n3 188.462
R6 a_711_307.n0 a_711_307.t7 176.733
R7 a_711_307.n2 a_711_307.n1 170.988
R8 a_711_307.n3 a_711_307.t4 147.495
R9 a_711_307.n1 a_711_307.t3 139.78
R10 a_711_307.n1 a_711_307.n0 137.298
R11 a_711_307.n4 a_711_307.n2 69.2216
R12 a_711_307.n5 a_711_307.t1 34.4755
R13 a_711_307.t0 a_711_307.n5 26.5955
R14 VGND.n4 VGND.t5 240.575
R15 VGND.n9 VGND.n7 205.748
R16 VGND.n28 VGND.n27 199.739
R17 VGND.n2 VGND.n1 198.964
R18 VGND.n13 VGND.n12 185
R19 VGND.n11 VGND.n10 185
R20 VGND.n12 VGND.n11 81.2313
R21 VGND.n7 VGND.t4 54.2862
R22 VGND.n1 VGND.t7 38.5719
R23 VGND.n1 VGND.t0 38.5719
R24 VGND.n27 VGND.t1 38.5719
R25 VGND.n27 VGND.t8 38.5719
R26 VGND.n15 VGND.n14 34.6358
R27 VGND.n20 VGND.n19 34.6358
R28 VGND.n21 VGND.n20 34.6358
R29 VGND.n26 VGND.n25 34.6358
R30 VGND.n7 VGND.t2 25.9346
R31 VGND.n14 VGND.n13 25.5411
R32 VGND.n11 VGND.t3 24.9236
R33 VGND.n12 VGND.t6 24.9236
R34 VGND.n21 VGND.n2 24.4711
R35 VGND.n28 VGND.n26 22.9652
R36 VGND.n15 VGND.n4 22.5887
R37 VGND.n19 VGND.n4 21.4593
R38 VGND.n25 VGND.n2 19.9534
R39 VGND.n10 VGND.n6 9.76892
R40 VGND.n8 VGND.n6 9.3005
R41 VGND.n14 VGND.n5 9.3005
R42 VGND.n16 VGND.n15 9.3005
R43 VGND.n17 VGND.n4 9.3005
R44 VGND.n19 VGND.n18 9.3005
R45 VGND.n20 VGND.n3 9.3005
R46 VGND.n22 VGND.n21 9.3005
R47 VGND.n23 VGND.n2 9.3005
R48 VGND.n25 VGND.n24 9.3005
R49 VGND.n26 VGND.n0 9.3005
R50 VGND.n10 VGND.n9 7.8135
R51 VGND.n29 VGND.n28 7.12063
R52 VGND.n9 VGND.n8 0.215935
R53 VGND.n29 VGND.n0 0.148519
R54 VGND.n8 VGND.n5 0.120292
R55 VGND.n16 VGND.n5 0.120292
R56 VGND.n17 VGND.n16 0.120292
R57 VGND.n18 VGND.n17 0.120292
R58 VGND.n18 VGND.n3 0.120292
R59 VGND.n22 VGND.n3 0.120292
R60 VGND.n23 VGND.n22 0.120292
R61 VGND.n24 VGND.n23 0.120292
R62 VGND.n24 VGND.n0 0.120292
R63 VGND VGND.n29 0.11354
R64 VGND.n13 VGND.n6 0.112781
R65 Q.n0 Q 591.4
R66 Q.n1 Q.n0 585
R67 Q.n2 Q.t0 209.923
R68 Q.n0 Q.t1 26.5955
R69 Q Q.n2 9.32621
R70 Q Q.n1 6.4005
R71 Q.n1 Q 6.03479
R72 Q.n2 Q 3.10907
R73 VNB.t5 VNB.t3 2677.02
R74 VNB.t4 VNB.t11 2677.02
R75 VNB.t1 VNB.t0 2677.02
R76 VNB.t6 VNB.t5 2449.19
R77 VNB.t8 VNB.t10 1395.47
R78 VNB.t3 VNB.t2 1352.75
R79 VNB.t10 VNB.t4 1352.75
R80 VNB.t7 VNB.t8 1352.75
R81 VNB.t11 VNB.t6 1267.31
R82 VNB.t0 VNB.t7 1196.12
R83 VNB.t9 VNB.t1 1196.12
R84 VNB VNB.t9 669.256
R85 D.n0 D.t0 327.644
R86 D.n0 D.t1 157.338
R87 D D.n0 154.595
R88 a_299_47.t1 a_299_47.n1 438.971
R89 a_299_47.n0 a_299_47.t3 373.283
R90 a_299_47.n1 a_299_47.t0 275.149
R91 a_299_47.n1 a_299_47.n0 156.462
R92 a_299_47.n0 a_299_47.t2 132.282
R93 VPWR.n17 VPWR.t9 853.981
R94 VPWR.n5 VPWR.t2 648.322
R95 VPWR.n30 VPWR.n1 604.394
R96 VPWR.n9 VPWR.n8 318.733
R97 VPWR.n3 VPWR.n2 311.356
R98 VPWR.n10 VPWR.n7 292.5
R99 VPWR.n12 VPWR.n11 292.5
R100 VPWR.n11 VPWR.n10 86.6805
R101 VPWR.n8 VPWR.t3 58.4849
R102 VPWR.n1 VPWR.t0 41.5552
R103 VPWR.n1 VPWR.t5 41.5552
R104 VPWR.n2 VPWR.t6 41.5552
R105 VPWR.n2 VPWR.t8 41.5552
R106 VPWR.n29 VPWR.n28 34.6358
R107 VPWR.n23 VPWR.n22 34.6358
R108 VPWR.n24 VPWR.n23 34.6358
R109 VPWR.n8 VPWR.t7 31.6057
R110 VPWR.n11 VPWR.t4 26.5955
R111 VPWR.n10 VPWR.t1 26.5955
R112 VPWR.n28 VPWR.n3 25.977
R113 VPWR.n22 VPWR.n5 24.5891
R114 VPWR.n16 VPWR.n7 24.2634
R115 VPWR.n30 VPWR.n29 22.9652
R116 VPWR.n17 VPWR.n16 21.6054
R117 VPWR.n24 VPWR.n3 19.577
R118 VPWR.n14 VPWR.n13 9.3005
R119 VPWR.n16 VPWR.n15 9.3005
R120 VPWR.n18 VPWR.n6 9.3005
R121 VPWR.n20 VPWR.n19 9.3005
R122 VPWR.n22 VPWR.n21 9.3005
R123 VPWR.n23 VPWR.n4 9.3005
R124 VPWR.n25 VPWR.n24 9.3005
R125 VPWR.n26 VPWR.n3 9.3005
R126 VPWR.n28 VPWR.n27 9.3005
R127 VPWR.n29 VPWR.n0 9.3005
R128 VPWR.n19 VPWR.n18 8.78856
R129 VPWR.n12 VPWR.n9 7.57306
R130 VPWR.n31 VPWR.n30 7.12063
R131 VPWR.n13 VPWR.n12 6.4005
R132 VPWR.n19 VPWR.n5 1.33781
R133 VPWR.n18 VPWR.n17 0.669157
R134 VPWR.n14 VPWR.n9 0.213951
R135 VPWR.n31 VPWR.n0 0.148519
R136 VPWR.n15 VPWR.n14 0.120292
R137 VPWR.n15 VPWR.n6 0.120292
R138 VPWR.n20 VPWR.n6 0.120292
R139 VPWR.n21 VPWR.n20 0.120292
R140 VPWR.n21 VPWR.n4 0.120292
R141 VPWR.n25 VPWR.n4 0.120292
R142 VPWR.n26 VPWR.n25 0.120292
R143 VPWR.n27 VPWR.n26 0.120292
R144 VPWR.n27 VPWR.n0 0.120292
R145 VPWR VPWR.n31 0.11354
R146 VPWR.n13 VPWR.n7 0.0740632
R147 VPB.t5 VPB.t11 583.023
R148 VPB.t4 VPB.t3 556.386
R149 VPB.t0 VPB.t10 556.386
R150 VPB.t1 VPB.t4 509.034
R151 VPB.t2 VPB.t5 284.113
R152 VPB.t8 VPB.t7 284.113
R153 VPB.t3 VPB.t9 281.154
R154 VPB.t11 VPB.t1 272.274
R155 VPB.t7 VPB.t2 248.599
R156 VPB.t10 VPB.t8 248.599
R157 VPB.t6 VPB.t0 248.599
R158 VPB VPB.t6 139.097
R159 a_193_47.t1 a_193_47.n1 366.837
R160 a_193_47.n0 a_193_47.t2 337.24
R161 a_193_47.n1 a_193_47.t0 322.567
R162 a_193_47.n0 a_193_47.t3 300.252
R163 a_193_47.n1 a_193_47.n0 25.0495
R164 a_465_47.n0 a_465_47.t1 66.6672
R165 a_465_47.n0 a_465_47.t0 26.3935
R166 a_465_47.n1 a_465_47.n0 14.4005
R167 a_560_47.n3 a_560_47.n2 699.951
R168 a_560_47.n2 a_560_47.n1 285.894
R169 a_560_47.n2 a_560_47.n0 247.619
R170 a_560_47.n0 a_560_47.t4 212.081
R171 a_560_47.n0 a_560_47.t5 141.971
R172 a_560_47.n1 a_560_47.t1 68.3338
R173 a_560_47.n3 a_560_47.t2 63.3219
R174 a_560_47.t0 a_560_47.n3 63.3219
R175 a_560_47.n1 a_560_47.t3 45.0005
R176 a_645_413.t0 a_645_413.t1 154.786
R177 RESET_B.n0 RESET_B.t1 241.536
R178 RESET_B.n0 RESET_B.t0 169.237
R179 RESET_B.n1 RESET_B.n0 152
R180 RESET_B.n1 RESET_B 10.8611
R181 RESET_B RESET_B.n1 6.98232
R182 a_941_47.t0 a_941_47.t1 54.462
R183 a_27_47.n2 a_27_47.t3 462.721
R184 a_27_47.t0 a_27_47.n3 411.32
R185 a_27_47.n1 a_27_47.t1 289.399
R186 a_27_47.n0 a_27_47.t5 263.173
R187 a_27_47.n2 a_27_47.t2 242.607
R188 a_27_47.n0 a_27_47.t4 227.826
R189 a_27_47.n3 a_27_47.n2 176.62
R190 a_27_47.n1 a_27_47.n0 152
R191 a_27_47.n3 a_27_47.n1 18.9713
R192 a_465_369.t0 a_465_369.t1 134.631
R193 GATE.n0 GATE.t0 272.062
R194 GATE.n0 GATE.t1 236.716
R195 GATE.n1 GATE.n0 152
R196 GATE GATE.n1 11.2005
R197 GATE.n1 GATE 6.93383
R198 a_658_47.t0 a_658_47.t1 93.0601
R199 a_1308_47.t1 a_1308_47.n1 669.563
R200 a_1308_47.n1 a_1308_47.t0 251.744
R201 a_1308_47.n0 a_1308_47.t2 238.59
R202 a_1308_47.n1 a_1308_47.n0 175.468
R203 a_1308_47.n0 a_1308_47.t3 166.291
R204 Q_N Q_N.n0 593.615
R205 Q_N.n2 Q_N.n0 585
R206 Q_N.n1 Q_N.t0 209.923
R207 Q_N Q_N.n1 97.7236
R208 Q_N.n0 Q_N.t1 26.5955
R209 Q_N.n2 Q_N 8.61589
R210 Q_N Q_N.n2 8.12358
R211 Q_N.n1 Q_N 0.246654
C0 VPB Q_N 0.01204f
C1 D VGND 0.018848f
C2 RESET_B VPWR 0.022807f
C3 RESET_B VGND 0.020733f
C4 RESET_B Q 3.58e-19
C5 VPWR VGND 0.11381f
C6 VPWR Q 0.09799f
C7 VPWR Q_N 0.093564f
C8 VGND Q 0.071859f
C9 VPB GATE 0.069428f
C10 VGND Q_N 0.057733f
C11 VPB D 0.062359f
C12 VPB RESET_B 0.032905f
C13 VPB VPWR 0.174768f
C14 GATE VPWR 0.017104f
C15 VPB VGND 0.017645f
C16 VPB Q 0.01158f
C17 D VPWR 0.014067f
C18 GATE VGND 0.016701f
C19 Q_N VNB 0.093502f
C20 Q VNB 0.012518f
C21 VGND VNB 0.881174f
C22 VPWR VNB 0.702185f
C23 RESET_B VNB 0.101527f
C24 D VNB 0.132433f
C25 GATE VNB 0.195339f
C26 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_1 VGND VPWR VPB VNB GATE_N D RESET_B Q
X0 VPWR.t5 D.t0 a_299_47.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_465_47.t1 a_299_47.t2 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_561_413.t1 a_27_47.t2 a_465_47.t0 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X3 a_561_413.t2 a_193_47.t2 a_465_369.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X4 a_724_21.t0 a_561_413.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND.t6 a_724_21.t3 a_659_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6 VPWR.t1 GATE_N.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_659_47.t1 a_193_47.t3 a_561_413.t3 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X8 VPWR.t3 a_724_21.t4 a_682_413.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 Q.t0 a_724_21.t5 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3825 ps=1.765 w=1 l=0.15
X10 a_193_47.t1 a_27_47.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_682_413.t0 a_27_47.t4 a_561_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X12 a_942_47.t0 a_561_413.t5 a_724_21.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47.t0 a_27_47.t5 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14 Q.t1 a_724_21.t6 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.248625 ps=1.415 w=0.65 l=0.15
X15 VPWR.t7 RESET_B.t0 a_724_21.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t4 D.t1 a_299_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t3 RESET_B.t1 a_942_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.248625 pd=1.415 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_465_369.t0 a_299_47.t3 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 VGND.t1 GATE_N.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 327.644
R1 D.n0 D.t1 157.338
R2 D D.n0 154.595
R3 a_299_47.t1 a_299_47.n1 438.971
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t0 275.149
R6 a_299_47.n1 a_299_47.n0 156.462
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n15 VPWR.t0 871.352
R9 VPWR.n16 VPWR.t3 666.86
R10 VPWR.n27 VPWR.n1 604.394
R11 VPWR.n11 VPWR.n10 585.15
R12 VPWR.n9 VPWR.n8 585
R13 VPWR.n22 VPWR.n4 311.356
R14 VPWR.n10 VPWR.n9 80.7705
R15 VPWR.n9 VPWR.t7 43.3405
R16 VPWR.n1 VPWR.t2 41.5552
R17 VPWR.n1 VPWR.t1 41.5552
R18 VPWR.n4 VPWR.t6 41.5552
R19 VPWR.n4 VPWR.t5 41.5552
R20 VPWR.n26 VPWR.n2 34.6358
R21 VPWR.n20 VPWR.n5 34.6358
R22 VPWR.n21 VPWR.n20 34.6358
R23 VPWR.n28 VPWR.n27 30.7593
R24 VPWR.n16 VPWR.n5 27.8593
R25 VPWR.n10 VPWR.t4 26.5955
R26 VPWR.n22 VPWR.n2 25.977
R27 VPWR.n14 VPWR.n7 24.5217
R28 VPWR.n27 VPWR.n26 22.9652
R29 VPWR.n22 VPWR.n21 19.577
R30 VPWR.n15 VPWR.n14 18.824
R31 VPWR.n16 VPWR.n15 14.3064
R32 VPWR.n12 VPWR.n7 9.3005
R33 VPWR.n14 VPWR.n13 9.3005
R34 VPWR.n15 VPWR.n6 9.3005
R35 VPWR.n17 VPWR.n16 9.3005
R36 VPWR.n18 VPWR.n5 9.3005
R37 VPWR.n20 VPWR.n19 9.3005
R38 VPWR.n21 VPWR.n3 9.3005
R39 VPWR.n23 VPWR.n22 9.3005
R40 VPWR.n24 VPWR.n2 9.3005
R41 VPWR.n26 VPWR.n25 9.3005
R42 VPWR.n27 VPWR.n0 9.3005
R43 VPWR.n11 VPWR.n8 7.68361
R44 VPWR.n12 VPWR.n11 7.39269
R45 VPWR.n8 VPWR.n7 1.14677
R46 VPWR.n13 VPWR.n12 0.120292
R47 VPWR.n13 VPWR.n6 0.120292
R48 VPWR.n17 VPWR.n6 0.120292
R49 VPWR.n18 VPWR.n17 0.120292
R50 VPWR.n19 VPWR.n18 0.120292
R51 VPWR.n19 VPWR.n3 0.120292
R52 VPWR.n23 VPWR.n3 0.120292
R53 VPWR.n24 VPWR.n23 0.120292
R54 VPWR.n25 VPWR.n24 0.120292
R55 VPWR.n25 VPWR.n0 0.120292
R56 VPWR.n0 VPWR 0.11899
R57 VPWR VPWR.n28 0.0213333
R58 VPWR.n28 VPWR 0.00180208
R59 VPB.t4 VPB.t0 556.386
R60 VPB.t3 VPB.t6 556.386
R61 VPB.t8 VPB.t5 541.59
R62 VPB.t9 VPB.t2 358.101
R63 VPB.t7 VPB.t9 284.113
R64 VPB.t0 VPB.t8 248.599
R65 VPB.t6 VPB.t7 248.599
R66 VPB.t1 VPB.t3 248.599
R67 VPB.t2 VPB.t4 213.084
R68 VPB VPB.t1 139.097
R69 VGND.n4 VGND.t6 240.833
R70 VGND.n26 VGND.n25 199.739
R71 VGND.n2 VGND.n1 198.964
R72 VGND.n9 VGND.n8 185.089
R73 VGND.n7 VGND.n6 185
R74 VGND.n8 VGND.n7 74.7697
R75 VGND.n7 VGND.t3 40.6159
R76 VGND.n1 VGND.t5 38.5719
R77 VGND.n1 VGND.t4 38.5719
R78 VGND.n25 VGND.t2 38.5719
R79 VGND.n25 VGND.t1 38.5719
R80 VGND.n13 VGND.n12 34.6358
R81 VGND.n18 VGND.n17 34.6358
R82 VGND.n19 VGND.n18 34.6358
R83 VGND.n24 VGND.n23 34.6358
R84 VGND.n8 VGND.t0 25.8467
R85 VGND.n19 VGND.n2 24.4711
R86 VGND.n12 VGND.n11 24.3324
R87 VGND.n26 VGND.n24 22.9652
R88 VGND.n13 VGND.n4 22.5887
R89 VGND.n17 VGND.n4 21.8358
R90 VGND.n23 VGND.n2 19.9534
R91 VGND.n11 VGND.n10 9.3005
R92 VGND.n12 VGND.n5 9.3005
R93 VGND.n14 VGND.n13 9.3005
R94 VGND.n15 VGND.n4 9.3005
R95 VGND.n17 VGND.n16 9.3005
R96 VGND.n18 VGND.n3 9.3005
R97 VGND.n20 VGND.n19 9.3005
R98 VGND.n21 VGND.n2 9.3005
R99 VGND.n23 VGND.n22 9.3005
R100 VGND.n24 VGND.n0 9.3005
R101 VGND.n9 VGND.n6 9.00713
R102 VGND.n10 VGND.n9 7.43627
R103 VGND.n27 VGND.n26 7.12063
R104 VGND.n11 VGND.n6 1.34787
R105 VGND.n27 VGND.n0 0.148519
R106 VGND.n10 VGND.n5 0.120292
R107 VGND.n14 VGND.n5 0.120292
R108 VGND.n15 VGND.n14 0.120292
R109 VGND.n16 VGND.n15 0.120292
R110 VGND.n16 VGND.n3 0.120292
R111 VGND.n20 VGND.n3 0.120292
R112 VGND.n21 VGND.n20 0.120292
R113 VGND.n22 VGND.n21 0.120292
R114 VGND.n22 VGND.n0 0.120292
R115 VGND VGND.n27 0.0927068
R116 a_465_47.n0 a_465_47.t0 88.3338
R117 a_465_47.n0 a_465_47.t1 26.3935
R118 a_465_47.n1 a_465_47.n0 14.4005
R119 VNB.t9 VNB.t0 2677.02
R120 VNB.t4 VNB.t6 2677.02
R121 VNB.t5 VNB.t2 2605.83
R122 VNB.t7 VNB.t1 1537.86
R123 VNB.t8 VNB.t9 1352.75
R124 VNB.t1 VNB.t8 1224.6
R125 VNB.t0 VNB.t5 1196.12
R126 VNB.t6 VNB.t7 1196.12
R127 VNB.t3 VNB.t4 1196.12
R128 VNB VNB.t3 669.256
R129 a_27_47.t0 a_27_47.n3 415.863
R130 a_27_47.n2 a_27_47.t4 316.111
R131 a_27_47.n2 a_27_47.t2 315.729
R132 a_27_47.n1 a_27_47.t1 294.873
R133 a_27_47.n0 a_27_47.t5 263.173
R134 a_27_47.n0 a_27_47.t3 227.826
R135 a_27_47.n1 a_27_47.n0 152
R136 a_27_47.n3 a_27_47.n2 20.5706
R137 a_27_47.n3 a_27_47.n1 18.9713
R138 a_561_413.n3 a_561_413.n2 747.072
R139 a_561_413.n2 a_561_413.n1 281.274
R140 a_561_413.n2 a_561_413.n0 253.439
R141 a_561_413.n0 a_561_413.t4 221.72
R142 a_561_413.n0 a_561_413.t5 149.421
R143 a_561_413.n3 a_561_413.t2 121.953
R144 a_561_413.t0 a_561_413.n3 91.4648
R145 a_561_413.n1 a_561_413.t3 46.6672
R146 a_561_413.n1 a_561_413.t1 46.6672
R147 a_193_47.n0 a_193_47.t3 464.327
R148 a_193_47.t0 a_193_47.n1 366.837
R149 a_193_47.n1 a_193_47.t1 322.567
R150 a_193_47.n0 a_193_47.t2 242.607
R151 a_193_47.n1 a_193_47.n0 187.469
R152 a_465_369.t0 a_465_369.t1 134.631
R153 a_724_21.n2 a_724_21.t3 368.329
R154 a_724_21.n4 a_724_21.n3 299.166
R155 a_724_21.n0 a_724_21.t5 235.471
R156 a_724_21.n1 a_724_21.t1 228.059
R157 a_724_21.n3 a_724_21.n2 187.685
R158 a_724_21.n0 a_724_21.t6 163.172
R159 a_724_21.n1 a_724_21.n0 152
R160 a_724_21.n2 a_724_21.t4 149.822
R161 a_724_21.n3 a_724_21.n1 50.6853
R162 a_724_21.n4 a_724_21.t2 26.5955
R163 a_724_21.t0 a_724_21.n4 26.5955
R164 a_659_47.t0 a_659_47.t1 93.0601
R165 GATE_N.n0 GATE_N.t0 269.921
R166 GATE_N.n0 GATE_N.t1 234.573
R167 GATE_N.n1 GATE_N.n0 152
R168 GATE_N GATE_N.n1 10.9719
R169 GATE_N.n1 GATE_N 6.79234
R170 a_682_413.t0 a_682_413.t1 98.5005
R171 Q.n0 Q.t0 374.618
R172 Q.n1 Q.t1 209.923
R173 Q Q.n1 9.10819
R174 Q Q.n0 8.95158
R175 Q.n0 Q 7.65628
R176 Q.n1 Q 7.63127
R177 a_942_47.t0 a_942_47.t1 49.8467
R178 RESET_B.n0 RESET_B.t0 241.536
R179 RESET_B.n0 RESET_B.t1 169.237
R180 RESET_B.n1 RESET_B.n0 152
R181 RESET_B.n1 RESET_B 10.6672
R182 RESET_B RESET_B.n1 7.17626
C0 RESET_B VGND 0.020525f
C1 VPB GATE_N 0.070092f
C2 VPWR VGND 0.083329f
C3 RESET_B Q 4.35e-19
C4 VPB D 0.062359f
C5 VPWR Q 0.068789f
C6 VPB RESET_B 0.032594f
C7 VGND Q 0.03582f
C8 VPB VPWR 0.146436f
C9 VPB VGND 0.013642f
C10 VPB Q 0.010449f
C11 GATE_N VPWR 0.019242f
C12 D VPWR 0.014067f
C13 GATE_N VGND 0.019085f
C14 D VGND 0.018848f
C15 RESET_B VPWR 0.020489f
C16 Q VNB 0.088693f
C17 VGND VNB 0.745621f
C18 VPWR VNB 0.58894f
C19 RESET_B VNB 0.102165f
C20 D VNB 0.132433f
C21 GATE_N VNB 0.195771f
C22 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_2 VGND VPWR VPB VNB Q RESET_B D GATE_N
X0 VPWR.t0 D.t0 a_299_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47.t3 a_27_47.t2 a_465_47.t1 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.0612 pd=0.7 as=0.066 ps=0.745 w=0.36 l=0.15
X2 a_645_413.t1 a_27_47.t3 a_560_47.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR.t1 a_711_307.t3 a_645_413.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.45 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_465_47.t0 a_299_47.t2 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VPWR.t6 RESET_B.t0 a_711_307.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6 a_560_47.t0 a_193_47.t2 a_465_369.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0968 ps=0.97 w=0.42 l=0.15
X7 VPWR.t8 GATE_N.t0 a_27_47.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 Q.t1 a_711_307.t4 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.165 ps=1.33 w=1 l=0.15
X9 VGND.t4 a_711_307.t5 a_658_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10 a_658_47.t0 a_193_47.t3 a_560_47.t1 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0612 ps=0.7 w=0.36 l=0.15
X11 VPWR.t4 a_711_307.t6 Q.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X12 a_193_47.t1 a_27_47.t4 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_711_307.t1 a_560_47.t4 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Q.t3 a_711_307.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15 a_941_47.t1 a_560_47.t5 a_711_307.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_193_47.t0 a_27_47.t5 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X17 VGND.t2 a_711_307.t8 Q.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t0 D.t1 a_299_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 VGND.t5 RESET_B.t1 a_941_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_465_369.t0 a_299_47.t3 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND.t7 GATE_N.t1 a_27_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 327.644
R1 D.n0 D.t1 157.338
R2 D D.n0 154.595
R3 a_299_47.t1 a_299_47.n1 435.498
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t0 273.433
R6 a_299_47.n1 a_299_47.n0 156.268
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n11 VPWR.t5 871.352
R9 VPWR.n5 VPWR.t1 685.12
R10 VPWR.n23 VPWR.n1 604.394
R11 VPWR.n7 VPWR.t4 410.932
R12 VPWR.n3 VPWR.n2 311.356
R13 VPWR.n9 VPWR.n8 307.866
R14 VPWR.n1 VPWR.t7 41.5552
R15 VPWR.n1 VPWR.t8 41.5552
R16 VPWR.n2 VPWR.t3 41.5552
R17 VPWR.n2 VPWR.t0 41.5552
R18 VPWR.n22 VPWR.n21 34.6358
R19 VPWR.n16 VPWR.n15 34.6358
R20 VPWR.n17 VPWR.n16 34.6358
R21 VPWR.n8 VPWR.t2 32.5055
R22 VPWR.n8 VPWR.t6 32.5055
R23 VPWR.n15 VPWR.n5 26.3534
R24 VPWR.n21 VPWR.n3 25.977
R25 VPWR.n23 VPWR.n22 22.9652
R26 VPWR.n11 VPWR.n10 20.3299
R27 VPWR.n17 VPWR.n3 19.577
R28 VPWR.n10 VPWR.n9 19.577
R29 VPWR.n11 VPWR.n5 12.8005
R30 VPWR.n10 VPWR.n6 9.3005
R31 VPWR.n12 VPWR.n11 9.3005
R32 VPWR.n13 VPWR.n5 9.3005
R33 VPWR.n15 VPWR.n14 9.3005
R34 VPWR.n16 VPWR.n4 9.3005
R35 VPWR.n18 VPWR.n17 9.3005
R36 VPWR.n19 VPWR.n3 9.3005
R37 VPWR.n21 VPWR.n20 9.3005
R38 VPWR.n22 VPWR.n0 9.3005
R39 VPWR.n24 VPWR.n23 7.12063
R40 VPWR.n9 VPWR.n7 6.56061
R41 VPWR.n7 VPWR.n6 0.621726
R42 VPWR.n24 VPWR.n0 0.148519
R43 VPWR.n12 VPWR.n6 0.120292
R44 VPWR.n13 VPWR.n12 0.120292
R45 VPWR.n14 VPWR.n13 0.120292
R46 VPWR.n14 VPWR.n4 0.120292
R47 VPWR.n18 VPWR.n4 0.120292
R48 VPWR.n19 VPWR.n18 0.120292
R49 VPWR.n20 VPWR.n19 0.120292
R50 VPWR.n20 VPWR.n0 0.120292
R51 VPWR VPWR.n24 0.0927068
R52 VPB.t2 VPB.t6 583.023
R53 VPB.t9 VPB.t0 556.386
R54 VPB.t7 VPB.t3 284.113
R55 VPB.t8 VPB.t2 284.113
R56 VPB.t4 VPB.t1 284.113
R57 VPB.t3 VPB.t5 269.315
R58 VPB.t6 VPB.t7 248.599
R59 VPB.t1 VPB.t8 248.599
R60 VPB.t0 VPB.t4 248.599
R61 VPB.t10 VPB.t9 248.599
R62 VPB VPB.t10 139.097
R63 a_27_47.t0 a_27_47.n3 415.863
R64 a_27_47.n2 a_27_47.t2 315.678
R65 a_27_47.n2 a_27_47.t3 308.158
R66 a_27_47.n1 a_27_47.t1 294.873
R67 a_27_47.n0 a_27_47.t5 263.173
R68 a_27_47.n0 a_27_47.t4 227.826
R69 a_27_47.n1 a_27_47.n0 152
R70 a_27_47.n3 a_27_47.n2 20.5706
R71 a_27_47.n3 a_27_47.n1 18.9713
R72 a_465_47.n0 a_465_47.t1 66.6672
R73 a_465_47.n0 a_465_47.t0 26.3935
R74 a_465_47.n1 a_465_47.n0 14.4005
R75 a_560_47.n3 a_560_47.n2 754.694
R76 a_560_47.n2 a_560_47.n1 281.12
R77 a_560_47.n0 a_560_47.t4 268.313
R78 a_560_47.n2 a_560_47.n0 252.797
R79 a_560_47.n0 a_560_47.t5 151.206
R80 a_560_47.n3 a_560_47.t2 63.3219
R81 a_560_47.t0 a_560_47.n3 63.3219
R82 a_560_47.n1 a_560_47.t3 60.0005
R83 a_560_47.n1 a_560_47.t1 53.3338
R84 VNB.t6 VNB.t2 2677.02
R85 VNB.t8 VNB.t0 2677.02
R86 VNB.t7 VNB.t3 1423.95
R87 VNB.t9 VNB.t1 1395.47
R88 VNB.t1 VNB.t6 1352.75
R89 VNB.t5 VNB.t9 1352.75
R90 VNB.t3 VNB.t4 1196.12
R91 VNB.t2 VNB.t7 1196.12
R92 VNB.t0 VNB.t5 1196.12
R93 VNB.t10 VNB.t8 1196.12
R94 VNB VNB.t10 669.256
R95 a_645_413.t0 a_645_413.t1 154.786
R96 a_711_307.n4 a_711_307.t5 366.002
R97 a_711_307.n6 a_711_307.n5 299.166
R98 a_711_307.n3 a_711_307.t0 224.123
R99 a_711_307.n2 a_711_307.t4 214.272
R100 a_711_307.n0 a_711_307.t6 212.081
R101 a_711_307.n5 a_711_307.n4 186.91
R102 a_711_307.n3 a_711_307.n2 152
R103 a_711_307.n4 a_711_307.t3 147.495
R104 a_711_307.n0 a_711_307.t8 139.78
R105 a_711_307.n1 a_711_307.t7 139.78
R106 a_711_307.n5 a_711_307.n3 71.1375
R107 a_711_307.n1 a_711_307.n0 61.346
R108 a_711_307.n6 a_711_307.t2 26.5955
R109 a_711_307.t1 a_711_307.n6 26.5955
R110 a_711_307.n2 a_711_307.n1 2.92171
R111 VGND.n6 VGND.t2 293.767
R112 VGND.n4 VGND.t4 240.575
R113 VGND.n23 VGND.n22 199.739
R114 VGND.n8 VGND.n7 198.964
R115 VGND.n2 VGND.n1 198.964
R116 VGND.n7 VGND.t3 39.6928
R117 VGND.n1 VGND.t1 38.5719
R118 VGND.n1 VGND.t0 38.5719
R119 VGND.n22 VGND.t6 38.5719
R120 VGND.n22 VGND.t7 38.5719
R121 VGND.n10 VGND.n9 34.6358
R122 VGND.n15 VGND.n14 34.6358
R123 VGND.n16 VGND.n15 34.6358
R124 VGND.n21 VGND.n20 34.6358
R125 VGND.n7 VGND.t5 24.9236
R126 VGND.n16 VGND.n2 24.4711
R127 VGND.n23 VGND.n21 22.9652
R128 VGND.n10 VGND.n4 22.5887
R129 VGND.n14 VGND.n4 21.4593
R130 VGND.n9 VGND.n8 19.9534
R131 VGND.n20 VGND.n2 19.9534
R132 VGND.n9 VGND.n5 9.3005
R133 VGND.n11 VGND.n10 9.3005
R134 VGND.n12 VGND.n4 9.3005
R135 VGND.n14 VGND.n13 9.3005
R136 VGND.n15 VGND.n3 9.3005
R137 VGND.n17 VGND.n16 9.3005
R138 VGND.n18 VGND.n2 9.3005
R139 VGND.n20 VGND.n19 9.3005
R140 VGND.n21 VGND.n0 9.3005
R141 VGND.n24 VGND.n23 7.12063
R142 VGND.n8 VGND.n6 6.73566
R143 VGND.n6 VGND.n5 0.589728
R144 VGND.n24 VGND.n0 0.148519
R145 VGND.n11 VGND.n5 0.120292
R146 VGND.n12 VGND.n11 0.120292
R147 VGND.n13 VGND.n12 0.120292
R148 VGND.n13 VGND.n3 0.120292
R149 VGND.n17 VGND.n3 0.120292
R150 VGND.n18 VGND.n17 0.120292
R151 VGND.n19 VGND.n18 0.120292
R152 VGND.n19 VGND.n0 0.120292
R153 VGND VGND.n24 0.0927068
R154 RESET_B.n0 RESET_B.t0 241.536
R155 RESET_B.n0 RESET_B.t1 169.237
R156 RESET_B RESET_B.n0 162.862
R157 a_193_47.n0 a_193_47.t3 462.721
R158 a_193_47.t0 a_193_47.n1 366.837
R159 a_193_47.n1 a_193_47.t1 322.567
R160 a_193_47.n0 a_193_47.t2 242.607
R161 a_193_47.n1 a_193_47.n0 187.469
R162 a_465_369.t0 a_465_369.t1 134.631
R163 GATE_N.n0 GATE_N.t0 269.921
R164 GATE_N.n0 GATE_N.t1 234.573
R165 GATE_N.n1 GATE_N.n0 152
R166 GATE_N GATE_N.n1 10.9719
R167 GATE_N.n1 GATE_N 6.79234
R168 Q Q.n2 593.297
R169 Q.n1 Q.n0 239.091
R170 Q.n2 Q.t0 30.5355
R171 Q.n2 Q.t1 29.5505
R172 Q.n0 Q.t2 24.9236
R173 Q.n0 Q.t3 24.9236
R174 Q.n1 Q 9.6005
R175 Q.n3 Q 4.82857
R176 Q Q.n3 2.80752
R177 Q.n1 Q 2.18853
R178 Q.n3 Q.n1 0.547509
R179 a_658_47.t1 a_658_47.t0 93.0601
R180 a_941_47.t0 a_941_47.t1 49.8467
C0 VPB D 0.062355f
C1 VPB RESET_B 0.027237f
C2 VPB VPWR 0.151945f
C3 VPB VGND 0.013535f
C4 GATE_N VPWR 0.019242f
C5 GATE_N VGND 0.019085f
C6 D VPWR 0.014067f
C7 VPB Q 0.006968f
C8 D VGND 0.018848f
C9 RESET_B VPWR 0.022024f
C10 RESET_B VGND 0.018162f
C11 RESET_B Q 0.001136f
C12 VPWR VGND 0.082133f
C13 VPWR Q 0.186248f
C14 VGND Q 0.130452f
C15 VPB GATE_N 0.070092f
C16 Q VNB 0.047486f
C17 VGND VNB 0.756611f
C18 VPWR VNB 0.619563f
C19 RESET_B VNB 0.091055f
C20 D VNB 0.132265f
C21 GATE_N VNB 0.195771f
C22 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbn_2 VNB VPB VPWR VGND D GATE_N Q RESET_B Q_N
X0 VPWR.t1 D.t0 a_299_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_465_47.t1 a_299_47.t2 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_561_413.t1 a_27_47.t2 a_465_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X3 Q_N.t0 a_1313_47# VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.149 ps=1.325 w=1 l=0.15
X4 Q_N.t1 a_1313_47# VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.097 ps=0.975 w=0.65 l=0.15
X5 a_561_413.t3 a_193_47.t2 a_465_369.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X6 a_724_21.t1 a_561_413.t4 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t8 a_724_21.t3 a_659_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8 VPWR.t5 GATE_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 VPWR a_1313_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X10 a_659_47.t0 a_193_47.t3 a_561_413.t2 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X11 VPWR.t9 a_724_21.t4 a_682_413.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 VGND a_1313_47# Q_N VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.089375 ps=0.925 w=0.65 l=0.15
X13 a_193_47.t1 a_27_47.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_682_413.t0 a_27_47.t4 a_561_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X15 Q.t3 a_724_21.t5 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_942_47.t1 a_561_413.t5 a_724_21.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VPWR.t7 a_724_21.t6 Q.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X18 a_193_47.t0 a_27_47.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 Q.t0 a_724_21.t7 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t2 RESET_B.t0 a_724_21.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND.t1 D.t1 a_299_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X22 VGND.t2 RESET_B.t1 a_942_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VGND.t6 a_724_21.t8 Q.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.105625 ps=0.975 w=0.65 l=0.15
X24 a_465_369.t1 a_299_47.t3 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 VGND.t5 GATE_N.t1 a_27_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 327.644
R1 D.n0 D.t1 157.338
R2 D D.n0 154.595
R3 a_299_47.t1 a_299_47.n1 438.971
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t0 275.149
R6 a_299_47.n1 a_299_47.n0 156.462
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n16 VPWR.t6 853.981
R9 VPWR.n5 VPWR.t9 648.322
R10 VPWR.n29 VPWR.n1 604.394
R11 VPWR.n9 VPWR.t3 349.832
R12 VPWR.n10 VPWR.t7 343.057
R13 VPWR.n8 VPWR.n7 315.221
R14 VPWR.n3 VPWR.n2 311.356
R15 VPWR.n1 VPWR.t0 41.5552
R16 VPWR.n1 VPWR.t5 41.5552
R17 VPWR.n2 VPWR.t4 41.5552
R18 VPWR.n2 VPWR.t1 41.5552
R19 VPWR.n28 VPWR.n27 34.6358
R20 VPWR.n22 VPWR.n21 34.6358
R21 VPWR.n23 VPWR.n22 34.6358
R22 VPWR.n11 VPWR.n8 30.1181
R23 VPWR.n21 VPWR.n5 29.4832
R24 VPWR.n7 VPWR.t8 26.5955
R25 VPWR.n7 VPWR.t2 26.5955
R26 VPWR.n27 VPWR.n3 25.977
R27 VPWR.n11 VPWR.n10 25.224
R28 VPWR.n29 VPWR.n28 22.9652
R29 VPWR.n16 VPWR.n15 21.2233
R30 VPWR.n15 VPWR.n8 20.3299
R31 VPWR.n23 VPWR.n3 19.577
R32 VPWR.n12 VPWR.n11 9.3005
R33 VPWR.n13 VPWR.n8 9.3005
R34 VPWR.n15 VPWR.n14 9.3005
R35 VPWR.n17 VPWR.n6 9.3005
R36 VPWR.n19 VPWR.n18 9.3005
R37 VPWR.n21 VPWR.n20 9.3005
R38 VPWR.n22 VPWR.n4 9.3005
R39 VPWR.n24 VPWR.n23 9.3005
R40 VPWR.n25 VPWR.n3 9.3005
R41 VPWR.n27 VPWR.n26 9.3005
R42 VPWR.n28 VPWR.n0 9.3005
R43 VPWR.n18 VPWR.n17 8.78856
R44 VPWR.n30 VPWR.n29 7.12063
R45 VPWR.n10 VPWR.n9 6.79261
R46 VPWR.n17 VPWR.n16 1.05125
R47 VPWR.n12 VPWR.n9 0.49177
R48 VPWR.n30 VPWR.n0 0.148519
R49 VPWR.n13 VPWR.n12 0.120292
R50 VPWR.n14 VPWR.n13 0.120292
R51 VPWR.n14 VPWR.n6 0.120292
R52 VPWR.n19 VPWR.n6 0.120292
R53 VPWR.n20 VPWR.n19 0.120292
R54 VPWR.n20 VPWR.n4 0.120292
R55 VPWR.n24 VPWR.n4 0.120292
R56 VPWR.n25 VPWR.n24 0.120292
R57 VPWR.n26 VPWR.n25 0.120292
R58 VPWR.n26 VPWR.n0 0.120292
R59 VPWR VPWR.n30 0.11354
R60 VPWR.n18 VPWR.n5 0.0960224
R61 VPB.t8 VPB.t4 843.458
R62 VPB.t11 VPB.t7 556.386
R63 VPB.t1 VPB.t2 556.386
R64 VPB.t10 VPB.t0 358.101
R65 VPB.t5 VPB.t10 284.113
R66 VPB.t9 VPB.t8 281.154
R67 VPB.t3 VPB.t9 248.599
R68 VPB.t7 VPB.t3 248.599
R69 VPB.t2 VPB.t5 248.599
R70 VPB.t6 VPB.t1 248.599
R71 VPB.t0 VPB.t11 213.084
R72 VPB VPB.t6 189.409
R73 VGND.n7 VGND.t6 283.015
R74 VGND.n4 VGND.t8 240.833
R75 VGND.n8 VGND.t3 232.448
R76 VGND.n28 VGND.n27 199.739
R77 VGND.n2 VGND.n1 198.964
R78 VGND.n13 VGND.n12 185
R79 VGND.n1 VGND.t4 38.5719
R80 VGND.n1 VGND.t1 38.5719
R81 VGND.n27 VGND.t0 38.5719
R82 VGND.n27 VGND.t5 38.5719
R83 VGND.n15 VGND.n14 34.6358
R84 VGND.n20 VGND.n19 34.6358
R85 VGND.n21 VGND.n20 34.6358
R86 VGND.n26 VGND.n25 34.6358
R87 VGND.n7 VGND.n6 25.224
R88 VGND.n12 VGND.t7 24.9236
R89 VGND.n12 VGND.t2 24.9236
R90 VGND.n11 VGND.n6 24.5966
R91 VGND.n21 VGND.n2 24.4711
R92 VGND.n14 VGND.n13 24.0352
R93 VGND.n28 VGND.n26 22.9652
R94 VGND.n15 VGND.n4 22.5887
R95 VGND.n19 VGND.n4 21.8358
R96 VGND.n25 VGND.n2 19.9534
R97 VGND.n26 VGND.n0 9.3005
R98 VGND.n25 VGND.n24 9.3005
R99 VGND.n23 VGND.n2 9.3005
R100 VGND.n22 VGND.n21 9.3005
R101 VGND.n20 VGND.n3 9.3005
R102 VGND.n19 VGND.n18 9.3005
R103 VGND.n17 VGND.n4 9.3005
R104 VGND.n9 VGND.n6 9.3005
R105 VGND.n11 VGND.n10 9.3005
R106 VGND.n14 VGND.n5 9.3005
R107 VGND.n16 VGND.n15 9.3005
R108 VGND.n29 VGND.n28 7.12063
R109 VGND.n8 VGND.n7 6.78446
R110 VGND.n13 VGND.n11 0.561904
R111 VGND.n9 VGND.n8 0.498094
R112 VGND.n29 VGND.n0 0.148519
R113 VGND.n10 VGND.n9 0.120292
R114 VGND.n10 VGND.n5 0.120292
R115 VGND.n16 VGND.n5 0.120292
R116 VGND.n17 VGND.n16 0.120292
R117 VGND.n18 VGND.n17 0.120292
R118 VGND.n18 VGND.n3 0.120292
R119 VGND.n22 VGND.n3 0.120292
R120 VGND.n23 VGND.n22 0.120292
R121 VGND.n24 VGND.n23 0.120292
R122 VGND.n24 VGND.n0 0.120292
R123 VGND VGND.n29 0.11354
R124 a_465_47.n0 a_465_47.t0 88.3338
R125 a_465_47.n0 a_465_47.t1 26.3935
R126 a_465_47.n1 a_465_47.n0 14.4005
R127 VNB.t9 VNB.t6 4058.25
R128 VNB.t11 VNB.t3 2677.02
R129 VNB.t1 VNB.t2 2677.02
R130 VNB.t7 VNB.t0 1537.86
R131 VNB.t10 VNB.t9 1352.75
R132 VNB.t5 VNB.t11 1352.75
R133 VNB.t0 VNB.t5 1224.6
R134 VNB.t4 VNB.t10 1196.12
R135 VNB.t3 VNB.t4 1196.12
R136 VNB.t2 VNB.t7 1196.12
R137 VNB.t8 VNB.t1 1196.12
R138 VNB VNB.t8 911.327
R139 a_27_47.t0 a_27_47.n3 410.19
R140 a_27_47.n2 a_27_47.t4 316.111
R141 a_27_47.n2 a_27_47.t2 315.729
R142 a_27_47.n1 a_27_47.t1 288.075
R143 a_27_47.n0 a_27_47.t5 263.173
R144 a_27_47.n0 a_27_47.t3 227.826
R145 a_27_47.n1 a_27_47.n0 152
R146 a_27_47.n3 a_27_47.n2 20.5706
R147 a_27_47.n3 a_27_47.n1 18.4963
R148 a_561_413.n3 a_561_413.n2 714.672
R149 a_561_413.n2 a_561_413.n1 282.507
R150 a_561_413.n2 a_561_413.n0 248.657
R151 a_561_413.n0 a_561_413.t4 212.081
R152 a_561_413.n0 a_561_413.t5 139.78
R153 a_561_413.n3 a_561_413.t3 121.953
R154 a_561_413.t0 a_561_413.n3 91.4648
R155 a_561_413.n1 a_561_413.t2 46.6672
R156 a_561_413.n1 a_561_413.t1 46.6672
R157 Q_N.n2 Q_N.t0 350.031
R158 Q_N.n0 Q_N.t1 209.923
R159 Q_N.n1 Q_N.n0 27.3215
R160 Q_N Q_N.n1 24.3815
R161 Q_N.n1 Q_N 15.882
R162 Q_N.n2 Q_N 9.28312
R163 Q_N Q_N.n2 7.62171
R164 Q_N.n0 Q_N 6.77697
R165 a_193_47.n0 a_193_47.t3 464.327
R166 a_193_47.t0 a_193_47.n1 366.837
R167 a_193_47.n1 a_193_47.t1 322.567
R168 a_193_47.n0 a_193_47.t2 242.607
R169 a_193_47.n1 a_193_47.n0 187.469
R170 a_465_369.t1 a_465_369.t0 134.631
R171 a_724_21.n7 a_724_21.t3 368.329
R172 a_724_21.n6 a_724_21.t2 301.716
R173 a_724_21.n9 a_724_21.n8 299.93
R174 a_724_21.n2 a_724_21.n0 247.542
R175 a_724_21.n3 a_724_21.t6 212.081
R176 a_724_21.n4 a_724_21.t7 212.081
R177 a_724_21.n8 a_724_21.n7 183.827
R178 a_724_21.n2 a_724_21.n1 154.356
R179 a_724_21.n6 a_724_21.n5 152
R180 a_724_21.n7 a_724_21.t4 149.822
R181 a_724_21.n3 a_724_21.t8 139.78
R182 a_724_21.n4 a_724_21.t5 139.78
R183 a_724_21.n3 a_724_21.n2 119.77
R184 a_724_21.n5 a_724_21.n3 60.6157
R185 a_724_21.n8 a_724_21.n6 57.5657
R186 a_724_21.t0 a_724_21.n9 26.5955
R187 a_724_21.n9 a_724_21.t1 26.5955
R188 a_724_21.n5 a_724_21.n4 8.76414
R189 a_659_47.t1 a_659_47.t0 93.0601
R190 GATE_N.n0 GATE_N.t0 269.921
R191 GATE_N.n0 GATE_N.t1 234.573
R192 GATE_N.n1 GATE_N.n0 152
R193 GATE_N GATE_N.n1 10.9719
R194 GATE_N.n1 GATE_N 6.79234
R195 a_682_413.t0 a_682_413.t1 98.5005
R196 Q.n0 Q 593.453
R197 Q.n1 Q.n0 585
R198 Q.n3 Q.n2 185
R199 Q Q.n1 37.7358
R200 Q.n0 Q.t0 36.4455
R201 Q.n2 Q.t3 34.1543
R202 Q.n0 Q.t1 27.5805
R203 Q.n2 Q.t2 25.8467
R204 Q Q.n3 19.1068
R205 Q.n1 Q 7.97031
R206 Q.n3 Q 7.63127
R207 a_942_47.t0 a_942_47.t1 49.8467
R208 RESET_B.n0 RESET_B.t0 241.536
R209 RESET_B.n0 RESET_B.t1 169.237
R210 RESET_B RESET_B.n0 162.28
C0 a_1313_47# VPB 0.079175f
C1 VPB GATE_N 0.069289f
C2 VGND Q_N 0.145594f
C3 VPB D 0.062359f
C4 VPB RESET_B 0.02634f
C5 VPB VPWR 0.197551f
C6 a_1313_47# VPWR 0.216142f
C7 GATE_N VPWR 0.017119f
C8 VPB VGND 0.01826f
C9 a_1313_47# VGND 0.160021f
C10 GATE_N VGND 0.016722f
C11 VPB Q 0.006988f
C12 D VPWR 0.014067f
C13 a_1313_47# Q 0.06653f
C14 RESET_B VPWR 0.022084f
C15 D VGND 0.018848f
C16 VPB Q_N 0.007371f
C17 a_1313_47# Q_N 0.124109f
C18 RESET_B VGND 0.018675f
C19 RESET_B Q 8.3e-19
C20 VPWR VGND 0.124166f
C21 VPWR Q 0.154624f
C22 VGND Q 0.078035f
C23 VPWR Q_N 0.20168f
C24 Q_N VNB 0.032932f
C25 Q VNB 0.010393f
C26 VGND VNB 0.964845f
C27 VPWR VNB 0.779022f
C28 RESET_B VNB 0.089508f
C29 D VNB 0.132433f
C30 GATE_N VNB 0.19496f
C31 VPB VNB 1.66792f
C32 a_1313_47# VNB 0.22538f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbp_2 VGND VPWR VPB VNB Q RESET_B Q_N D GATE
X0 VPWR.t11 D.t0 a_299_47.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 Q_N.t1 a_1316_47.t2 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2 a_645_413.t0 a_193_47.t2 a_561_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR.t0 a_711_307.t3 a_645_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_465_47.t1 a_299_47.t2 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_561_413.t1 a_193_47.t3 a_465_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X6 VGND.t1 a_711_307.t4 a_1316_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR.t1 a_711_307.t5 a_1316_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_561_413.t2 a_27_47.t2 a_465_369.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0968 ps=0.97 w=0.42 l=0.15
X9 a_711_307.t2 a_561_413.t4 VPWR.t8 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND.t2 a_711_307.t6 a_659_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11 VPWR.t4 GATE.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12 VPWR.t6 RESET_B.t0 a_711_307.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND.t3 a_711_307.t7 Q.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.09425 ps=0.94 w=0.65 l=0.15
X14 a_659_47.t1 a_27_47.t3 a_561_413.t3 VNB.t13 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X15 VGND.t5 a_1316_47.t3 Q_N.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_193_47.t0 a_27_47.t4 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR.t9 a_711_307.t8 Q.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.145 ps=1.29 w=1 l=0.15
X18 VPWR.t3 a_1316_47.t4 Q_N.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 a_942_47.t1 a_561_413.t5 a_711_307.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X20 Q.t0 a_711_307.t9 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.104 ps=0.97 w=0.65 l=0.15
X21 Q_N.t2 a_1316_47.t5 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X22 a_193_47.t1 a_27_47.t5 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND.t10 RESET_B.t1 a_942_47.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VGND.t9 D.t1 a_299_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 Q.t2 a_711_307.t10 VPWR.t10 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.16 ps=1.32 w=1 l=0.15
X26 a_465_369.t0 a_299_47.t3 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 VGND.t0 GATE.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 327.644
R1 D.n0 D.t1 157.338
R2 D D.n0 154.595
R3 a_299_47.t0 a_299_47.n1 438.971
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t1 275.149
R6 a_299_47.n1 a_299_47.n0 156.462
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n21 VPWR.t8 853.981
R9 VPWR.n5 VPWR.t0 648.322
R10 VPWR.n34 VPWR.n1 604.394
R11 VPWR.n15 VPWR.t9 341.93
R12 VPWR.n11 VPWR.n10 312.632
R13 VPWR.n3 VPWR.n2 311.356
R14 VPWR.n8 VPWR.n7 307.464
R15 VPWR.n12 VPWR.t3 256.253
R16 VPWR.n10 VPWR.t1 56.9458
R17 VPWR.n1 VPWR.t5 41.5552
R18 VPWR.n1 VPWR.t4 41.5552
R19 VPWR.n2 VPWR.t7 41.5552
R20 VPWR.n2 VPWR.t11 41.5552
R21 VPWR.n7 VPWR.t10 36.4455
R22 VPWR.n33 VPWR.n32 34.6358
R23 VPWR.n27 VPWR.n26 34.6358
R24 VPWR.n28 VPWR.n27 34.6358
R25 VPWR.n10 VPWR.t2 33.1448
R26 VPWR.n14 VPWR.n11 28.2358
R27 VPWR.n7 VPWR.t6 26.5955
R28 VPWR.n16 VPWR.n15 26.3534
R29 VPWR.n32 VPWR.n3 25.977
R30 VPWR.n26 VPWR.n5 24.5891
R31 VPWR.n15 VPWR.n14 23.3417
R32 VPWR.n34 VPWR.n33 22.9652
R33 VPWR.n20 VPWR.n8 21.0829
R34 VPWR.n21 VPWR.n20 20.6614
R35 VPWR.n28 VPWR.n3 19.577
R36 VPWR.n16 VPWR.n8 19.577
R37 VPWR.n14 VPWR.n13 9.3005
R38 VPWR.n15 VPWR.n9 9.3005
R39 VPWR.n17 VPWR.n16 9.3005
R40 VPWR.n18 VPWR.n8 9.3005
R41 VPWR.n20 VPWR.n19 9.3005
R42 VPWR.n22 VPWR.n6 9.3005
R43 VPWR.n24 VPWR.n23 9.3005
R44 VPWR.n26 VPWR.n25 9.3005
R45 VPWR.n27 VPWR.n4 9.3005
R46 VPWR.n29 VPWR.n28 9.3005
R47 VPWR.n30 VPWR.n3 9.3005
R48 VPWR.n32 VPWR.n31 9.3005
R49 VPWR.n33 VPWR.n0 9.3005
R50 VPWR.n23 VPWR.n22 8.78856
R51 VPWR.n35 VPWR.n34 7.12063
R52 VPWR.n12 VPWR.n11 6.32884
R53 VPWR.n23 VPWR.n5 1.33781
R54 VPWR.n22 VPWR.n21 1.05125
R55 VPWR.n13 VPWR.n12 0.664094
R56 VPWR.n35 VPWR.n0 0.148519
R57 VPWR.n13 VPWR.n9 0.120292
R58 VPWR.n17 VPWR.n9 0.120292
R59 VPWR.n18 VPWR.n17 0.120292
R60 VPWR.n19 VPWR.n18 0.120292
R61 VPWR.n19 VPWR.n6 0.120292
R62 VPWR.n24 VPWR.n6 0.120292
R63 VPWR.n25 VPWR.n24 0.120292
R64 VPWR.n25 VPWR.n4 0.120292
R65 VPWR.n29 VPWR.n4 0.120292
R66 VPWR.n30 VPWR.n29 0.120292
R67 VPWR.n31 VPWR.n30 0.120292
R68 VPWR.n31 VPWR.n0 0.120292
R69 VPWR VPWR.n35 0.11354
R70 VPB.t1 VPB.t9 594.861
R71 VPB.t10 VPB.t2 556.386
R72 VPB.t6 VPB.t12 556.386
R73 VPB.t0 VPB.t1 284.113
R74 VPB.t8 VPB.t13 284.113
R75 VPB.t2 VPB.t3 281.154
R76 VPB.t7 VPB.t11 278.193
R77 VPB.t11 VPB.t10 260.437
R78 VPB.t9 VPB.t7 254.518
R79 VPB.t3 VPB.t4 248.599
R80 VPB.t13 VPB.t0 248.599
R81 VPB.t12 VPB.t8 248.599
R82 VPB.t5 VPB.t6 248.599
R83 VPB VPB.t5 139.097
R84 a_1316_47.t1 a_1316_47.n2 392.175
R85 a_1316_47.n0 a_1316_47.t5 300.447
R86 a_1316_47.n2 a_1316_47.t0 248.689
R87 a_1316_47.n0 a_1316_47.t2 228.148
R88 a_1316_47.n1 a_1316_47.t4 221.72
R89 a_1316_47.n2 a_1316_47.n0 170.231
R90 a_1316_47.n1 a_1316_47.t3 149.421
R91 a_1316_47.n0 a_1316_47.n1 84.7968
R92 VGND.n12 VGND.t3 282.384
R93 VGND.n4 VGND.t2 240.833
R94 VGND.n10 VGND.n9 200.948
R95 VGND.n33 VGND.n32 199.739
R96 VGND.n2 VGND.n1 198.964
R97 VGND.n18 VGND.n17 185
R98 VGND.n8 VGND.t5 161.489
R99 VGND.n9 VGND.t1 52.8576
R100 VGND.n1 VGND.t7 38.5719
R101 VGND.n1 VGND.t9 38.5719
R102 VGND.n32 VGND.t4 38.5719
R103 VGND.n32 VGND.t0 38.5719
R104 VGND.n20 VGND.n19 34.6358
R105 VGND.n25 VGND.n24 34.6358
R106 VGND.n26 VGND.n25 34.6358
R107 VGND.n31 VGND.n30 34.6358
R108 VGND.n17 VGND.t8 34.1543
R109 VGND.n11 VGND.n10 27.4829
R110 VGND.n9 VGND.t6 27.3631
R111 VGND.n17 VGND.t10 24.9236
R112 VGND.n19 VGND.n18 24.7881
R113 VGND.n26 VGND.n2 24.4711
R114 VGND.n16 VGND.n6 24.0682
R115 VGND.n12 VGND.n11 23.3417
R116 VGND.n33 VGND.n31 22.9652
R117 VGND.n20 VGND.n4 22.5887
R118 VGND.n24 VGND.n4 21.8358
R119 VGND.n12 VGND.n6 20.3299
R120 VGND.n30 VGND.n2 19.9534
R121 VGND.n31 VGND.n0 9.3005
R122 VGND.n30 VGND.n29 9.3005
R123 VGND.n28 VGND.n2 9.3005
R124 VGND.n27 VGND.n26 9.3005
R125 VGND.n25 VGND.n3 9.3005
R126 VGND.n24 VGND.n23 9.3005
R127 VGND.n22 VGND.n4 9.3005
R128 VGND.n21 VGND.n20 9.3005
R129 VGND.n19 VGND.n5 9.3005
R130 VGND.n16 VGND.n15 9.3005
R131 VGND.n14 VGND.n6 9.3005
R132 VGND.n13 VGND.n12 9.3005
R133 VGND.n11 VGND.n7 9.3005
R134 VGND.n34 VGND.n33 7.12063
R135 VGND.n10 VGND.n8 6.32884
R136 VGND.n8 VGND.n7 0.664094
R137 VGND.n18 VGND.n16 0.337342
R138 VGND.n34 VGND.n0 0.148519
R139 VGND.n13 VGND.n7 0.120292
R140 VGND.n14 VGND.n13 0.120292
R141 VGND.n15 VGND.n14 0.120292
R142 VGND.n15 VGND.n5 0.120292
R143 VGND.n21 VGND.n5 0.120292
R144 VGND.n22 VGND.n21 0.120292
R145 VGND.n23 VGND.n22 0.120292
R146 VGND.n23 VGND.n3 0.120292
R147 VGND.n27 VGND.n3 0.120292
R148 VGND.n28 VGND.n27 0.120292
R149 VGND.n29 VGND.n28 0.120292
R150 VGND.n29 VGND.n0 0.120292
R151 VGND VGND.n34 0.11354
R152 Q_N Q_N.n0 586.793
R153 Q_N.n4 Q_N.n0 585
R154 Q_N.n2 Q_N.n1 185
R155 Q_N.n3 Q_N.n2 30.8861
R156 Q_N Q_N.n3 30.2989
R157 Q_N.n0 Q_N.t3 26.5955
R158 Q_N.n0 Q_N.t2 26.5955
R159 Q_N.n1 Q_N.t0 24.9236
R160 Q_N.n1 Q_N.t1 24.9236
R161 Q_N Q_N.n4 15.6165
R162 Q_N.n3 Q_N 14.9338
R163 Q_N.n2 Q_N 6.9125
R164 Q_N.n4 Q_N 1.7925
R165 VNB.t4 VNB.t2 2677.02
R166 VNB.t3 VNB.t9 2677.02
R167 VNB.t5 VNB.t11 2677.02
R168 VNB.t8 VNB.t0 1537.86
R169 VNB.t2 VNB.t7 1352.75
R170 VNB.t13 VNB.t3 1352.75
R171 VNB.t12 VNB.t10 1338.51
R172 VNB.t10 VNB.t4 1253.07
R173 VNB.t9 VNB.t12 1224.6
R174 VNB.t0 VNB.t13 1224.6
R175 VNB.t7 VNB.t6 1196.12
R176 VNB.t11 VNB.t8 1196.12
R177 VNB.t1 VNB.t5 1196.12
R178 VNB VNB.t1 669.256
R179 a_193_47.t1 a_193_47.n1 366.837
R180 a_193_47.n0 a_193_47.t3 329.659
R181 a_193_47.n1 a_193_47.t0 322.567
R182 a_193_47.n0 a_193_47.t2 300.252
R183 a_193_47.n1 a_193_47.n0 25.054
R184 a_561_413.n3 a_561_413.n2 699.951
R185 a_561_413.n2 a_561_413.n1 280.625
R186 a_561_413.n2 a_561_413.n0 250.541
R187 a_561_413.n0 a_561_413.t4 212.081
R188 a_561_413.n0 a_561_413.t5 139.78
R189 a_561_413.t0 a_561_413.n3 63.3219
R190 a_561_413.n3 a_561_413.t2 63.3219
R191 a_561_413.n1 a_561_413.t3 46.6672
R192 a_561_413.n1 a_561_413.t1 46.6672
R193 a_645_413.t0 a_645_413.t1 154.786
R194 a_711_307.n4 a_711_307.t6 366.002
R195 a_711_307.n6 a_711_307.n5 299.93
R196 a_711_307.n3 a_711_307.t1 297.44
R197 a_711_307.n0 a_711_307.t5 269.921
R198 a_711_307.n2 a_711_307.t10 212.081
R199 a_711_307.n1 a_711_307.t8 212.081
R200 a_711_307.n5 a_711_307.n4 188.073
R201 a_711_307.n0 a_711_307.t4 176.733
R202 a_711_307.n3 a_711_307.n2 152
R203 a_711_307.n4 a_711_307.t3 147.495
R204 a_711_307.n2 a_711_307.t9 139.78
R205 a_711_307.n1 a_711_307.t7 139.78
R206 a_711_307.n1 a_711_307.n0 137.298
R207 a_711_307.n2 a_711_307.n1 64.2672
R208 a_711_307.n5 a_711_307.n3 58.8229
R209 a_711_307.n6 a_711_307.t2 28.5655
R210 a_711_307.t0 a_711_307.n6 26.5955
R211 a_465_47.n0 a_465_47.t0 88.3338
R212 a_465_47.n0 a_465_47.t1 26.3935
R213 a_465_47.n1 a_465_47.n0 14.4005
R214 a_27_47.n2 a_27_47.t3 464.327
R215 a_27_47.t1 a_27_47.n3 411.32
R216 a_27_47.n1 a_27_47.t0 289.399
R217 a_27_47.n0 a_27_47.t5 263.173
R218 a_27_47.n2 a_27_47.t2 242.607
R219 a_27_47.n0 a_27_47.t4 227.826
R220 a_27_47.n3 a_27_47.n2 176.62
R221 a_27_47.n1 a_27_47.n0 152
R222 a_27_47.n3 a_27_47.n1 18.9713
R223 a_465_369.t0 a_465_369.t1 134.631
R224 a_659_47.t0 a_659_47.t1 93.0601
R225 GATE.n0 GATE.t0 269.921
R226 GATE.n0 GATE.t1 234.573
R227 GATE.n1 GATE.n0 152
R228 GATE GATE.n1 10.9719
R229 GATE.n1 GATE 6.79234
R230 RESET_B.n0 RESET_B.t0 241.536
R231 RESET_B.n0 RESET_B.t1 169.237
R232 RESET_B RESET_B.n0 161.892
R233 Q.n0 Q 593.961
R234 Q.n1 Q.n0 585
R235 Q.n3 Q.n2 185
R236 Q Q.n1 33.6993
R237 Q.n0 Q.t2 30.5355
R238 Q.n2 Q.t0 28.6159
R239 Q Q.n3 28.5539
R240 Q.n0 Q.t3 26.5955
R241 Q.n2 Q.t1 24.9236
R242 Q.n3 Q 11.6711
R243 Q.n1 Q 8.4485
R244 a_942_47.t0 a_942_47.t1 51.6928
C0 VPWR Q 0.161686f
C1 VPWR Q_N 0.198775f
C2 VGND Q 0.086355f
C3 VPB GATE 0.069313f
C4 VGND Q_N 0.143042f
C5 VPB D 0.062359f
C6 VPB RESET_B 0.027283f
C7 VPB VPWR 0.196624f
C8 VPB VGND 0.018879f
C9 GATE VPWR 0.017119f
C10 GATE VGND 0.016722f
C11 D VPWR 0.014067f
C12 VPB Q 0.006615f
C13 VPB Q_N 0.006804f
C14 RESET_B VPWR 0.022129f
C15 D VGND 0.018848f
C16 RESET_B VGND 0.018755f
C17 VPWR VGND 0.123907f
C18 RESET_B Q 7.19e-19
C19 Q_N VNB 0.032678f
C20 Q VNB 0.011117f
C21 VGND VNB 0.960417f
C22 VPWR VNB 0.777038f
C23 RESET_B VNB 0.090182f
C24 D VNB 0.132433f
C25 GATE VNB 0.194986f
C26 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_4 VPWR VGND VPB VNB Q RESET_B D GATE_N
X0 VPWR.t3 RESET_B.t0 a_725_21.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_466_47.t1 a_300_47.t2 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_562_413.t1 a_27_47.t2 a_466_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X3 VGND.t6 a_725_21.t3 a_660_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4 VGND.t8 a_725_21.t4 Q.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.099125 ps=0.955 w=0.65 l=0.15
X5 a_466_369.t1 a_300_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 VPWR.t2 GATE_N.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 VPWR.t4 D.t0 a_300_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 VPWR.t6 a_725_21.t5 Q.t5 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.1525 ps=1.305 w=1 l=0.15
X9 VGND.t7 a_725_21.t6 Q.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X10 a_562_413.t0 a_193_47.t2 a_466_369.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X11 a_725_21.t2 a_562_413.t4 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47.t0 a_27_47.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VPWR.t7 a_725_21.t7 a_683_413.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 a_943_47.t0 a_562_413.t5 a_725_21.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 Q.t4 a_725_21.t8 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1425 ps=1.285 w=1 l=0.15
X16 a_683_413.t0 a_27_47.t4 a_562_413.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X17 a_193_47.t1 a_27_47.t5 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X18 a_660_47.t0 a_193_47.t3 a_562_413.t3 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X19 Q.t0 a_725_21.t9 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.092625 ps=0.935 w=0.65 l=0.15
X20 VGND.t4 D.t1 a_300_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VGND.t2 RESET_B.t1 a_943_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t8 a_725_21.t10 Q.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X23 VGND.t1 GATE_N.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 RESET_B.n0 RESET_B.t0 241.536
R1 RESET_B.n0 RESET_B.t1 169.237
R2 RESET_B RESET_B.n0 162.28
R3 a_725_21.n7 a_725_21.t3 368.329
R4 a_725_21.n9 a_725_21.n8 299.166
R5 a_725_21.n6 a_725_21.t1 231.212
R6 a_725_21.n5 a_725_21.n1 212.081
R7 a_725_21.n2 a_725_21.t10 212.081
R8 a_725_21.n3 a_725_21.t8 212.081
R9 a_725_21.n4 a_725_21.t5 212.081
R10 a_725_21.n8 a_725_21.n7 187.685
R11 a_725_21.n6 a_725_21.n5 152
R12 a_725_21.n7 a_725_21.t7 149.822
R13 a_725_21.n5 a_725_21.n0 139.78
R14 a_725_21.n2 a_725_21.t6 139.78
R15 a_725_21.n3 a_725_21.t9 139.78
R16 a_725_21.n4 a_725_21.t4 139.78
R17 a_725_21.n8 a_725_21.n6 76.7206
R18 a_725_21.n3 a_725_21.n2 67.1884
R19 a_725_21.n5 a_725_21.n4 66.4581
R20 a_725_21.n4 a_725_21.n3 63.5369
R21 a_725_21.t0 a_725_21.n9 26.5955
R22 a_725_21.n9 a_725_21.t2 26.5955
R23 VPWR.n15 VPWR.t5 871.352
R24 VPWR.n5 VPWR.t7 666.86
R25 VPWR.n27 VPWR.n1 604.394
R26 VPWR.n13 VPWR.t3 340.372
R27 VPWR.n3 VPWR.n2 311.356
R28 VPWR.n10 VPWR.t8 250.055
R29 VPWR.n9 VPWR.n8 221.748
R30 VPWR.n1 VPWR.t1 41.5552
R31 VPWR.n1 VPWR.t2 41.5552
R32 VPWR.n2 VPWR.t0 41.5552
R33 VPWR.n2 VPWR.t4 41.5552
R34 VPWR.n26 VPWR.n25 34.6358
R35 VPWR.n20 VPWR.n19 34.6358
R36 VPWR.n21 VPWR.n20 34.6358
R37 VPWR.n8 VPWR.t6 29.5505
R38 VPWR.n12 VPWR.n9 28.9887
R39 VPWR.n19 VPWR.n5 28.2358
R40 VPWR.n8 VPWR.t9 26.5955
R41 VPWR.n25 VPWR.n3 26.3534
R42 VPWR.n27 VPWR.n26 22.9652
R43 VPWR.n14 VPWR.n13 21.4593
R44 VPWR.n13 VPWR.n12 19.9534
R45 VPWR.n21 VPWR.n3 19.2005
R46 VPWR.n15 VPWR.n14 18.4476
R47 VPWR.n15 VPWR.n5 14.3064
R48 VPWR.n12 VPWR.n11 9.3005
R49 VPWR.n13 VPWR.n7 9.3005
R50 VPWR.n14 VPWR.n6 9.3005
R51 VPWR.n16 VPWR.n15 9.3005
R52 VPWR.n17 VPWR.n5 9.3005
R53 VPWR.n19 VPWR.n18 9.3005
R54 VPWR.n20 VPWR.n4 9.3005
R55 VPWR.n22 VPWR.n21 9.3005
R56 VPWR.n23 VPWR.n3 9.3005
R57 VPWR.n25 VPWR.n24 9.3005
R58 VPWR.n26 VPWR.n0 9.3005
R59 VPWR.n28 VPWR.n27 7.12063
R60 VPWR.n10 VPWR.n9 6.33298
R61 VPWR.n11 VPWR.n10 0.717924
R62 VPWR.n28 VPWR.n0 0.148519
R63 VPWR.n11 VPWR.n7 0.120292
R64 VPWR.n7 VPWR.n6 0.120292
R65 VPWR.n16 VPWR.n6 0.120292
R66 VPWR.n17 VPWR.n16 0.120292
R67 VPWR.n18 VPWR.n17 0.120292
R68 VPWR.n18 VPWR.n4 0.120292
R69 VPWR.n22 VPWR.n4 0.120292
R70 VPWR.n23 VPWR.n22 0.120292
R71 VPWR.n24 VPWR.n23 0.120292
R72 VPWR.n24 VPWR.n0 0.120292
R73 VPWR VPWR.n28 0.0927068
R74 VPB.t2 VPB.t6 559.346
R75 VPB.t10 VPB.t7 556.386
R76 VPB.t4 VPB.t11 553.428
R77 VPB.t5 VPB.t1 358.101
R78 VPB.t0 VPB.t5 284.113
R79 VPB.t9 VPB.t8 272.274
R80 VPB.t11 VPB.t9 257.478
R81 VPB.t7 VPB.t4 248.599
R82 VPB.t6 VPB.t0 248.599
R83 VPB.t3 VPB.t2 248.599
R84 VPB.t1 VPB.t10 213.084
R85 VPB VPB.t3 139.097
R86 a_300_47.t0 a_300_47.n1 438.971
R87 a_300_47.n0 a_300_47.t3 373.283
R88 a_300_47.n1 a_300_47.t1 275.149
R89 a_300_47.n1 a_300_47.n0 156.462
R90 a_300_47.n0 a_300_47.t2 132.282
R91 VGND.n9 VGND.t7 289.36
R92 VGND.n12 VGND.t2 271.281
R93 VGND.n4 VGND.t6 240.833
R94 VGND.n8 VGND.n7 203.016
R95 VGND.n27 VGND.n26 199.739
R96 VGND.n2 VGND.n1 198.964
R97 VGND.n1 VGND.t3 38.5719
R98 VGND.n1 VGND.t4 38.5719
R99 VGND.n26 VGND.t0 38.5719
R100 VGND.n26 VGND.t1 38.5719
R101 VGND.n14 VGND.n13 34.6358
R102 VGND.n19 VGND.n18 34.6358
R103 VGND.n20 VGND.n19 34.6358
R104 VGND.n25 VGND.n24 34.6358
R105 VGND.n8 VGND.n6 28.9887
R106 VGND.n7 VGND.t8 27.6928
R107 VGND.n7 VGND.t5 24.9236
R108 VGND.n20 VGND.n2 24.0946
R109 VGND.n12 VGND.n6 23.3417
R110 VGND.n27 VGND.n25 22.9652
R111 VGND.n14 VGND.n4 22.2123
R112 VGND.n18 VGND.n4 22.2123
R113 VGND.n13 VGND.n12 20.3299
R114 VGND.n24 VGND.n2 20.3299
R115 VGND.n10 VGND.n6 9.3005
R116 VGND.n12 VGND.n11 9.3005
R117 VGND.n13 VGND.n5 9.3005
R118 VGND.n15 VGND.n14 9.3005
R119 VGND.n16 VGND.n4 9.3005
R120 VGND.n18 VGND.n17 9.3005
R121 VGND.n19 VGND.n3 9.3005
R122 VGND.n21 VGND.n20 9.3005
R123 VGND.n22 VGND.n2 9.3005
R124 VGND.n24 VGND.n23 9.3005
R125 VGND.n25 VGND.n0 9.3005
R126 VGND.n28 VGND.n27 7.12063
R127 VGND.n9 VGND.n8 6.33298
R128 VGND.n10 VGND.n9 0.717924
R129 VGND.n28 VGND.n0 0.148519
R130 VGND.n11 VGND.n10 0.120292
R131 VGND.n11 VGND.n5 0.120292
R132 VGND.n15 VGND.n5 0.120292
R133 VGND.n16 VGND.n15 0.120292
R134 VGND.n17 VGND.n16 0.120292
R135 VGND.n17 VGND.n3 0.120292
R136 VGND.n21 VGND.n3 0.120292
R137 VGND.n22 VGND.n21 0.120292
R138 VGND.n23 VGND.n22 0.120292
R139 VGND.n23 VGND.n0 0.120292
R140 VGND VGND.n28 0.11354
R141 a_466_47.n0 a_466_47.t0 88.3338
R142 a_466_47.n0 a_466_47.t1 26.3935
R143 a_466_47.n1 a_466_47.n0 14.4005
R144 VNB.t1 VNB.t7 2691.26
R145 VNB.t11 VNB.t5 2677.02
R146 VNB.t3 VNB.t10 2662.78
R147 VNB.t4 VNB.t0 1537.86
R148 VNB.t6 VNB.t11 1352.75
R149 VNB.t8 VNB.t9 1310.03
R150 VNB.t10 VNB.t8 1238.83
R151 VNB.t0 VNB.t6 1224.6
R152 VNB.t5 VNB.t3 1196.12
R153 VNB.t7 VNB.t4 1196.12
R154 VNB.t2 VNB.t1 1196.12
R155 VNB VNB.t2 911.327
R156 Q Q.t5 796.319
R157 Q.n3 Q.n0 338.481
R158 Q.n2 Q.t2 289.279
R159 Q.n3 Q.n1 202.601
R160 Q.n2 Q 52.6403
R161 Q.n0 Q.t3 30.5355
R162 Q.n0 Q.t4 30.5355
R163 Q.n1 Q.t1 28.6159
R164 Q.n1 Q.t0 28.6159
R165 Q Q.n3 9.6005
R166 Q Q.n2 6.74336
R167 Q.n3 Q 0.914786
R168 a_27_47.t0 a_27_47.n3 415.863
R169 a_27_47.n2 a_27_47.t4 316.111
R170 a_27_47.n2 a_27_47.t2 315.729
R171 a_27_47.n1 a_27_47.t1 294.873
R172 a_27_47.n0 a_27_47.t5 263.173
R173 a_27_47.n0 a_27_47.t3 227.826
R174 a_27_47.n1 a_27_47.n0 152
R175 a_27_47.n3 a_27_47.n2 20.5751
R176 a_27_47.n3 a_27_47.n1 18.9713
R177 a_562_413.n3 a_562_413.n2 745.471
R178 a_562_413.n2 a_562_413.n1 280.692
R179 a_562_413.n2 a_562_413.n0 254.02
R180 a_562_413.n0 a_562_413.t4 221.72
R181 a_562_413.n0 a_562_413.t5 149.421
R182 a_562_413.t0 a_562_413.n3 121.953
R183 a_562_413.n3 a_562_413.t2 91.4648
R184 a_562_413.n1 a_562_413.t3 46.6672
R185 a_562_413.n1 a_562_413.t1 46.6672
R186 a_660_47.t1 a_660_47.t0 93.0601
R187 a_466_369.t1 a_466_369.t0 134.631
R188 GATE_N.n0 GATE_N.t0 269.921
R189 GATE_N.n0 GATE_N.t1 234.573
R190 GATE_N.n1 GATE_N.n0 152
R191 GATE_N GATE_N.n1 10.9719
R192 GATE_N.n1 GATE_N 6.79234
R193 D.n0 D.t0 327.644
R194 D.n0 D.t1 157.338
R195 D D.n0 154.595
R196 a_193_47.n0 a_193_47.t3 464.327
R197 a_193_47.t1 a_193_47.n1 366.837
R198 a_193_47.n1 a_193_47.t0 322.567
R199 a_193_47.n0 a_193_47.t2 242.607
R200 a_193_47.n1 a_193_47.n0 187.472
R201 a_683_413.t0 a_683_413.t1 98.5005
R202 a_943_47.t0 a_943_47.t1 49.8467
C0 VPB D 0.062421f
C1 VPWR VPB 0.17189f
C2 VPB RESET_B 0.027079f
C3 VGND VPB 0.014587f
C4 VPWR GATE_N 0.019242f
C5 VPWR D 0.014068f
C6 Q VPB 0.011077f
C7 VGND GATE_N 0.019085f
C8 VGND D 0.018841f
C9 VPWR RESET_B 0.021845f
C10 VPWR VGND 0.101051f
C11 VGND RESET_B 0.017916f
C12 VPWR Q 0.432995f
C13 Q RESET_B 0.001091f
C14 VGND Q 0.275622f
C15 VPB GATE_N 0.070092f
C16 Q VNB 0.046058f
C17 VGND VNB 0.846722f
C18 VPWR VNB 0.69903f
C19 RESET_B VNB 0.091276f
C20 D VNB 0.132563f
C21 GATE_N VNB 0.195771f
C22 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_1 VGND VPWR VPB VNB Q RESET_B D GATE
X0 a_929_47.t1 a_560_425.t4 a_711_21.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR.t1 D.t0 a_299_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 Q.t0 a_711_21.t3 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3 a_465_47.t0 a_299_47.t2 VGND.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VGND.t4 a_711_21.t4 a_654_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.05985 ps=0.705 w=0.42 l=0.15
X5 VPWR.t5 GATE.t0 a_27_47.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 Q.t1 a_711_21.t5 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X7 a_560_425.t1 a_27_47.t2 a_465_369.t1 VPB.t3 sky130_fd_pr__special_pfet_01v8_hvt ad=0.0666 pd=0.73 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 VPWR.t4 a_711_21.t6 a_664_425.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2006 pd=1.61 as=0.0822 ps=0.835 w=0.42 l=0.15
X9 a_654_47.t0 a_27_47.t3 a_560_425.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_193_47.t1 a_27_47.t4 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_711_21.t1 a_560_425.t5 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2006 ps=1.61 w=1 l=0.15
X12 VPWR.t7 RESET_B.t0 a_711_21.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.165 ps=1.33 w=1 l=0.15
X13 a_193_47.t0 a_27_47.t5 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14 a_560_425.t3 a_193_47.t2 a_465_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07665 ps=0.785 w=0.42 l=0.15
X15 a_664_425.t0 a_193_47.t3 a_560_425.t0 VPB.t2 sky130_fd_pr__special_pfet_01v8_hvt ad=0.0822 pd=0.835 as=0.0666 ps=0.73 w=0.36 l=0.15
X16 VGND.t1 D.t1 a_299_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t2 RESET_B.t1 a_929_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X18 a_465_369.t0 a_299_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0935 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X19 VGND.t5 GATE.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_560_425.n2 a_560_425.n0 719.566
R1 a_560_425.n3 a_560_425.n2 282.507
R2 a_560_425.n2 a_560_425.n1 242.815
R3 a_560_425.n1 a_560_425.t5 212.081
R4 a_560_425.n1 a_560_425.t4 139.78
R5 a_560_425.n0 a_560_425.t0 106.709
R6 a_560_425.n0 a_560_425.t1 95.7644
R7 a_560_425.t2 a_560_425.n3 40.0005
R8 a_560_425.n3 a_560_425.t3 40.0005
R9 a_711_21.n1 a_711_21.t4 358.182
R10 a_711_21.n4 a_711_21.n3 296.087
R11 a_711_21.n0 a_711_21.t3 241.536
R12 a_711_21.n3 a_711_21.n0 196.675
R13 a_711_21.n2 a_711_21.t0 176.216
R14 a_711_21.n2 a_711_21.n1 173.351
R15 a_711_21.n0 a_711_21.t5 169.237
R16 a_711_21.n1 a_711_21.t6 149.822
R17 a_711_21.t1 a_711_21.n4 33.4905
R18 a_711_21.n4 a_711_21.t2 31.5205
R19 a_711_21.n3 a_711_21.n2 12.272
R20 a_929_47.t0 a_929_47.t1 60.9236
R21 VNB.t6 VNB.t4 2677.02
R22 VNB.t8 VNB.t3 2677.02
R23 VNB.t9 VNB.t2 1466.67
R24 VNB.t4 VNB.t0 1366.99
R25 VNB.t0 VNB.t5 1310.03
R26 VNB.t1 VNB.t6 1238.83
R27 VNB.t2 VNB.t1 1224.6
R28 VNB.t3 VNB.t9 1196.12
R29 VNB.t7 VNB.t8 1196.12
R30 VNB VNB.t7 683.495
R31 D.n0 D.t0 332.983
R32 D.n0 D.t1 156.249
R33 D D.n0 154.595
R34 a_299_47.t1 a_299_47.n1 435.738
R35 a_299_47.n0 a_299_47.t3 373.283
R36 a_299_47.n1 a_299_47.t0 271.432
R37 a_299_47.n1 a_299_47.n0 157.237
R38 a_299_47.n0 a_299_47.t2 132.282
R39 VPWR.n22 VPWR.n1 604.394
R40 VPWR.n8 VPWR.n7 585
R41 VPWR.n10 VPWR.n9 585
R42 VPWR.n11 VPWR.n6 316.12
R43 VPWR.n3 VPWR.n2 312.978
R44 VPWR.n9 VPWR.n8 159.476
R45 VPWR.n8 VPWR.t4 63.3219
R46 VPWR.n1 VPWR.t6 41.5552
R47 VPWR.n1 VPWR.t5 41.5552
R48 VPWR.n2 VPWR.t0 41.5552
R49 VPWR.n2 VPWR.t1 41.5552
R50 VPWR.n21 VPWR.n20 34.6358
R51 VPWR.n14 VPWR.n5 34.6358
R52 VPWR.n15 VPWR.n14 34.6358
R53 VPWR.n16 VPWR.n15 34.6358
R54 VPWR.n6 VPWR.t7 34.4755
R55 VPWR.n9 VPWR.t2 29.316
R56 VPWR.n6 VPWR.t3 26.5955
R57 VPWR.n20 VPWR.n3 25.977
R58 VPWR.n22 VPWR.n21 22.9652
R59 VPWR.n16 VPWR.n3 21.4593
R60 VPWR.n12 VPWR.n5 9.3005
R61 VPWR.n14 VPWR.n13 9.3005
R62 VPWR.n15 VPWR.n4 9.3005
R63 VPWR.n17 VPWR.n16 9.3005
R64 VPWR.n18 VPWR.n3 9.3005
R65 VPWR.n20 VPWR.n19 9.3005
R66 VPWR.n21 VPWR.n0 9.3005
R67 VPWR.n11 VPWR.n10 7.28759
R68 VPWR.n23 VPWR.n22 7.12063
R69 VPWR.n10 VPWR.n7 6.49602
R70 VPWR.n7 VPWR.n5 3.22579
R71 VPWR.n12 VPWR.n11 0.483236
R72 VPWR.n23 VPWR.n0 0.148519
R73 VPWR.n13 VPWR.n12 0.120292
R74 VPWR.n13 VPWR.n4 0.120292
R75 VPWR.n17 VPWR.n4 0.120292
R76 VPWR.n18 VPWR.n17 0.120292
R77 VPWR.n19 VPWR.n18 0.120292
R78 VPWR.n19 VPWR.n0 0.120292
R79 VPWR VPWR.n23 0.114842
R80 VPB.t8 VPB.t1 556.386
R81 VPB.t5 VPB.t4 449.844
R82 VPB.t2 VPB.t5 334.425
R83 VPB.t3 VPB.t2 307.788
R84 VPB.t4 VPB.t9 284.113
R85 VPB.t0 VPB.t3 281.154
R86 VPB.t9 VPB.t6 272.274
R87 VPB.t1 VPB.t0 248.599
R88 VPB.t7 VPB.t8 248.599
R89 VPB VPB.t7 142.056
R90 Q.n0 Q.t0 374.618
R91 Q.n1 Q.t1 209.923
R92 Q Q.n1 82.7196
R93 Q Q.n0 8.95158
R94 Q.n0 Q 7.65628
R95 Q.n1 Q 6.9619
R96 VGND.n4 VGND.t4 244.668
R97 VGND.n6 VGND.n5 215.827
R98 VGND.n17 VGND.n16 199.739
R99 VGND.n2 VGND.n1 198.964
R100 VGND.n1 VGND.t0 38.5719
R101 VGND.n1 VGND.t1 38.5719
R102 VGND.n16 VGND.t6 38.5719
R103 VGND.n16 VGND.t5 38.5719
R104 VGND.n9 VGND.n8 34.6358
R105 VGND.n10 VGND.n9 34.6358
R106 VGND.n15 VGND.n14 34.6358
R107 VGND.n5 VGND.t2 32.3082
R108 VGND.n5 VGND.t3 24.9236
R109 VGND.n10 VGND.n2 24.4711
R110 VGND.n8 VGND.n4 22.9652
R111 VGND.n17 VGND.n15 22.9652
R112 VGND.n14 VGND.n2 19.9534
R113 VGND.n15 VGND.n0 9.3005
R114 VGND.n14 VGND.n13 9.3005
R115 VGND.n12 VGND.n2 9.3005
R116 VGND.n11 VGND.n10 9.3005
R117 VGND.n9 VGND.n3 9.3005
R118 VGND.n8 VGND.n7 9.3005
R119 VGND.n6 VGND.n4 7.194
R120 VGND.n18 VGND.n17 7.12063
R121 VGND.n7 VGND.n6 0.216848
R122 VGND.n18 VGND.n0 0.148519
R123 VGND.n7 VGND.n3 0.120292
R124 VGND.n11 VGND.n3 0.120292
R125 VGND.n12 VGND.n11 0.120292
R126 VGND.n13 VGND.n12 0.120292
R127 VGND.n13 VGND.n0 0.120292
R128 VGND VGND.n18 0.114842
R129 a_465_47.t0 a_465_47.t1 104.287
R130 a_654_47.t0 a_654_47.t1 81.4291
R131 GATE.n0 GATE.t0 272.062
R132 GATE.n0 GATE.t1 236.716
R133 GATE.n1 GATE.n0 152
R134 GATE GATE.n1 11.2005
R135 GATE.n1 GATE 6.93383
R136 a_27_47.n2 a_27_47.t3 426.659
R137 a_27_47.t0 a_27_47.n3 410.943
R138 a_27_47.n1 a_27_47.t1 294.043
R139 a_27_47.n0 a_27_47.t5 262.945
R140 a_27_47.n2 a_27_47.t2 228.631
R141 a_27_47.n0 a_27_47.t4 227.597
R142 a_27_47.n3 a_27_47.n2 177.572
R143 a_27_47.n1 a_27_47.n0 152
R144 a_27_47.n3 a_27_47.n1 18.9713
R145 a_465_369.t0 a_465_369.t1 147.922
R146 a_664_425.n0 a_664_425.t0 158.695
R147 a_664_425.n0 a_664_425.t1 43.3289
R148 a_664_425.n1 a_664_425.n0 23.6405
R149 a_193_47.t0 a_193_47.n1 367.062
R150 a_193_47.n0 a_193_47.t2 334.781
R151 a_193_47.n1 a_193_47.t1 322.807
R152 a_193_47.n0 a_193_47.t3 290.613
R153 a_193_47.n1 a_193_47.n0 23.606
R154 RESET_B.n0 RESET_B.t0 241.536
R155 RESET_B.n0 RESET_B.t1 169.237
R156 RESET_B.n1 RESET_B.n0 157.042
R157 RESET_B RESET_B.n1 12.8005
R158 RESET_B.n1 RESET_B 4.46111
C0 RESET_B Q 0.009647f
C1 D VGND 0.018889f
C2 RESET_B VGND 0.07767f
C3 VPWR Q 0.083402f
C4 VPWR VGND 0.071358f
C5 Q VGND 0.065713f
C6 VPB GATE 0.06938f
C7 VPB D 0.072383f
C8 VPB RESET_B 0.027185f
C9 VPB VPWR 0.130924f
C10 GATE VPWR 0.017104f
C11 VPB Q 0.010797f
C12 D VPWR 0.014303f
C13 VPB VGND 0.012927f
C14 GATE VGND 0.018932f
C15 RESET_B VPWR 0.02126f
C16 VGND VNB 0.700745f
C17 Q VNB 0.090048f
C18 VPWR VNB 0.555865f
C19 RESET_B VNB 0.09197f
C20 D VNB 0.136397f
C21 GATE VNB 0.196004f
C22 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_2 VGND VPWR VPB VNB Q RESET_B D GATE
X0 VPWR.t1 D.t0 a_299_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47.t1 a_193_47.t2 a_465_47.t0 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0603 pd=0.695 as=0.066 ps=0.745 w=0.36 l=0.15
X2 VPWR.t4 a_711_307.t3 a_644_413.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3 a_465_47.t1 a_299_47.t2 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR.t8 GATE.t0 a_27_47.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 Q.t1 a_711_307.t4 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t5 a_711_307.t5 a_657_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7 VPWR.t6 a_711_307.t6 Q.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X8 a_657_47.t0 a_27_47.t2 a_560_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0603 ps=0.695 w=0.36 l=0.15
X9 a_193_47.t0 a_27_47.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 Q.t3 a_711_307.t7 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X11 VPWR.t3 RESET_B.t0 a_711_307.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.32 w=1 l=0.15
X12 a_940_47.t0 a_560_47.t4 a_711_307.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47.t1 a_27_47.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14 VGND.t4 a_711_307.t8 Q.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_711_307.t0 a_560_47.t5 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.27 ps=2.54 w=1 l=0.15
X16 VGND.t2 D.t1 a_299_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 a_644_413.t0 a_193_47.t3 a_560_47.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VGND.t1 RESET_B.t1 a_940_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.104 ps=0.97 w=0.65 l=0.15
X19 a_465_369.t0 a_299_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_560_47.t3 a_27_47.t5 a_465_369.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X21 VGND.t7 GATE.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 326.764
R1 D.n0 D.t1 156.457
R2 D D.n0 154.595
R3 a_299_47.t0 a_299_47.n1 436.368
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t1 272.137
R6 a_299_47.n1 a_299_47.n0 157.042
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n12 VPWR.t7 861.39
R9 VPWR.n13 VPWR.t4 662.628
R10 VPWR.n24 VPWR.n1 604.394
R11 VPWR.n9 VPWR.t6 410.901
R12 VPWR.n19 VPWR.n4 312.632
R13 VPWR.n8 VPWR.n7 308.978
R14 VPWR.n1 VPWR.t0 41.5552
R15 VPWR.n1 VPWR.t8 41.5552
R16 VPWR.n4 VPWR.t2 41.5552
R17 VPWR.n4 VPWR.t1 41.5552
R18 VPWR.n23 VPWR.n2 34.6358
R19 VPWR.n17 VPWR.n5 34.6358
R20 VPWR.n18 VPWR.n17 34.6358
R21 VPWR.n25 VPWR.n24 30.7593
R22 VPWR.n7 VPWR.t5 26.5955
R23 VPWR.n7 VPWR.t3 26.5955
R24 VPWR.n19 VPWR.n2 25.977
R25 VPWR.n11 VPWR.n8 23.3417
R26 VPWR.n24 VPWR.n23 22.9652
R27 VPWR.n13 VPWR.n5 22.5887
R28 VPWR.n19 VPWR.n18 21.0829
R29 VPWR.n12 VPWR.n11 20.3299
R30 VPWR.n13 VPWR.n12 14.3064
R31 VPWR.n11 VPWR.n10 9.3005
R32 VPWR.n12 VPWR.n6 9.3005
R33 VPWR.n14 VPWR.n13 9.3005
R34 VPWR.n15 VPWR.n5 9.3005
R35 VPWR.n17 VPWR.n16 9.3005
R36 VPWR.n18 VPWR.n3 9.3005
R37 VPWR.n20 VPWR.n19 9.3005
R38 VPWR.n21 VPWR.n2 9.3005
R39 VPWR.n23 VPWR.n22 9.3005
R40 VPWR.n24 VPWR.n0 9.3005
R41 VPWR.n9 VPWR.n8 6.4202
R42 VPWR.n10 VPWR.n9 0.647392
R43 VPWR.n10 VPWR.n6 0.120292
R44 VPWR.n14 VPWR.n6 0.120292
R45 VPWR.n15 VPWR.n14 0.120292
R46 VPWR.n16 VPWR.n15 0.120292
R47 VPWR.n16 VPWR.n3 0.120292
R48 VPWR.n20 VPWR.n3 0.120292
R49 VPWR.n21 VPWR.n20 0.120292
R50 VPWR.n22 VPWR.n21 0.120292
R51 VPWR.n22 VPWR.n0 0.120292
R52 VPWR.n0 VPWR 0.11899
R53 VPWR VPWR.n25 0.0213333
R54 VPWR.n25 VPWR 0.00180208
R55 VPB.t5 VPB.t8 588.942
R56 VPB.t0 VPB.t1 556.386
R57 VPB.t10 VPB.t5 287.072
R58 VPB.t2 VPB.t3 281.154
R59 VPB.t8 VPB.t4 278.193
R60 VPB.t6 VPB.t7 269.315
R61 VPB.t4 VPB.t6 248.599
R62 VPB.t3 VPB.t10 248.599
R63 VPB.t1 VPB.t2 248.599
R64 VPB.t9 VPB.t0 248.599
R65 VPB VPB.t9 139.097
R66 a_193_47.t1 a_193_47.n1 366.837
R67 a_193_47.n0 a_193_47.t2 343.087
R68 a_193_47.n1 a_193_47.t0 322.567
R69 a_193_47.n0 a_193_47.t3 298.646
R70 a_193_47.n1 a_193_47.n0 24.9193
R71 a_465_47.n0 a_465_47.t0 66.6672
R72 a_465_47.n0 a_465_47.t1 26.3935
R73 a_465_47.n1 a_465_47.n0 14.4005
R74 a_560_47.n3 a_560_47.n2 708.375
R75 a_560_47.n2 a_560_47.n0 263.329
R76 a_560_47.n2 a_560_47.n1 256.486
R77 a_560_47.n0 a_560_47.t5 221.72
R78 a_560_47.n0 a_560_47.t4 149.421
R79 a_560_47.n1 a_560_47.t0 66.6672
R80 a_560_47.t2 a_560_47.n3 63.3219
R81 a_560_47.n3 a_560_47.t3 63.3219
R82 a_560_47.n1 a_560_47.t1 45.0005
R83 VNB.t8 VNB.t4 2677.02
R84 VNB.t1 VNB.t5 2677.02
R85 VNB.t2 VNB.t0 1381.23
R86 VNB.t0 VNB.t8 1352.75
R87 VNB.t6 VNB.t2 1352.75
R88 VNB.t4 VNB.t3 1338.51
R89 VNB.t3 VNB.t9 1295.79
R90 VNB.t9 VNB.t10 1196.12
R91 VNB.t5 VNB.t6 1196.12
R92 VNB.t7 VNB.t1 1196.12
R93 VNB VNB.t7 911.327
R94 a_711_307.n4 a_711_307.t5 368.329
R95 a_711_307.n6 a_711_307.n5 299.93
R96 a_711_307.n3 a_711_307.t1 222.536
R97 a_711_307.n2 a_711_307.t4 214.272
R98 a_711_307.n0 a_711_307.t6 212.081
R99 a_711_307.n5 a_711_307.n4 191.758
R100 a_711_307.n3 a_711_307.n2 152
R101 a_711_307.n4 a_711_307.t3 149.822
R102 a_711_307.n0 a_711_307.t8 139.78
R103 a_711_307.n1 a_711_307.t7 139.78
R104 a_711_307.n5 a_711_307.n3 69.5751
R105 a_711_307.n1 a_711_307.n0 61.346
R106 a_711_307.t0 a_711_307.n6 36.4455
R107 a_711_307.n6 a_711_307.t2 26.5955
R108 a_711_307.n2 a_711_307.n1 2.92171
R109 a_644_413.t0 a_644_413.t1 157.131
R110 VGND.n8 VGND.t4 292.26
R111 VGND.n4 VGND.t5 240.325
R112 VGND.n7 VGND.n6 205.707
R113 VGND.n25 VGND.n24 199.739
R114 VGND.n2 VGND.n1 198.964
R115 VGND.n1 VGND.t3 38.5719
R116 VGND.n1 VGND.t2 38.5719
R117 VGND.n24 VGND.t0 38.5719
R118 VGND.n24 VGND.t7 38.5719
R119 VGND.n8 VGND.n7 36.2765
R120 VGND.n11 VGND.n10 34.6358
R121 VGND.n12 VGND.n11 34.6358
R122 VGND.n17 VGND.n16 34.6358
R123 VGND.n18 VGND.n17 34.6358
R124 VGND.n23 VGND.n22 34.6358
R125 VGND.n6 VGND.t1 31.3851
R126 VGND.n6 VGND.t6 24.9236
R127 VGND.n18 VGND.n2 24.4711
R128 VGND.n12 VGND.n4 23.3417
R129 VGND.n25 VGND.n23 22.9652
R130 VGND.n16 VGND.n4 20.3299
R131 VGND.n22 VGND.n2 19.9534
R132 VGND.n10 VGND.n9 9.3005
R133 VGND.n11 VGND.n5 9.3005
R134 VGND.n13 VGND.n12 9.3005
R135 VGND.n14 VGND.n4 9.3005
R136 VGND.n16 VGND.n15 9.3005
R137 VGND.n17 VGND.n3 9.3005
R138 VGND.n19 VGND.n18 9.3005
R139 VGND.n20 VGND.n2 9.3005
R140 VGND.n22 VGND.n21 9.3005
R141 VGND.n23 VGND.n0 9.3005
R142 VGND.n26 VGND.n25 7.12063
R143 VGND.n10 VGND.n7 3.76521
R144 VGND.n9 VGND.n8 2.08078
R145 VGND.n26 VGND.n0 0.148519
R146 VGND.n9 VGND.n5 0.120292
R147 VGND.n13 VGND.n5 0.120292
R148 VGND.n14 VGND.n13 0.120292
R149 VGND.n15 VGND.n14 0.120292
R150 VGND.n15 VGND.n3 0.120292
R151 VGND.n19 VGND.n3 0.120292
R152 VGND.n20 VGND.n19 0.120292
R153 VGND.n21 VGND.n20 0.120292
R154 VGND.n21 VGND.n0 0.120292
R155 VGND VGND.n26 0.11354
R156 GATE.n0 GATE.t0 270.457
R157 GATE.n0 GATE.t1 235.109
R158 GATE.n1 GATE.n0 152
R159 GATE GATE.n1 11.2005
R160 GATE.n1 GATE 6.93383
R161 a_27_47.n2 a_27_47.t2 453.743
R162 a_27_47.t0 a_27_47.n3 415.863
R163 a_27_47.n1 a_27_47.t1 289.399
R164 a_27_47.n0 a_27_47.t4 263.173
R165 a_27_47.n2 a_27_47.t5 236.369
R166 a_27_47.n0 a_27_47.t3 227.826
R167 a_27_47.n3 a_27_47.n2 177.379
R168 a_27_47.n1 a_27_47.n0 152
R169 a_27_47.n3 a_27_47.n1 18.9713
R170 Q Q.n2 593.297
R171 Q.n1 Q.n0 239.091
R172 Q.n2 Q.t0 30.5355
R173 Q.n2 Q.t1 29.5505
R174 Q.n0 Q.t2 24.9236
R175 Q.n0 Q.t3 24.9236
R176 Q.n1 Q 11.5205
R177 Q.n3 Q 4.82857
R178 Q Q.n3 2.80752
R179 Q.n1 Q 2.18853
R180 Q.n3 Q.n1 0.547509
R181 a_657_47.t1 a_657_47.t0 93.0601
R182 RESET_B.n0 RESET_B.t0 241
R183 RESET_B.n0 RESET_B.t1 168.701
R184 RESET_B.n1 RESET_B.n0 162.373
R185 RESET_B.n1 RESET_B 2.86617
R186 RESET_B RESET_B.n1 1.98671
R187 a_940_47.t0 a_940_47.t1 59.0774
R188 a_465_369.t0 a_465_369.t1 132.286
C0 VPWR VGND 0.081538f
C1 VPWR Q 0.189666f
C2 VPWR VPB 0.153112f
C3 VGND Q 0.132663f
C4 VGND VPB 0.014088f
C5 VPWR GATE 0.019079f
C6 Q VPB 0.006968f
C7 VPWR D 0.014099f
C8 VGND GATE 0.016666f
C9 VPWR RESET_B 0.02147f
C10 VGND D 0.019078f
C11 VPB GATE 0.069748f
C12 VGND RESET_B 0.01688f
C13 VPB D 0.063192f
C14 Q RESET_B 0.001182f
C15 VPB RESET_B 0.027589f
C16 Q VNB 0.047407f
C17 VGND VNB 0.758809f
C18 VPWR VNB 0.619736f
C19 RESET_B VNB 0.092088f
C20 D VNB 0.134235f
C21 GATE VNB 0.194444f
C22 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_4 VGND VPWR VPB VNB Q GATE D RESET_B
X0 VPWR.t1 RESET_B.t0 a_725_21.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_466_47.t1 a_300_47.t2 VGND.t8 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_562_413.t0 a_193_47.t2 a_466_47.t0 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X3 VGND.t3 a_725_21.t3 a_660_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4 VGND.t6 a_725_21.t4 Q.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.099125 ps=0.955 w=0.65 l=0.15
X5 a_466_369.t1 a_300_47.t3 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X6 VPWR.t0 GATE.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 VPWR.t7 D.t0 a_300_47.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 VPWR.t6 a_725_21.t5 Q.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.1525 ps=1.305 w=1 l=0.15
X9 VGND.t5 a_725_21.t6 Q.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X10 a_562_413.t2 a_27_47.t2 a_466_369.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X11 a_725_21.t1 a_562_413.t4 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47.t0 a_27_47.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VPWR.t3 a_725_21.t7 a_683_413.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X14 a_943_47.t1 a_562_413.t5 a_725_21.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 Q.t1 a_725_21.t8 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1425 ps=1.285 w=1 l=0.15
X16 a_683_413.t0 a_193_47.t3 a_562_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X17 a_193_47.t1 a_27_47.t4 VPWR.t9 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X18 a_660_47.t1 a_27_47.t5 a_562_413.t3 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X19 Q.t3 a_725_21.t9 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.092625 ps=0.935 w=0.65 l=0.15
X20 VGND.t7 D.t1 a_300_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VGND.t1 RESET_B.t1 a_943_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t4 a_725_21.t10 Q.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X23 VGND.t0 GATE.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 RESET_B.n0 RESET_B.t0 241.536
R1 RESET_B.n0 RESET_B.t1 169.237
R2 RESET_B RESET_B.n0 162.28
R3 a_725_21.n7 a_725_21.t3 368.329
R4 a_725_21.n9 a_725_21.n8 299.166
R5 a_725_21.n6 a_725_21.t2 231.398
R6 a_725_21.n5 a_725_21.n1 212.081
R7 a_725_21.n2 a_725_21.t10 212.081
R8 a_725_21.n3 a_725_21.t8 212.081
R9 a_725_21.n4 a_725_21.t5 212.081
R10 a_725_21.n8 a_725_21.n7 187.685
R11 a_725_21.n6 a_725_21.n5 152
R12 a_725_21.n7 a_725_21.t7 149.822
R13 a_725_21.n5 a_725_21.n0 139.78
R14 a_725_21.n2 a_725_21.t6 139.78
R15 a_725_21.n3 a_725_21.t9 139.78
R16 a_725_21.n4 a_725_21.t4 139.78
R17 a_725_21.n8 a_725_21.n6 76.7206
R18 a_725_21.n3 a_725_21.n2 67.1884
R19 a_725_21.n5 a_725_21.n4 66.4581
R20 a_725_21.n4 a_725_21.n3 63.5369
R21 a_725_21.t0 a_725_21.n9 26.5955
R22 a_725_21.n9 a_725_21.t1 26.5955
R23 VPWR.n15 VPWR.t2 871.352
R24 VPWR.n5 VPWR.t3 666.86
R25 VPWR.n27 VPWR.n1 604.394
R26 VPWR.n13 VPWR.t1 340.372
R27 VPWR.n3 VPWR.n2 311.356
R28 VPWR.n10 VPWR.t4 250.055
R29 VPWR.n9 VPWR.n8 221.748
R30 VPWR.n1 VPWR.t9 41.5552
R31 VPWR.n1 VPWR.t0 41.5552
R32 VPWR.n2 VPWR.t8 41.5552
R33 VPWR.n2 VPWR.t7 41.5552
R34 VPWR.n26 VPWR.n25 34.6358
R35 VPWR.n20 VPWR.n19 34.6358
R36 VPWR.n21 VPWR.n20 34.6358
R37 VPWR.n8 VPWR.t6 29.5505
R38 VPWR.n12 VPWR.n9 28.9887
R39 VPWR.n19 VPWR.n5 28.2358
R40 VPWR.n8 VPWR.t5 26.5955
R41 VPWR.n25 VPWR.n3 26.3534
R42 VPWR.n27 VPWR.n26 22.9652
R43 VPWR.n14 VPWR.n13 21.4593
R44 VPWR.n13 VPWR.n12 19.9534
R45 VPWR.n21 VPWR.n3 19.2005
R46 VPWR.n15 VPWR.n14 18.4476
R47 VPWR.n15 VPWR.n5 14.3064
R48 VPWR.n12 VPWR.n11 9.3005
R49 VPWR.n13 VPWR.n7 9.3005
R50 VPWR.n14 VPWR.n6 9.3005
R51 VPWR.n16 VPWR.n15 9.3005
R52 VPWR.n17 VPWR.n5 9.3005
R53 VPWR.n19 VPWR.n18 9.3005
R54 VPWR.n20 VPWR.n4 9.3005
R55 VPWR.n22 VPWR.n21 9.3005
R56 VPWR.n23 VPWR.n3 9.3005
R57 VPWR.n25 VPWR.n24 9.3005
R58 VPWR.n26 VPWR.n0 9.3005
R59 VPWR.n28 VPWR.n27 7.12063
R60 VPWR.n10 VPWR.n9 6.33298
R61 VPWR.n11 VPWR.n10 0.717924
R62 VPWR.n28 VPWR.n0 0.148519
R63 VPWR.n11 VPWR.n7 0.120292
R64 VPWR.n7 VPWR.n6 0.120292
R65 VPWR.n16 VPWR.n6 0.120292
R66 VPWR.n17 VPWR.n16 0.120292
R67 VPWR.n18 VPWR.n17 0.120292
R68 VPWR.n18 VPWR.n4 0.120292
R69 VPWR.n22 VPWR.n4 0.120292
R70 VPWR.n23 VPWR.n22 0.120292
R71 VPWR.n24 VPWR.n23 0.120292
R72 VPWR.n24 VPWR.n0 0.120292
R73 VPWR VPWR.n28 0.0927068
R74 VPB.t11 VPB.t9 559.346
R75 VPB.t7 VPB.t3 556.386
R76 VPB.t2 VPB.t8 553.428
R77 VPB.t4 VPB.t1 358.101
R78 VPB.t10 VPB.t4 284.113
R79 VPB.t6 VPB.t5 272.274
R80 VPB.t8 VPB.t6 257.478
R81 VPB.t3 VPB.t2 248.599
R82 VPB.t9 VPB.t10 248.599
R83 VPB.t0 VPB.t11 248.599
R84 VPB.t1 VPB.t7 213.084
R85 VPB VPB.t0 139.097
R86 a_300_47.t0 a_300_47.n1 438.971
R87 a_300_47.n0 a_300_47.t3 373.283
R88 a_300_47.n1 a_300_47.t1 275.149
R89 a_300_47.n1 a_300_47.n0 156.462
R90 a_300_47.n0 a_300_47.t2 132.282
R91 VGND.n9 VGND.t5 289.36
R92 VGND.n12 VGND.t1 271.281
R93 VGND.n4 VGND.t3 240.833
R94 VGND.n8 VGND.n7 203.016
R95 VGND.n27 VGND.n26 199.739
R96 VGND.n2 VGND.n1 198.964
R97 VGND.n1 VGND.t8 38.5719
R98 VGND.n1 VGND.t7 38.5719
R99 VGND.n26 VGND.t2 38.5719
R100 VGND.n26 VGND.t0 38.5719
R101 VGND.n14 VGND.n13 34.6358
R102 VGND.n19 VGND.n18 34.6358
R103 VGND.n20 VGND.n19 34.6358
R104 VGND.n25 VGND.n24 34.6358
R105 VGND.n8 VGND.n6 28.9887
R106 VGND.n7 VGND.t6 27.6928
R107 VGND.n7 VGND.t4 24.9236
R108 VGND.n20 VGND.n2 24.0946
R109 VGND.n12 VGND.n6 23.3417
R110 VGND.n27 VGND.n25 22.9652
R111 VGND.n14 VGND.n4 22.2123
R112 VGND.n18 VGND.n4 22.2123
R113 VGND.n13 VGND.n12 20.3299
R114 VGND.n24 VGND.n2 20.3299
R115 VGND.n10 VGND.n6 9.3005
R116 VGND.n12 VGND.n11 9.3005
R117 VGND.n13 VGND.n5 9.3005
R118 VGND.n15 VGND.n14 9.3005
R119 VGND.n16 VGND.n4 9.3005
R120 VGND.n18 VGND.n17 9.3005
R121 VGND.n19 VGND.n3 9.3005
R122 VGND.n21 VGND.n20 9.3005
R123 VGND.n22 VGND.n2 9.3005
R124 VGND.n24 VGND.n23 9.3005
R125 VGND.n25 VGND.n0 9.3005
R126 VGND.n28 VGND.n27 7.12063
R127 VGND.n9 VGND.n8 6.33298
R128 VGND.n10 VGND.n9 0.717924
R129 VGND.n28 VGND.n0 0.148519
R130 VGND.n11 VGND.n10 0.120292
R131 VGND.n11 VGND.n5 0.120292
R132 VGND.n15 VGND.n5 0.120292
R133 VGND.n16 VGND.n15 0.120292
R134 VGND.n17 VGND.n16 0.120292
R135 VGND.n17 VGND.n3 0.120292
R136 VGND.n21 VGND.n3 0.120292
R137 VGND.n22 VGND.n21 0.120292
R138 VGND.n23 VGND.n22 0.120292
R139 VGND.n23 VGND.n0 0.120292
R140 VGND VGND.n28 0.11354
R141 a_466_47.n0 a_466_47.t0 88.3338
R142 a_466_47.n0 a_466_47.t1 26.3935
R143 a_466_47.n1 a_466_47.n0 14.4005
R144 VNB.t3 VNB.t9 2691.26
R145 VNB.t7 VNB.t2 2677.02
R146 VNB.t1 VNB.t6 2662.78
R147 VNB.t11 VNB.t8 1537.86
R148 VNB.t10 VNB.t7 1352.75
R149 VNB.t4 VNB.t5 1310.03
R150 VNB.t6 VNB.t4 1238.83
R151 VNB.t8 VNB.t10 1224.6
R152 VNB.t2 VNB.t1 1196.12
R153 VNB.t9 VNB.t11 1196.12
R154 VNB.t0 VNB.t3 1196.12
R155 VNB VNB.t0 911.327
R156 Q Q.t2 796.319
R157 Q.n2 Q.n0 338.481
R158 Q.n3 Q.t5 289.279
R159 Q.n2 Q.n1 202.601
R160 Q.n3 Q 52.6403
R161 Q.n0 Q.t0 30.5355
R162 Q.n0 Q.t1 30.5355
R163 Q.n1 Q.t4 28.6159
R164 Q.n1 Q.t3 28.6159
R165 Q.n2 Q 9.6005
R166 Q Q.n3 6.74336
R167 Q Q.n2 0.914786
R168 a_193_47.t1 a_193_47.n1 366.837
R169 a_193_47.n0 a_193_47.t2 329.659
R170 a_193_47.n1 a_193_47.t0 322.567
R171 a_193_47.n0 a_193_47.t3 308.204
R172 a_193_47.n1 a_193_47.n0 25.0585
R173 a_562_413.n3 a_562_413.n2 715.871
R174 a_562_413.n2 a_562_413.n1 283.635
R175 a_562_413.n2 a_562_413.n0 261.31
R176 a_562_413.n0 a_562_413.t4 221.72
R177 a_562_413.n0 a_562_413.t5 149.421
R178 a_562_413.n3 a_562_413.t2 121.953
R179 a_562_413.t1 a_562_413.n3 91.4648
R180 a_562_413.n1 a_562_413.t3 46.6672
R181 a_562_413.n1 a_562_413.t0 46.6672
R182 a_660_47.t0 a_660_47.t1 93.0601
R183 a_466_369.t1 a_466_369.t0 134.631
R184 GATE.n0 GATE.t0 269.921
R185 GATE.n0 GATE.t1 234.573
R186 GATE.n1 GATE.n0 152
R187 GATE GATE.n1 10.9719
R188 GATE.n1 GATE 6.79234
R189 a_27_47.n2 a_27_47.t5 464.327
R190 a_27_47.t0 a_27_47.n3 415.863
R191 a_27_47.n1 a_27_47.t1 294.873
R192 a_27_47.n0 a_27_47.t4 263.173
R193 a_27_47.n2 a_27_47.t2 242.607
R194 a_27_47.n0 a_27_47.t3 227.826
R195 a_27_47.n3 a_27_47.n2 176.625
R196 a_27_47.n1 a_27_47.n0 152
R197 a_27_47.n3 a_27_47.n1 18.9713
R198 D.n0 D.t0 327.644
R199 D.n0 D.t1 157.338
R200 D D.n0 154.595
R201 a_683_413.t0 a_683_413.t1 98.5005
R202 a_943_47.t0 a_943_47.t1 49.8467
C0 VPB RESET_B 0.027109f
C1 VPB VPWR 0.172518f
C2 VPB VGND 0.015263f
C3 GATE VPWR 0.019242f
C4 VPB Q 0.011077f
C5 D VPWR 0.014068f
C6 GATE VGND 0.019085f
C7 RESET_B VPWR 0.021845f
C8 D VGND 0.018841f
C9 RESET_B VGND 0.017916f
C10 VPWR VGND 0.101051f
C11 RESET_B Q 0.001091f
C12 VPWR Q 0.432995f
C13 VGND Q 0.275622f
C14 VPB GATE 0.070092f
C15 VPB D 0.062421f
C16 Q VNB 0.046058f
C17 VGND VNB 0.846901f
C18 VPWR VNB 0.69959f
C19 RESET_B VNB 0.091013f
C20 D VNB 0.132563f
C21 GATE VNB 0.195771f
C22 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxbn_1 VGND VPWR VPB VNB Q_N Q D GATE_N
X0 a_560_47.t2 a_193_47.t2 a_470_369.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0968 ps=0.97 w=0.42 l=0.15
X1 a_560_47.t0 a_27_47.t2 a_465_47.t1 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0549 pd=0.665 as=0.066 ps=0.745 w=0.36 l=0.15
X2 a_465_47.t0 a_299_47.t2 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_674_413.t1 a_27_47.t3 a_560_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X4 VPWR.t3 a_716_21.t2 a_1124_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t6 GATE_N.t0 a_27_47.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 VGND.t2 a_560_47.t4 a_716_21.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Q.t1 a_716_21.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_193_47.t0 a_27_47.t4 VGND.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_651_47.t1 a_193_47.t3 a_560_47.t3 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0549 ps=0.665 w=0.36 l=0.15
X10 Q.t0 a_716_21.t4 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Q_N.t1 a_1124_47.t2 VPWR.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X12 a_193_47.t1 a_27_47.t5 VPWR.t8 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 VPWR.t5 a_560_47.t5 a_716_21.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Q_N.t0 a_1124_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15 a_470_369.t1 a_299_47.t3 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 VGND.t6 D.t0 a_299_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t5 a_716_21.t5 a_1124_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 VPWR.t0 D.t1 a_299_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X19 VPWR.t1 a_716_21.t6 a_674_413.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X20 VGND.t7 a_716_21.t7 a_651_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X21 VGND.t3 GATE_N.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_193_47.n0 a_193_47.t3 562.716
R1 a_193_47.t1 a_193_47.n1 366.837
R2 a_193_47.n1 a_193_47.t0 322.567
R3 a_193_47.n0 a_193_47.t2 219.042
R4 a_193_47.n1 a_193_47.n0 187.49
R5 a_470_369.t1 a_470_369.t0 134.631
R6 a_560_47.n3 a_560_47.n2 728.84
R7 a_560_47.n2 a_560_47.n1 286.272
R8 a_560_47.n2 a_560_47.n0 241.047
R9 a_560_47.n0 a_560_47.t5 212.081
R10 a_560_47.n0 a_560_47.t4 139.78
R11 a_560_47.n3 a_560_47.t2 119.608
R12 a_560_47.t1 a_560_47.n3 63.3219
R13 a_560_47.n1 a_560_47.t0 51.6672
R14 a_560_47.n1 a_560_47.t3 50.0005
R15 VPB.t4 VPB.t0 571.184
R16 VPB.t2 VPB.t1 556.386
R17 VPB.t10 VPB.t8 556.386
R18 VPB.t6 VPB.t3 319.627
R19 VPB.t7 VPB.t6 284.113
R20 VPB.t1 VPB.t5 281.154
R21 VPB.t8 VPB.t2 248.599
R22 VPB.t0 VPB.t7 248.599
R23 VPB.t9 VPB.t4 248.599
R24 VPB.t3 VPB.t10 213.084
R25 VPB VPB.t9 139.097
R26 a_27_47.t0 a_27_47.n3 415.863
R27 a_27_47.n2 a_27_47.t2 371.238
R28 a_27_47.n2 a_27_47.t3 303.087
R29 a_27_47.n1 a_27_47.t1 294.873
R30 a_27_47.n0 a_27_47.t5 263.173
R31 a_27_47.n0 a_27_47.t4 227.826
R32 a_27_47.n1 a_27_47.n0 152
R33 a_27_47.n3 a_27_47.n2 20.5929
R34 a_27_47.n3 a_27_47.n1 18.9713
R35 a_465_47.n0 a_465_47.t1 66.6672
R36 a_465_47.n0 a_465_47.t0 26.3935
R37 a_465_47.n1 a_465_47.n0 14.4005
R38 VNB.t5 VNB.t6 2677.02
R39 VNB.t8 VNB.t2 2677.02
R40 VNB.t9 VNB.t7 2677.02
R41 VNB.t6 VNB.t0 1352.75
R42 VNB.t1 VNB.t8 1352.75
R43 VNB.t4 VNB.t10 1352.75
R44 VNB.t10 VNB.t1 1295.79
R45 VNB.t2 VNB.t5 1196.12
R46 VNB.t7 VNB.t4 1196.12
R47 VNB.t3 VNB.t9 1196.12
R48 VNB VNB.t3 669.256
R49 a_299_47.n0 a_299_47.t2 464.685
R50 a_299_47.t0 a_299_47.n1 421.714
R51 a_299_47.n0 a_299_47.t3 328.296
R52 a_299_47.n1 a_299_47.t1 280.856
R53 a_299_47.n1 a_299_47.n0 152
R54 VGND.n11 VGND.t7 240.833
R55 VGND.n8 VGND.n7 207.585
R56 VGND.n6 VGND.n5 199.739
R57 VGND.n23 VGND.n1 199.739
R58 VGND.n18 VGND.n17 197.981
R59 VGND.n7 VGND.t5 54.2862
R60 VGND.n17 VGND.t1 38.5719
R61 VGND.n17 VGND.t6 38.5719
R62 VGND.n1 VGND.t8 38.5719
R63 VGND.n1 VGND.t3 38.5719
R64 VGND.n12 VGND.n3 34.6358
R65 VGND.n16 VGND.n3 34.6358
R66 VGND.n19 VGND.n0 34.6358
R67 VGND.n24 VGND.n23 30.7593
R68 VGND.n7 VGND.t0 25.9346
R69 VGND.n5 VGND.t4 24.9236
R70 VGND.n5 VGND.t2 24.9236
R71 VGND.n12 VGND.n11 23.7181
R72 VGND.n23 VGND.n0 22.9652
R73 VGND.n18 VGND.n16 22.5887
R74 VGND.n11 VGND.n10 20.7064
R75 VGND.n10 VGND.n6 20.3299
R76 VGND.n19 VGND.n18 19.9534
R77 VGND.n23 VGND.n22 9.3005
R78 VGND.n21 VGND.n0 9.3005
R79 VGND.n20 VGND.n19 9.3005
R80 VGND.n18 VGND.n2 9.3005
R81 VGND.n16 VGND.n15 9.3005
R82 VGND.n14 VGND.n3 9.3005
R83 VGND.n13 VGND.n12 9.3005
R84 VGND.n11 VGND.n4 9.3005
R85 VGND.n10 VGND.n9 9.3005
R86 VGND.n8 VGND.n6 7.10028
R87 VGND.n9 VGND.n8 0.218617
R88 VGND.n9 VGND.n4 0.120292
R89 VGND.n13 VGND.n4 0.120292
R90 VGND.n14 VGND.n13 0.120292
R91 VGND.n15 VGND.n14 0.120292
R92 VGND.n15 VGND.n2 0.120292
R93 VGND.n20 VGND.n2 0.120292
R94 VGND.n21 VGND.n20 0.120292
R95 VGND.n22 VGND.n21 0.120292
R96 VGND.n22 VGND 0.11899
R97 VGND VGND.n24 0.0213333
R98 VGND.n24 VGND 0.00180208
R99 a_674_413.t0 a_674_413.t1 98.5005
R100 a_716_21.t1 a_716_21.n5 406.075
R101 a_716_21.n4 a_716_21.t7 368.329
R102 a_716_21.n0 a_716_21.t2 268.365
R103 a_716_21.n3 a_716_21.t0 234.9
R104 a_716_21.n1 a_716_21.t3 212.081
R105 a_716_21.n0 a_716_21.t5 175.179
R106 a_716_21.n3 a_716_21.n2 174.109
R107 a_716_21.n5 a_716_21.n4 167.151
R108 a_716_21.n4 a_716_21.t6 149.822
R109 a_716_21.n1 a_716_21.t4 139.78
R110 a_716_21.n2 a_716_21.n0 130.725
R111 a_716_21.n5 a_716_21.n3 61.2126
R112 a_716_21.n2 a_716_21.n1 5.84292
R113 a_1124_47.t1 a_1124_47.n1 669.563
R114 a_1124_47.n1 a_1124_47.t0 248.404
R115 a_1124_47.n0 a_1124_47.t2 241.536
R116 a_1124_47.n1 a_1124_47.n0 174.691
R117 a_1124_47.n0 a_1124_47.t3 169.237
R118 VPWR.n12 VPWR.t1 670.534
R119 VPWR.n24 VPWR.n1 604.394
R120 VPWR.n8 VPWR.n7 318.728
R121 VPWR.n10 VPWR.n9 316.502
R122 VPWR.n19 VPWR.n4 311.356
R123 VPWR.n7 VPWR.t3 58.4849
R124 VPWR.n1 VPWR.t8 41.5552
R125 VPWR.n1 VPWR.t6 41.5552
R126 VPWR.n4 VPWR.t4 41.5552
R127 VPWR.n4 VPWR.t0 41.5552
R128 VPWR.n23 VPWR.n2 34.6358
R129 VPWR.n13 VPWR.n11 34.6358
R130 VPWR.n17 VPWR.n5 34.6358
R131 VPWR.n18 VPWR.n17 34.6358
R132 VPWR.n7 VPWR.t7 31.6057
R133 VPWR.n12 VPWR.n5 31.2476
R134 VPWR.n25 VPWR.n24 30.7593
R135 VPWR.n19 VPWR.n2 27.8593
R136 VPWR.n9 VPWR.t2 26.5955
R137 VPWR.n9 VPWR.t5 26.5955
R138 VPWR.n11 VPWR.n10 26.3534
R139 VPWR.n24 VPWR.n23 22.9652
R140 VPWR.n19 VPWR.n18 17.6946
R141 VPWR.n11 VPWR.n6 9.3005
R142 VPWR.n14 VPWR.n13 9.3005
R143 VPWR.n15 VPWR.n5 9.3005
R144 VPWR.n17 VPWR.n16 9.3005
R145 VPWR.n18 VPWR.n3 9.3005
R146 VPWR.n20 VPWR.n19 9.3005
R147 VPWR.n21 VPWR.n2 9.3005
R148 VPWR.n23 VPWR.n22 9.3005
R149 VPWR.n24 VPWR.n0 9.3005
R150 VPWR.n10 VPWR.n8 7.10028
R151 VPWR.n13 VPWR.n12 3.38874
R152 VPWR.n8 VPWR.n6 0.218617
R153 VPWR.n14 VPWR.n6 0.120292
R154 VPWR.n15 VPWR.n14 0.120292
R155 VPWR.n16 VPWR.n15 0.120292
R156 VPWR.n16 VPWR.n3 0.120292
R157 VPWR.n20 VPWR.n3 0.120292
R158 VPWR.n21 VPWR.n20 0.120292
R159 VPWR.n22 VPWR.n21 0.120292
R160 VPWR.n22 VPWR.n0 0.120292
R161 VPWR.n0 VPWR 0.11899
R162 VPWR VPWR.n25 0.0213333
R163 VPWR.n25 VPWR 0.00180208
R164 GATE_N.n0 GATE_N.t0 270.457
R165 GATE_N.n0 GATE_N.t1 235.109
R166 GATE_N.n1 GATE_N.n0 152
R167 GATE_N GATE_N.n1 11.2005
R168 GATE_N.n1 GATE_N 6.93383
R169 Q.n0 Q.t1 375.036
R170 Q.n1 Q.t0 209.923
R171 Q Q.n1 80.1887
R172 Q Q.n0 6.86263
R173 Q.n0 Q 5.86156
R174 Q.n1 Q 5.83579
R175 a_651_47.t0 a_651_47.t1 93.0601
R176 Q_N.n1 Q_N.t1 353.606
R177 Q_N.n0 Q_N.t0 209.923
R178 Q_N Q_N.n0 72.6418
R179 Q_N.n1 Q_N 9.10538
R180 Q_N Q_N.n1 7.47898
R181 Q_N.n0 Q_N 6.64665
R182 D.n0 D.t1 314.3
R183 D.n0 D.t0 157.544
R184 D D.n0 154.447
C0 VPB GATE_N 0.069748f
C1 VPB D 0.067771f
C2 VPB VPWR 0.163712f
C3 VPB VGND 0.016779f
C4 GATE_N VPWR 0.019079f
C5 D VPWR 0.014857f
C6 VPB Q 0.012499f
C7 GATE_N VGND 0.018898f
C8 D VGND 0.019229f
C9 VPB Q_N 0.011972f
C10 VPWR VGND 0.092294f
C11 VPWR Q 0.104256f
C12 VGND Q 0.043733f
C13 VPWR Q_N 0.093184f
C14 VGND Q_N 0.06408f
C15 Q_N VNB 0.095041f
C16 Q VNB 0.01145f
C17 VGND VNB 0.795325f
C18 VPWR VNB 0.639789f
C19 D VNB 0.136483f
C20 GATE_N VNB 0.19517f
C21 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxbn_2 VNB VPB VPWR VGND Q_N Q D GATE_N
X0 VPWR.t4 a_728_21.t2 Q.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t5 a_728_21.t3 a_663_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2 VPWR.t5 a_728_21.t4 a_686_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 Q_N.t1 a_1223_47.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.149 ps=1.325 w=1 l=0.15
X4 VPWR.t10 GATE_N.t0 a_27_47.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_686_413.t1 a_27_47.t2 a_565_413.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X6 VPWR.t1 a_1223_47.t3 Q_N.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X7 VGND.t4 a_728_21.t5 Q.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Q.t2 a_728_21.t6 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X9 VGND.t7 a_565_413.t4 a_728_21.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_193_47.t1 a_27_47.t3 VGND.t10 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 Q_N.t3 a_1223_47.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.097 ps=0.975 w=0.65 l=0.15
X12 VPWR.t2 a_728_21.t7 a_1223_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X13 a_663_47.t1 a_193_47.t2 a_565_413.t0 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X14 VGND.t2 a_728_21.t8 a_1223_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_469_369.t1 a_303_47.t2 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 VGND.t6 D.t0 a_303_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 a_193_47.t0 a_27_47.t4 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X18 VPWR.t6 D.t1 a_303_47.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X19 VGND.t1 a_1223_47.t5 Q_N.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.089375 ps=0.925 w=0.65 l=0.15
X20 a_565_413.t1 a_193_47.t3 a_469_369.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X21 VPWR.t9 a_565_413.t5 a_728_21.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X22 a_469_47.t1 a_303_47.t3 VGND.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 VGND.t8 GATE_N.t1 a_27_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_565_413.t2 a_27_47.t5 a_469_47.t0 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X25 Q.t0 a_728_21.t9 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
R0 a_728_21.t1 a_728_21.n0 395.272
R1 a_728_21.n5 a_728_21.t3 368.329
R2 a_728_21.n1 a_728_21.t7 247.542
R3 a_728_21.n4 a_728_21.t0 236.978
R4 a_728_21.n2 a_728_21.t2 212.081
R5 a_728_21.n3 a_728_21.t6 212.081
R6 a_728_21.n4 a_728_21.n3 176.689
R7 a_728_21.n0 a_728_21.n5 171.394
R8 a_728_21.n1 a_728_21.t8 154.356
R9 a_728_21.n5 a_728_21.t4 149.822
R10 a_728_21.n2 a_728_21.t5 139.78
R11 a_728_21.n3 a_728_21.t9 139.78
R12 a_728_21.n2 a_728_21.n1 118.309
R13 a_728_21.n3 a_728_21.n2 61.346
R14 a_728_21.n0 a_728_21.n4 17.7517
R15 Q.n0 Q 593.448
R16 Q.n1 Q.n0 585
R17 Q.n3 Q.n2 185
R18 Q Q.n3 26.7557
R19 Q.n0 Q.t3 26.5955
R20 Q.n0 Q.t2 26.5955
R21 Q.n2 Q.t1 24.9236
R22 Q.n2 Q.t0 24.9236
R23 Q.n1 Q 14.8485
R24 Q.n3 Q 7.9365
R25 Q Q.n1 2.5605
R26 VPWR.n5 VPWR.t5 666.241
R27 VPWR.n30 VPWR.n1 604.394
R28 VPWR.n8 VPWR.t4 341.087
R29 VPWR.n17 VPWR.n7 316.377
R30 VPWR.n11 VPWR.n10 312.632
R31 VPWR.n3 VPWR.n2 311.356
R32 VPWR.n9 VPWR.t1 256.253
R33 VPWR.n10 VPWR.t2 58.4849
R34 VPWR.n1 VPWR.t8 41.5552
R35 VPWR.n1 VPWR.t10 41.5552
R36 VPWR.n2 VPWR.t7 41.5552
R37 VPWR.n2 VPWR.t6 41.5552
R38 VPWR.n29 VPWR.n28 34.6358
R39 VPWR.n23 VPWR.n22 34.6358
R40 VPWR.n24 VPWR.n23 34.6358
R41 VPWR.n10 VPWR.t0 31.6057
R42 VPWR.n7 VPWR.t9 29.5505
R43 VPWR.n22 VPWR.n5 29.3652
R44 VPWR.n18 VPWR.n17 29.3652
R45 VPWR.n12 VPWR.n11 28.2358
R46 VPWR.n28 VPWR.n3 27.4829
R47 VPWR.n7 VPWR.t3 26.5955
R48 VPWR.n16 VPWR.n8 25.977
R49 VPWR.n30 VPWR.n29 22.9652
R50 VPWR.n12 VPWR.n8 22.9652
R51 VPWR.n17 VPWR.n16 18.4476
R52 VPWR.n24 VPWR.n3 18.0711
R53 VPWR.n18 VPWR.n5 17.3181
R54 VPWR.n13 VPWR.n12 9.3005
R55 VPWR.n14 VPWR.n8 9.3005
R56 VPWR.n16 VPWR.n15 9.3005
R57 VPWR.n17 VPWR.n6 9.3005
R58 VPWR.n19 VPWR.n18 9.3005
R59 VPWR.n20 VPWR.n5 9.3005
R60 VPWR.n22 VPWR.n21 9.3005
R61 VPWR.n23 VPWR.n4 9.3005
R62 VPWR.n25 VPWR.n24 9.3005
R63 VPWR.n26 VPWR.n3 9.3005
R64 VPWR.n28 VPWR.n27 9.3005
R65 VPWR.n29 VPWR.n0 9.3005
R66 VPWR.n31 VPWR.n30 7.12063
R67 VPWR.n11 VPWR.n9 6.32884
R68 VPWR.n13 VPWR.n9 0.664094
R69 VPWR.n31 VPWR.n0 0.148519
R70 VPWR.n14 VPWR.n13 0.120292
R71 VPWR.n15 VPWR.n14 0.120292
R72 VPWR.n15 VPWR.n6 0.120292
R73 VPWR.n19 VPWR.n6 0.120292
R74 VPWR.n20 VPWR.n19 0.120292
R75 VPWR.n21 VPWR.n20 0.120292
R76 VPWR.n21 VPWR.n4 0.120292
R77 VPWR.n25 VPWR.n4 0.120292
R78 VPWR.n26 VPWR.n25 0.120292
R79 VPWR.n27 VPWR.n26 0.120292
R80 VPWR.n27 VPWR.n0 0.120292
R81 VPWR VPWR.n31 0.114842
R82 VPB.t10 VPB.t7 568.225
R83 VPB.t5 VPB.t2 556.386
R84 VPB.t4 VPB.t11 556.386
R85 VPB.t6 VPB.t9 358.101
R86 VPB.t8 VPB.t6 284.113
R87 VPB.t2 VPB.t0 281.154
R88 VPB.t11 VPB.t3 257.478
R89 VPB.t0 VPB.t1 251.559
R90 VPB.t3 VPB.t5 248.599
R91 VPB.t7 VPB.t8 248.599
R92 VPB.t12 VPB.t10 248.599
R93 VPB.t9 VPB.t4 213.084
R94 VPB VPB.t12 192.369
R95 a_663_47.t0 a_663_47.t1 93.0601
R96 VGND.n6 VGND.t4 286.092
R97 VGND.n4 VGND.t5 240.833
R98 VGND.n16 VGND.n15 209.702
R99 VGND.n9 VGND.n8 201.488
R100 VGND.n30 VGND.n29 199.739
R101 VGND.n2 VGND.n1 198.964
R102 VGND.n7 VGND.t1 161.489
R103 VGND.n8 VGND.t2 54.2862
R104 VGND.n1 VGND.t9 38.5719
R105 VGND.n1 VGND.t6 38.5719
R106 VGND.n29 VGND.t10 38.5719
R107 VGND.n29 VGND.t8 38.5719
R108 VGND.n22 VGND.n21 34.6358
R109 VGND.n23 VGND.n22 34.6358
R110 VGND.n28 VGND.n27 34.6358
R111 VGND.n17 VGND.n16 29.3652
R112 VGND.n10 VGND.n9 28.2358
R113 VGND.n15 VGND.t7 27.6928
R114 VGND.n14 VGND.n6 25.977
R115 VGND.n8 VGND.t0 25.9346
R116 VGND.n15 VGND.t3 24.9236
R117 VGND.n21 VGND.n4 23.3417
R118 VGND.n10 VGND.n6 22.9652
R119 VGND.n23 VGND.n2 22.9652
R120 VGND.n30 VGND.n28 22.9652
R121 VGND.n27 VGND.n2 21.4593
R122 VGND.n17 VGND.n4 21.0829
R123 VGND.n16 VGND.n14 18.4476
R124 VGND.n28 VGND.n0 9.3005
R125 VGND.n27 VGND.n26 9.3005
R126 VGND.n25 VGND.n2 9.3005
R127 VGND.n24 VGND.n23 9.3005
R128 VGND.n22 VGND.n3 9.3005
R129 VGND.n21 VGND.n20 9.3005
R130 VGND.n19 VGND.n4 9.3005
R131 VGND.n11 VGND.n10 9.3005
R132 VGND.n12 VGND.n6 9.3005
R133 VGND.n14 VGND.n13 9.3005
R134 VGND.n16 VGND.n5 9.3005
R135 VGND.n18 VGND.n17 9.3005
R136 VGND.n31 VGND.n30 7.12063
R137 VGND.n9 VGND.n7 6.32884
R138 VGND.n11 VGND.n7 0.664094
R139 VGND.n31 VGND.n0 0.148519
R140 VGND.n12 VGND.n11 0.120292
R141 VGND.n13 VGND.n12 0.120292
R142 VGND.n13 VGND.n5 0.120292
R143 VGND.n18 VGND.n5 0.120292
R144 VGND.n19 VGND.n18 0.120292
R145 VGND.n20 VGND.n19 0.120292
R146 VGND.n20 VGND.n3 0.120292
R147 VGND.n24 VGND.n3 0.120292
R148 VGND.n25 VGND.n24 0.120292
R149 VGND.n26 VGND.n25 0.120292
R150 VGND.n26 VGND.n0 0.120292
R151 VGND VGND.n31 0.114842
R152 VNB.t11 VNB.t7 2733.98
R153 VNB.t4 VNB.t3 2677.02
R154 VNB.t5 VNB.t8 2677.02
R155 VNB.t10 VNB.t12 1537.86
R156 VNB.t3 VNB.t0 1352.75
R157 VNB.t6 VNB.t5 1352.75
R158 VNB.t8 VNB.t2 1238.83
R159 VNB.t12 VNB.t6 1224.6
R160 VNB.t0 VNB.t1 1210.36
R161 VNB.t2 VNB.t4 1196.12
R162 VNB.t7 VNB.t10 1196.12
R163 VNB.t9 VNB.t11 1196.12
R164 VNB VNB.t9 925.567
R165 a_686_413.t0 a_686_413.t1 98.5005
R166 a_1223_47.t0 a_1223_47.n2 386.31
R167 a_1223_47.n2 a_1223_47.t1 242.385
R168 a_1223_47.n1 a_1223_47.t2 239.04
R169 a_1223_47.n0 a_1223_47.t3 221.72
R170 a_1223_47.n2 a_1223_47.n1 175.274
R171 a_1223_47.n1 a_1223_47.t4 166.739
R172 a_1223_47.n0 a_1223_47.t5 149.421
R173 a_1223_47.n1 a_1223_47.n0 62.482
R174 Q_N Q_N.n0 586.758
R175 Q_N.n4 Q_N.n0 585
R176 Q_N.n2 Q_N.n1 185
R177 Q_N.n0 Q_N.t0 27.5805
R178 Q_N.n3 Q_N.n2 27.3215
R179 Q_N.n0 Q_N.t1 26.5955
R180 Q_N.n1 Q_N.t2 25.8467
R181 Q_N.n1 Q_N.t3 24.9236
R182 Q_N Q_N.n3 24.3815
R183 Q_N.n3 Q_N 16.8301
R184 Q_N Q_N.n4 15.3103
R185 Q_N.n2 Q_N 6.77697
R186 Q_N.n4 Q_N 1.75736
R187 GATE_N.n0 GATE_N.t0 270.457
R188 GATE_N.n0 GATE_N.t1 235.109
R189 GATE_N.n1 GATE_N.n0 152
R190 GATE_N GATE_N.n1 10.9719
R191 GATE_N.n1 GATE_N 6.79234
R192 a_27_47.t0 a_27_47.n3 415.863
R193 a_27_47.n2 a_27_47.t2 316.111
R194 a_27_47.n2 a_27_47.t5 315.729
R195 a_27_47.n1 a_27_47.t1 294.873
R196 a_27_47.n0 a_27_47.t4 263.173
R197 a_27_47.n0 a_27_47.t3 227.826
R198 a_27_47.n1 a_27_47.n0 152
R199 a_27_47.n3 a_27_47.n2 20.5885
R200 a_27_47.n3 a_27_47.n1 18.9713
R201 a_565_413.n3 a_565_413.n2 714.672
R202 a_565_413.n2 a_565_413.n1 282.507
R203 a_565_413.n2 a_565_413.n0 248.657
R204 a_565_413.n0 a_565_413.t5 212.081
R205 a_565_413.n0 a_565_413.t4 139.78
R206 a_565_413.t1 a_565_413.n3 121.953
R207 a_565_413.n3 a_565_413.t3 91.4648
R208 a_565_413.n1 a_565_413.t0 46.6672
R209 a_565_413.n1 a_565_413.t2 46.6672
R210 a_193_47.n0 a_193_47.t2 464.327
R211 a_193_47.t0 a_193_47.n1 366.837
R212 a_193_47.n1 a_193_47.t1 322.567
R213 a_193_47.n0 a_193_47.t3 242.607
R214 a_193_47.n1 a_193_47.n0 187.487
R215 a_303_47.t1 a_303_47.n1 438.971
R216 a_303_47.n0 a_303_47.t2 373.283
R217 a_303_47.n1 a_303_47.t0 275.149
R218 a_303_47.n1 a_303_47.n0 156.462
R219 a_303_47.n0 a_303_47.t3 132.282
R220 a_469_369.t1 a_469_369.t0 134.631
R221 D.n0 D.t1 327.644
R222 D.n0 D.t0 157.338
R223 D D.n0 154.595
R224 a_469_47.n0 a_469_47.t0 88.3338
R225 a_469_47.n0 a_469_47.t1 26.3935
R226 a_469_47.n1 a_469_47.n0 14.4005
C0 VPB VPWR 0.193155f
C1 GATE_N VPWR 0.019233f
C2 VPB VGND 0.018479f
C3 GATE_N VGND 0.019072f
C4 D VPWR 0.01407f
C5 VPB Q 0.007435f
C6 VPB Q_N 0.007306f
C7 D VGND 0.018822f
C8 VPWR VGND 0.115399f
C9 VPWR Q 0.190021f
C10 VPWR Q_N 0.200715f
C11 VGND Q 0.098487f
C12 VGND Q_N 0.144624f
C13 VPB GATE_N 0.069861f
C14 VPB D 0.062606f
C15 Q_N VNB 0.032832f
C16 Q VNB 0.00752f
C17 VGND VNB 0.921025f
C18 VPWR VNB 0.74275f
C19 D VNB 0.132945f
C20 GATE_N VNB 0.195334f
C21 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxbp_1 VGND VPWR VPB VNB Q_N Q D GATE
X0 a_560_47.t1 a_193_47.t2 a_465_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0549 pd=0.665 as=0.066 ps=0.745 w=0.36 l=0.15
X1 a_465_47.t1 a_299_47.t2 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR.t3 a_716_21.t2 a_1124_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 VPWR.t4 GATE.t0 a_27_47.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_467_369.t1 a_299_47.t3 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 a_560_47.t3 a_27_47.t2 a_467_369.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.09575 ps=0.965 w=0.42 l=0.15
X6 VGND.t6 a_560_47.t4 a_716_21.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR.t8 D.t0 a_299_47.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 Q.t1 a_716_21.t3 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_193_47.t1 a_27_47.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_651_47.t1 a_27_47.t4 a_560_47.t2 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0549 ps=0.665 w=0.36 l=0.15
X11 a_648_413.t0 a_193_47.t3 a_560_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 Q.t0 a_716_21.t4 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Q_N.t1 a_1124_47.t2 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X14 a_193_47.t0 a_27_47.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 VPWR.t7 a_560_47.t5 a_716_21.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 Q_N.t0 a_1124_47.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X17 VGND.t1 D.t1 a_299_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 VGND.t8 a_716_21.t5 a_1124_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 VPWR.t1 a_716_21.t6 a_648_413.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X20 VGND.t0 a_716_21.t7 a_651_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X21 VGND.t4 GATE.t1 a_27_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_193_47.n0 a_193_47.t2 383.005
R1 a_193_47.t0 a_193_47.n1 366.837
R2 a_193_47.n1 a_193_47.t1 322.567
R3 a_193_47.n0 a_193_47.t3 286.067
R4 a_193_47.n1 a_193_47.n0 25.1142
R5 a_465_47.n0 a_465_47.t0 66.6672
R6 a_465_47.n0 a_465_47.t1 26.3935
R7 a_465_47.n1 a_465_47.n0 14.4005
R8 a_560_47.n3 a_560_47.n2 709.649
R9 a_560_47.n2 a_560_47.n1 283.26
R10 a_560_47.n2 a_560_47.n0 246.466
R11 a_560_47.n0 a_560_47.t5 212.081
R12 a_560_47.n0 a_560_47.t4 139.78
R13 a_560_47.t0 a_560_47.n3 65.6672
R14 a_560_47.n3 a_560_47.t3 65.6672
R15 a_560_47.n1 a_560_47.t1 56.6672
R16 a_560_47.n1 a_560_47.t2 45.0005
R17 VNB.t9 VNB.t10 2677.02
R18 VNB.t2 VNB.t8 2677.02
R19 VNB.t5 VNB.t3 2677.02
R20 VNB.t10 VNB.t4 1352.75
R21 VNB.t1 VNB.t2 1352.75
R22 VNB.t7 VNB.t0 1352.75
R23 VNB.t0 VNB.t1 1295.79
R24 VNB.t8 VNB.t9 1196.12
R25 VNB.t3 VNB.t7 1196.12
R26 VNB.t6 VNB.t5 1196.12
R27 VNB VNB.t6 669.256
R28 a_299_47.t1 a_299_47.n1 400.163
R29 a_299_47.n0 a_299_47.t3 328.296
R30 a_299_47.n1 a_299_47.t0 260.538
R31 a_299_47.n0 a_299_47.t2 177.269
R32 a_299_47.n1 a_299_47.n0 152
R33 VGND.n4 VGND.t0 240.083
R34 VGND.n8 VGND.n7 213.161
R35 VGND.n6 VGND.n5 207.585
R36 VGND.n22 VGND.n21 199.739
R37 VGND.n2 VGND.n1 198.964
R38 VGND.n5 VGND.t8 54.2862
R39 VGND.n1 VGND.t5 38.5719
R40 VGND.n1 VGND.t1 38.5719
R41 VGND.n21 VGND.t3 38.5719
R42 VGND.n21 VGND.t4 38.5719
R43 VGND.n14 VGND.n13 34.6358
R44 VGND.n15 VGND.n14 34.6358
R45 VGND.n20 VGND.n19 34.6358
R46 VGND.n9 VGND.n8 26.3534
R47 VGND.n5 VGND.t2 25.9346
R48 VGND.n7 VGND.t7 24.9236
R49 VGND.n7 VGND.t6 24.9236
R50 VGND.n9 VGND.n4 24.4711
R51 VGND.n15 VGND.n2 24.4711
R52 VGND.n22 VGND.n20 22.9652
R53 VGND.n19 VGND.n2 19.9534
R54 VGND.n13 VGND.n4 18.824
R55 VGND.n20 VGND.n0 9.3005
R56 VGND.n19 VGND.n18 9.3005
R57 VGND.n17 VGND.n2 9.3005
R58 VGND.n16 VGND.n15 9.3005
R59 VGND.n14 VGND.n3 9.3005
R60 VGND.n13 VGND.n12 9.3005
R61 VGND.n11 VGND.n4 9.3005
R62 VGND.n10 VGND.n9 9.3005
R63 VGND.n23 VGND.n22 7.12063
R64 VGND.n8 VGND.n6 7.10028
R65 VGND.n10 VGND.n6 0.218617
R66 VGND.n23 VGND.n0 0.148519
R67 VGND.n11 VGND.n10 0.120292
R68 VGND.n12 VGND.n11 0.120292
R69 VGND.n12 VGND.n3 0.120292
R70 VGND.n16 VGND.n3 0.120292
R71 VGND.n17 VGND.n16 0.120292
R72 VGND.n18 VGND.n17 0.120292
R73 VGND.n18 VGND.n0 0.120292
R74 VGND VGND.n23 0.11354
R75 a_716_21.t0 a_716_21.n0 395.036
R76 a_716_21.n5 a_716_21.t7 367.543
R77 a_716_21.n1 a_716_21.t2 261.887
R78 a_716_21.n4 a_716_21.t1 233.504
R79 a_716_21.n2 a_716_21.t3 212.081
R80 a_716_21.n4 a_716_21.n3 176.048
R81 a_716_21.n0 a_716_21.n5 170.619
R82 a_716_21.n1 a_716_21.t5 168.701
R83 a_716_21.n5 a_716_21.t6 149.036
R84 a_716_21.n2 a_716_21.t4 139.78
R85 a_716_21.n3 a_716_21.n1 125.612
R86 a_716_21.n0 a_716_21.n4 18.1395
R87 a_716_21.n3 a_716_21.n2 7.30353
R88 a_1124_47.t0 a_1124_47.n1 669.563
R89 a_1124_47.n1 a_1124_47.t1 248.404
R90 a_1124_47.n0 a_1124_47.t2 239.04
R91 a_1124_47.n1 a_1124_47.n0 173.721
R92 a_1124_47.n0 a_1124_47.t3 166.739
R93 VPWR.n5 VPWR.t1 672.641
R94 VPWR.n22 VPWR.n1 604.394
R95 VPWR.n7 VPWR.n6 318.728
R96 VPWR.n9 VPWR.n8 316.377
R97 VPWR.n3 VPWR.n2 313.707
R98 VPWR.n6 VPWR.t3 58.4849
R99 VPWR.n1 VPWR.t0 41.5552
R100 VPWR.n1 VPWR.t4 41.5552
R101 VPWR.n2 VPWR.t5 41.5552
R102 VPWR.n2 VPWR.t8 41.5552
R103 VPWR.n21 VPWR.n20 34.6358
R104 VPWR.n15 VPWR.n14 34.6358
R105 VPWR.n16 VPWR.n15 34.6358
R106 VPWR.n6 VPWR.t6 31.6057
R107 VPWR.n10 VPWR.n5 29.3652
R108 VPWR.n20 VPWR.n3 26.7299
R109 VPWR.n8 VPWR.t2 26.5955
R110 VPWR.n8 VPWR.t7 26.5955
R111 VPWR.n14 VPWR.n5 24.8476
R112 VPWR.n10 VPWR.n9 23.7181
R113 VPWR.n22 VPWR.n21 22.9652
R114 VPWR.n16 VPWR.n3 21.4593
R115 VPWR.n11 VPWR.n10 9.3005
R116 VPWR.n12 VPWR.n5 9.3005
R117 VPWR.n14 VPWR.n13 9.3005
R118 VPWR.n15 VPWR.n4 9.3005
R119 VPWR.n17 VPWR.n16 9.3005
R120 VPWR.n18 VPWR.n3 9.3005
R121 VPWR.n20 VPWR.n19 9.3005
R122 VPWR.n21 VPWR.n0 9.3005
R123 VPWR.n23 VPWR.n22 7.12063
R124 VPWR.n9 VPWR.n7 7.10028
R125 VPWR.n11 VPWR.n7 0.218617
R126 VPWR.n23 VPWR.n0 0.148519
R127 VPWR.n12 VPWR.n11 0.120292
R128 VPWR.n13 VPWR.n12 0.120292
R129 VPWR.n13 VPWR.n4 0.120292
R130 VPWR.n17 VPWR.n4 0.120292
R131 VPWR.n18 VPWR.n17 0.120292
R132 VPWR.n19 VPWR.n18 0.120292
R133 VPWR.n19 VPWR.n0 0.120292
R134 VPWR VPWR.n23 0.11354
R135 VPB.t1 VPB.t10 562.306
R136 VPB.t3 VPB.t4 556.386
R137 VPB.t2 VPB.t9 556.386
R138 VPB.t0 VPB.t2 290.031
R139 VPB.t4 VPB.t8 281.154
R140 VPB.t7 VPB.t5 281.154
R141 VPB.t5 VPB.t0 254.518
R142 VPB.t9 VPB.t3 248.599
R143 VPB.t10 VPB.t7 248.599
R144 VPB.t6 VPB.t1 248.599
R145 VPB VPB.t6 139.097
R146 GATE.n0 GATE.t0 269.921
R147 GATE.n0 GATE.t1 234.573
R148 GATE.n1 GATE.n0 152
R149 GATE GATE.n1 10.9719
R150 GATE.n1 GATE 6.79234
R151 a_27_47.n2 a_27_47.t4 522.033
R152 a_27_47.t1 a_27_47.n3 415.863
R153 a_27_47.n1 a_27_47.t0 294.873
R154 a_27_47.n0 a_27_47.t5 263.173
R155 a_27_47.n0 a_27_47.t3 227.826
R156 a_27_47.n2 a_27_47.t2 219.042
R157 a_27_47.n3 a_27_47.n2 173.787
R158 a_27_47.n1 a_27_47.n0 152
R159 a_27_47.n3 a_27_47.n1 18.9713
R160 a_467_369.t1 a_467_369.t0 132.286
R161 D.n0 D.t0 393.534
R162 D.n0 D.t1 215.792
R163 D D.n0 154.595
R164 Q.n0 Q.t1 375.075
R165 Q Q.t0 249.798
R166 Q Q.n0 6.66813
R167 Q.n0 Q 5.6947
R168 a_651_47.t0 a_651_47.t1 93.0601
R169 a_648_413.t0 a_648_413.t1 159.476
R170 Q_N.n1 Q_N.t1 353.606
R171 Q_N.n0 Q_N.t0 209.923
R172 Q_N Q_N.n0 66.6967
R173 Q_N.n1 Q_N 9.10538
R174 Q_N Q_N.n1 7.47898
R175 Q_N.n0 Q_N 6.64665
C0 VPB GATE 0.070092f
C1 VPB D 0.079103f
C2 VPB VPWR 0.163405f
C3 GATE VPWR 0.019242f
C4 VPB VGND 0.016561f
C5 VPB Q 0.012712f
C6 GATE VGND 0.019085f
C7 D VPWR 0.015919f
C8 D VGND 0.021092f
C9 VPB Q_N 0.012f
C10 VPWR VGND 0.091033f
C11 VPWR Q 0.121666f
C12 VPWR Q_N 0.093352f
C13 VGND Q 0.089189f
C14 VGND Q_N 0.064368f
C15 Q_N VNB 0.094915f
C16 Q VNB 0.010388f
C17 VGND VNB 0.793185f
C18 VPWR VNB 0.631364f
C19 D VNB 0.152238f
C20 GATE VNB 0.195771f
C21 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtn_1 VGND VPWR VPB VNB Q D GATE_N
X0 VPWR.t0 D.t0 a_299_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47.t3 a_27_47.t2 a_465_47.t1 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.054 pd=0.66 as=0.066 ps=0.745 w=0.36 l=0.15
X2 a_465_47.t0 a_299_47.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR.t2 GATE_N.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VGND.t5 a_560_47.t4 a_715_21.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_193_47.t1 a_27_47.t3 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR.t3 a_560_47.t5 a_715_21.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7 a_650_47.t0 a_193_47.t2 a_560_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.054 ps=0.66 w=0.36 l=0.15
X8 Q.t0 a_715_21.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X9 a_193_47.t0 a_27_47.t4 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 VPWR.t5 a_715_21.t3 a_644_413.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 VGND.t0 D.t1 a_299_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 Q.t1 a_715_21.t4 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13 a_644_413.t1 a_27_47.t5 a_560_47.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_465_369.t0 a_299_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_560_47.t1 a_193_47.t3 a_465_369.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X16 VGND.t2 GATE_N.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t4 a_715_21.t5 a_650_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R0 D.n0 D.t0 344.363
R1 D.n0 D.t1 161.582
R2 D D.n0 154.595
R3 a_299_47.n0 a_299_47.t2 464.685
R4 a_299_47.t1 a_299_47.n1 430.467
R5 a_299_47.n0 a_299_47.t3 328.296
R6 a_299_47.n1 a_299_47.t0 276.702
R7 a_299_47.n1 a_299_47.n0 154.724
R8 VPWR.n5 VPWR.t5 663.521
R9 VPWR.n17 VPWR.n1 604.394
R10 VPWR.n7 VPWR.n6 322.038
R11 VPWR.n3 VPWR.n2 312.978
R12 VPWR.n1 VPWR.t6 41.5552
R13 VPWR.n1 VPWR.t2 41.5552
R14 VPWR.n2 VPWR.t1 41.5552
R15 VPWR.n2 VPWR.t0 41.5552
R16 VPWR.n16 VPWR.n15 34.6358
R17 VPWR.n10 VPWR.n9 34.6358
R18 VPWR.n11 VPWR.n10 34.6358
R19 VPWR.n6 VPWR.t3 34.4755
R20 VPWR.n6 VPWR.t4 26.5955
R21 VPWR.n15 VPWR.n3 25.977
R22 VPWR.n9 VPWR.n5 24.4711
R23 VPWR.n17 VPWR.n16 22.9652
R24 VPWR.n11 VPWR.n3 21.4593
R25 VPWR.n9 VPWR.n8 9.3005
R26 VPWR.n10 VPWR.n4 9.3005
R27 VPWR.n12 VPWR.n11 9.3005
R28 VPWR.n13 VPWR.n3 9.3005
R29 VPWR.n15 VPWR.n14 9.3005
R30 VPWR.n16 VPWR.n0 9.3005
R31 VPWR.n18 VPWR.n17 7.12063
R32 VPWR.n7 VPWR.n5 6.5678
R33 VPWR.n8 VPWR.n7 0.542133
R34 VPWR.n18 VPWR.n0 0.148519
R35 VPWR.n8 VPWR.n4 0.120292
R36 VPWR.n12 VPWR.n4 0.120292
R37 VPWR.n13 VPWR.n12 0.120292
R38 VPWR.n14 VPWR.n13 0.120292
R39 VPWR.n14 VPWR.n0 0.120292
R40 VPWR VPWR.n18 0.11354
R41 VPB.t5 VPB.t3 556.386
R42 VPB.t7 VPB.t0 556.386
R43 VPB.t8 VPB.t5 298.911
R44 VPB.t1 VPB.t6 281.154
R45 VPB.t3 VPB.t4 272.274
R46 VPB.t6 VPB.t8 248.599
R47 VPB.t0 VPB.t1 248.599
R48 VPB.t2 VPB.t7 248.599
R49 VPB VPB.t2 139.097
R50 a_27_47.t0 a_27_47.n3 415.863
R51 a_27_47.n2 a_27_47.t2 361.195
R52 a_27_47.n2 a_27_47.t5 297.034
R53 a_27_47.n1 a_27_47.t1 294.873
R54 a_27_47.n0 a_27_47.t4 263.173
R55 a_27_47.n0 a_27_47.t3 227.826
R56 a_27_47.n1 a_27_47.n0 152
R57 a_27_47.n3 a_27_47.n2 20.5885
R58 a_27_47.n3 a_27_47.n1 18.9713
R59 a_465_47.n0 a_465_47.t1 66.6672
R60 a_465_47.n0 a_465_47.t0 26.3935
R61 a_465_47.n1 a_465_47.n0 14.4005
R62 a_560_47.n3 a_560_47.n2 730.726
R63 a_560_47.n2 a_560_47.n1 264.459
R64 a_560_47.n2 a_560_47.n0 243.683
R65 a_560_47.n0 a_560_47.t5 212.081
R66 a_560_47.n0 a_560_47.t4 139.78
R67 a_560_47.n3 a_560_47.t2 63.3219
R68 a_560_47.t1 a_560_47.n3 63.3219
R69 a_560_47.n1 a_560_47.t0 55.0005
R70 a_560_47.n1 a_560_47.t3 45.0005
R71 VNB.t5 VNB.t6 2677.02
R72 VNB.t7 VNB.t1 2677.02
R73 VNB.t0 VNB.t5 1352.75
R74 VNB.t2 VNB.t8 1352.75
R75 VNB.t6 VNB.t4 1310.03
R76 VNB.t8 VNB.t0 1281.55
R77 VNB.t1 VNB.t2 1196.12
R78 VNB.t3 VNB.t7 1196.12
R79 VNB VNB.t3 669.256
R80 VGND.n4 VGND.t4 241.587
R81 VGND.n6 VGND.n5 222.159
R82 VGND.n17 VGND.n16 199.739
R83 VGND.n2 VGND.n1 198.964
R84 VGND.n1 VGND.t1 38.5719
R85 VGND.n1 VGND.t0 38.5719
R86 VGND.n16 VGND.t6 38.5719
R87 VGND.n16 VGND.t2 38.5719
R88 VGND.n9 VGND.n8 34.6358
R89 VGND.n10 VGND.n9 34.6358
R90 VGND.n15 VGND.n14 34.6358
R91 VGND.n5 VGND.t5 32.3082
R92 VGND.n5 VGND.t3 24.9236
R93 VGND.n8 VGND.n4 24.4711
R94 VGND.n10 VGND.n2 24.4711
R95 VGND.n17 VGND.n15 22.9652
R96 VGND.n14 VGND.n2 19.9534
R97 VGND.n15 VGND.n0 9.3005
R98 VGND.n14 VGND.n13 9.3005
R99 VGND.n12 VGND.n2 9.3005
R100 VGND.n11 VGND.n10 9.3005
R101 VGND.n9 VGND.n3 9.3005
R102 VGND.n8 VGND.n7 9.3005
R103 VGND.n18 VGND.n17 7.12063
R104 VGND.n6 VGND.n4 6.84171
R105 VGND.n7 VGND.n6 0.485732
R106 VGND.n18 VGND.n0 0.148519
R107 VGND.n7 VGND.n3 0.120292
R108 VGND.n11 VGND.n3 0.120292
R109 VGND.n12 VGND.n11 0.120292
R110 VGND.n13 VGND.n12 0.120292
R111 VGND.n13 VGND.n0 0.120292
R112 VGND VGND.n18 0.11354
R113 GATE_N.n0 GATE_N.t0 269.921
R114 GATE_N.n0 GATE_N.t1 234.573
R115 GATE_N.n1 GATE_N.n0 152
R116 GATE_N GATE_N.n1 10.9719
R117 GATE_N.n1 GATE_N 6.79234
R118 a_715_21.t0 a_715_21.n2 822.102
R119 a_715_21.t0 a_715_21.n4 759.269
R120 a_715_21.n3 a_715_21.t5 367.543
R121 a_715_21.n1 a_715_21.t1 246.042
R122 a_715_21.n0 a_715_21.t2 239.04
R123 a_715_21.n1 a_715_21.n0 173.528
R124 a_715_21.n4 a_715_21.n3 170.619
R125 a_715_21.n0 a_715_21.t4 166.739
R126 a_715_21.n3 a_715_21.t3 149.036
R127 a_715_21.n2 a_715_21.n1 17.3638
R128 a_715_21.n4 a_715_21.n2 1.35808
R129 a_193_47.n0 a_193_47.t2 562.716
R130 a_193_47.t0 a_193_47.n1 366.837
R131 a_193_47.n1 a_193_47.t1 322.567
R132 a_193_47.n0 a_193_47.t3 219.042
R133 a_193_47.n1 a_193_47.n0 185.101
R134 a_650_47.t1 a_650_47.t0 93.0601
R135 Q.n0 Q.t0 374.618
R136 Q.n1 Q.t1 209.923
R137 Q Q.n1 83.4322
R138 Q Q.n0 8.95158
R139 Q.n0 Q 7.65628
R140 Q.n1 Q 7.63127
R141 a_644_413.t0 a_644_413.t1 166.512
R142 a_465_369.t0 a_465_369.t1 132.286
C0 VPB GATE_N 0.070092f
C1 VPB D 0.071941f
C2 VPB VPWR 0.13016f
C3 GATE_N VPWR 0.019242f
C4 VPB VGND 0.012776f
C5 GATE_N VGND 0.019085f
C6 D VPWR 0.014335f
C7 VPB Q 0.011547f
C8 D VGND 0.018418f
C9 VPWR VGND 0.062945f
C10 VPWR Q 0.111042f
C11 VGND Q 0.053341f
C12 Q VNB 0.085917f
C13 VGND VNB 0.659055f
C14 VPWR VNB 0.518511f
C15 D VNB 0.140732f
C16 GATE_N VNB 0.195771f
C17 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtn_2 VNB VPB VPWR VGND Q D GATE_N
X0 VPWR.t4 a_728_21.t2 Q.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t5 a_728_21.t3 a_663_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2 VPWR.t5 a_728_21.t4 a_686_413.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR.t7 GATE_N.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_686_413.t0 a_27_47.t2 a_565_413.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X5 VGND.t4 a_728_21.t5 Q.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Q.t0 a_728_21.t6 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X7 VGND.t7 a_565_413.t4 a_728_21.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_193_47.t0 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_663_47.t1 a_193_47.t2 a_565_413.t1 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X10 a_469_369.t1 a_303_47.t2 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VGND.t2 D.t0 a_303_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_193_47.t1 a_27_47.t4 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 VPWR.t2 D.t1 a_303_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14 a_565_413.t0 a_193_47.t3 a_469_369.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X15 VPWR.t6 a_565_413.t5 a_728_21.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X16 a_469_47.t0 a_303_47.t3 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND.t6 GATE_N.t1 a_27_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_565_413.t2 a_27_47.t5 a_469_47.t1 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X19 Q.t2 a_728_21.t7 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
R0 a_728_21.t0 a_728_21.n0 395.272
R1 a_728_21.n4 a_728_21.t3 368.329
R2 a_728_21.n3 a_728_21.t1 236.978
R3 a_728_21.n1 a_728_21.t2 212.081
R4 a_728_21.n2 a_728_21.t6 212.081
R5 a_728_21.n3 a_728_21.n2 176.689
R6 a_728_21.n0 a_728_21.n4 171.394
R7 a_728_21.n4 a_728_21.t4 149.822
R8 a_728_21.n1 a_728_21.t5 139.78
R9 a_728_21.n2 a_728_21.t7 139.78
R10 a_728_21.n2 a_728_21.n1 61.346
R11 a_728_21.n0 a_728_21.n3 17.7517
R12 Q.n0 Q 593.448
R13 Q.n1 Q.n0 585
R14 Q.n3 Q.n2 185
R15 Q Q.n3 26.9563
R16 Q.n0 Q.t1 26.5955
R17 Q.n0 Q.t0 26.5955
R18 Q.n2 Q.t3 24.9236
R19 Q.n2 Q.t2 24.9236
R20 Q.n1 Q 14.8485
R21 Q.n3 Q 7.9365
R22 Q Q.n1 2.5605
R23 VPWR.n5 VPWR.t5 666.241
R24 VPWR.n21 VPWR.n1 604.394
R25 VPWR.n6 VPWR.t4 348.813
R26 VPWR.n8 VPWR.n7 316.377
R27 VPWR.n3 VPWR.n2 311.356
R28 VPWR.n1 VPWR.t0 41.5552
R29 VPWR.n1 VPWR.t7 41.5552
R30 VPWR.n2 VPWR.t1 41.5552
R31 VPWR.n2 VPWR.t2 41.5552
R32 VPWR.n20 VPWR.n19 34.6358
R33 VPWR.n14 VPWR.n13 34.6358
R34 VPWR.n15 VPWR.n14 34.6358
R35 VPWR.n7 VPWR.t6 29.5505
R36 VPWR.n13 VPWR.n5 29.3652
R37 VPWR.n9 VPWR.n8 29.3652
R38 VPWR.n19 VPWR.n3 27.4829
R39 VPWR.n7 VPWR.t3 26.5955
R40 VPWR.n21 VPWR.n20 22.9652
R41 VPWR.n15 VPWR.n3 18.0711
R42 VPWR.n9 VPWR.n5 17.3181
R43 VPWR.n10 VPWR.n9 9.3005
R44 VPWR.n11 VPWR.n5 9.3005
R45 VPWR.n13 VPWR.n12 9.3005
R46 VPWR.n14 VPWR.n4 9.3005
R47 VPWR.n16 VPWR.n15 9.3005
R48 VPWR.n17 VPWR.n3 9.3005
R49 VPWR.n19 VPWR.n18 9.3005
R50 VPWR.n20 VPWR.n0 9.3005
R51 VPWR.n22 VPWR.n21 7.12063
R52 VPWR.n8 VPWR.n6 6.29708
R53 VPWR.n10 VPWR.n6 0.669899
R54 VPWR.n22 VPWR.n0 0.148519
R55 VPWR.n11 VPWR.n10 0.120292
R56 VPWR.n12 VPWR.n11 0.120292
R57 VPWR.n12 VPWR.n4 0.120292
R58 VPWR.n16 VPWR.n4 0.120292
R59 VPWR.n17 VPWR.n16 0.120292
R60 VPWR.n18 VPWR.n17 0.120292
R61 VPWR.n18 VPWR.n0 0.120292
R62 VPWR VPWR.n22 0.11354
R63 VPB.t1 VPB.t3 568.225
R64 VPB.t5 VPB.t7 556.386
R65 VPB.t8 VPB.t0 358.101
R66 VPB.t2 VPB.t8 284.113
R67 VPB.t7 VPB.t4 257.478
R68 VPB.t4 VPB.t6 248.599
R69 VPB.t3 VPB.t2 248.599
R70 VPB.t9 VPB.t1 248.599
R71 VPB.t0 VPB.t5 213.084
R72 VPB VPB.t9 189.409
R73 a_663_47.t0 a_663_47.t1 93.0601
R74 VGND.n5 VGND.t4 293.67
R75 VGND.n4 VGND.t5 240.833
R76 VGND.n7 VGND.n6 209.702
R77 VGND.n21 VGND.n20 199.739
R78 VGND.n2 VGND.n1 198.964
R79 VGND.n1 VGND.t1 38.5719
R80 VGND.n1 VGND.t2 38.5719
R81 VGND.n20 VGND.t0 38.5719
R82 VGND.n20 VGND.t6 38.5719
R83 VGND.n13 VGND.n12 34.6358
R84 VGND.n14 VGND.n13 34.6358
R85 VGND.n19 VGND.n18 34.6358
R86 VGND.n8 VGND.n7 29.3652
R87 VGND.n6 VGND.t7 27.6928
R88 VGND.n6 VGND.t3 24.9236
R89 VGND.n12 VGND.n4 23.3417
R90 VGND.n14 VGND.n2 22.9652
R91 VGND.n21 VGND.n19 22.9652
R92 VGND.n18 VGND.n2 21.4593
R93 VGND.n8 VGND.n4 21.0829
R94 VGND.n19 VGND.n0 9.3005
R95 VGND.n18 VGND.n17 9.3005
R96 VGND.n16 VGND.n2 9.3005
R97 VGND.n15 VGND.n14 9.3005
R98 VGND.n13 VGND.n3 9.3005
R99 VGND.n12 VGND.n11 9.3005
R100 VGND.n10 VGND.n4 9.3005
R101 VGND.n9 VGND.n8 9.3005
R102 VGND.n22 VGND.n21 7.12063
R103 VGND.n7 VGND.n5 6.29708
R104 VGND.n9 VGND.n5 0.669899
R105 VGND.n22 VGND.n0 0.148519
R106 VGND.n10 VGND.n9 0.120292
R107 VGND.n11 VGND.n10 0.120292
R108 VGND.n11 VGND.n3 0.120292
R109 VGND.n15 VGND.n3 0.120292
R110 VGND.n16 VGND.n15 0.120292
R111 VGND.n17 VGND.n16 0.120292
R112 VGND.n17 VGND.n0 0.120292
R113 VGND VGND.n22 0.11354
R114 VNB.t0 VNB.t3 2733.98
R115 VNB.t6 VNB.t9 2677.02
R116 VNB.t2 VNB.t1 1537.86
R117 VNB.t7 VNB.t6 1352.75
R118 VNB.t9 VNB.t4 1238.83
R119 VNB.t1 VNB.t7 1224.6
R120 VNB.t4 VNB.t5 1196.12
R121 VNB.t3 VNB.t2 1196.12
R122 VNB.t8 VNB.t0 1196.12
R123 VNB VNB.t8 911.327
R124 a_686_413.t0 a_686_413.t1 98.5005
R125 GATE_N.n0 GATE_N.t0 269.921
R126 GATE_N.n0 GATE_N.t1 234.573
R127 GATE_N.n1 GATE_N.n0 152
R128 GATE_N GATE_N.n1 10.9719
R129 GATE_N.n1 GATE_N 6.79234
R130 a_27_47.t1 a_27_47.n3 415.863
R131 a_27_47.n2 a_27_47.t2 316.111
R132 a_27_47.n2 a_27_47.t5 315.729
R133 a_27_47.n1 a_27_47.t0 294.873
R134 a_27_47.n0 a_27_47.t4 263.173
R135 a_27_47.n0 a_27_47.t3 227.826
R136 a_27_47.n1 a_27_47.n0 152
R137 a_27_47.n3 a_27_47.n2 20.5885
R138 a_27_47.n3 a_27_47.n1 18.9713
R139 a_565_413.n3 a_565_413.n2 714.672
R140 a_565_413.n2 a_565_413.n1 282.507
R141 a_565_413.n2 a_565_413.n0 248.657
R142 a_565_413.n0 a_565_413.t5 212.081
R143 a_565_413.n0 a_565_413.t4 139.78
R144 a_565_413.t0 a_565_413.n3 121.953
R145 a_565_413.n3 a_565_413.t3 91.4648
R146 a_565_413.n1 a_565_413.t1 46.6672
R147 a_565_413.n1 a_565_413.t2 46.6672
R148 a_193_47.n0 a_193_47.t2 464.327
R149 a_193_47.t1 a_193_47.n1 366.837
R150 a_193_47.n1 a_193_47.t0 322.567
R151 a_193_47.n0 a_193_47.t3 242.607
R152 a_193_47.n1 a_193_47.n0 187.487
R153 a_303_47.t1 a_303_47.n1 438.971
R154 a_303_47.n0 a_303_47.t2 373.283
R155 a_303_47.n1 a_303_47.t0 275.149
R156 a_303_47.n1 a_303_47.n0 156.462
R157 a_303_47.n0 a_303_47.t3 132.282
R158 a_469_369.t1 a_469_369.t0 134.631
R159 D.n0 D.t1 327.644
R160 D.n0 D.t0 157.338
R161 D D.n0 154.595
R162 a_469_47.n0 a_469_47.t1 88.3338
R163 a_469_47.n0 a_469_47.t0 26.3935
R164 a_469_47.n1 a_469_47.n0 14.4005
C0 VPWR VGND 0.074005f
C1 VPWR Q 0.196602f
C2 VGND Q 0.098344f
C3 VPB VPWR 0.145747f
C4 GATE_N VPWR 0.019242f
C5 VPB VGND 0.013536f
C6 D VPWR 0.01407f
C7 GATE_N VGND 0.019085f
C8 VPB Q 0.007933f
C9 D VGND 0.018822f
C10 VPB GATE_N 0.070092f
C11 VPB D 0.062606f
C12 Q VNB 0.050004f
C13 VGND VNB 0.716623f
C14 VPWR VNB 0.582914f
C15 D VNB 0.132945f
C16 GATE_N VNB 0.195771f
C17 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtn_4 VNB VPB VPWR VGND Q D GATE_N
X0 VPWR.t2 D.t0 a_299_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 Q.t3 a_724_21.t2 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.1525 ps=1.305 w=1 l=0.15
X2 a_465_47.t0 a_299_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_561_413.t1 a_27_47.t2 a_465_47.t1 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X4 a_561_413.t2 a_193_47.t2 a_465_369.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X5 VGND.t9 a_724_21.t3 a_659_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6 Q.t7 a_724_21.t4 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.099125 ps=0.955 w=0.65 l=0.15
X7 VPWR.t4 GATE_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 Q.t2 a_724_21.t5 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X9 a_659_47.t0 a_193_47.t3 a_561_413.t3 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X10 VPWR.t7 a_724_21.t6 a_682_413.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 a_193_47.t1 a_27_47.t3 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_682_413.t0 a_27_47.t4 a_561_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X13 VPWR.t8 a_724_21.t7 Q.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.145 ps=1.29 w=1 l=0.15
X14 VGND.t7 a_724_21.t8 Q.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_193_47.t0 a_27_47.t5 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 VPWR.t1 a_561_413.t4 a_724_21.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X17 VGND.t2 a_561_413.t5 a_724_21.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VGND.t6 a_724_21.t9 Q.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.09425 ps=0.94 w=0.65 l=0.15
X19 Q.t4 a_724_21.t10 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X20 VGND.t1 D.t1 a_299_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VPWR.t9 a_724_21.t11 Q.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X22 a_465_369.t0 a_299_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND.t4 GATE_N.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 327.644
R1 D.n0 D.t1 157.338
R2 D D.n0 154.595
R3 a_299_47.t1 a_299_47.n1 438.971
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t0 275.149
R6 a_299_47.n1 a_299_47.n0 156.462
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n5 VPWR.t7 666.241
R9 VPWR.n26 VPWR.n1 604.394
R10 VPWR.n10 VPWR.t8 410.901
R11 VPWR.n9 VPWR.n8 320.228
R12 VPWR.n13 VPWR.n7 316.377
R13 VPWR.n3 VPWR.n2 311.356
R14 VPWR.n1 VPWR.t3 41.5552
R15 VPWR.n1 VPWR.t4 41.5552
R16 VPWR.n2 VPWR.t0 41.5552
R17 VPWR.n2 VPWR.t2 41.5552
R18 VPWR.n25 VPWR.n24 34.6358
R19 VPWR.n19 VPWR.n18 34.6358
R20 VPWR.n20 VPWR.n19 34.6358
R21 VPWR.n8 VPWR.t9 33.4905
R22 VPWR.n14 VPWR.n13 31.2476
R23 VPWR.n12 VPWR.n9 30.4946
R24 VPWR.n7 VPWR.t1 29.5505
R25 VPWR.n18 VPWR.n5 27.8593
R26 VPWR.n7 VPWR.t6 26.5955
R27 VPWR.n8 VPWR.t5 26.5955
R28 VPWR.n24 VPWR.n3 25.977
R29 VPWR.n26 VPWR.n25 22.9652
R30 VPWR.n20 VPWR.n3 19.577
R31 VPWR.n14 VPWR.n5 18.824
R32 VPWR.n13 VPWR.n12 16.5652
R33 VPWR.n12 VPWR.n11 9.3005
R34 VPWR.n13 VPWR.n6 9.3005
R35 VPWR.n15 VPWR.n14 9.3005
R36 VPWR.n16 VPWR.n5 9.3005
R37 VPWR.n18 VPWR.n17 9.3005
R38 VPWR.n19 VPWR.n4 9.3005
R39 VPWR.n21 VPWR.n20 9.3005
R40 VPWR.n22 VPWR.n3 9.3005
R41 VPWR.n24 VPWR.n23 9.3005
R42 VPWR.n25 VPWR.n0 9.3005
R43 VPWR.n27 VPWR.n26 7.12063
R44 VPWR.n10 VPWR.n9 6.4202
R45 VPWR.n11 VPWR.n10 0.647392
R46 VPWR.n27 VPWR.n0 0.148519
R47 VPWR.n11 VPWR.n6 0.120292
R48 VPWR.n15 VPWR.n6 0.120292
R49 VPWR.n16 VPWR.n15 0.120292
R50 VPWR.n17 VPWR.n16 0.120292
R51 VPWR.n17 VPWR.n4 0.120292
R52 VPWR.n21 VPWR.n4 0.120292
R53 VPWR.n22 VPWR.n21 0.120292
R54 VPWR.n23 VPWR.n22 0.120292
R55 VPWR.n23 VPWR.n0 0.120292
R56 VPWR VPWR.n27 0.114842
R57 VPB.t9 VPB.t1 583.023
R58 VPB.t5 VPB.t2 556.386
R59 VPB.t3 VPB.t4 358.101
R60 VPB.t0 VPB.t3 284.113
R61 VPB.t11 VPB.t7 269.315
R62 VPB.t7 VPB.t10 260.437
R63 VPB.t1 VPB.t8 257.478
R64 VPB.t8 VPB.t11 248.599
R65 VPB.t2 VPB.t0 248.599
R66 VPB.t6 VPB.t5 248.599
R67 VPB.t4 VPB.t9 213.084
R68 VPB VPB.t6 192.369
R69 a_724_21.t0 a_724_21.n0 395.272
R70 a_724_21.n6 a_724_21.t3 368.329
R71 a_724_21.n5 a_724_21.t1 238.347
R72 a_724_21.n1 a_724_21.t7 212.081
R73 a_724_21.n2 a_724_21.t2 212.081
R74 a_724_21.n3 a_724_21.t11 212.081
R75 a_724_21.n4 a_724_21.t5 212.081
R76 a_724_21.n5 a_724_21.n4 176.689
R77 a_724_21.n0 a_724_21.n6 173.139
R78 a_724_21.n6 a_724_21.t6 149.822
R79 a_724_21.n1 a_724_21.t9 139.78
R80 a_724_21.n2 a_724_21.t4 139.78
R81 a_724_21.n3 a_724_21.t8 139.78
R82 a_724_21.n4 a_724_21.t10 139.78
R83 a_724_21.n3 a_724_21.n2 66.4581
R84 a_724_21.n2 a_724_21.n1 64.2672
R85 a_724_21.n4 a_724_21.n3 61.346
R86 a_724_21.n0 a_724_21.n5 17.7517
R87 Q.n0 Q 592.412
R88 Q.n1 Q.n0 585
R89 Q.n5 Q.n4 291.046
R90 Q.n3 Q.n2 185
R91 Q.n7 Q.n6 185
R92 Q.n4 Q.t1 30.5355
R93 Q.n6 Q.t5 28.6159
R94 Q.n0 Q.t0 26.5955
R95 Q.n0 Q.t2 26.5955
R96 Q.n4 Q.t3 26.5955
R97 Q.n9 Q.n3 26.2346
R98 Q Q.n9 25.8251
R99 Q.n2 Q.t6 24.9236
R100 Q.n2 Q.t4 24.9236
R101 Q.n6 Q.t7 24.9236
R102 Q.n8 Q 21.8079
R103 Q.n8 Q 14.352
R104 Q.n1 Q 13.0251
R105 Q.n8 Q 10.9042
R106 Q Q.n7 10.1931
R107 Q.n9 Q 10.0853
R108 Q Q.n5 9.12101
R109 Q.n3 Q 6.9619
R110 Q.n5 Q 6.84089
R111 Q.n7 Q 5.92643
R112 Q Q.n8 3.49141
R113 Q Q.n1 2.24611
R114 VGND.n8 VGND.t6 243.911
R115 VGND.n4 VGND.t9 240.833
R116 VGND.n7 VGND.n6 213.161
R117 VGND.n12 VGND.n11 209.702
R118 VGND.n26 VGND.n25 199.739
R119 VGND.n2 VGND.n1 198.964
R120 VGND.n1 VGND.t0 38.5719
R121 VGND.n1 VGND.t1 38.5719
R122 VGND.n25 VGND.t3 38.5719
R123 VGND.n25 VGND.t4 38.5719
R124 VGND.n18 VGND.n17 34.6358
R125 VGND.n19 VGND.n18 34.6358
R126 VGND.n24 VGND.n23 34.6358
R127 VGND.n6 VGND.t7 31.3851
R128 VGND.n13 VGND.n12 31.2476
R129 VGND.n10 VGND.n7 30.4946
R130 VGND.n11 VGND.t2 27.6928
R131 VGND.n6 VGND.t8 24.9236
R132 VGND.n11 VGND.t5 24.9236
R133 VGND.n19 VGND.n2 24.4711
R134 VGND.n26 VGND.n24 22.9652
R135 VGND.n13 VGND.n4 22.5887
R136 VGND.n17 VGND.n4 21.8358
R137 VGND.n23 VGND.n2 19.9534
R138 VGND.n12 VGND.n10 16.5652
R139 VGND.n24 VGND.n0 9.3005
R140 VGND.n23 VGND.n22 9.3005
R141 VGND.n21 VGND.n2 9.3005
R142 VGND.n20 VGND.n19 9.3005
R143 VGND.n18 VGND.n3 9.3005
R144 VGND.n17 VGND.n16 9.3005
R145 VGND.n15 VGND.n4 9.3005
R146 VGND.n14 VGND.n13 9.3005
R147 VGND.n12 VGND.n5 9.3005
R148 VGND.n10 VGND.n9 9.3005
R149 VGND.n27 VGND.n26 7.12063
R150 VGND.n8 VGND.n7 6.4202
R151 VGND.n9 VGND.n8 0.647392
R152 VGND.n27 VGND.n0 0.148519
R153 VGND.n9 VGND.n5 0.120292
R154 VGND.n14 VGND.n5 0.120292
R155 VGND.n15 VGND.n14 0.120292
R156 VGND.n16 VGND.n15 0.120292
R157 VGND.n16 VGND.n3 0.120292
R158 VGND.n20 VGND.n3 0.120292
R159 VGND.n21 VGND.n20 0.120292
R160 VGND.n22 VGND.n21 0.120292
R161 VGND.n22 VGND.n0 0.120292
R162 VGND VGND.n27 0.114842
R163 a_465_47.n0 a_465_47.t1 88.3338
R164 a_465_47.n0 a_465_47.t0 26.3935
R165 a_465_47.n1 a_465_47.n0 14.4005
R166 VNB.t11 VNB.t3 2805.18
R167 VNB.t5 VNB.t1 2677.02
R168 VNB.t0 VNB.t4 1537.86
R169 VNB.t2 VNB.t11 1352.75
R170 VNB.t9 VNB.t10 1295.79
R171 VNB.t10 VNB.t8 1253.07
R172 VNB.t3 VNB.t7 1238.83
R173 VNB.t4 VNB.t2 1224.6
R174 VNB.t7 VNB.t9 1196.12
R175 VNB.t1 VNB.t0 1196.12
R176 VNB.t6 VNB.t5 1196.12
R177 VNB VNB.t6 925.567
R178 a_27_47.t0 a_27_47.n3 415.863
R179 a_27_47.n2 a_27_47.t4 316.111
R180 a_27_47.n2 a_27_47.t2 315.729
R181 a_27_47.n1 a_27_47.t1 294.873
R182 a_27_47.n0 a_27_47.t5 263.173
R183 a_27_47.n0 a_27_47.t3 227.826
R184 a_27_47.n1 a_27_47.n0 152
R185 a_27_47.n3 a_27_47.n2 20.5706
R186 a_27_47.n3 a_27_47.n1 18.9713
R187 a_561_413.n3 a_561_413.n2 714.672
R188 a_561_413.n2 a_561_413.n1 282.507
R189 a_561_413.n2 a_561_413.n0 255.231
R190 a_561_413.n0 a_561_413.t4 212.081
R191 a_561_413.n0 a_561_413.t5 139.78
R192 a_561_413.n3 a_561_413.t2 121.953
R193 a_561_413.t0 a_561_413.n3 91.4648
R194 a_561_413.n1 a_561_413.t3 46.6672
R195 a_561_413.n1 a_561_413.t1 46.6672
R196 a_193_47.n0 a_193_47.t3 464.327
R197 a_193_47.t0 a_193_47.n1 366.837
R198 a_193_47.n1 a_193_47.t1 322.567
R199 a_193_47.n0 a_193_47.t2 242.607
R200 a_193_47.n1 a_193_47.n0 187.469
R201 a_465_369.t0 a_465_369.t1 134.631
R202 a_659_47.t1 a_659_47.t0 93.0601
R203 GATE_N.n0 GATE_N.t0 269.921
R204 GATE_N.n0 GATE_N.t1 234.573
R205 GATE_N.n1 GATE_N.n0 152
R206 GATE_N GATE_N.n1 10.9719
R207 GATE_N.n1 GATE_N 6.79234
R208 a_682_413.t0 a_682_413.t1 98.5005
C0 GATE_N VGND 0.019085f
C1 D VPWR 0.014067f
C2 VPB Q 0.011781f
C3 D VGND 0.018848f
C4 VPWR VGND 0.09333f
C5 VPWR Q 0.460724f
C6 VGND Q 0.251721f
C7 VPB GATE_N 0.070092f
C8 VPB D 0.062359f
C9 VPB VPWR 0.164758f
C10 VPB VGND 0.014125f
C11 GATE_N VPWR 0.019242f
C12 Q VNB 0.042422f
C13 VGND VNB 0.813516f
C14 VPWR VNB 0.666829f
C15 D VNB 0.132433f
C16 GATE_N VNB 0.195771f
C17 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtp_1 VGND VPWR VPB VNB Q D GATE
X0 VPWR.t4 D.t0 a_299_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47.t1 a_193_47.t2 a_465_47.t0 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.066 ps=0.745 w=0.36 l=0.15
X2 VGND.t1 a_713_21.t2 a_659_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0936 pd=1.24 as=0.0486 ps=0.63 w=0.36 l=0.15
X3 Q.t0 a_713_21.t3 VGND.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.092625 ps=0.935 w=0.65 l=0.15
X4 a_465_47.t1 a_299_47.t2 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VPWR.t2 GATE.t0 a_27_47.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_659_47.t1 a_27_47.t2 a_560_47.t2 VNB.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0486 pd=0.63 as=0.0621 ps=0.705 w=0.36 l=0.15
X7 VGND.t6 a_560_47.t4 a_713_21.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR.t6 a_713_21.t4 a_644_413.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.07245 ps=0.765 w=0.42 l=0.15
X9 a_193_47.t0 a_27_47.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR.t5 a_560_47.t5 a_713_21.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X11 a_193_47.t1 a_27_47.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 Q.t1 a_713_21.t5 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.1425 ps=1.285 w=1 l=0.15
X13 VGND.t5 D.t1 a_299_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14 a_644_413.t1 a_193_47.t3 a_560_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_465_369.t1 a_299_47.t3 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X16 a_560_47.t3 a_27_47.t5 a_465_369.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X17 VGND.t3 GATE.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 D.n0 D.t0 327.644
R1 D.n0 D.t1 157.338
R2 D D.n0 154.595
R3 a_299_47.t1 a_299_47.n1 438.971
R4 a_299_47.n0 a_299_47.t3 373.283
R5 a_299_47.n1 a_299_47.t0 275.149
R6 a_299_47.n1 a_299_47.n0 156.462
R7 a_299_47.n0 a_299_47.t2 132.282
R8 VPWR.n5 VPWR.t6 678.236
R9 VPWR.n17 VPWR.n1 604.394
R10 VPWR.n7 VPWR.n6 331.558
R11 VPWR.n3 VPWR.n2 311.356
R12 VPWR.n1 VPWR.t0 41.5552
R13 VPWR.n1 VPWR.t2 41.5552
R14 VPWR.n2 VPWR.t1 41.5552
R15 VPWR.n2 VPWR.t4 41.5552
R16 VPWR.n16 VPWR.n15 34.6358
R17 VPWR.n10 VPWR.n9 34.6358
R18 VPWR.n11 VPWR.n10 34.6358
R19 VPWR.n9 VPWR.n5 30.8711
R20 VPWR.n6 VPWR.t5 29.5505
R21 VPWR.n6 VPWR.t3 26.5955
R22 VPWR.n15 VPWR.n3 25.977
R23 VPWR.n17 VPWR.n16 22.9652
R24 VPWR.n11 VPWR.n3 19.577
R25 VPWR.n7 VPWR.n5 11.0462
R26 VPWR.n9 VPWR.n8 9.3005
R27 VPWR.n10 VPWR.n4 9.3005
R28 VPWR.n12 VPWR.n11 9.3005
R29 VPWR.n13 VPWR.n3 9.3005
R30 VPWR.n15 VPWR.n14 9.3005
R31 VPWR.n16 VPWR.n0 9.3005
R32 VPWR.n18 VPWR.n17 7.12063
R33 VPWR.n8 VPWR.n7 0.453238
R34 VPWR.n18 VPWR.n0 0.148519
R35 VPWR.n8 VPWR.n4 0.120292
R36 VPWR.n12 VPWR.n4 0.120292
R37 VPWR.n13 VPWR.n12 0.120292
R38 VPWR.n14 VPWR.n13 0.120292
R39 VPWR.n14 VPWR.n0 0.120292
R40 VPWR VPWR.n18 0.114842
R41 VPB.t7 VPB.t6 562.306
R42 VPB.t0 VPB.t5 556.386
R43 VPB.t8 VPB.t7 292.991
R44 VPB.t2 VPB.t1 281.154
R45 VPB.t6 VPB.t4 257.478
R46 VPB.t1 VPB.t8 248.599
R47 VPB.t5 VPB.t2 248.599
R48 VPB.t3 VPB.t0 248.599
R49 VPB VPB.t3 142.056
R50 a_193_47.t1 a_193_47.n1 366.837
R51 a_193_47.n0 a_193_47.t2 328.108
R52 a_193_47.n1 a_193_47.t0 322.567
R53 a_193_47.n0 a_193_47.t3 300.252
R54 a_193_47.n1 a_193_47.n0 25.054
R55 a_465_47.n0 a_465_47.t0 66.6672
R56 a_465_47.n0 a_465_47.t1 26.3935
R57 a_465_47.n1 a_465_47.n0 14.4005
R58 a_560_47.n3 a_560_47.n2 721.871
R59 a_560_47.n2 a_560_47.n1 279.872
R60 a_560_47.n2 a_560_47.n0 246.489
R61 a_560_47.n0 a_560_47.t5 212.081
R62 a_560_47.n0 a_560_47.t4 139.78
R63 a_560_47.n1 a_560_47.t1 68.3338
R64 a_560_47.t0 a_560_47.n3 63.3219
R65 a_560_47.n3 a_560_47.t3 63.3219
R66 a_560_47.n1 a_560_47.t2 46.6672
R67 VNB.t0 VNB.t7 2705.5
R68 VNB.t3 VNB.t6 2677.02
R69 VNB.t1 VNB.t2 1409.71
R70 VNB.t5 VNB.t1 1352.75
R71 VNB.t7 VNB.t8 1238.83
R72 VNB.t2 VNB.t0 1196.12
R73 VNB.t6 VNB.t5 1196.12
R74 VNB.t4 VNB.t3 1196.12
R75 VNB VNB.t4 683.495
R76 a_713_21.t1 a_713_21.n0 395.272
R77 a_713_21.n3 a_713_21.t2 375.961
R78 a_713_21.n1 a_713_21.t5 241.536
R79 a_713_21.n2 a_713_21.t0 238.347
R80 a_713_21.n2 a_713_21.n1 174.498
R81 a_713_21.n0 a_713_21.n3 169.649
R82 a_713_21.n1 a_713_21.t3 169.237
R83 a_713_21.n3 a_713_21.t4 147.814
R84 a_713_21.n0 a_713_21.n2 17.7517
R85 a_659_47.t0 a_659_47.t1 90.0005
R86 VGND.n4 VGND.t1 247.262
R87 VGND.n6 VGND.n5 225.21
R88 VGND.n17 VGND.n16 199.739
R89 VGND.n2 VGND.n1 198.964
R90 VGND.n1 VGND.t4 38.5719
R91 VGND.n1 VGND.t5 38.5719
R92 VGND.n16 VGND.t2 38.5719
R93 VGND.n16 VGND.t3 38.5719
R94 VGND.n9 VGND.n8 34.6358
R95 VGND.n10 VGND.n9 34.6358
R96 VGND.n15 VGND.n14 34.6358
R97 VGND.n5 VGND.t6 27.6928
R98 VGND.n5 VGND.t0 24.9236
R99 VGND.n10 VGND.n2 24.4711
R100 VGND.n17 VGND.n15 22.9652
R101 VGND.n14 VGND.n2 19.9534
R102 VGND.n8 VGND.n4 17.6946
R103 VGND.n15 VGND.n0 9.3005
R104 VGND.n14 VGND.n13 9.3005
R105 VGND.n12 VGND.n2 9.3005
R106 VGND.n11 VGND.n10 9.3005
R107 VGND.n9 VGND.n3 9.3005
R108 VGND.n8 VGND.n7 9.3005
R109 VGND.n18 VGND.n17 7.12063
R110 VGND.n6 VGND.n4 6.91327
R111 VGND.n7 VGND.n6 0.513852
R112 VGND.n18 VGND.n0 0.148519
R113 VGND.n7 VGND.n3 0.120292
R114 VGND.n11 VGND.n3 0.120292
R115 VGND.n12 VGND.n11 0.120292
R116 VGND.n13 VGND.n12 0.120292
R117 VGND.n13 VGND.n0 0.120292
R118 VGND VGND.n18 0.114842
R119 Q.n0 Q 592.412
R120 Q.n1 Q.n0 585
R121 Q.n2 Q.t0 214.538
R122 Q Q.n2 82.223
R123 Q.n0 Q.t1 31.5205
R124 Q.n1 Q 13.0251
R125 Q.n2 Q 6.9619
R126 Q Q.n1 2.24611
R127 GATE.n0 GATE.t0 270.457
R128 GATE.n0 GATE.t1 235.109
R129 GATE.n1 GATE.n0 152
R130 GATE GATE.n1 11.2005
R131 GATE.n1 GATE 6.93383
R132 a_27_47.n2 a_27_47.t2 425.945
R133 a_27_47.t1 a_27_47.n3 415.863
R134 a_27_47.n1 a_27_47.t0 294.873
R135 a_27_47.n0 a_27_47.t4 263.173
R136 a_27_47.n0 a_27_47.t3 227.826
R137 a_27_47.n2 a_27_47.t5 219.042
R138 a_27_47.n3 a_27_47.n2 176.62
R139 a_27_47.n1 a_27_47.n0 152
R140 a_27_47.n3 a_27_47.n1 18.9713
R141 a_644_413.t0 a_644_413.t1 161.821
R142 a_465_369.t1 a_465_369.t0 132.286
C0 VPB VGND 0.013865f
C1 GATE VPWR 0.019079f
C2 GATE VGND 0.018898f
C3 D VPWR 0.014067f
C4 VPB Q 0.011783f
C5 D VGND 0.018848f
C6 VPWR VGND 0.062839f
C7 VPWR Q 0.100486f
C8 VGND Q 0.052621f
C9 VPB GATE 0.069748f
C10 VPB D 0.062359f
C11 VPB VPWR 0.131202f
C12 Q VNB 0.08476f
C13 VGND VNB 0.659888f
C14 VPWR VNB 0.523436f
C15 D VNB 0.132433f
C16 GATE VNB 0.19517f
C17 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd1_1 VPWR VGND VPB VNB X A
X0 X.t1 a_299_93.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1 VPWR.t1 a_193_47.t2 a_299_93.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t2 A.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_193_47.t0 a_27_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_193_47.t1 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND.t2 a_193_47.t3 a_299_93.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X.t0 a_299_93.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_299_93.t0 a_299_93.n1 716.485
R1 a_299_93.n1 a_299_93.t1 271.241
R2 a_299_93.n0 a_299_93.t3 238.59
R3 a_299_93.n0 a_299_93.t2 166.291
R4 a_299_93.n1 a_299_93.n0 152
R5 VGND.n2 VGND.n0 213.603
R6 VGND.n2 VGND.n1 208.339
R7 VGND.n1 VGND.t2 58.5719
R8 VGND.n0 VGND.t0 38.5719
R9 VGND.n0 VGND.t1 38.5719
R10 VGND.n1 VGND.t3 24.0005
R11 VGND VGND.n2 0.197535
R12 X X.n0 589.186
R13 X.n2 X.n0 585
R14 X.n1 X.t1 209.923
R15 X X.n1 78.6279
R16 X.n0 X.t0 26.5955
R17 X X.n2 12.5543
R18 X.n2 X 4.18512
R19 X.n1 X 3.75222
R20 VNB.t0 VNB.t2 2677.02
R21 VNB.t2 VNB.t3 1381.23
R22 VNB.t1 VNB.t0 1196.12
R23 VNB VNB.t1 939.807
R24 a_193_47.n1 a_193_47.t1 721.572
R25 a_193_47.t0 a_193_47.n1 268.964
R26 a_193_47.n0 a_193_47.t2 206.69
R27 a_193_47.n1 a_193_47.n0 177.28
R28 a_193_47.n0 a_193_47.t3 119.93
R29 VPWR.n2 VPWR.n0 616.504
R30 VPWR.n2 VPWR.n1 613.605
R31 VPWR.n0 VPWR.t1 89.1195
R32 VPWR.n1 VPWR.t0 63.3219
R33 VPWR.n1 VPWR.t2 63.3219
R34 VPWR.n0 VPWR.t3 37.3146
R35 VPWR VPWR.n2 0.196563
R36 VPB.t0 VPB.t1 562.306
R37 VPB.t1 VPB.t3 281.154
R38 VPB.t2 VPB.t0 248.599
R39 VPB VPB.t2 195.327
R40 A.n0 A.t0 326.762
R41 A.n0 A.t1 198.228
R42 A.n1 A.n0 152
R43 A.n1 A 7.7622
R44 A A.n1 1.49837
R45 a_27_47.t0 a_27_47.n1 729.926
R46 a_27_47.n0 a_27_47.t3 334.723
R47 a_27_47.n1 a_27_47.t1 285.538
R48 a_27_47.n0 a_27_47.t2 206.19
R49 a_27_47.n1 a_27_47.n0 152
C0 VPB A 0.07869f
C1 VPB VPWR 0.08957f
C2 VPB X 0.019387f
C3 A VPWR 0.017834f
C4 VPB VGND 0.015112f
C5 VPWR X 0.085284f
C6 A VGND 0.018684f
C7 VPWR VGND 0.066675f
C8 X VGND 0.06793f
C9 VGND VNB 0.408705f
C10 X VNB 0.084601f
C11 VPWR VNB 0.335714f
C12 A VNB 0.182357f
C13 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd2_1 VPB VNB VGND VPWR X A
X0 VPWR.t3 A.t0 a_49_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR.t2 a_221_47.t2 a_327_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.18
X2 X.t1 a_327_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3 VGND.t3 A.t1 a_49_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X.t0 a_327_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X5 a_221_47.t1 a_49_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.18
X6 a_221_47.t0 a_49_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.18
X7 VGND.t2 a_221_47.t3 a_327_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.18
R0 A.n0 A.t0 322.188
R1 A.n0 A.t1 193.655
R2 A.n1 A.n0 152
R3 A.n1 A 6.75606
R4 A A.n1 1.3042
R5 a_49_47.t0 a_49_47.n1 714.768
R6 a_49_47.n0 a_49_47.t3 283.844
R7 a_49_47.n1 a_49_47.t1 274.098
R8 a_49_47.n0 a_49_47.t2 176.733
R9 a_49_47.n1 a_49_47.n0 152
R10 VPWR.n2 VPWR.n1 608.726
R11 VPWR.n2 VPWR.n0 605.726
R12 VPWR.n0 VPWR.t2 75.0481
R13 VPWR.n1 VPWR.t1 63.3219
R14 VPWR.n1 VPWR.t3 63.3219
R15 VPWR.n0 VPWR.t0 43.3874
R16 VPWR VPWR.n2 0.207476
R17 VPB.t1 VPB.t2 574.144
R18 VPB.t2 VPB.t0 290.031
R19 VPB.t3 VPB.t1 257.478
R20 VPB VPB.t3 257.478
R21 a_221_47.t0 a_221_47.n1 702.812
R22 a_221_47.n0 a_221_47.t2 272.062
R23 a_221_47.n1 a_221_47.t1 268.517
R24 a_221_47.n0 a_221_47.t3 164.952
R25 a_221_47.n1 a_221_47.n0 152
R26 a_327_47.t0 a_327_47.n1 724.922
R27 a_327_47.n1 a_327_47.t1 281.724
R28 a_327_47.n0 a_327_47.t3 241.536
R29 a_327_47.n0 a_327_47.t2 169.237
R30 a_327_47.n1 a_327_47.n0 152
R31 VGND.n2 VGND.n0 208.726
R32 VGND.n2 VGND.n1 205.726
R33 VGND.n1 VGND.t2 45.7148
R34 VGND.n0 VGND.t0 38.5719
R35 VGND.n0 VGND.t3 38.5719
R36 VGND.n1 VGND.t1 34.506
R37 VGND VGND.n2 0.207671
R38 X.n0 X 586.927
R39 X.n1 X.n0 585
R40 X.n3 X.t1 209.923
R41 X.n0 X.t0 26.5955
R42 X X.n4 7.7918
R43 X.n2 X 6.57041
R44 X.n1 X 5.77749
R45 X X.n3 5.77749
R46 X X.n1 1.92616
R47 X.n3 X 1.92616
R48 X.n4 X 1.67007
R49 X X.n2 1.3918
R50 X.n4 X 1.35979
R51 X.n2 X 1.13324
R52 VNB.t0 VNB.t2 2762.46
R53 VNB.t2 VNB.t1 1395.47
R54 VNB.t3 VNB.t0 1238.83
R55 VNB VNB.t3 1238.83
C0 VPB VGND 0.007731f
C1 A VGND 0.018415f
C2 VPWR X 0.105065f
C3 VPWR VGND 0.062504f
C4 X VGND 0.104492f
C5 VPB A 0.087159f
C6 VPB VPWR 0.073796f
C7 VPB X 0.023807f
C8 A VPWR 0.017617f
C9 VGND VNB 0.397454f
C10 X VNB 0.103025f
C11 VPWR VNB 0.330896f
C12 A VNB 0.1896f
C13 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR.t0 A.t0 a_49_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND.t0 a_285_47.t2 a_391_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X.t0 a_391_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND.t1 A.t1 a_49_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR.t2 a_285_47.t3 a_391_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47.t1 a_49_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47.t0 a_49_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X.t1 a_391_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
R0 A.n0 A.t0 331.777
R1 A.n0 A.t1 203.244
R2 A.n1 A.n0 152
R3 A A.n1 7.88621
R4 A.n1 A 2.62907
R5 a_49_47.n1 a_49_47.t1 733.438
R6 a_49_47.t0 a_49_47.n1 293.175
R7 a_49_47.n1 a_49_47.n0 152
R8 a_49_47.n0 a_49_47.t3 107.487
R9 a_49_47.n0 a_49_47.t2 68.9265
R10 VPWR.n2 VPWR.n1 608.769
R11 VPWR.n2 VPWR.n0 606.074
R12 VPWR.n0 VPWR.t2 75.0481
R13 VPWR.n1 VPWR.t1 63.3219
R14 VPWR.n1 VPWR.t0 63.3219
R15 VPWR.n0 VPWR.t3 43.3874
R16 VPWR VPWR.n2 0.163864
R17 VPB.t1 VPB.t2 763.552
R18 VPB.t2 VPB.t3 384.736
R19 VPB.t0 VPB.t1 352.182
R20 VPB VPB.t0 257.478
R21 a_285_47.t0 a_285_47.n1 672.681
R22 a_285_47.n1 a_285_47.t1 242.239
R23 a_285_47.n1 a_285_47.n0 171.719
R24 a_285_47.n0 a_285_47.t3 107.487
R25 a_285_47.n0 a_285_47.t2 68.9265
R26 a_391_47.t0 a_391_47.n1 706.611
R27 a_391_47.n1 a_391_47.t1 276.81
R28 a_391_47.n0 a_391_47.t2 241.536
R29 a_391_47.n0 a_391_47.t3 169.237
R30 a_391_47.n1 a_391_47.n0 152.776
R31 VGND.n2 VGND.n1 208.769
R32 VGND.n2 VGND.n0 206.075
R33 VGND.n0 VGND.t0 45.7148
R34 VGND.n1 VGND.t3 38.5719
R35 VGND.n1 VGND.t1 38.5719
R36 VGND.n0 VGND.t2 34.506
R37 VGND VGND.n2 0.164057
R38 VNB.t3 VNB.t0 3673.79
R39 VNB.t0 VNB.t2 1851.13
R40 VNB.t1 VNB.t3 1694.5
R41 VNB VNB.t1 1238.83
R42 X X.t0 758.308
R43 X.n0 X.t1 209.923
R44 X X.n1 12.8005
R45 X.n2 X 9.64206
R46 X X.n0 8.47842
R47 X.n0 X 2.82647
R48 X.n1 X 2.74336
R49 X.n2 X 2.28621
R50 X.n1 X 1.99531
R51 X X.n2 1.66284
C0 VPB A 0.082837f
C1 VPB VPWR 0.0787f
C2 VPB X 0.015496f
C3 A VPWR 0.020643f
C4 VPB VGND 0.007167f
C5 A VGND 0.021393f
C6 VPWR X 0.080229f
C7 VPWR VGND 0.071507f
C8 X VGND 0.07961f
C9 VGND VNB 0.43965f
C10 X VNB 0.095447f
C11 VPWR VNB 0.367348f
C12 A VNB 0.178652f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlymetal6s2s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB X A
X0 a_558_47.t0 a_381_47.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND.t2 X.t2 a_381_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47.t1 a_664_47.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR.t2 A.t0 a_62_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND.t5 A.t1 a_62_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47.t1 a_381_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X.t0 a_62_47.t2 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR.t5 X.t3 a_381_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47.t0 a_664_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X.t1 a_62_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR.t3 a_558_47.t2 a_664_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND.t4 a_558_47.t3 a_664_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_381_47.n1 a_381_47.t1 705.896
R1 a_381_47.t0 a_381_47.n1 269.426
R2 a_381_47.n0 a_381_47.t2 241.536
R3 a_381_47.n0 a_381_47.t3 169.237
R4 a_381_47.n1 a_381_47.n0 152
R5 VPWR.n5 VPWR.n4 591.333
R6 VPWR.n11 VPWR.n10 585
R7 VPWR.n3 VPWR.n2 585
R8 VPWR.n4 VPWR.t3 77.3934
R9 VPWR.n2 VPWR.t5 77.3934
R10 VPWR.n10 VPWR.t2 77.3934
R11 VPWR.n4 VPWR.t1 41.0422
R12 VPWR.n2 VPWR.t0 41.0422
R13 VPWR.n10 VPWR.t4 41.0422
R14 VPWR.n8 VPWR.n1 34.6358
R15 VPWR.n9 VPWR.n8 34.6358
R16 VPWR.n3 VPWR.n1 20.3837
R17 VPWR.n12 VPWR.n11 11.8541
R18 VPWR.n11 VPWR.n9 9.73495
R19 VPWR.n6 VPWR.n1 9.3005
R20 VPWR.n8 VPWR.n7 9.3005
R21 VPWR.n9 VPWR.n0 9.3005
R22 VPWR.n5 VPWR.n3 8.3181
R23 VPWR.n6 VPWR.n5 0.219762
R24 VPWR.n12 VPWR.n0 0.141672
R25 VPWR VPWR.n12 0.128288
R26 VPWR.n7 VPWR.n6 0.120292
R27 VPWR.n7 VPWR.n0 0.120292
R28 a_558_47.t0 a_558_47.n1 364.868
R29 a_558_47.n0 a_558_47.t2 323.55
R30 a_558_47.n1 a_558_47.t1 246.088
R31 a_558_47.n0 a_558_47.t3 195.017
R32 a_558_47.n1 a_558_47.n0 152
R33 VPB.t3 VPB.t4 662.928
R34 VPB.t0 VPB.t5 556.386
R35 VPB VPB.t2 310.748
R36 VPB.t5 VPB.t1 281.154
R37 VPB.t4 VPB.t0 281.154
R38 VPB.t2 VPB.t3 281.154
R39 X.n0 X 590.271
R40 X.n1 X.n0 585
R41 X.n2 X.t3 323.55
R42 X.n5 X.t1 209.923
R43 X.n2 X.t2 195.017
R44 X X.n2 153.409
R45 X.n0 X.t0 26.5955
R46 X.n3 X 16.7116
R47 X.n3 X 16.0005
R48 X X.n5 9.78874
R49 X.n4 X 6.34564
R50 X X.n3 6.0165
R51 X.n3 X 5.7605
R52 X X.n1 5.27109
R53 X.n1 X 4.96991
R54 X.n4 X 2.19479
R55 X X.n4 1.80756
R56 X.n5 X 0.452265
R57 VGND.n5 VGND.n4 191.421
R58 VGND.n3 VGND.n2 185
R59 VGND.n11 VGND.n10 185
R60 VGND.n10 VGND.t5 45.7148
R61 VGND.n2 VGND.t2 45.7148
R62 VGND.n4 VGND.t4 45.7148
R63 VGND.n8 VGND.n1 34.6358
R64 VGND.n9 VGND.n8 34.6358
R65 VGND.n10 VGND.t3 34.506
R66 VGND.n2 VGND.t0 34.506
R67 VGND.n4 VGND.t1 34.506
R68 VGND.n3 VGND.n1 20.4554
R69 VGND.n12 VGND.n11 11.9258
R70 VGND.n11 VGND.n9 10.0265
R71 VGND.n6 VGND.n1 9.3005
R72 VGND.n8 VGND.n7 9.3005
R73 VGND.n9 VGND.n0 9.3005
R74 VGND.n5 VGND.n3 8.4829
R75 VGND.n6 VGND.n5 0.220277
R76 VGND.n12 VGND.n0 0.141672
R77 VGND VGND.n12 0.128288
R78 VGND.n7 VGND.n6 0.120292
R79 VGND.n7 VGND.n0 0.120292
R80 VNB.t3 VNB.t2 3189.64
R81 VNB.t0 VNB.t4 2677.02
R82 VNB VNB.t5 1495.15
R83 VNB.t4 VNB.t1 1352.75
R84 VNB.t2 VNB.t0 1352.75
R85 VNB.t5 VNB.t3 1352.75
R86 a_664_47.n1 a_664_47.t1 707.12
R87 a_664_47.t0 a_664_47.n1 269.426
R88 a_664_47.n0 a_664_47.t2 241.536
R89 a_664_47.n0 a_664_47.t3 169.237
R90 a_664_47.n1 a_664_47.n0 152
R91 a_841_47.t1 a_841_47.t0 621.348
R92 A.n0 A.t0 323.55
R93 A.n0 A.t1 195.017
R94 A.n1 A.n0 152
R95 A.n1 A 7.52215
R96 A A.n1 1.45205
R97 a_62_47.n1 a_62_47.t1 704.678
R98 a_62_47.t0 a_62_47.n1 264.865
R99 a_62_47.n0 a_62_47.t2 241.536
R100 a_62_47.n0 a_62_47.t3 169.237
R101 a_62_47.n1 a_62_47.n0 152
C0 A VPWR 0.017441f
C1 VPB VGND 0.008004f
C2 A VGND 0.017615f
C3 VPB A 0.104964f
C4 X VPWR 0.107956f
C5 X VGND 0.106174f
C6 VPWR VGND 0.090191f
C7 VPB X 0.1257f
C8 A X 0.014223f
C9 VPB VPWR 0.102518f
C10 VGND VNB 0.536721f
C11 VPWR VNB 0.439129f
C12 X VNB 0.162711f
C13 A VNB 0.198339f
C14 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlymetal6s4s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlymetal6s4s_1 VPWR VGND VPB VNB X A
X0 X.t1 a_345_47.t2 VGND.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 VPWR.t1 a_239_47.t2 a_345_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47.t0 a_664_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND.t1 a_239_47.t3 a_345_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR.t0 A.t0 a_62_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t0 A.t1 a_62_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X.t0 a_345_47.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 a_239_47.t0 a_62_47.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8 a_841_47.t1 a_664_47.t3 VGND.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 a_239_47.t1 a_62_47.t3 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR.t5 X.t2 a_664_47.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND.t2 X.t3 a_664_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_345_47.n1 a_345_47.t1 707.457
R1 a_345_47.t0 a_345_47.n1 269.728
R2 a_345_47.n0 a_345_47.t3 241.536
R3 a_345_47.n0 a_345_47.t2 169.237
R4 a_345_47.n1 a_345_47.n0 152
R5 VGND.n5 VGND.n4 191.435
R6 VGND.n3 VGND.n2 185
R7 VGND.n11 VGND.n10 185
R8 VGND.n10 VGND.t0 45.7148
R9 VGND.n2 VGND.t1 45.7148
R10 VGND.n4 VGND.t2 45.7148
R11 VGND.n8 VGND.n1 34.6358
R12 VGND.n9 VGND.n8 34.6358
R13 VGND.n10 VGND.t3 34.506
R14 VGND.n2 VGND.t5 34.506
R15 VGND.n4 VGND.t4 34.506
R16 VGND.n5 VGND.n3 14.9325
R17 VGND.n12 VGND.n11 11.9258
R18 VGND.n11 VGND.n9 10.0265
R19 VGND.n6 VGND.n1 9.3005
R20 VGND.n8 VGND.n7 9.3005
R21 VGND.n9 VGND.n0 9.3005
R22 VGND.n3 VGND.n1 6.90246
R23 VGND.n6 VGND.n5 0.206034
R24 VGND.n12 VGND.n0 0.141672
R25 VGND VGND.n12 0.128288
R26 VGND.n7 VGND.n6 0.120292
R27 VGND.n7 VGND.n0 0.120292
R28 X.n0 X 590.034
R29 X.n1 X.n0 585
R30 X.n2 X.t2 323.55
R31 X.n6 X.t1 209.923
R32 X.n2 X.t3 195.017
R33 X X.n2 153.792
R34 X.n0 X.t0 26.5955
R35 X.n3 X 17.7783
R36 X.n3 X 14.9338
R37 X X.n6 9.34881
R38 X.n4 X.n3 5.8885
R39 X.n5 X.n4 5.88158
R40 X.n3 X 5.3765
R41 X X.n1 5.03421
R42 X.n1 X 4.74657
R43 X.n5 X 2.07618
R44 X X.n5 1.72634
R45 X.n4 X 0.5125
R46 X.n6 X 0.431961
R47 VNB.t4 VNB.t5 3189.64
R48 VNB.t2 VNB.t1 2677.02
R49 VNB VNB.t0 1495.15
R50 VNB.t5 VNB.t3 1352.75
R51 VNB.t1 VNB.t4 1352.75
R52 VNB.t0 VNB.t2 1352.75
R53 a_239_47.t0 a_239_47.n1 362.024
R54 a_239_47.n0 a_239_47.t2 323.55
R55 a_239_47.n1 a_239_47.t1 242.583
R56 a_239_47.n0 a_239_47.t3 195.017
R57 a_239_47.n1 a_239_47.n0 152
R58 VPWR.n5 VPWR.n4 591.348
R59 VPWR.n11 VPWR.n10 585
R60 VPWR.n3 VPWR.n2 585
R61 VPWR.n4 VPWR.t5 77.3934
R62 VPWR.n2 VPWR.t1 77.3934
R63 VPWR.n10 VPWR.t0 77.3934
R64 VPWR.n4 VPWR.t3 41.0422
R65 VPWR.n2 VPWR.t4 41.0422
R66 VPWR.n10 VPWR.t2 41.0422
R67 VPWR.n8 VPWR.n1 34.6358
R68 VPWR.n9 VPWR.n8 34.6358
R69 VPWR.n5 VPWR.n3 14.6416
R70 VPWR.n12 VPWR.n11 11.8541
R71 VPWR.n11 VPWR.n9 9.73495
R72 VPWR.n6 VPWR.n1 9.3005
R73 VPWR.n8 VPWR.n7 9.3005
R74 VPWR.n9 VPWR.n0 9.3005
R75 VPWR.n3 VPWR.n1 6.83075
R76 VPWR.n6 VPWR.n5 0.205339
R77 VPWR.n12 VPWR.n0 0.141672
R78 VPWR VPWR.n12 0.128288
R79 VPWR.n7 VPWR.n6 0.120292
R80 VPWR.n7 VPWR.n0 0.120292
R81 VPB.t4 VPB.t5 662.928
R82 VPB.t2 VPB.t1 556.386
R83 VPB VPB.t0 310.748
R84 VPB.t5 VPB.t3 281.154
R85 VPB.t1 VPB.t4 281.154
R86 VPB.t0 VPB.t2 281.154
R87 a_664_47.t0 a_664_47.n1 707.12
R88 a_664_47.n1 a_664_47.t1 269.426
R89 a_664_47.n0 a_664_47.t2 241.536
R90 a_664_47.n0 a_664_47.t3 169.237
R91 a_664_47.n1 a_664_47.n0 152
R92 a_841_47.t0 a_841_47.t1 621.348
R93 A.n0 A.t0 323.55
R94 A.n0 A.t1 195.017
R95 A.n1 A.n0 152
R96 A.n1 A 7.52215
R97 A A.n1 1.45205
R98 a_62_47.t0 a_62_47.n1 704.678
R99 a_62_47.n1 a_62_47.t1 264.865
R100 a_62_47.n0 a_62_47.t2 241.536
R101 a_62_47.n0 a_62_47.t3 169.237
R102 a_62_47.n1 a_62_47.n0 152
C0 X VPWR 0.111451f
C1 A VGND 0.017615f
C2 X VGND 0.109054f
C3 VPWR VGND 0.090168f
C4 VPB A 0.104121f
C5 VPB X 0.124968f
C6 VPB VPWR 0.100625f
C7 A VPWR 0.017441f
C8 VPB VGND 0.007842f
C9 VGND VNB 0.538104f
C10 VPWR VNB 0.442872f
C11 X VNB 0.174165f
C12 A VNB 0.198004f
C13 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlymetal6s6s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND VPB VNB X A
X0 X.t0 a_629_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 a_523_47.t0 a_346_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2 VGND.t5 a_240_47.t2 a_346_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_240_47.t0 a_63_47.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VPWR.t0 a_240_47.t3 a_346_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t2 A.t0 a_63_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR.t5 A.t1 a_63_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR.t4 a_523_47.t2 a_629_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND.t0 a_523_47.t3 a_629_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_523_47.t1 a_346_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X10 a_240_47.t1 a_63_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X11 X.t1 a_629_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
R0 a_629_47.t0 a_629_47.n1 706.186
R1 a_629_47.n1 a_629_47.t1 268.589
R2 a_629_47.n0 a_629_47.t3 241.536
R3 a_629_47.n0 a_629_47.t2 169.237
R4 a_629_47.n1 a_629_47.n0 152
R5 VGND.n6 VGND.n5 192.263
R6 VGND.n4 VGND.n3 185
R7 VGND.n1 VGND.n0 185
R8 VGND.n0 VGND.t2 45.7148
R9 VGND.n3 VGND.t5 45.7148
R10 VGND.n5 VGND.t0 45.7148
R11 VGND.n9 VGND.n8 34.6358
R12 VGND.n10 VGND.n9 34.6358
R13 VGND.n0 VGND.t4 34.506
R14 VGND.n3 VGND.t3 34.506
R15 VGND.n5 VGND.t1 34.506
R16 VGND.n6 VGND.n4 14.4956
R17 VGND.n12 VGND.n1 12.3022
R18 VGND.n10 VGND.n1 9.65004
R19 VGND.n8 VGND.n7 9.3005
R20 VGND.n9 VGND.n2 9.3005
R21 VGND.n11 VGND.n10 9.3005
R22 VGND.n8 VGND.n4 7.27893
R23 VGND.n7 VGND.n6 0.265833
R24 VGND.n12 VGND.n11 0.141672
R25 VGND VGND.n12 0.126986
R26 VGND.n7 VGND.n2 0.120292
R27 VGND.n11 VGND.n2 0.120292
R28 X.n0 X 590.149
R29 X.n1 X.n0 585
R30 X.n4 X.t0 209.923
R31 X.n0 X.t1 26.5955
R32 X.n3 X 9.95606
R33 X.n4 X 9.56372
R34 X.n2 X 8.53383
R35 X X.n1 5.14993
R36 X.n1 X 4.85567
R37 X.n3 X 2.13383
R38 X X.n2 1.77828
R39 X X.n3 1.76602
R40 X.n2 X 1.47176
R41 X X.n4 0.441879
R42 VNB.t3 VNB.t0 2677.02
R43 VNB.t4 VNB.t5 2677.02
R44 VNB VNB.t2 1495.15
R45 VNB.t0 VNB.t1 1352.75
R46 VNB.t5 VNB.t3 1352.75
R47 VNB.t2 VNB.t4 1352.75
R48 a_346_47.t0 a_346_47.n1 707.457
R49 a_346_47.n1 a_346_47.t1 269.728
R50 a_346_47.n0 a_346_47.t3 241.536
R51 a_346_47.n0 a_346_47.t2 169.237
R52 a_346_47.n1 a_346_47.n0 152
R53 a_523_47.t1 a_523_47.n1 364.13
R54 a_523_47.n0 a_523_47.t2 323.55
R55 a_523_47.n1 a_523_47.t0 245.32
R56 a_523_47.n0 a_523_47.t3 195.017
R57 a_523_47.n1 a_523_47.n0 152
R58 a_240_47.t1 a_240_47.n1 362.024
R59 a_240_47.n0 a_240_47.t3 323.55
R60 a_240_47.n1 a_240_47.t0 242.583
R61 a_240_47.n0 a_240_47.t2 195.017
R62 a_240_47.n1 a_240_47.n0 152
R63 a_63_47.n1 a_63_47.t1 704.572
R64 a_63_47.t0 a_63_47.n1 264.767
R65 a_63_47.n0 a_63_47.t3 241.536
R66 a_63_47.n0 a_63_47.t2 169.237
R67 a_63_47.n1 a_63_47.n0 152
R68 VPWR.n5 VPWR.n4 592.152
R69 VPWR.n11 VPWR.n10 585
R70 VPWR.n3 VPWR.n2 585
R71 VPWR.n4 VPWR.t4 77.3934
R72 VPWR.n2 VPWR.t0 77.3934
R73 VPWR.n10 VPWR.t5 77.3934
R74 VPWR.n4 VPWR.t2 41.0422
R75 VPWR.n2 VPWR.t3 41.0422
R76 VPWR.n10 VPWR.t1 41.0422
R77 VPWR.n8 VPWR.n1 34.6358
R78 VPWR.n9 VPWR.n8 34.6358
R79 VPWR.n5 VPWR.n3 14.2054
R80 VPWR.n12 VPWR.n11 12.2305
R81 VPWR.n11 VPWR.n9 9.35848
R82 VPWR.n6 VPWR.n1 9.3005
R83 VPWR.n8 VPWR.n7 9.3005
R84 VPWR.n9 VPWR.n0 9.3005
R85 VPWR.n3 VPWR.n1 7.20722
R86 VPWR.n6 VPWR.n5 0.264419
R87 VPWR.n12 VPWR.n0 0.141672
R88 VPWR VPWR.n12 0.126986
R89 VPWR.n7 VPWR.n6 0.120292
R90 VPWR.n7 VPWR.n0 0.120292
R91 VPB.t3 VPB.t4 556.386
R92 VPB.t1 VPB.t0 556.386
R93 VPB VPB.t5 310.748
R94 VPB.t4 VPB.t2 281.154
R95 VPB.t0 VPB.t3 281.154
R96 VPB.t5 VPB.t1 281.154
R97 A.n0 A.t1 323.55
R98 A.n0 A.t0 195.017
R99 A.n1 A.n0 152
R100 A.n1 A 7.4454
R101 A A.n1 1.43723
C0 VPWR X 0.086118f
C1 A VGND 0.017536f
C2 VPWR VGND 0.090168f
C3 X VGND 0.083173f
C4 VPB A 0.104303f
C5 VPB VPWR 0.098471f
C6 A VPWR 0.017356f
C7 VPB X 0.01886f
C8 VPB VGND 0.007892f
C9 VGND VNB 0.538855f
C10 X VNB 0.100265f
C11 VPWR VNB 0.446134f
C12 A VNB 0.197984f
C13 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_1 VNB VPB VPWR VGND Z TE_B A
X0 Z.t1 a_27_47.t2 a_383_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.475 ps=1.95 w=1 l=0.15
X1 a_193_369.t1 TE_B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.2583 pd=2.07 as=0.098125 ps=1.005 w=0.42 l=0.15
X2 a_383_297.t0 TE_B.t1 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=1.95 as=0.27 ps=2.54 w=1 l=0.15
X3 VPWR.t2 A.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_531_47.t0 a_193_369.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.2275 ps=2 w=0.65 l=0.15
X5 Z.t0 a_27_47.t3 a_531_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.286 pd=2.18 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 a_193_369.t0 TE_B.t2 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7 VGND.t2 A.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.098125 pd=1.005 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t1 a_27_47.n1 722.542
R1 a_27_47.n1 a_27_47.n0 329.921
R2 a_27_47.n1 a_27_47.t0 248.082
R3 a_27_47.n0 a_27_47.t2 241.536
R4 a_27_47.n0 a_27_47.t3 169.237
R5 a_383_297.t0 a_383_297.t1 187.15
R6 Z.n3 Z.t1 329.93
R7 Z.n0 Z 186.77
R8 Z.n1 Z.n0 185
R9 Z.n0 Z.t0 50.7697
R10 Z Z.n2 10.5417
R11 Z.n1 Z 7.48986
R12 Z Z.n3 3.89328
R13 Z.n2 Z 2.25932
R14 Z.n3 Z 2.17782
R15 Z Z.n1 1.77071
R16 Z.n2 Z 1.63454
R17 VPB.t0 VPB.t3 651.091
R18 VPB.t2 VPB.t0 562.306
R19 VPB.t1 VPB.t2 248.599
R20 VPB VPB.t1 189.409
R21 TE_B.n1 TE_B.t1 323.817
R22 TE_B.n0 TE_B.t2 282.336
R23 TE_B.n2 TE_B.n1 152
R24 TE_B.n0 TE_B.t0 102.828
R25 TE_B.n1 TE_B.n0 14.6066
R26 TE_B.n2 TE_B 11.055
R27 TE_B TE_B.n2 2.13383
R28 VGND.n1 VGND.t1 233.887
R29 VGND.n1 VGND.n0 205.831
R30 VGND.n0 VGND.t0 88.798
R31 VGND.n0 VGND.t2 38.5724
R32 VGND VGND.n1 0.167388
R33 a_193_369.t0 a_193_369.n0 676.302
R34 a_193_369.n0 a_193_369.t2 351.382
R35 a_193_369.n0 a_193_369.t1 337.998
R36 VNB.t0 VNB.t2 4570.87
R37 VNB.t1 VNB.t0 1438.19
R38 VNB.t2 VNB.t3 1025.24
R39 VNB VNB.t1 911.327
R40 VPWR.n1 VPWR.t1 807.249
R41 VPWR.n1 VPWR.n0 604.366
R42 VPWR.n0 VPWR.t0 41.5552
R43 VPWR.n0 VPWR.t2 41.5552
R44 VPWR VPWR.n1 0.471431
R45 A.n0 A.t0 289.318
R46 A.n0 A.t1 196.131
R47 A.n1 A.n0 152
R48 A.n1 A 13.5116
R49 A A.n1 2.60791
R50 a_531_47.t0 a_531_47.t1 38.7697
C0 VPB VGND 0.007748f
C1 VPB A 0.064652f
C2 A VGND 0.01737f
C3 VPB TE_B 0.127958f
C4 TE_B VGND 0.0199f
C5 VPB VPWR 0.082415f
C6 A TE_B 0.064835f
C7 VPWR VGND 0.070492f
C8 A VPWR 0.017206f
C9 TE_B VPWR 0.04252f
C10 VPB Z 0.029612f
C11 Z VGND 0.101739f
C12 A Z 1.04e-19
C13 TE_B Z 0.00859f
C14 VPWR Z 0.243182f
C15 VGND VNB 0.442579f
C16 Z VNB 0.097664f
C17 VPWR VNB 0.361695f
C18 TE_B VNB 0.22258f
C19 A VNB 0.195718f
C20 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_2 VNB VPB VGND VPWR A TE_B Z
X0 a_320_309.t3 a_27_47.t2 Z.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Z.t0 a_27_47.t3 a_320_309.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37025 ps=1.745 w=1 l=0.15
X2 VPWR.t3 A.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.015 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 VGND.t3 a_214_47.t2 a_392_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_214_47.t1 TE_B.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12 ps=1.015 w=0.64 l=0.15
X5 a_320_309.t1 TE_B.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.37025 pd=1.745 as=0.1269 ps=1.21 w=0.94 l=0.15
X6 a_392_47.t2 a_214_47.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR.t0 TE_B.t2 a_320_309.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.2444 ps=2.4 w=0.94 l=0.15
X8 Z.t3 a_27_47.t4 a_392_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X9 a_214_47.t0 TE_B.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07875 ps=0.795 w=0.42 l=0.15
X10 a_392_47.t0 a_27_47.t5 Z.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t1 A.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.07875 pd=0.795 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t0 a_27_47.n3 680.693
R1 a_27_47.n3 a_27_47.t1 263.26
R2 a_27_47.n0 a_27_47.t2 221.72
R3 a_27_47.n1 a_27_47.t3 221.72
R4 a_27_47.n3 a_27_47.n2 174.32
R5 a_27_47.n0 a_27_47.t5 149.421
R6 a_27_47.n1 a_27_47.t4 149.421
R7 a_27_47.n2 a_27_47.n0 37.4894
R8 a_27_47.n2 a_27_47.n1 37.4894
R9 Z.n0 Z 593.145
R10 Z.n1 Z.n0 585
R11 Z Z.n2 207.35
R12 Z.n0 Z.t1 26.5955
R13 Z.n0 Z.t0 26.5955
R14 Z.n2 Z.t2 24.9236
R15 Z.n2 Z.t3 24.9236
R16 Z.n3 Z 21.9466
R17 Z Z.n3 15.0005
R18 Z.n1 Z 5.04292
R19 Z.n3 Z.n1 1.93989
R20 a_320_309.n2 a_320_309.t0 871.958
R21 a_320_309.n1 a_320_309.n0 590.778
R22 a_320_309.n3 a_320_309.n2 585
R23 a_320_309.n1 a_320_309.t3 381.471
R24 a_320_309.n4 a_320_309.n3 45.059
R25 a_320_309.n3 a_320_309.t1 40.8675
R26 a_320_309.n0 a_320_309.t2 28.5298
R27 a_320_309.n4 a_320_309.n0 16.9824
R28 a_320_309.n5 a_320_309.n4 8.8214
R29 a_320_309.n2 a_320_309.n1 8.21182
R30 VPB.t2 VPB.t0 556.386
R31 VPB.t3 VPB.t4 529.751
R32 VPB.t1 VPB.t2 310.748
R33 VPB.t4 VPB.t5 248.599
R34 VPB.t0 VPB.t3 248.599
R35 VPB VPB.t1 189.409
R36 A.n0 A.t0 295.168
R37 A.n0 A.t1 201.982
R38 A.n1 A.n0 152
R39 A.n1 A 17.435
R40 A A.n1 12.5798
R41 VPWR.n2 VPWR.n0 604.86
R42 VPWR.n2 VPWR.n1 310.899
R43 VPWR.n1 VPWR.t3 58.4849
R44 VPWR.n1 VPWR.t1 56.9458
R45 VPWR.n0 VPWR.t2 28.2931
R46 VPWR.n0 VPWR.t0 28.2931
R47 VPWR VPWR.n2 0.216573
R48 a_214_47.t1 a_214_47.n1 672.888
R49 a_214_47.n1 a_214_47.t0 263.337
R50 a_214_47.n0 a_214_47.t2 237.787
R51 a_214_47.n1 a_214_47.n0 224.786
R52 a_214_47.n0 a_214_47.t3 139.488
R53 a_392_47.n0 a_392_47.t0 327.474
R54 a_392_47.n0 a_392_47.t3 270.805
R55 a_392_47.n1 a_392_47.n0 185
R56 a_392_47.t1 a_392_47.n1 36.0005
R57 a_392_47.n1 a_392_47.t2 35.0774
R58 VGND.n2 VGND.n0 205.097
R59 VGND.n2 VGND.n1 204.48
R60 VGND.n1 VGND.t0 68.5719
R61 VGND.n1 VGND.t1 38.5719
R62 VGND.n0 VGND.t2 24.9236
R63 VGND.n0 VGND.t3 24.9236
R64 VGND VGND.n2 0.158598
R65 VNB.t0 VNB.t5 3702.27
R66 VNB.t4 VNB.t2 1523.62
R67 VNB.t3 VNB.t0 1495.15
R68 VNB.t2 VNB.t1 1196.12
R69 VNB.t5 VNB.t4 1196.12
R70 VNB VNB.t3 911.327
R71 TE_B.n0 TE_B.t1 284.38
R72 TE_B.n1 TE_B.t0 233.369
R73 TE_B.n1 TE_B.n0 210.474
R74 TE_B.n2 TE_B.t3 204.448
R75 TE_B.n0 TE_B.t2 175.127
R76 TE_B TE_B.n2 167.321
R77 TE_B.n2 TE_B.n1 31.4644
C0 A TE_B 0.124986f
C1 VPWR Z 0.023178f
C2 VPWR VGND 0.016998f
C3 Z VGND 0.011142f
C4 VPB VPWR 0.088255f
C5 A VPWR 0.044881f
C6 VPB Z 0.012981f
C7 TE_B VPWR 0.053172f
C8 VPB VGND 0.004366f
C9 A VGND 0.042829f
C10 TE_B Z 0.023743f
C11 TE_B VGND 0.020636f
C12 VPB A 0.063734f
C13 VPB TE_B 0.163644f
C14 VGND VNB 0.486559f
C15 Z VNB 0.054717f
C16 VPWR VNB 0.398468f
C17 TE_B VNB 0.245427f
C18 A VNB 0.156127f
C19 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_4 VNB VPB VGND VPWR TE_B Z A
X0 a_214_47.t1 TE_B.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1875 ps=1.375 w=1 l=0.15
X1 Z.t5 a_27_47.t2 a_320_309.t7 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37525 ps=1.755 w=1 l=0.15
X2 VGND.t5 a_214_47.t2 a_393_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_320_309.t3 TE_B.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.37525 pd=1.755 as=0.1269 ps=1.21 w=0.94 l=0.15
X4 VGND.t4 a_214_47.t3 a_393_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t2 TE_B.t2 a_320_309.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X6 a_320_309.t1 TE_B.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X7 a_393_47.t1 a_214_47.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Z.t7 a_27_47.t3 a_393_47.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X9 VPWR.t0 TE_B.t4 a_320_309.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.2444 ps=2.4 w=0.94 l=0.15
X10 a_393_47.t0 a_214_47.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Z.t6 a_27_47.t4 a_393_47.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_393_47.t5 a_27_47.t5 Z.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_214_47.t0 TE_B.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.121875 ps=1.025 w=0.65 l=0.15
X14 Z.t4 a_27_47.t6 a_320_309.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_320_309.t5 a_27_47.t7 Z.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X16 a_393_47.t4 a_27_47.t8 Z.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_320_309.t4 a_27_47.t9 Z.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR.t5 A.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1875 pd=1.375 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND.t1 A.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.169 ps=1.82 w=0.65 l=0.15
R0 TE_B.n4 TE_B.t5 365.813
R1 TE_B.n0 TE_B.t1 310.087
R2 TE_B.n3 TE_B.t0 194.28
R3 TE_B.n3 TE_B.n2 186.603
R4 TE_B.n0 TE_B.t2 175.127
R5 TE_B.n1 TE_B.t3 175.127
R6 TE_B.n2 TE_B.t4 175.127
R7 TE_B TE_B.n4 167.321
R8 TE_B.n1 TE_B.n0 134.96
R9 TE_B.n2 TE_B.n1 134.96
R10 TE_B.n4 TE_B.n3 22.1979
R11 VPWR.n5 VPWR.n4 604.323
R12 VPWR.n3 VPWR.n2 598.965
R13 VPWR.n9 VPWR.n1 306.202
R14 VPWR.n1 VPWR.t4 39.4005
R15 VPWR.n8 VPWR.n7 34.6358
R16 VPWR.n1 VPWR.t5 34.4755
R17 VPWR.n2 VPWR.t1 28.2931
R18 VPWR.n2 VPWR.t0 28.2931
R19 VPWR.n4 VPWR.t3 28.2931
R20 VPWR.n4 VPWR.t2 28.2931
R21 VPWR.n7 VPWR.n3 27.8593
R22 VPWR.n9 VPWR.n8 16.5652
R23 VPWR.n7 VPWR.n6 9.3005
R24 VPWR.n8 VPWR.n0 9.3005
R25 VPWR.n10 VPWR.n9 7.12063
R26 VPWR.n5 VPWR.n3 6.15486
R27 VPWR.n6 VPWR.n5 0.648523
R28 VPWR.n10 VPWR.n0 0.148519
R29 VPWR.n6 VPWR.n0 0.120292
R30 VPWR VPWR.n10 0.11354
R31 a_214_47.t1 a_214_47.n3 369.178
R32 a_214_47.n3 a_214_47.n2 268.562
R33 a_214_47.n0 a_214_47.t2 263.493
R34 a_214_47.n3 a_214_47.t0 250.062
R35 a_214_47.n2 a_214_47.t5 139.488
R36 a_214_47.n1 a_214_47.n0 134.96
R37 a_214_47.n0 a_214_47.t4 128.534
R38 a_214_47.n1 a_214_47.t3 128.534
R39 a_214_47.n2 a_214_47.n1 109.254
R40 VPB.t4 VPB.t0 556.386
R41 VPB.t3 VPB.t6 535.67
R42 VPB.t5 VPB.t4 310.748
R43 VPB.t7 VPB.t8 248.599
R44 VPB.t9 VPB.t7 248.599
R45 VPB.t6 VPB.t9 248.599
R46 VPB.t2 VPB.t3 248.599
R47 VPB.t1 VPB.t2 248.599
R48 VPB.t0 VPB.t1 248.599
R49 VPB VPB.t5 189.409
R50 a_27_47.t1 a_27_47.n11 364.142
R51 a_27_47.n11 a_27_47.t0 249.351
R52 a_27_47.n2 a_27_47.t7 221.72
R53 a_27_47.n1 a_27_47.t6 221.72
R54 a_27_47.n7 a_27_47.t9 221.72
R55 a_27_47.n8 a_27_47.t2 221.72
R56 a_27_47.n4 a_27_47.n3 169.409
R57 a_27_47.n10 a_27_47.n9 159.424
R58 a_27_47.n6 a_27_47.n0 152
R59 a_27_47.n5 a_27_47.n4 152
R60 a_27_47.n2 a_27_47.t5 149.421
R61 a_27_47.n1 a_27_47.t4 149.421
R62 a_27_47.n7 a_27_47.t8 149.421
R63 a_27_47.n8 a_27_47.t3 149.421
R64 a_27_47.n6 a_27_47.n5 60.6968
R65 a_27_47.n3 a_27_47.n1 58.9116
R66 a_27_47.n9 a_27_47.n7 48.2005
R67 a_27_47.n9 a_27_47.n8 26.7783
R68 a_27_47.n11 a_27_47.n10 22.2135
R69 a_27_47.n4 a_27_47.n0 17.4085
R70 a_27_47.n3 a_27_47.n2 16.0672
R71 a_27_47.n7 a_27_47.n6 12.4968
R72 a_27_47.n10 a_27_47.n0 9.9845
R73 a_27_47.n5 a_27_47.n1 1.78569
R74 a_320_309.n3 a_320_309.t0 862.809
R75 a_320_309.n3 a_320_309.n2 599.683
R76 a_320_309.n1 a_320_309.t5 337.959
R77 a_320_309.n1 a_320_309.n0 292.5
R78 a_320_309.n5 a_320_309.n4 146.25
R79 a_320_309.t3 a_320_309.n5 82.7824
R80 a_320_309.n4 a_320_309.n3 53.7669
R81 a_320_309.n5 a_320_309.t7 49.8979
R82 a_320_309.n2 a_320_309.t2 28.2931
R83 a_320_309.n2 a_320_309.t1 28.2931
R84 a_320_309.n0 a_320_309.t6 26.5955
R85 a_320_309.n0 a_320_309.t4 26.5955
R86 a_320_309.n4 a_320_309.n1 23.9163
R87 Z.n6 Z.n5 585
R88 Z.n4 Z.n3 585
R89 Z.n2 Z.n0 229.8
R90 Z.n2 Z.n1 185
R91 Z Z.n2 28.8005
R92 Z.n3 Z.t2 26.5955
R93 Z.n3 Z.t5 26.5955
R94 Z.n5 Z.t3 26.5955
R95 Z.n5 Z.t4 26.5955
R96 Z.n0 Z.t0 24.9236
R97 Z.n0 Z.t7 24.9236
R98 Z.n1 Z.t1 24.9236
R99 Z.n1 Z.t6 24.9236
R100 Z Z.n4 21.0291
R101 Z.n4 Z 21.0291
R102 Z.n6 Z 17.3719
R103 Z.n7 Z 14.546
R104 Z Z.n7 5.23686
R105 Z.n7 Z 5.06717
R106 Z Z.n6 3.65764
R107 a_393_47.n4 a_393_47.t5 327.305
R108 a_393_47.n1 a_393_47.t3 267.158
R109 a_393_47.n1 a_393_47.n0 192.154
R110 a_393_47.n3 a_393_47.n2 185
R111 a_393_47.n5 a_393_47.n4 185
R112 a_393_47.n4 a_393_47.n3 60.1326
R113 a_393_47.n3 a_393_47.n1 56.9274
R114 a_393_47.n2 a_393_47.t7 36.0005
R115 a_393_47.n2 a_393_47.t0 36.0005
R116 a_393_47.n0 a_393_47.t2 24.9236
R117 a_393_47.n0 a_393_47.t1 24.9236
R118 a_393_47.t6 a_393_47.n5 24.9236
R119 a_393_47.n5 a_393_47.t4 24.9236
R120 VGND.n3 VGND.n2 204.149
R121 VGND.n5 VGND.n4 198.964
R122 VGND.n13 VGND.n12 185
R123 VGND.n12 VGND.t0 44.3082
R124 VGND.n6 VGND.n1 34.6358
R125 VGND.n10 VGND.n1 34.6358
R126 VGND.n14 VGND.n13 33.8652
R127 VGND.n12 VGND.t1 24.9236
R128 VGND.n2 VGND.t2 24.9236
R129 VGND.n2 VGND.t4 24.9236
R130 VGND.n4 VGND.t3 24.9236
R131 VGND.n4 VGND.t5 24.9236
R132 VGND.n11 VGND.n10 21.0829
R133 VGND.n6 VGND.n5 20.7064
R134 VGND.n11 VGND.n0 9.3005
R135 VGND.n7 VGND.n6 9.3005
R136 VGND.n8 VGND.n1 9.3005
R137 VGND.n10 VGND.n9 9.3005
R138 VGND.n5 VGND.n3 6.5713
R139 VGND.n7 VGND.n3 0.671755
R140 VGND.n13 VGND.n11 0.188735
R141 VGND.n8 VGND.n7 0.120292
R142 VGND.n9 VGND.n8 0.120292
R143 VGND.n9 VGND.n0 0.120292
R144 VGND.n14 VGND.n0 0.120292
R145 VGND VGND.n14 0.0213333
R146 VNB.t0 VNB.t5 3716.5
R147 VNB.t2 VNB.t9 1537.86
R148 VNB.t1 VNB.t0 1495.15
R149 VNB.t8 VNB.t7 1196.12
R150 VNB.t6 VNB.t8 1196.12
R151 VNB.t9 VNB.t6 1196.12
R152 VNB.t4 VNB.t2 1196.12
R153 VNB.t3 VNB.t4 1196.12
R154 VNB.t5 VNB.t3 1196.12
R155 VNB VNB.t1 911.327
R156 A.n0 A.t0 237.328
R157 A.n0 A.t1 165.029
R158 A.n1 A.n0 152
R159 A.n1 A 17.435
R160 A A.n1 12.5798
C0 TE_B Z 0.04535f
C1 A VGND 0.045825f
C2 VPWR Z 0.03233f
C3 TE_B VGND 0.026659f
C4 VPWR VGND 0.034204f
C5 Z VGND 0.0312f
C6 VPB A 0.035325f
C7 VPB TE_B 0.199796f
C8 VPB VPWR 0.115876f
C9 A TE_B 0.107483f
C10 A VPWR 0.049404f
C11 VPB Z 0.019538f
C12 TE_B VPWR 0.080073f
C13 VPB VGND 0.004931f
C14 VGND VNB 0.663671f
C15 Z VNB 0.062428f
C16 VPWR VNB 0.547045f
C17 TE_B VNB 0.285072f
C18 A VNB 0.123613f
C19 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_0 VPWR VGND VPB VNB A Z TE_B
X0 VGND.t1 TE_B.t0 a_30_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Z.t0 A.t0 a_215_369.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X2 a_215_369.t1 TE_B.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.10855 ps=1.005 w=0.64 l=0.15
X3 a_215_47.t1 a_30_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.07665 ps=0.785 w=0.42 l=0.15
X4 Z.t1 A.t1 a_215_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR.t0 TE_B.t2 a_30_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 TE_B.n0 TE_B.t1 292.413
R1 TE_B.n1 TE_B.t0 206.19
R2 TE_B.n0 TE_B.t2 162.274
R3 TE_B.n2 TE_B.n1 152
R4 TE_B.n1 TE_B.n0 124.249
R5 TE_B.n2 TE_B 6.45714
R6 TE_B TE_B.n2 1.24652
R7 a_30_47.t0 a_30_47.n0 753.674
R8 a_30_47.n0 a_30_47.t2 354.81
R9 a_30_47.n0 a_30_47.t1 303.562
R10 VGND VGND.n0 191.477
R11 VGND.n0 VGND.t0 52.8576
R12 VGND.n0 VGND.t1 51.4291
R13 VNB.t1 VNB.t0 1466.67
R14 VNB.t0 VNB.t2 1025.24
R15 VNB VNB.t1 968.285
R16 A.n0 A.t0 288.204
R17 A.n0 A.t1 195.017
R18 A.n1 A.n0 152
R19 A.n1 A 14.3064
R20 A A.n1 2.76128
R21 a_215_369.t0 a_215_369.t1 64.6411
R22 Z Z.t0 628.25
R23 Z Z.t1 225.267
R24 VPB.t1 VPB.t2 304.829
R25 VPB.t2 VPB.t0 213.084
R26 VPB VPB.t1 201.246
R27 VPWR VPWR.n0 591.583
R28 VPWR.n0 VPWR.t0 86.7743
R29 VPWR.n0 VPWR.t1 61.05
R30 a_215_47.t0 a_215_47.t1 60.0005
C0 VPWR VPB 0.042411f
C1 VPB TE_B 0.136539f
C2 Z VPB 0.010484f
C3 VPWR TE_B 0.034405f
C4 VPWR Z 0.094759f
C5 VPB A 0.073348f
C6 VGND VPB 0.005482f
C7 VPWR A 0.012311f
C8 Z TE_B 0.007676f
C9 VPWR VGND 0.037578f
C10 TE_B A 0.034031f
C11 Z A 0.188537f
C12 VGND TE_B 0.020448f
C13 Z VGND 0.094442f
C14 VGND A 0.012693f
C15 VGND VNB 0.251746f
C16 Z VNB 0.044696f
C17 VPWR VNB 0.213824f
C18 A VNB 0.206932f
C19 TE_B VNB 0.220088f
C20 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_1 VGND VPWR VPB VNB Z A TE_B
X0 VPWR.t1 TE_B.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_204_297.t0 TE_B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.149 ps=1.325 w=1 l=0.15
X2 Z.t0 A.t0 a_204_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3675 ps=1.735 w=1 l=0.15
X3 Z.t1 A.t1 a_286_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_286_47.t1 a_27_47.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.23025 ps=1.385 w=0.65 l=0.15
X5 VGND.t0 TE_B.t2 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.23025 pd=1.385 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 TE_B.n0 TE_B.t1 313.3
R1 TE_B.n0 TE_B.t0 266.707
R2 TE_B.n1 TE_B.t2 229.754
R3 TE_B.n2 TE_B.n1 152
R4 TE_B.n1 TE_B.n0 56.2338
R5 TE_B.n2 TE_B 8.58403
R6 TE_B TE_B.n2 1.65697
R7 a_27_47.t0 a_27_47.n0 691.448
R8 a_27_47.n0 a_27_47.t2 317.029
R9 a_27_47.n0 a_27_47.t1 266.438
R10 VPWR VPWR.n0 604.854
R11 VPWR.n0 VPWR.t1 49.2505
R12 VPWR.n0 VPWR.t0 40.8401
R13 VPB.t0 VPB.t2 523.832
R14 VPB.t1 VPB.t0 281.154
R15 VPB VPB.t1 192.369
R16 a_204_297.t0 a_204_297.t1 144.796
R17 A.n0 A.t0 230.363
R18 A.n0 A.t1 158.064
R19 A.n1 A.n0 152
R20 A.n1 A 14.8903
R21 A A.n1 2.87397
R22 Z Z.t0 320.224
R23 Z Z.t1 212.183
R24 Z.n0 Z 94.7874
R25 Z.n0 Z 5.08285
R26 Z Z.n0 3.57697
R27 a_286_47.t0 a_286_47.t1 60.0005
R28 VNB.t0 VNB.t2 2520.39
R29 VNB.t2 VNB.t1 1352.75
R30 VNB VNB.t0 925.567
R31 VGND VGND.n0 83.5196
R32 VGND.n0 VGND.t0 70.4693
R33 VGND.n0 VGND.t1 63.8192
C0 VPB TE_B 0.110791f
C1 VPB A 0.045045f
C2 VPB VPWR 0.048834f
C3 TE_B A 0.006508f
C4 VPB Z 0.011362f
C5 TE_B VPWR 0.035386f
C6 A VPWR 0.009185f
C7 TE_B Z 0.008978f
C8 VPB VGND 0.004335f
C9 A Z 0.161437f
C10 TE_B VGND 0.021622f
C11 VPWR Z 0.173614f
C12 A VGND 0.011807f
C13 VPWR VGND 0.044838f
C14 Z VGND 0.09749f
C15 VGND VNB 0.293412f
C16 Z VNB 0.054798f
C17 VPWR VNB 0.247318f
C18 A VNB 0.166607f
C19 TE_B VNB 0.252019f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_2 VPWR VGND VPB VNB Z TE_B A
X0 Z.t2 A.t0 a_204_309.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t1 a_27_47.t2 a_214_120.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.16535 ps=1.82 w=0.65 l=0.15
X2 a_204_309.t1 A.t1 Z.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2593 ps=2.56 w=1 l=0.15
X3 Z.t0 A.t2 a_214_120.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VPWR.t0 TE_B.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1415 pd=1.265 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 VPWR.t2 TE_B.t1 a_204_309.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.241375 pd=2.4 as=0.1269 ps=1.21 w=0.94 l=0.15
X6 a_204_309.t3 TE_B.t2 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1415 ps=1.265 w=0.94 l=0.15
X7 a_214_120.t0 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_214_120.t2 A.t3 Z.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t2 TE_B.t3 a_27_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1079 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A.n1 A.t0 234.038
R1 A.n0 A.t1 221.72
R2 A.n1 A.t3 161.738
R3 A A.n1 154.012
R4 A.n0 A.t2 149.421
R5 A.n1 A.n0 61.5894
R6 a_204_309.n1 a_204_309.n0 950.731
R7 a_204_309.n0 a_204_309.t0 28.2931
R8 a_204_309.n0 a_204_309.t3 28.2931
R9 a_204_309.n1 a_204_309.t2 26.5955
R10 a_204_309.t1 a_204_309.n1 26.5955
R11 Z.n3 Z.t1 785.784
R12 Z.n1 Z.t2 354.366
R13 Z.n5 Z.n0 187.048
R14 Z.n0 Z.t3 24.9236
R15 Z.n0 Z.t0 24.9236
R16 Z Z.n4 17.4085
R17 Z Z.n3 17.1525
R18 Z.n4 Z.n2 15.1045
R19 Z.n5 Z 13.3125
R20 Z.n2 Z 7.86336
R21 Z Z.n1 6.71777
R22 Z.n3 Z 6.4005
R23 Z.n1 Z 5.62926
R24 Z.n2 Z 4.57193
R25 Z Z.n5 4.0965
R26 Z.n4 Z 2.3045
R27 Z.n5 Z 2.3045
R28 VPB.t1 VPB.t2 565.265
R29 VPB.t0 VPB.t4 281.154
R30 VPB.t2 VPB.t3 248.599
R31 VPB.t4 VPB.t1 248.599
R32 VPB VPB.t0 192.369
R33 a_27_47.t0 a_27_47.n1 679.856
R34 a_27_47.n1 a_27_47.t1 263.329
R35 a_27_47.n1 a_27_47.n0 227.47
R36 a_27_47.n0 a_27_47.t2 224.934
R37 a_27_47.n0 a_27_47.t3 147.072
R38 a_214_120.t2 a_214_120.n1 282.295
R39 a_214_120.n1 a_214_120.t1 274.048
R40 a_214_120.n1 a_214_120.n0 185
R41 a_214_120.n0 a_214_120.t0 32.3082
R42 a_214_120.n0 a_214_120.t3 31.3851
R43 VGND.n1 VGND.t2 245
R44 VGND.n1 VGND.n0 204.536
R45 VGND.n0 VGND.t0 24.9236
R46 VGND.n0 VGND.t1 24.9236
R47 VGND VGND.n1 0.470326
R48 VNB.t4 VNB.t1 2662.78
R49 VNB.t0 VNB.t3 1409.71
R50 VNB.t3 VNB.t2 1196.12
R51 VNB.t1 VNB.t0 1196.12
R52 VNB VNB.t4 925.567
R53 TE_B.n0 TE_B.t1 310.087
R54 TE_B.n1 TE_B.t0 247.428
R55 TE_B.n2 TE_B.t3 229.754
R56 TE_B TE_B.n2 177.757
R57 TE_B.n0 TE_B.t2 175.127
R58 TE_B.n1 TE_B.n0 128.534
R59 TE_B.n2 TE_B.n1 75.5138
R60 VPWR.n1 VPWR.t2 786.087
R61 VPWR.n1 VPWR.n0 312.692
R62 VPWR.n0 VPWR.t0 49.2505
R63 VPWR.n0 VPWR.t1 42.2041
R64 VPWR VPWR.n1 0.496779
C0 Z VGND 0.011904f
C1 VPB TE_B 0.14929f
C2 VPB A 0.074895f
C3 TE_B A 0.006099f
C4 VPB VPWR 0.069241f
C5 TE_B VPWR 0.056442f
C6 VPB Z 0.017924f
C7 TE_B Z 0.001958f
C8 A VPWR 0.02752f
C9 VPB VGND 0.006524f
C10 A Z 0.11699f
C11 TE_B VGND 0.021297f
C12 A VGND 0.018859f
C13 VPWR Z 0.062474f
C14 VPWR VGND 0.062256f
C15 VGND VNB 0.390245f
C16 Z VNB 0.058262f
C17 VPWR VNB 0.322944f
C18 A VNB 0.23366f
C19 TE_B VNB 0.294504f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_4 VGND VPWR VPB VNB TE_B Z A
X0 VGND.t4 a_27_47.t2 a_215_47.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_204_309.t5 A.t0 Z.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t3 a_27_47.t3 a_215_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t3 TE_B.t0 a_204_309.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2444 pd=2.4 as=0.1269 ps=1.21 w=0.94 l=0.15
X4 Z.t5 A.t1 a_215_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X5 a_204_309.t0 TE_B.t1 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X6 a_215_47.t4 a_27_47.t4 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Z.t4 A.t2 a_215_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Z.t0 A.t3 a_204_309.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VPWR.t1 TE_B.t2 a_204_309.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X10 a_204_309.t6 TE_B.t3 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.16025 ps=1.325 w=0.94 l=0.15
X11 a_215_47.t0 A.t4 Z.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_215_47.t7 A.t5 Z.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_215_47.t3 a_27_47.t5 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_204_309.t3 A.t6 Z.t7 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t4 TE_B.t4 a_27_47.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.16025 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X16 Z.t6 A.t7 a_204_309.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t0 TE_B.t5 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t1 a_27_47.n3 395.301
R1 a_27_47.n0 a_27_47.t2 263.493
R2 a_27_47.n3 a_27_47.t0 241.476
R3 a_27_47.n3 a_27_47.n2 227.442
R4 a_27_47.n1 a_27_47.n0 134.96
R5 a_27_47.n2 a_27_47.t4 134.476
R6 a_27_47.n0 a_27_47.t5 128.534
R7 a_27_47.n1 a_27_47.t3 128.534
R8 a_27_47.n2 a_27_47.n1 94.9479
R9 a_215_47.n4 a_215_47.t7 323.711
R10 a_215_47.n1 a_215_47.t6 275.303
R11 a_215_47.n1 a_215_47.n0 192.154
R12 a_215_47.n3 a_215_47.n2 185
R13 a_215_47.n5 a_215_47.n4 185
R14 a_215_47.n3 a_215_47.n1 72.6593
R15 a_215_47.n4 a_215_47.n3 65.0623
R16 a_215_47.n2 a_215_47.t4 30.462
R17 a_215_47.n2 a_215_47.t1 29.539
R18 a_215_47.n0 a_215_47.t5 24.9236
R19 a_215_47.n0 a_215_47.t3 24.9236
R20 a_215_47.n5 a_215_47.t2 24.9236
R21 a_215_47.t0 a_215_47.n5 24.9236
R22 VGND.n6 VGND.t0 282.817
R23 VGND.n2 VGND.n1 204.238
R24 VGND.n4 VGND.n3 198.964
R25 VGND.n1 VGND.t2 24.9236
R26 VGND.n1 VGND.t3 24.9236
R27 VGND.n3 VGND.t1 24.9236
R28 VGND.n3 VGND.t4 24.9236
R29 VGND.n5 VGND.n4 22.9652
R30 VGND.n6 VGND.n5 22.9652
R31 VGND.n5 VGND.n0 9.3005
R32 VGND.n7 VGND.n6 7.12063
R33 VGND.n4 VGND.n2 6.46197
R34 VGND.n2 VGND.n0 0.660443
R35 VGND.n7 VGND.n0 0.148519
R36 VGND VGND.n7 0.11354
R37 VNB.t0 VNB.t7 2677.02
R38 VNB.t5 VNB.t2 1352.75
R39 VNB.t3 VNB.t8 1196.12
R40 VNB.t1 VNB.t3 1196.12
R41 VNB.t2 VNB.t1 1196.12
R42 VNB.t6 VNB.t5 1196.12
R43 VNB.t4 VNB.t6 1196.12
R44 VNB.t7 VNB.t4 1196.12
R45 VNB VNB.t0 911.327
R46 A A.n3 214.197
R47 A.n3 A.t6 212.081
R48 A.n2 A.t7 212.081
R49 A.n1 A.t0 212.081
R50 A.n0 A.t3 212.081
R51 A.n3 A.t5 139.78
R52 A.n2 A.t2 139.78
R53 A.n1 A.t4 139.78
R54 A.n0 A.t1 139.78
R55 A.n3 A.n2 61.346
R56 A.n2 A.n1 61.346
R57 A.n1 A.n0 61.346
R58 Z.n5 Z.n3 300.805
R59 Z.n2 Z.n0 300.803
R60 Z.n2 Z.n1 185
R61 Z.n5 Z.n4 185
R62 Z.n3 Z.t1 26.5955
R63 Z.n3 Z.t0 26.5955
R64 Z.n0 Z.t7 26.5955
R65 Z.n0 Z.t6 26.5955
R66 Z.n4 Z.t3 24.9236
R67 Z.n4 Z.t5 24.9236
R68 Z.n1 Z.t2 24.9236
R69 Z.n1 Z.t4 24.9236
R70 Z Z.n2 5.43306
R71 Z Z.n5 0.223756
R72 a_204_309.n4 a_204_309.t3 422.652
R73 a_204_309.n2 a_204_309.n1 367.474
R74 a_204_309.n3 a_204_309.t4 351.798
R75 a_204_309.n2 a_204_309.n0 310.058
R76 a_204_309.n5 a_204_309.n4 309.305
R77 a_204_309.n3 a_204_309.n2 85.9032
R78 a_204_309.n4 a_204_309.n3 80.776
R79 a_204_309.n1 a_204_309.t1 28.2931
R80 a_204_309.n1 a_204_309.t6 28.2931
R81 a_204_309.n0 a_204_309.t7 28.2931
R82 a_204_309.n0 a_204_309.t0 28.2931
R83 a_204_309.n5 a_204_309.t2 26.5955
R84 a_204_309.t5 a_204_309.n5 26.5955
R85 VPB.t8 VPB.t4 556.386
R86 VPB.t6 VPB.t7 281.154
R87 VPB.t2 VPB.t3 248.599
R88 VPB.t5 VPB.t2 248.599
R89 VPB.t4 VPB.t5 248.599
R90 VPB.t0 VPB.t8 248.599
R91 VPB.t1 VPB.t0 248.599
R92 VPB.t7 VPB.t1 248.599
R93 VPB VPB.t6 189.409
R94 TE_B.n0 TE_B.t0 310.087
R95 TE_B.n3 TE_B.t4 220.391
R96 TE_B.n2 TE_B.t3 199.227
R97 TE_B.n0 TE_B.t1 175.127
R98 TE_B.n1 TE_B.t2 175.127
R99 TE_B.n4 TE_B.t5 158.064
R100 TE_B TE_B.n4 155.685
R101 TE_B.n3 TE_B.n2 151.028
R102 TE_B.n1 TE_B.n0 134.96
R103 TE_B.n2 TE_B.n1 110.861
R104 TE_B.n4 TE_B.n3 9.97291
R105 VPWR.n2 VPWR.t3 341.065
R106 VPWR.n4 VPWR.n3 309.726
R107 VPWR.n6 VPWR.n1 309.724
R108 VPWR.n1 VPWR.t0 39.8196
R109 VPWR.n3 VPWR.t2 28.2931
R110 VPWR.n3 VPWR.t1 28.2931
R111 VPWR.n1 VPWR.t4 26.4528
R112 VPWR.n6 VPWR.n5 22.9652
R113 VPWR.n5 VPWR.n4 19.577
R114 VPWR.n5 VPWR.n0 9.3005
R115 VPWR.n7 VPWR.n6 7.12063
R116 VPWR.n4 VPWR.n2 6.62798
R117 VPWR.n2 VPWR.n0 0.669349
R118 VPWR.n7 VPWR.n0 0.148519
R119 VPWR VPWR.n7 0.11354
C0 VPB A 0.148061f
C1 VPB VPWR 0.103727f
C2 TE_B A 0.005873f
C3 TE_B VPWR 0.104251f
C4 VPB Z 0.010561f
C5 A VPWR 0.032294f
C6 TE_B Z 0.001725f
C7 VPB VGND 0.007414f
C8 TE_B VGND 0.025611f
C9 A Z 0.194222f
C10 VPWR Z 0.02172f
C11 A VGND 0.036773f
C12 VPWR VGND 0.097631f
C13 Z VGND 0.029046f
C14 VPB TE_B 0.183389f
C15 VGND VNB 0.566134f
C16 Z VNB 0.013739f
C17 VPWR VNB 0.468984f
C18 A VNB 0.456615f
C19 TE_B VNB 0.321488f
C20 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_8 VNB VPB VGND VPWR A TE_B Z
X0 VPWR.t9 TE_B.t0 a_407_309.t15 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.2444 ps=2.4 w=0.94 l=0.15
X1 a_455_47.t15 a_301_47.t2 VGND.t7 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Z.t15 a_116_47.t4 a_407_309.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Z.t7 a_116_47.t5 a_455_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.18 w=0.65 l=0.15
X4 a_116_47.t2 A.t0 VPWR.t10 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5 a_407_309.t1 a_116_47.t6 Z.t14 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t8 TE_B.t1 a_407_309.t14 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X7 a_407_309.t13 TE_B.t2 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.38275 pd=1.77 as=0.1269 ps=1.21 w=0.94 l=0.15
X8 VGND.t6 a_301_47.t3 a_455_47.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VGND.t5 a_301_47.t4 a_455_47.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Z.t13 a_116_47.t7 a_407_309.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_116_47.t3 A.t1 VGND.t10 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19175 ps=1.89 w=0.65 l=0.15
X12 VGND.t4 a_301_47.t5 a_455_47.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_407_309.t12 TE_B.t3 VPWR.t6 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X14 VGND.t3 a_301_47.t6 a_455_47.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_455_47.t1 a_116_47.t8 Z.t6 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t5 TE_B.t4 a_407_309.t11 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X17 a_455_47.t2 a_116_47.t9 Z.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_455_47.t3 a_116_47.t10 Z.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_301_47.t0 TE_B.t5 VGND.t9 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.115375 ps=1.005 w=0.65 l=0.15
X20 a_455_47.t10 a_301_47.t7 VGND.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.18 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_301_47.t1 TE_B.t6 VPWR.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1775 ps=1.355 w=1 l=0.15
X22 a_455_47.t9 a_301_47.t8 VGND.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_455_47.t8 a_301_47.t9 VGND.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_407_309.t3 a_116_47.t11 Z.t12 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Z.t3 a_116_47.t12 a_455_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Z.t2 a_116_47.t13 a_455_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR.t0 A.t2 a_116_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.135 ps=1.27 w=1 l=0.15
X28 Z.t11 a_116_47.t14 a_407_309.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.38275 ps=1.77 w=1 l=0.15
X29 Z.t1 a_116_47.t15 a_455_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_407_309.t10 TE_B.t7 VPWR.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X31 VGND.t8 A.t3 a_116_47.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 VPWR.t3 TE_B.t8 a_407_309.t9 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X33 a_407_309.t5 a_116_47.t16 Z.t10 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X34 Z.t9 a_116_47.t17 a_407_309.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_407_309.t8 TE_B.t9 VPWR.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X36 a_455_47.t7 a_116_47.t18 Z.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 a_407_309.t7 a_116_47.t19 Z.t8 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 TE_B.n0 TE_B.t2 310.087
R1 TE_B.n7 TE_B.n6 243.483
R2 TE_B.n7 TE_B.t6 212.081
R3 TE_B.n0 TE_B.t1 175.127
R4 TE_B.n1 TE_B.t3 175.127
R5 TE_B.n2 TE_B.t4 175.127
R6 TE_B.n3 TE_B.t7 175.127
R7 TE_B.n4 TE_B.t8 175.127
R8 TE_B.n5 TE_B.t9 175.127
R9 TE_B.n6 TE_B.t0 175.127
R10 TE_B.n8 TE_B.n7 165.968
R11 TE_B.n7 TE_B.t5 139.78
R12 TE_B.n1 TE_B.n0 134.96
R13 TE_B.n2 TE_B.n1 134.96
R14 TE_B.n3 TE_B.n2 134.96
R15 TE_B.n4 TE_B.n3 134.96
R16 TE_B.n5 TE_B.n4 134.96
R17 TE_B.n6 TE_B.n5 134.96
R18 TE_B.n8 TE_B 15.093
R19 TE_B TE_B.n8 10.8901
R20 a_407_309.n6 a_407_309.t15 874.173
R21 a_407_309.n8 a_407_309.n3 602.694
R22 a_407_309.n7 a_407_309.n4 602.694
R23 a_407_309.n6 a_407_309.n5 602.694
R24 a_407_309.n12 a_407_309.n11 591.52
R25 a_407_309.n10 a_407_309.n9 585
R26 a_407_309.n1 a_407_309.t5 337.959
R27 a_407_309.n1 a_407_309.n0 292.5
R28 a_407_309.n13 a_407_309.n2 292.5
R29 a_407_309.n15 a_407_309.n14 292.5
R30 a_407_309.n8 a_407_309.n7 63.2476
R31 a_407_309.n7 a_407_309.n6 63.2476
R32 a_407_309.n9 a_407_309.n8 60.6651
R33 a_407_309.n11 a_407_309.n10 60.3907
R34 a_407_309.n10 a_407_309.t13 46.1069
R35 a_407_309.n3 a_407_309.t14 28.2931
R36 a_407_309.n3 a_407_309.t12 28.2931
R37 a_407_309.n4 a_407_309.t11 28.2931
R38 a_407_309.n4 a_407_309.t10 28.2931
R39 a_407_309.n5 a_407_309.t9 28.2931
R40 a_407_309.n5 a_407_309.t8 28.2931
R41 a_407_309.n11 a_407_309.t4 27.7133
R42 a_407_309.n2 a_407_309.t2 26.5955
R43 a_407_309.n2 a_407_309.t3 26.5955
R44 a_407_309.n0 a_407_309.t6 26.5955
R45 a_407_309.n0 a_407_309.t7 26.5955
R46 a_407_309.t0 a_407_309.n15 26.5955
R47 a_407_309.n15 a_407_309.t1 26.5955
R48 a_407_309.n13 a_407_309.n12 20.5479
R49 a_407_309.n14 a_407_309.n1 18.8637
R50 a_407_309.n14 a_407_309.n13 18.8637
R51 a_407_309.n12 a_407_309.n9 7.63559
R52 VPWR.n11 VPWR.n10 604.301
R53 VPWR.n16 VPWR.n5 598.965
R54 VPWR.n14 VPWR.n7 598.965
R55 VPWR.n9 VPWR.n8 598.965
R56 VPWR.n23 VPWR.t10 337.841
R57 VPWR.n21 VPWR.n2 309.469
R58 VPWR.n2 VPWR.t1 43.3405
R59 VPWR.n20 VPWR.n3 34.6358
R60 VPWR.n5 VPWR.t2 28.2931
R61 VPWR.n5 VPWR.t9 28.2931
R62 VPWR.n7 VPWR.t4 28.2931
R63 VPWR.n7 VPWR.t3 28.2931
R64 VPWR.n8 VPWR.t6 28.2931
R65 VPWR.n8 VPWR.t5 28.2931
R66 VPWR.n10 VPWR.t7 28.2931
R67 VPWR.n10 VPWR.t8 28.2931
R68 VPWR.n2 VPWR.t0 26.5955
R69 VPWR.n16 VPWR.n3 25.977
R70 VPWR.n14 VPWR.n13 24.4711
R71 VPWR.n21 VPWR.n20 22.9652
R72 VPWR.n22 VPWR.n21 21.0829
R73 VPWR.n15 VPWR.n14 19.9534
R74 VPWR.n23 VPWR.n22 18.4476
R75 VPWR.n16 VPWR.n15 18.4476
R76 VPWR.n13 VPWR.n9 13.9299
R77 VPWR.n13 VPWR.n12 9.3005
R78 VPWR.n14 VPWR.n6 9.3005
R79 VPWR.n15 VPWR.n4 9.3005
R80 VPWR.n17 VPWR.n16 9.3005
R81 VPWR.n18 VPWR.n3 9.3005
R82 VPWR.n20 VPWR.n19 9.3005
R83 VPWR.n21 VPWR.n1 9.3005
R84 VPWR.n22 VPWR.n0 9.3005
R85 VPWR.n24 VPWR.n23 9.3005
R86 VPWR.n11 VPWR.n9 6.72135
R87 VPWR.n12 VPWR.n11 0.819886
R88 VPWR.n12 VPWR.n6 0.120292
R89 VPWR.n6 VPWR.n4 0.120292
R90 VPWR.n17 VPWR.n4 0.120292
R91 VPWR.n18 VPWR.n17 0.120292
R92 VPWR.n19 VPWR.n18 0.120292
R93 VPWR.n19 VPWR.n1 0.120292
R94 VPWR.n1 VPWR.n0 0.120292
R95 VPWR.n24 VPWR.n0 0.120292
R96 VPWR VPWR.n24 0.0226354
R97 VPB.t12 VPB.t17 556.386
R98 VPB.t15 VPB.t4 544.548
R99 VPB.t8 VPB.t12 298.911
R100 VPB.t6 VPB.t5 248.599
R101 VPB.t7 VPB.t6 248.599
R102 VPB.t0 VPB.t7 248.599
R103 VPB.t1 VPB.t0 248.599
R104 VPB.t2 VPB.t1 248.599
R105 VPB.t3 VPB.t2 248.599
R106 VPB.t4 VPB.t3 248.599
R107 VPB.t16 VPB.t15 248.599
R108 VPB.t14 VPB.t16 248.599
R109 VPB.t13 VPB.t14 248.599
R110 VPB.t11 VPB.t13 248.599
R111 VPB.t10 VPB.t11 248.599
R112 VPB.t9 VPB.t10 248.599
R113 VPB.t17 VPB.t9 248.599
R114 VPB.t18 VPB.t8 248.599
R115 VPB VPB.t18 213.084
R116 a_301_47.n7 a_301_47.n6 376.656
R117 a_301_47.n0 a_301_47.t3 263.493
R118 a_301_47.t1 a_301_47.n7 249.98
R119 a_301_47.n7 a_301_47.t0 227.38
R120 a_301_47.n5 a_301_47.n4 134.96
R121 a_301_47.n4 a_301_47.n3 134.96
R122 a_301_47.n3 a_301_47.n2 134.96
R123 a_301_47.n2 a_301_47.n1 134.96
R124 a_301_47.n1 a_301_47.n0 134.96
R125 a_301_47.n6 a_301_47.n5 132.942
R126 a_301_47.n0 a_301_47.t2 128.534
R127 a_301_47.n1 a_301_47.t5 128.534
R128 a_301_47.n2 a_301_47.t8 128.534
R129 a_301_47.n3 a_301_47.t6 128.534
R130 a_301_47.n4 a_301_47.t9 128.534
R131 a_301_47.n5 a_301_47.t4 128.534
R132 a_301_47.n6 a_301_47.t7 126.612
R133 VGND.n6 VGND.n5 204.291
R134 VGND.n8 VGND.n7 198.964
R135 VGND.n10 VGND.n9 198.964
R136 VGND.n17 VGND.n16 198.964
R137 VGND.n23 VGND.n2 198.756
R138 VGND.n25 VGND.t10 135.921
R139 VGND.n2 VGND.t9 40.6159
R140 VGND.n15 VGND.n4 34.6358
R141 VGND.n19 VGND.n18 34.6358
R142 VGND.n19 VGND.n1 34.6358
R143 VGND.n11 VGND.n8 32.0005
R144 VGND.n5 VGND.t2 24.9236
R145 VGND.n5 VGND.t5 24.9236
R146 VGND.n7 VGND.t0 24.9236
R147 VGND.n7 VGND.t3 24.9236
R148 VGND.n9 VGND.t1 24.9236
R149 VGND.n9 VGND.t4 24.9236
R150 VGND.n16 VGND.t7 24.9236
R151 VGND.n16 VGND.t6 24.9236
R152 VGND.n2 VGND.t8 24.9236
R153 VGND.n23 VGND.n1 22.9652
R154 VGND.n24 VGND.n23 21.0829
R155 VGND.n25 VGND.n24 18.4476
R156 VGND.n18 VGND.n17 9.41227
R157 VGND.n26 VGND.n25 9.3005
R158 VGND.n12 VGND.n11 9.3005
R159 VGND.n13 VGND.n4 9.3005
R160 VGND.n15 VGND.n14 9.3005
R161 VGND.n18 VGND.n3 9.3005
R162 VGND.n20 VGND.n19 9.3005
R163 VGND.n21 VGND.n1 9.3005
R164 VGND.n23 VGND.n22 9.3005
R165 VGND.n24 VGND.n0 9.3005
R166 VGND.n11 VGND.n10 6.4005
R167 VGND.n8 VGND.n6 5.79899
R168 VGND.n10 VGND.n4 3.38874
R169 VGND.n12 VGND.n6 0.650401
R170 VGND.n17 VGND.n15 0.376971
R171 VGND.n13 VGND.n12 0.120292
R172 VGND.n14 VGND.n13 0.120292
R173 VGND.n14 VGND.n3 0.120292
R174 VGND.n20 VGND.n3 0.120292
R175 VGND.n21 VGND.n20 0.120292
R176 VGND.n22 VGND.n21 0.120292
R177 VGND.n22 VGND.n0 0.120292
R178 VGND.n26 VGND.n0 0.120292
R179 VGND VGND.n26 0.0226354
R180 a_455_47.n4 a_455_47.t7 327.305
R181 a_455_47.t14 a_455_47.n13 265.808
R182 a_455_47.n13 a_455_47.n0 192.154
R183 a_455_47.n12 a_455_47.n1 192.154
R184 a_455_47.n11 a_455_47.n2 192.154
R185 a_455_47.n4 a_455_47.n3 185
R186 a_455_47.n6 a_455_47.n5 185
R187 a_455_47.n8 a_455_47.n7 185
R188 a_455_47.n10 a_455_47.n9 185
R189 a_455_47.n6 a_455_47.n4 56.59
R190 a_455_47.n8 a_455_47.n6 56.59
R191 a_455_47.n10 a_455_47.n8 55.3437
R192 a_455_47.n12 a_455_47.n11 53.7605
R193 a_455_47.n13 a_455_47.n12 53.7605
R194 a_455_47.n11 a_455_47.n10 53.0138
R195 a_455_47.n9 a_455_47.t10 49.8467
R196 a_455_47.n9 a_455_47.t0 48.0005
R197 a_455_47.n7 a_455_47.t4 24.9236
R198 a_455_47.n7 a_455_47.t1 24.9236
R199 a_455_47.n5 a_455_47.t5 24.9236
R200 a_455_47.n5 a_455_47.t2 24.9236
R201 a_455_47.n3 a_455_47.t6 24.9236
R202 a_455_47.n3 a_455_47.t3 24.9236
R203 a_455_47.n0 a_455_47.t12 24.9236
R204 a_455_47.n0 a_455_47.t15 24.9236
R205 a_455_47.n1 a_455_47.t11 24.9236
R206 a_455_47.n1 a_455_47.t9 24.9236
R207 a_455_47.n2 a_455_47.t13 24.9236
R208 a_455_47.n2 a_455_47.t8 24.9236
R209 VNB.t17 VNB.t14 3360.52
R210 VNB.t10 VNB.t0 1936.57
R211 VNB.t16 VNB.t17 1438.19
R212 VNB.t6 VNB.t7 1196.12
R213 VNB.t3 VNB.t6 1196.12
R214 VNB.t5 VNB.t3 1196.12
R215 VNB.t2 VNB.t5 1196.12
R216 VNB.t4 VNB.t2 1196.12
R217 VNB.t1 VNB.t4 1196.12
R218 VNB.t0 VNB.t1 1196.12
R219 VNB.t13 VNB.t10 1196.12
R220 VNB.t8 VNB.t13 1196.12
R221 VNB.t11 VNB.t8 1196.12
R222 VNB.t9 VNB.t11 1196.12
R223 VNB.t12 VNB.t9 1196.12
R224 VNB.t15 VNB.t12 1196.12
R225 VNB.t14 VNB.t15 1196.12
R226 VNB.t18 VNB.t16 1196.12
R227 VNB VNB.t18 1025.24
R228 a_116_47.n23 a_116_47.n22 654.059
R229 a_116_47.n22 a_116_47.n0 235.535
R230 a_116_47.n5 a_116_47.t16 221.72
R231 a_116_47.n6 a_116_47.t17 221.72
R232 a_116_47.n4 a_116_47.t19 221.72
R233 a_116_47.n10 a_116_47.t4 221.72
R234 a_116_47.n12 a_116_47.t6 221.72
R235 a_116_47.n2 a_116_47.t7 221.72
R236 a_116_47.n18 a_116_47.t11 221.72
R237 a_116_47.n19 a_116_47.t14 221.72
R238 a_116_47.n21 a_116_47.n20 167.617
R239 a_116_47.n17 a_116_47.n1 152
R240 a_116_47.n16 a_116_47.n15 152
R241 a_116_47.n14 a_116_47.n13 152
R242 a_116_47.n11 a_116_47.n3 152
R243 a_116_47.n9 a_116_47.n8 152
R244 a_116_47.n5 a_116_47.t18 149.421
R245 a_116_47.n6 a_116_47.t15 149.421
R246 a_116_47.n4 a_116_47.t10 149.421
R247 a_116_47.n10 a_116_47.t13 149.421
R248 a_116_47.n12 a_116_47.t9 149.421
R249 a_116_47.n2 a_116_47.t12 149.421
R250 a_116_47.n18 a_116_47.t8 149.421
R251 a_116_47.n19 a_116_47.t5 149.421
R252 a_116_47.n8 a_116_47.n7 84.799
R253 a_116_47.n6 a_116_47.n5 74.9783
R254 a_116_47.n17 a_116_47.n16 60.6968
R255 a_116_47.n13 a_116_47.n2 55.3412
R256 a_116_47.n20 a_116_47.n18 51.7709
R257 a_116_47.n9 a_116_47.n4 48.2005
R258 a_116_47.n12 a_116_47.n11 41.0598
R259 a_116_47.n7 a_116_47.n4 36.6421
R260 a_116_47.n11 a_116_47.n10 33.919
R261 a_116_47.n7 a_116_47.n6 28.6962
R262 a_116_47.n10 a_116_47.n9 26.7783
R263 a_116_47.t0 a_116_47.n23 26.5955
R264 a_116_47.n23 a_116_47.t2 26.5955
R265 a_116_47.n0 a_116_47.t1 24.9236
R266 a_116_47.n0 a_116_47.t3 24.9236
R267 a_116_47.n22 a_116_47.n21 23.834
R268 a_116_47.n20 a_116_47.n19 23.2079
R269 a_116_47.n13 a_116_47.n12 19.6375
R270 a_116_47.n8 a_116_47.n3 17.4085
R271 a_116_47.n14 a_116_47.n3 17.4085
R272 a_116_47.n15 a_116_47.n14 17.4085
R273 a_116_47.n15 a_116_47.n1 17.4085
R274 a_116_47.n18 a_116_47.n17 8.92643
R275 a_116_47.n16 a_116_47.n2 5.35606
R276 a_116_47.n21 a_116_47.n1 1.7925
R277 Z.n7 Z.n6 585
R278 Z.n5 Z.n4 585
R279 Z.n3 Z.n2 585
R280 Z.n1 Z.n0 585
R281 Z.n10 Z.n8 229.8
R282 Z.n14 Z.n13 185
R283 Z.n12 Z.n11 185
R284 Z.n10 Z.n9 185
R285 Z.n14 Z.n12 44.8005
R286 Z.n12 Z.n10 44.8005
R287 Z Z.n1 27.4291
R288 Z.n0 Z.t12 26.5955
R289 Z.n0 Z.t11 26.5955
R290 Z.n2 Z.t14 26.5955
R291 Z.n2 Z.t13 26.5955
R292 Z.n4 Z.t8 26.5955
R293 Z.n4 Z.t15 26.5955
R294 Z.n6 Z.t10 26.5955
R295 Z.n6 Z.t9 26.5955
R296 Z.n8 Z.t6 24.9236
R297 Z.n8 Z.t7 24.9236
R298 Z.n9 Z.t5 24.9236
R299 Z.n9 Z.t3 24.9236
R300 Z.n11 Z.t4 24.9236
R301 Z.n11 Z.t2 24.9236
R302 Z.n13 Z.t0 24.9236
R303 Z.n13 Z.t1 24.9236
R304 Z Z.n14 21.0032
R305 Z Z.n7 17.3719
R306 Z.n1 Z 14.6291
R307 Z Z.n5 13.7148
R308 Z.n3 Z 10.9719
R309 Z Z.n3 10.0576
R310 Z.n5 Z 7.31479
R311 Z.n7 Z 3.65764
R312 A.n1 A.t0 231.017
R313 A.n0 A.t2 221.72
R314 A.n1 A.t1 158.716
R315 A.n2 A.n1 152
R316 A.n0 A.t3 149.421
R317 A.n1 A.n0 61.5894
R318 A.n2 A 10.5744
R319 A A.n2 2.04108
C0 VPB A 0.072814f
C1 VPB TE_B 0.340703f
C2 VGND VPB 0.005681f
C3 A TE_B 0.065637f
C4 VPB VPWR 0.179256f
C5 VGND A 0.073719f
C6 VPB Z 0.027454f
C7 A VPWR 0.080343f
C8 VGND TE_B 0.060461f
C9 TE_B VPWR 0.167153f
C10 VGND VPWR 0.068364f
C11 TE_B Z 0.101783f
C12 VGND Z 0.045623f
C13 VPWR Z 0.062136f
C14 VGND VNB 1.04398f
C15 Z VNB 0.063938f
C16 VPWR VNB 0.867196f
C17 TE_B VNB 0.42661f
C18 A VNB 0.246447f
C19 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__edfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__edfxbp_1 VPWR VGND CLK DE Q D Q_N VPB VNB
X0 a_381_369.t0 D.t0 a_299_47.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 Q.t1 a_1591_413# VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR.t10 DE.t0 a_423_343.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 VPWR.t6 CLK.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q_N.t1 a_791_264.t2 VPWR.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_986_413.t3 a_193_47.t2 a_299_47.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.15985 ps=1.265 w=0.42 l=0.15
X6 VGND.t8 DE.t1 a_423_343.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_1500_413.t0 a_1150_159.t2 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_1101_47# a_193_47.t3 a_986_413.t2 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X9 a_1514_47.t0 a_1150_159.t3 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 Q.t0 a_1591_413# VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.154 ps=1.335 w=1 l=0.15
X11 VPWR.t1 a_1591_413# a_791_264.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1728 ps=1.82 w=0.64 l=0.15
X12 a_193_47.t0 a_27_47.t2 VGND.t10 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_729_47.t1 a_423_343.t2 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X14 a_729_369.t1 DE.t2 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X15 a_1077_413.t1 a_27_47.t3 a_986_413.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X16 VPWR.t4 a_791_264.t3 a_1675_413.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0882 ps=0.84 w=0.42 l=0.15
X17 a_299_47.t0 a_791_264.t4 a_729_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1446 pd=1.18 as=0.0756 ps=0.78 w=0.42 l=0.15
X18 VGND.t0 a_791_264.t5 a_1717_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.066 ps=0.745 w=0.42 l=0.15
X19 a_193_47.t1 a_27_47.t4 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VPWR.t0 a_1150_159.t4 a_1077_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X21 a_1717_47.t1 a_27_47.t5 a_1591_413# VNB.t13 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X22 a_1150_159.t1 a_986_413.t4 VPWR.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X23 a_986_413.t1 a_27_47.t6 a_299_47.t5 VNB.t14 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.1446 ps=1.18 w=0.36 l=0.15
X24 a_299_47.t1 a_791_264.t6 a_729_369.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.15985 pd=1.265 as=0.1152 ps=1 w=0.64 l=0.15
X25 VGND.t7 a_1591_413# a_791_264.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 a_381_47.t0 D.t1 a_299_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR.t8 a_423_343.t3 a_381_369.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X28 VGND.t5 CLK.t1 a_27_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VGND.t2 DE.t3 a_381_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 a_1150_159.t0 a_986_413.t5 VGND.t9 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
X31 Q_N.t0 a_791_264.t7 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
R0 D.n0 D.t1 220.367
R1 D.n0 D.t0 216.796
R2 D D.n0 71.33
R3 a_299_47.n1 a_299_47.t3 467.892
R4 a_299_47.n3 a_299_47.n2 391.748
R5 a_299_47.n1 a_299_47.t2 232.434
R6 a_299_47.n3 a_299_47.t4 230.97
R7 a_299_47.n0 a_299_47.t5 208.333
R8 a_299_47.n2 a_299_47.n0 188.082
R9 a_299_47.t1 a_299_47.n3 34.992
R10 a_299_47.n0 a_299_47.t0 28.3186
R11 a_299_47.n2 a_299_47.n1 20.4743
R12 a_381_369.t0 a_381_369.t1 64.6411
R13 VPB.t10 VPB.t9 855.297
R14 VPB.t8 VPB.t5 787.227
R15 VPB.t12 VPB.t10 556.386
R16 VPB.t2 VPB.t7 556.386
R17 VPB.t13 VPB.t1 556.386
R18 VPB.t0 VPB.t3 458.724
R19 VPB.t4 VPB.t12 390.654
R20 VPB.t15 VPB.t4 304.829
R21 VPB.t14 VPB.t0 301.87
R22 VPB.t5 VPB.t6 287.072
R23 VPB.t9 VPB.t8 287.072
R24 VPB.t3 VPB.t15 269.315
R25 VPB.t7 VPB.t14 260.437
R26 VPB.t11 VPB.t13 248.599
R27 VPB.t1 VPB.t2 213.084
R28 VPB VPB.t11 142.056
R29 VGND.n24 VGND.t9 273.476
R30 VGND.n8 VGND.t4 244.518
R31 VGND.n36 VGND.t2 238.311
R32 VGND.n34 VGND.n4 202.262
R33 VGND.n43 VGND.n42 199.739
R34 VGND.n14 VGND.n11 123.651
R35 VGND.n13 VGND.n12 117.118
R36 VGND.n12 VGND.t0 57.819
R37 VGND.n11 VGND.t7 57.8184
R38 VGND.n4 VGND.t3 41.4291
R39 VGND.n4 VGND.t8 41.4291
R40 VGND.n42 VGND.t10 38.5719
R41 VGND.n42 VGND.t5 38.5719
R42 VGND.n17 VGND.n10 34.6358
R43 VGND.n18 VGND.n17 34.6358
R44 VGND.n19 VGND.n18 34.6358
R45 VGND.n23 VGND.n22 34.6358
R46 VGND.n28 VGND.n6 34.6358
R47 VGND.n29 VGND.n28 34.6358
R48 VGND.n30 VGND.n29 34.6358
R49 VGND.n30 VGND.n3 34.6358
R50 VGND.n40 VGND.n1 34.6358
R51 VGND.n41 VGND.n40 34.6358
R52 VGND.n36 VGND.n35 32.0005
R53 VGND.n34 VGND.n3 29.7417
R54 VGND.n24 VGND.n23 24.8476
R55 VGND.n11 VGND.t6 24.7498
R56 VGND.n12 VGND.t1 24.7492
R57 VGND.n43 VGND.n41 22.9652
R58 VGND.n24 VGND.n6 14.6829
R59 VGND.n35 VGND.n34 14.6829
R60 VGND.n14 VGND.n13 13.9614
R61 VGND.n36 VGND.n1 12.424
R62 VGND.n19 VGND.n8 11.2946
R63 VGND.n13 VGND.n10 9.41227
R64 VGND.n41 VGND.n0 9.3005
R65 VGND.n40 VGND.n39 9.3005
R66 VGND.n38 VGND.n1 9.3005
R67 VGND.n37 VGND.n36 9.3005
R68 VGND.n35 VGND.n2 9.3005
R69 VGND.n34 VGND.n33 9.3005
R70 VGND.n32 VGND.n3 9.3005
R71 VGND.n31 VGND.n30 9.3005
R72 VGND.n29 VGND.n5 9.3005
R73 VGND.n28 VGND.n27 9.3005
R74 VGND.n26 VGND.n6 9.3005
R75 VGND.n25 VGND.n24 9.3005
R76 VGND.n23 VGND.n7 9.3005
R77 VGND.n22 VGND.n21 9.3005
R78 VGND.n20 VGND.n19 9.3005
R79 VGND.n18 VGND.n9 9.3005
R80 VGND.n17 VGND.n16 9.3005
R81 VGND.n15 VGND.n10 9.3005
R82 VGND.n44 VGND.n43 7.12063
R83 VGND.n22 VGND.n8 2.63579
R84 VGND.n15 VGND.n14 0.186831
R85 VGND.n44 VGND.n0 0.148519
R86 VGND.n16 VGND.n15 0.120292
R87 VGND.n16 VGND.n9 0.120292
R88 VGND.n20 VGND.n9 0.120292
R89 VGND.n21 VGND.n20 0.120292
R90 VGND.n21 VGND.n7 0.120292
R91 VGND.n25 VGND.n7 0.120292
R92 VGND.n26 VGND.n25 0.120292
R93 VGND.n27 VGND.n26 0.120292
R94 VGND.n27 VGND.n5 0.120292
R95 VGND.n31 VGND.n5 0.120292
R96 VGND.n32 VGND.n31 0.120292
R97 VGND.n33 VGND.n32 0.120292
R98 VGND.n33 VGND.n2 0.120292
R99 VGND.n37 VGND.n2 0.120292
R100 VGND.n38 VGND.n37 0.120292
R101 VGND.n39 VGND.n38 0.120292
R102 VGND.n39 VGND.n0 0.120292
R103 VGND VGND.n44 0.114842
R104 Q Q.t0 251.107
R105 Q Q.t1 146.542
R106 VNB.t2 VNB.t9 3460.19
R107 VNB.t6 VNB.t12 3203.88
R108 VNB.t7 VNB.t13 2890.61
R109 VNB.t12 VNB.t7 2677.02
R110 VNB.t4 VNB.t11 2677.02
R111 VNB.t15 VNB.t3 2677.02
R112 VNB.t0 VNB.t14 2591.59
R113 VNB.t5 VNB.t0 1452.43
R114 VNB.t9 VNB.t10 1381.23
R115 VNB.t1 VNB.t2 1381.23
R116 VNB.t13 VNB.t1 1352.75
R117 VNB.t14 VNB.t6 1253.07
R118 VNB.t11 VNB.t5 1253.07
R119 VNB.t8 VNB.t15 1196.12
R120 VNB.t3 VNB.t4 1025.24
R121 VNB VNB.t8 683.495
R122 DE.n0 DE.t2 319.728
R123 DE.n2 DE.n1 238.69
R124 DE.n0 DE.t0 178.34
R125 DE DE.n2 158.893
R126 DE.n1 DE.n0 147.814
R127 DE.n2 DE.t3 130.387
R128 DE.n1 DE.t1 130.141
R129 a_423_343.t0 a_423_343.n1 376.974
R130 a_423_343.n1 a_423_343.t3 375.568
R131 a_423_343.n0 a_423_343.t2 334.038
R132 a_423_343.n0 a_423_343.t1 244.181
R133 a_423_343.n1 a_423_343.n0 11.1343
R134 VPWR.n23 VPWR.t5 667.963
R135 VPWR.n43 VPWR.n1 604.394
R136 VPWR.n37 VPWR.t8 374.937
R137 VPWR.n35 VPWR.n5 323.079
R138 VPWR.n9 VPWR.n8 317.757
R139 VPWR.n15 VPWR.n14 245.905
R140 VPWR.n16 VPWR.n13 231.042
R141 VPWR.n8 VPWR.t0 106.1
R142 VPWR.n13 VPWR.t4 95.3126
R143 VPWR.n14 VPWR.t1 61.9802
R144 VPWR.n5 VPWR.t9 44.6333
R145 VPWR.n5 VPWR.t10 44.6333
R146 VPWR.n8 VPWR.t7 43.3405
R147 VPWR.n1 VPWR.t11 41.5552
R148 VPWR.n1 VPWR.t6 41.5552
R149 VPWR.n41 VPWR.n2 34.6358
R150 VPWR.n42 VPWR.n41 34.6358
R151 VPWR.n29 VPWR.n28 34.6358
R152 VPWR.n30 VPWR.n29 34.6358
R153 VPWR.n30 VPWR.n6 34.6358
R154 VPWR.n34 VPWR.n6 34.6358
R155 VPWR.n18 VPWR.n17 34.6358
R156 VPWR.n18 VPWR.n11 34.6358
R157 VPWR.n22 VPWR.n11 34.6358
R158 VPWR.n35 VPWR.n34 33.8829
R159 VPWR.n37 VPWR.n36 32.0005
R160 VPWR.n14 VPWR.t2 30.1762
R161 VPWR.n24 VPWR.n23 30.1181
R162 VPWR.n16 VPWR.n15 29.0203
R163 VPWR.n28 VPWR.n9 28.2358
R164 VPWR.n13 VPWR.t3 26.4482
R165 VPWR.n24 VPWR.n9 23.3417
R166 VPWR.n43 VPWR.n42 22.9652
R167 VPWR.n36 VPWR.n35 20.7064
R168 VPWR.n23 VPWR.n22 17.3181
R169 VPWR.n17 VPWR.n16 13.177
R170 VPWR.n37 VPWR.n2 12.424
R171 VPWR.n17 VPWR.n12 9.3005
R172 VPWR.n19 VPWR.n18 9.3005
R173 VPWR.n20 VPWR.n11 9.3005
R174 VPWR.n22 VPWR.n21 9.3005
R175 VPWR.n23 VPWR.n10 9.3005
R176 VPWR.n25 VPWR.n24 9.3005
R177 VPWR.n26 VPWR.n9 9.3005
R178 VPWR.n28 VPWR.n27 9.3005
R179 VPWR.n29 VPWR.n7 9.3005
R180 VPWR.n31 VPWR.n30 9.3005
R181 VPWR.n32 VPWR.n6 9.3005
R182 VPWR.n34 VPWR.n33 9.3005
R183 VPWR.n35 VPWR.n4 9.3005
R184 VPWR.n36 VPWR.n3 9.3005
R185 VPWR.n38 VPWR.n37 9.3005
R186 VPWR.n39 VPWR.n2 9.3005
R187 VPWR.n41 VPWR.n40 9.3005
R188 VPWR.n42 VPWR.n0 9.3005
R189 VPWR.n44 VPWR.n43 7.12063
R190 VPWR.n15 VPWR.n12 0.186831
R191 VPWR.n44 VPWR.n0 0.148519
R192 VPWR.n19 VPWR.n12 0.120292
R193 VPWR.n20 VPWR.n19 0.120292
R194 VPWR.n21 VPWR.n20 0.120292
R195 VPWR.n21 VPWR.n10 0.120292
R196 VPWR.n25 VPWR.n10 0.120292
R197 VPWR.n26 VPWR.n25 0.120292
R198 VPWR.n27 VPWR.n26 0.120292
R199 VPWR.n27 VPWR.n7 0.120292
R200 VPWR.n31 VPWR.n7 0.120292
R201 VPWR.n32 VPWR.n31 0.120292
R202 VPWR.n33 VPWR.n32 0.120292
R203 VPWR.n33 VPWR.n4 0.120292
R204 VPWR.n4 VPWR.n3 0.120292
R205 VPWR.n38 VPWR.n3 0.120292
R206 VPWR.n39 VPWR.n38 0.120292
R207 VPWR.n40 VPWR.n39 0.120292
R208 VPWR.n40 VPWR.n0 0.120292
R209 VPWR VPWR.n44 0.114842
R210 CLK.n0 CLK.t0 292.95
R211 CLK.n0 CLK.t1 209.403
R212 CLK CLK.n0 154.069
R213 a_27_47.n3 a_27_47.t5 443.44
R214 a_27_47.t1 a_27_47.n6 390.443
R215 a_27_47.n4 a_27_47.t6 344.428
R216 a_27_47.n4 a_27_47.t3 296.969
R217 a_27_47.n1 a_27_47.t0 288.373
R218 a_27_47.n0 a_27_47.t4 263.406
R219 a_27_47.n3 a_27_47.n2 254.389
R220 a_27_47.n0 a_27_47.t2 228.06
R221 a_27_47.n5 a_27_47.n3 194.501
R222 a_27_47.n1 a_27_47.n0 152
R223 a_27_47.n6 a_27_47.n1 35.3396
R224 a_27_47.n6 a_27_47.n5 13.284
R225 a_27_47.n5 a_27_47.n4 12.879
R226 a_193_47.t1 a_193_47.n5 395.625
R227 a_193_47.n3 a_193_47.t3 389.545
R228 a_193_47.n2 a_193_47.n0 308.651
R229 a_193_47.n5 a_193_47.t0 300.372
R230 a_193_47.n2 a_193_47.n1 298.373
R231 a_193_47.n3 a_193_47.t2 273.572
R232 a_193_47.n4 a_193_47.n3 173.755
R233 a_193_47.n5 a_193_47.n4 12.5786
R234 a_193_47.n4 a_193_47.n2 12.2528
R235 a_1514_47.n0 a_1514_47.t0 45.1697
R236 a_791_264.t1 a_791_264.n5 394.808
R237 a_791_264.n0 a_791_264.t3 368.969
R238 a_791_264.n3 a_791_264.t4 310.623
R239 a_791_264.n5 a_791_264.n2 308.443
R240 a_791_264.n1 a_791_264.t2 245.821
R241 a_791_264.n4 a_791_264.t0 241.077
R242 a_791_264.n4 a_791_264.n3 219.524
R243 a_791_264.n3 a_791_264.t6 194.942
R244 a_791_264.n0 a_791_264.t5 189.588
R245 a_791_264.n2 a_791_264.t7 152.633
R246 a_791_264.n1 a_791_264.n0 96.4005
R247 a_791_264.n2 a_791_264.n1 29.9627
R248 a_791_264.n5 a_791_264.n4 7.71815
R249 Q_N Q_N.t1 246.079
R250 Q_N Q_N.t0 148.946
R251 a_986_413.n3 a_986_413.n2 680.737
R252 a_986_413.n2 a_986_413.n1 276.272
R253 a_986_413.n0 a_986_413.t5 230.484
R254 a_986_413.n0 a_986_413.t4 196.013
R255 a_986_413.n2 a_986_413.n0 171.939
R256 a_986_413.t0 a_986_413.n3 72.7029
R257 a_986_413.n3 a_986_413.t3 70.3576
R258 a_986_413.n1 a_986_413.t2 51.6672
R259 a_986_413.n1 a_986_413.t1 45.0005
R260 a_1150_159.t1 a_1150_159.n4 408.848
R261 a_1150_159.n2 a_1150_159.t4 406.401
R262 a_1150_159.n0 a_1150_159.t2 318.12
R263 a_1150_159.n0 a_1150_159.t3 194.477
R264 a_1150_159.n3 a_1150_159.n2 176.534
R265 a_1150_159.n4 a_1150_159.n0 168.486
R266 a_1150_159.n3 a_1150_159.t0 140.249
R267 a_1150_159.n2 a_1150_159.n1 130.054
R268 a_1150_159.n4 a_1150_159.n3 9.32396
R269 a_729_47.t0 a_729_47.t1 102.858
R270 a_729_369.t0 a_729_369.t1 110.812
R271 a_1077_413.t0 a_1077_413.t1 171.202
R272 a_1717_47.t0 a_1717_47.t1 93.0601
R273 a_381_47.t0 a_381_47.t1 60.0005
C0 VPB VGND 0.015827f
C1 D DE 0.099354f
C2 CLK VPWR 0.019263f
C3 VPB Q_N 0.015582f
C4 CLK VGND 0.019296f
C5 D VPWR 0.01674f
C6 VPB Q 0.016876f
C7 D VGND 0.014495f
C8 DE VPWR 0.046893f
C9 a_1591_413# VPB 0.21251f
C10 DE VGND 0.057232f
C11 VPWR VGND 0.078008f
C12 VPWR Q_N 0.124307f
C13 VPWR Q 0.122443f
C14 VGND Q_N 0.097568f
C15 a_1591_413# VPWR 0.336655f
C16 a_1101_47# VGND 0.004436f
C17 VPB CLK 0.069635f
C18 VGND Q 0.100622f
C19 a_1591_413# VGND 0.18479f
C20 VPB D 0.068631f
C21 a_1591_413# Q_N 0.102624f
C22 VPB DE 0.114449f
C23 a_1591_413# Q 0.0374f
C24 VPB VPWR 0.275237f
C25 Q VNB 0.083148f
C26 Q_N VNB 0.012608f
C27 VGND VNB 1.33164f
C28 VPWR VNB 1.07887f
C29 DE VNB 0.282831f
C30 D VNB 0.122269f
C31 CLK VNB 0.195128f
C32 VPB VNB 2.37668f
C33 a_1591_413# VNB 0.287613f
.ends

* NGSPICE file created from sky130_fd_sc_hd__edfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__edfxtp_1 VPWR VGND CLK DE Q D VPB VNB
X0 a_381_369.t0 D.t0 a_299_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 VGND.t2 a_1591_413# a_791_264.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t1 DE.t0 a_423_343.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 VPWR.t8 CLK.t0 a_27_47.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_986_413.t2 a_193_47.t2 a_299_47.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.15985 ps=1.265 w=0.42 l=0.15
X5 Q.t1 a_1591_413# VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.154 ps=1.335 w=1 l=0.15
X6 VGND.t7 DE.t1 a_423_343.t0 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_1500_413.t0 a_1150_159.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_1101_47# a_193_47.t3 a_986_413.t3 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0759 pd=0.8 as=0.0522 ps=0.65 w=0.36 l=0.15
X9 a_1514_47.t0 a_1150_159.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0678 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 a_193_47.t0 a_27_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_729_47.t0 a_423_343.t2 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0609 ps=0.71 w=0.42 l=0.15
X12 a_729_369.t0 DE.t2 VPWR.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1152 pd=1 as=0.0928 ps=0.93 w=0.64 l=0.15
X13 a_1077_413.t1 a_27_47.t3 a_986_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06405 ps=0.725 w=0.42 l=0.15
X14 VPWR.t10 a_791_264.t2 a_1675_413# VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15 Q.t0 a_1591_413# VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10025 ps=0.985 w=0.65 l=0.15
X16 a_299_47.t4 a_791_264.t3 a_729_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1446 pd=1.18 as=0.0756 ps=0.78 w=0.42 l=0.15
X17 VPWR.t4 a_1591_413# a_791_264.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1728 ps=1.82 w=0.64 l=0.15
X18 VGND.t9 a_791_264.t4 a_1717_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X19 a_193_47.t1 a_27_47.t4 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VPWR.t5 a_1150_159.t4 a_1077_413.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X21 a_1717_47.t0 a_27_47.t5 a_1591_413# VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X22 a_1150_159.t1 a_986_413.t4 VPWR.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=2.02 as=0.178875 ps=1.26 w=0.75 l=0.15
X23 a_986_413.t1 a_27_47.t6 a_299_47.t3 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.0522 pd=0.65 as=0.1446 ps=1.18 w=0.36 l=0.15
X24 a_299_47.t5 a_791_264.t5 a_729_369.t1 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.15985 pd=1.265 as=0.1152 ps=1 w=0.64 l=0.15
X25 a_381_47.t1 D.t1 a_299_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 VPWR.t0 a_423_343.t3 a_381_369.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X27 VGND.t8 CLK.t1 a_27_47.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 VGND.t6 DE.t3 a_381_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X29 a_1150_159.t0 a_986_413.t5 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.12095 ps=1.085 w=0.64 l=0.15
R0 D.n0 D.t1 220.367
R1 D.n0 D.t0 216.796
R2 D D.n0 71.33
R3 a_299_47.t1 a_299_47.n3 467.892
R4 a_299_47.n2 a_299_47.n0 380.805
R5 a_299_47.n3 a_299_47.t0 232.434
R6 a_299_47.n0 a_299_47.t2 231.013
R7 a_299_47.n1 a_299_47.t3 208.333
R8 a_299_47.n2 a_299_47.n1 188.082
R9 a_299_47.n0 a_299_47.t5 41.1785
R10 a_299_47.n1 a_299_47.t4 28.3186
R11 a_299_47.n3 a_299_47.n2 20.4743
R12 a_381_369.t0 a_381_369.t1 64.6411
R13 VPB.t6 VPB.t11 855.297
R14 VPB.t11 VPB.t1 624.456
R15 VPB.t14 VPB.t6 556.386
R16 VPB.t5 VPB.t12 556.386
R17 VPB.t8 VPB.t4 556.386
R18 VPB.t10 VPB.t7 458.724
R19 VPB.t3 VPB.t14 390.654
R20 VPB.t0 VPB.t3 304.829
R21 VPB.t9 VPB.t10 301.87
R22 VPB.t1 VPB.t2 287.072
R23 VPB.t7 VPB.t0 269.315
R24 VPB.t12 VPB.t9 260.437
R25 VPB.t13 VPB.t8 248.599
R26 VPB.t4 VPB.t5 213.084
R27 VPB VPB.t13 142.056
R28 a_791_264.n2 a_791_264.t4 382.745
R29 a_791_264.t1 a_791_264.n3 362.808
R30 a_791_264.n0 a_791_264.t3 310.623
R31 a_791_264.n1 a_791_264.t0 242.322
R32 a_791_264.n1 a_791_264.n0 218.909
R33 a_791_264.n0 a_791_264.t5 194.942
R34 a_791_264.n3 a_791_264.n2 174.017
R35 a_791_264.n2 a_791_264.t2 138.53
R36 a_791_264.n3 a_791_264.n1 48.371
R37 VGND.n23 VGND.t4 273.476
R38 VGND.n8 VGND.t0 244.518
R39 VGND.n11 VGND.t9 241.857
R40 VGND.n35 VGND.t6 238.311
R41 VGND.n33 VGND.n4 202.262
R42 VGND.n42 VGND.n41 199.739
R43 VGND.n13 VGND.n12 124.519
R44 VGND.n12 VGND.t2 57.8184
R45 VGND.n4 VGND.t5 41.4291
R46 VGND.n4 VGND.t7 41.4291
R47 VGND.n41 VGND.t1 38.5719
R48 VGND.n41 VGND.t8 38.5719
R49 VGND.n16 VGND.n10 34.6358
R50 VGND.n17 VGND.n16 34.6358
R51 VGND.n18 VGND.n17 34.6358
R52 VGND.n22 VGND.n21 34.6358
R53 VGND.n27 VGND.n6 34.6358
R54 VGND.n28 VGND.n27 34.6358
R55 VGND.n29 VGND.n28 34.6358
R56 VGND.n29 VGND.n3 34.6358
R57 VGND.n39 VGND.n1 34.6358
R58 VGND.n40 VGND.n39 34.6358
R59 VGND.n35 VGND.n34 32.0005
R60 VGND.n33 VGND.n3 29.7417
R61 VGND.n23 VGND.n22 24.8476
R62 VGND.n12 VGND.t3 24.7498
R63 VGND.n42 VGND.n40 22.9652
R64 VGND.n23 VGND.n6 14.6829
R65 VGND.n34 VGND.n33 14.6829
R66 VGND.n35 VGND.n1 12.424
R67 VGND.n13 VGND.n11 11.8579
R68 VGND.n18 VGND.n8 11.2946
R69 VGND.n40 VGND.n0 9.3005
R70 VGND.n39 VGND.n38 9.3005
R71 VGND.n37 VGND.n1 9.3005
R72 VGND.n36 VGND.n35 9.3005
R73 VGND.n34 VGND.n2 9.3005
R74 VGND.n33 VGND.n32 9.3005
R75 VGND.n31 VGND.n3 9.3005
R76 VGND.n30 VGND.n29 9.3005
R77 VGND.n28 VGND.n5 9.3005
R78 VGND.n27 VGND.n26 9.3005
R79 VGND.n25 VGND.n6 9.3005
R80 VGND.n24 VGND.n23 9.3005
R81 VGND.n22 VGND.n7 9.3005
R82 VGND.n21 VGND.n20 9.3005
R83 VGND.n19 VGND.n18 9.3005
R84 VGND.n17 VGND.n9 9.3005
R85 VGND.n16 VGND.n15 9.3005
R86 VGND.n14 VGND.n10 9.3005
R87 VGND.n43 VGND.n42 7.12063
R88 VGND.n11 VGND.n10 6.02403
R89 VGND.n21 VGND.n8 2.63579
R90 VGND.n14 VGND.n13 0.754043
R91 VGND.n43 VGND.n0 0.148519
R92 VGND.n15 VGND.n14 0.120292
R93 VGND.n15 VGND.n9 0.120292
R94 VGND.n19 VGND.n9 0.120292
R95 VGND.n20 VGND.n19 0.120292
R96 VGND.n20 VGND.n7 0.120292
R97 VGND.n24 VGND.n7 0.120292
R98 VGND.n25 VGND.n24 0.120292
R99 VGND.n26 VGND.n25 0.120292
R100 VGND.n26 VGND.n5 0.120292
R101 VGND.n30 VGND.n5 0.120292
R102 VGND.n31 VGND.n30 0.120292
R103 VGND.n32 VGND.n31 0.120292
R104 VGND.n32 VGND.n2 0.120292
R105 VGND.n36 VGND.n2 0.120292
R106 VGND.n37 VGND.n36 0.120292
R107 VGND.n38 VGND.n37 0.120292
R108 VGND.n38 VGND.n0 0.120292
R109 VGND VGND.n43 0.114842
R110 VNB.t7 VNB.t5 3203.88
R111 VNB.t0 VNB.t8 2890.61
R112 VNB.t13 VNB.t3 2677.02
R113 VNB.t5 VNB.t0 2677.02
R114 VNB.t10 VNB.t11 2677.02
R115 VNB.t1 VNB.t4 2677.02
R116 VNB.t14 VNB.t9 2591.59
R117 VNB.t6 VNB.t14 1452.43
R118 VNB.t3 VNB.t2 1381.23
R119 VNB.t8 VNB.t13 1352.75
R120 VNB.t9 VNB.t7 1253.07
R121 VNB.t11 VNB.t6 1253.07
R122 VNB.t12 VNB.t1 1196.12
R123 VNB.t4 VNB.t10 1025.24
R124 VNB VNB.t12 683.495
R125 DE.n0 DE.t2 319.728
R126 DE.n2 DE.n1 238.69
R127 DE.n0 DE.t0 178.34
R128 DE DE.n2 158.893
R129 DE.n1 DE.n0 147.814
R130 DE.n2 DE.t3 130.387
R131 DE.n1 DE.t1 130.141
R132 a_423_343.t1 a_423_343.n1 376.974
R133 a_423_343.n1 a_423_343.t3 375.568
R134 a_423_343.n0 a_423_343.t2 334.038
R135 a_423_343.n0 a_423_343.t0 244.181
R136 a_423_343.n1 a_423_343.n0 11.1343
R137 VPWR.n15 VPWR.t10 671.345
R138 VPWR.n22 VPWR.t6 667.963
R139 VPWR.n42 VPWR.n1 604.394
R140 VPWR.n36 VPWR.t0 374.937
R141 VPWR.n34 VPWR.n5 323.079
R142 VPWR.n9 VPWR.n8 317.757
R143 VPWR.n14 VPWR.n13 246.773
R144 VPWR.n8 VPWR.t5 106.1
R145 VPWR.n13 VPWR.t4 61.9802
R146 VPWR.n5 VPWR.t2 44.6333
R147 VPWR.n5 VPWR.t1 44.6333
R148 VPWR.n8 VPWR.t9 43.3405
R149 VPWR.n1 VPWR.t7 41.5552
R150 VPWR.n1 VPWR.t8 41.5552
R151 VPWR.n40 VPWR.n2 34.6358
R152 VPWR.n41 VPWR.n40 34.6358
R153 VPWR.n28 VPWR.n27 34.6358
R154 VPWR.n29 VPWR.n28 34.6358
R155 VPWR.n29 VPWR.n6 34.6358
R156 VPWR.n33 VPWR.n6 34.6358
R157 VPWR.n17 VPWR.n16 34.6358
R158 VPWR.n17 VPWR.n11 34.6358
R159 VPWR.n21 VPWR.n11 34.6358
R160 VPWR.n34 VPWR.n33 33.8829
R161 VPWR.n36 VPWR.n35 32.0005
R162 VPWR.n13 VPWR.t3 30.1762
R163 VPWR.n23 VPWR.n22 30.1181
R164 VPWR.n27 VPWR.n9 28.2358
R165 VPWR.n23 VPWR.n9 23.3417
R166 VPWR.n42 VPWR.n41 22.9652
R167 VPWR.n15 VPWR.n14 21.2697
R168 VPWR.n35 VPWR.n34 20.7064
R169 VPWR.n22 VPWR.n21 17.3181
R170 VPWR.n36 VPWR.n2 12.424
R171 VPWR.n16 VPWR.n12 9.3005
R172 VPWR.n18 VPWR.n17 9.3005
R173 VPWR.n19 VPWR.n11 9.3005
R174 VPWR.n21 VPWR.n20 9.3005
R175 VPWR.n22 VPWR.n10 9.3005
R176 VPWR.n24 VPWR.n23 9.3005
R177 VPWR.n25 VPWR.n9 9.3005
R178 VPWR.n27 VPWR.n26 9.3005
R179 VPWR.n28 VPWR.n7 9.3005
R180 VPWR.n30 VPWR.n29 9.3005
R181 VPWR.n31 VPWR.n6 9.3005
R182 VPWR.n33 VPWR.n32 9.3005
R183 VPWR.n34 VPWR.n4 9.3005
R184 VPWR.n35 VPWR.n3 9.3005
R185 VPWR.n37 VPWR.n36 9.3005
R186 VPWR.n38 VPWR.n2 9.3005
R187 VPWR.n40 VPWR.n39 9.3005
R188 VPWR.n41 VPWR.n0 9.3005
R189 VPWR.n43 VPWR.n42 7.12063
R190 VPWR.n14 VPWR.n12 0.754043
R191 VPWR.n16 VPWR.n15 0.753441
R192 VPWR.n43 VPWR.n0 0.148519
R193 VPWR.n18 VPWR.n12 0.120292
R194 VPWR.n19 VPWR.n18 0.120292
R195 VPWR.n20 VPWR.n19 0.120292
R196 VPWR.n20 VPWR.n10 0.120292
R197 VPWR.n24 VPWR.n10 0.120292
R198 VPWR.n25 VPWR.n24 0.120292
R199 VPWR.n26 VPWR.n25 0.120292
R200 VPWR.n26 VPWR.n7 0.120292
R201 VPWR.n30 VPWR.n7 0.120292
R202 VPWR.n31 VPWR.n30 0.120292
R203 VPWR.n32 VPWR.n31 0.120292
R204 VPWR.n32 VPWR.n4 0.120292
R205 VPWR.n4 VPWR.n3 0.120292
R206 VPWR.n37 VPWR.n3 0.120292
R207 VPWR.n38 VPWR.n37 0.120292
R208 VPWR.n39 VPWR.n38 0.120292
R209 VPWR.n39 VPWR.n0 0.120292
R210 VPWR VPWR.n43 0.114842
R211 CLK.n0 CLK.t0 292.95
R212 CLK.n0 CLK.t1 209.403
R213 CLK CLK.n0 154.069
R214 a_27_47.n3 a_27_47.t5 443.44
R215 a_27_47.t1 a_27_47.n6 390.443
R216 a_27_47.n4 a_27_47.t6 344.428
R217 a_27_47.n4 a_27_47.t3 296.969
R218 a_27_47.n1 a_27_47.t0 288.373
R219 a_27_47.n0 a_27_47.t4 263.406
R220 a_27_47.n3 a_27_47.n2 254.389
R221 a_27_47.n0 a_27_47.t2 228.06
R222 a_27_47.n5 a_27_47.n3 194.501
R223 a_27_47.n1 a_27_47.n0 152
R224 a_27_47.n6 a_27_47.n1 35.3396
R225 a_27_47.n6 a_27_47.n5 13.284
R226 a_27_47.n5 a_27_47.n4 12.879
R227 a_193_47.t1 a_193_47.n5 395.625
R228 a_193_47.n3 a_193_47.t3 389.545
R229 a_193_47.n2 a_193_47.n0 308.651
R230 a_193_47.n5 a_193_47.t0 300.372
R231 a_193_47.n2 a_193_47.n1 298.373
R232 a_193_47.n3 a_193_47.t2 273.572
R233 a_193_47.n4 a_193_47.n3 173.755
R234 a_193_47.n5 a_193_47.n4 12.5786
R235 a_193_47.n4 a_193_47.n2 12.2528
R236 a_1514_47.n0 a_1514_47.t0 45.1697
R237 a_986_413.n3 a_986_413.n2 680.737
R238 a_986_413.n2 a_986_413.n1 276.272
R239 a_986_413.n0 a_986_413.t5 230.484
R240 a_986_413.n0 a_986_413.t4 196.013
R241 a_986_413.n2 a_986_413.n0 171.939
R242 a_986_413.t0 a_986_413.n3 72.7029
R243 a_986_413.n3 a_986_413.t2 70.3576
R244 a_986_413.n1 a_986_413.t3 51.6672
R245 a_986_413.n1 a_986_413.t1 45.0005
R246 Q Q.t1 251.107
R247 Q Q.t0 146.542
R248 a_1150_159.t1 a_1150_159.n4 408.848
R249 a_1150_159.n2 a_1150_159.t4 406.401
R250 a_1150_159.n0 a_1150_159.t2 318.12
R251 a_1150_159.n0 a_1150_159.t3 194.477
R252 a_1150_159.n3 a_1150_159.n2 176.534
R253 a_1150_159.n4 a_1150_159.n0 168.486
R254 a_1150_159.n3 a_1150_159.t0 140.249
R255 a_1150_159.n2 a_1150_159.n1 130.054
R256 a_1150_159.n4 a_1150_159.n3 9.32396
R257 a_729_47.t0 a_729_47.t1 102.858
R258 a_729_369.t0 a_729_369.t1 110.812
R259 a_1077_413.t0 a_1077_413.t1 171.202
R260 a_1717_47.t1 a_1717_47.t0 93.0601
R261 a_381_47.t0 a_381_47.t1 60.0005
C0 VPB VPWR 0.25415f
C1 CLK VPWR 0.019263f
C2 D DE 0.099354f
C3 VPB VGND 0.013019f
C4 VPB Q 0.013891f
C5 CLK VGND 0.019296f
C6 D VPWR 0.01674f
C7 VPB a_1591_413# 0.147526f
C8 D VGND 0.014495f
C9 DE VPWR 0.046893f
C10 DE VGND 0.057232f
C11 VPWR VGND 0.061718f
C12 a_1675_413# VPWR 0.004673f
C13 VPWR Q 0.122606f
C14 VPWR a_1591_413# 0.160369f
C15 VGND Q 0.092175f
C16 VGND a_1591_413# 0.173214f
C17 VPB CLK 0.069635f
C18 a_1101_47# VGND 0.004436f
C19 a_1675_413# a_1591_413# 0.008717f
C20 Q a_1591_413# 0.036123f
C21 VPB D 0.068631f
C22 VPB DE 0.114449f
C23 Q VNB 0.084065f
C24 VGND VNB 1.23098f
C25 VPWR VNB 0.992377f
C26 DE VNB 0.282831f
C27 D VNB 0.122269f
C28 CLK VNB 0.195128f
C29 VPB VNB 2.19949f
C30 a_1591_413# VNB 0.312829f
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_8 VGND VPWR VPB VNB A Z TE_B
X0 a_204_309.t8 A.t0 Z.t10 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t7 a_27_47.t2 a_215_47.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_215_47.t7 A.t1 Z.t13 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Z.t9 A.t2 a_204_309.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t6 a_27_47.t3 a_215_47.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t5 a_27_47.t4 a_215_47.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_204_309.t13 TE_B.t0 VPWR.t7 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X7 a_204_309.t6 A.t3 Z.t8 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t4 a_27_47.t5 a_215_47.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR.t6 TE_B.t1 a_204_309.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X10 Z.t7 A.t4 a_204_309.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_204_309.t11 TE_B.t2 VPWR.t5 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X12 a_215_47.t11 a_27_47.t6 VGND.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Z.t12 A.t5 a_215_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X14 a_215_47.t10 a_27_47.t7 VGND.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_215_47.t9 a_27_47.t8 VGND.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t4 TE_B.t3 a_204_309.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X17 a_215_47.t5 A.t6 Z.t11 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_204_309.t15 TE_B.t4 VPWR.t3 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.16025 ps=1.325 w=0.94 l=0.15
X19 a_215_47.t4 A.t7 Z.t14 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_215_47.t3 A.t8 Z.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_204_309.t4 A.t9 Z.t6 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR.t2 TE_B.t5 a_204_309.t14 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.2444 pd=2.4 as=0.1269 ps=1.21 w=0.94 l=0.15
X23 a_204_309.t0 TE_B.t6 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X24 Z.t5 A.t10 a_204_309.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Z.t1 A.t11 a_215_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Z.t4 A.t12 a_204_309.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 a_204_309.t1 A.t13 Z.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Z.t15 A.t14 a_215_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VPWR.t0 TE_B.t7 a_204_309.t12 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1269 pd=1.21 as=0.1269 ps=1.21 w=0.94 l=0.15
X30 Z.t2 A.t15 a_215_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_215_47.t8 a_27_47.t9 VGND.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 VPWR.t8 TE_B.t8 a_27_47.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.16025 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X33 VGND.t8 TE_B.t9 a_27_47.t1 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A.n3 A.t0 212.081
R1 A.n2 A.t2 212.081
R2 A.n1 A.t3 212.081
R3 A.n11 A.t4 212.081
R4 A.n13 A.t9 212.081
R5 A.n22 A.t10 212.081
R6 A.n15 A.t13 212.081
R7 A.n16 A.t12 212.081
R8 A A.n4 157.518
R9 A.n6 A.n5 152
R10 A.n8 A.n7 152
R11 A.n10 A.n9 152
R12 A.n12 A.n0 152
R13 A.n24 A.n23 152
R14 A.n21 A.n20 152
R15 A.n19 A.n14 152
R16 A.n18 A.n17 152
R17 A.n3 A.t1 139.78
R18 A.n2 A.t15 139.78
R19 A.n1 A.t8 139.78
R20 A.n11 A.t14 139.78
R21 A.n13 A.t7 139.78
R22 A.n22 A.t11 139.78
R23 A.n15 A.t6 139.78
R24 A.n16 A.t5 139.78
R25 A.n7 A.n6 49.6611
R26 A.n21 A.n14 49.6611
R27 A.n17 A.n15 48.2005
R28 A.n10 A.n1 45.2793
R29 A.n4 A.n2 42.3581
R30 A.n23 A.n22 39.4369
R31 A.n12 A.n11 33.5944
R32 A.n13 A.n12 27.752
R33 A.n23 A.n13 21.9096
R34 A.n4 A.n3 18.9884
R35 A.n11 A.n10 16.0672
R36 A.n9 A.n8 15.0074
R37 A.n20 A.n19 15.0074
R38 A A.n0 13.9039
R39 A.n17 A.n16 13.146
R40 A A.n18 13.0212
R41 A.n24 A 11.6971
R42 A.n5 A 10.8143
R43 A.n22 A.n21 10.2247
R44 A.n5 A 9.49016
R45 A A.n24 8.6074
R46 A.n6 A.n2 7.30353
R47 A.n18 A 7.28326
R48 A A.n0 6.4005
R49 A.n7 A.n1 4.38232
R50 A.n8 A 4.1936
R51 A.n20 A 3.31084
R52 A.n19 A 1.98671
R53 A.n15 A.n14 1.46111
R54 A.n9 A 1.10395
R55 Z.n2 Z.n0 340.368
R56 Z.n2 Z.n1 301.966
R57 Z.n15 Z.n14 294.132
R58 Z.n11 Z.n10 294.132
R59 Z.n5 Z.n3 237.45
R60 Z.n9 Z.n8 185
R61 Z.n7 Z.n6 185
R62 Z.n5 Z.n4 185
R63 Z.n9 Z.n7 52.4493
R64 Z.n7 Z.n5 52.4493
R65 Z.n12 Z 43.5707
R66 Z.n13 Z.n2 38.4005
R67 Z.n13 Z.n12 38.4005
R68 Z Z.n9 28.4727
R69 Z.n10 Z.t10 26.5955
R70 Z.n10 Z.t9 26.5955
R71 Z.n0 Z.t3 26.5955
R72 Z.n0 Z.t4 26.5955
R73 Z.n1 Z.t6 26.5955
R74 Z.n1 Z.t5 26.5955
R75 Z.n14 Z.t8 26.5955
R76 Z.n14 Z.t7 26.5955
R77 Z.n3 Z.t11 24.9236
R78 Z.n3 Z.t12 24.9236
R79 Z.n4 Z.t14 24.9236
R80 Z.n4 Z.t1 24.9236
R81 Z.n6 Z.t0 24.9236
R82 Z.n6 Z.t15 24.9236
R83 Z.n8 Z.t13 24.9236
R84 Z.n8 Z.t2 24.9236
R85 Z.n15 Z.n13 7.83717
R86 Z.n12 Z.n11 7.83717
R87 Z Z.n15 1.65867
R88 Z.n11 Z 1.65867
R89 a_204_309.t8 a_204_309.n13 382.825
R90 a_204_309.n7 a_204_309.n6 367.474
R91 a_204_309.n10 a_204_309.t2 352.606
R92 a_204_309.n9 a_204_309.n3 310.058
R93 a_204_309.n8 a_204_309.n4 310.058
R94 a_204_309.n7 a_204_309.n5 310.058
R95 a_204_309.n11 a_204_309.n2 298.673
R96 a_204_309.n12 a_204_309.n1 298.673
R97 a_204_309.n13 a_204_309.n0 298.673
R98 a_204_309.n10 a_204_309.n9 78.9851
R99 a_204_309.n11 a_204_309.n10 76.9672
R100 a_204_309.n9 a_204_309.n8 63.2476
R101 a_204_309.n8 a_204_309.n7 63.2476
R102 a_204_309.n13 a_204_309.n12 63.2476
R103 a_204_309.n12 a_204_309.n11 63.2476
R104 a_204_309.n6 a_204_309.t9 28.2931
R105 a_204_309.n6 a_204_309.t15 28.2931
R106 a_204_309.n3 a_204_309.t14 28.2931
R107 a_204_309.n3 a_204_309.t0 28.2931
R108 a_204_309.n4 a_204_309.t12 28.2931
R109 a_204_309.n4 a_204_309.t13 28.2931
R110 a_204_309.n5 a_204_309.t10 28.2931
R111 a_204_309.n5 a_204_309.t11 28.2931
R112 a_204_309.n2 a_204_309.t3 26.5955
R113 a_204_309.n2 a_204_309.t1 26.5955
R114 a_204_309.n1 a_204_309.t5 26.5955
R115 a_204_309.n1 a_204_309.t4 26.5955
R116 a_204_309.n0 a_204_309.t7 26.5955
R117 a_204_309.n0 a_204_309.t6 26.5955
R118 VPB.t15 VPB.t2 556.386
R119 VPB.t12 VPB.t16 281.154
R120 VPB.t7 VPB.t8 248.599
R121 VPB.t6 VPB.t7 248.599
R122 VPB.t5 VPB.t6 248.599
R123 VPB.t4 VPB.t5 248.599
R124 VPB.t3 VPB.t4 248.599
R125 VPB.t1 VPB.t3 248.599
R126 VPB.t2 VPB.t1 248.599
R127 VPB.t0 VPB.t15 248.599
R128 VPB.t13 VPB.t0 248.599
R129 VPB.t14 VPB.t13 248.599
R130 VPB.t10 VPB.t14 248.599
R131 VPB.t11 VPB.t10 248.599
R132 VPB.t9 VPB.t11 248.599
R133 VPB.t16 VPB.t9 248.599
R134 VPB VPB.t12 189.409
R135 a_27_47.t0 a_27_47.n7 395.608
R136 a_27_47.n7 a_27_47.n6 292.606
R137 a_27_47.n0 a_27_47.t2 263.493
R138 a_27_47.n7 a_27_47.t1 241.649
R139 a_27_47.n5 a_27_47.n4 134.96
R140 a_27_47.n4 a_27_47.n3 134.96
R141 a_27_47.n3 a_27_47.n2 134.96
R142 a_27_47.n2 a_27_47.n1 134.96
R143 a_27_47.n1 a_27_47.n0 134.96
R144 a_27_47.n6 a_27_47.t8 134.476
R145 a_27_47.n0 a_27_47.t9 128.534
R146 a_27_47.n1 a_27_47.t3 128.534
R147 a_27_47.n2 a_27_47.t6 128.534
R148 a_27_47.n3 a_27_47.t4 128.534
R149 a_27_47.n4 a_27_47.t7 128.534
R150 a_27_47.n5 a_27_47.t5 128.534
R151 a_27_47.n6 a_27_47.n5 94.9479
R152 a_215_47.t7 a_215_47.n13 323.711
R153 a_215_47.n3 a_215_47.t15 275.303
R154 a_215_47.n3 a_215_47.n2 192.154
R155 a_215_47.n4 a_215_47.n1 192.154
R156 a_215_47.n5 a_215_47.n0 192.154
R157 a_215_47.n7 a_215_47.n6 185
R158 a_215_47.n13 a_215_47.n12 185
R159 a_215_47.n11 a_215_47.n10 185
R160 a_215_47.n9 a_215_47.n8 185
R161 a_215_47.n7 a_215_47.n5 68.3168
R162 a_215_47.n5 a_215_47.n4 63.2476
R163 a_215_47.n4 a_215_47.n3 63.2476
R164 a_215_47.n9 a_215_47.n7 62.0618
R165 a_215_47.n13 a_215_47.n11 55.139
R166 a_215_47.n11 a_215_47.n9 55.139
R167 a_215_47.n6 a_215_47.t9 30.462
R168 a_215_47.n6 a_215_47.t6 29.539
R169 a_215_47.n8 a_215_47.t2 24.9236
R170 a_215_47.n8 a_215_47.t5 24.9236
R171 a_215_47.n10 a_215_47.t1 24.9236
R172 a_215_47.n10 a_215_47.t4 24.9236
R173 a_215_47.n12 a_215_47.t0 24.9236
R174 a_215_47.n12 a_215_47.t3 24.9236
R175 a_215_47.n2 a_215_47.t14 24.9236
R176 a_215_47.n2 a_215_47.t8 24.9236
R177 a_215_47.n1 a_215_47.t13 24.9236
R178 a_215_47.n1 a_215_47.t11 24.9236
R179 a_215_47.n0 a_215_47.t12 24.9236
R180 a_215_47.n0 a_215_47.t10 24.9236
R181 VGND.n16 VGND.t8 282.817
R182 VGND.n5 VGND.n4 203.927
R183 VGND.n7 VGND.n6 198.964
R184 VGND.n10 VGND.n9 198.964
R185 VGND.n14 VGND.n2 198.964
R186 VGND.n10 VGND.n8 27.4829
R187 VGND.n4 VGND.t1 24.9236
R188 VGND.n4 VGND.t4 24.9236
R189 VGND.n6 VGND.t2 24.9236
R190 VGND.n6 VGND.t5 24.9236
R191 VGND.n9 VGND.t3 24.9236
R192 VGND.n9 VGND.t6 24.9236
R193 VGND.n2 VGND.t0 24.9236
R194 VGND.n2 VGND.t7 24.9236
R195 VGND.n15 VGND.n14 22.9652
R196 VGND.n16 VGND.n15 22.9652
R197 VGND.n14 VGND.n1 21.4593
R198 VGND.n10 VGND.n1 16.9417
R199 VGND.n8 VGND.n7 10.9181
R200 VGND.n8 VGND.n3 9.3005
R201 VGND.n11 VGND.n10 9.3005
R202 VGND.n12 VGND.n1 9.3005
R203 VGND.n14 VGND.n13 9.3005
R204 VGND.n15 VGND.n0 9.3005
R205 VGND.n17 VGND.n16 7.12063
R206 VGND.n7 VGND.n5 6.70383
R207 VGND.n5 VGND.n3 0.949634
R208 VGND.n17 VGND.n0 0.148519
R209 VGND.n11 VGND.n3 0.120292
R210 VGND.n12 VGND.n11 0.120292
R211 VGND.n13 VGND.n12 0.120292
R212 VGND.n13 VGND.n0 0.120292
R213 VGND VGND.n17 0.11354
R214 VNB.t16 VNB.t15 2677.02
R215 VNB.t9 VNB.t6 1352.75
R216 VNB.t0 VNB.t7 1196.12
R217 VNB.t3 VNB.t0 1196.12
R218 VNB.t1 VNB.t3 1196.12
R219 VNB.t4 VNB.t1 1196.12
R220 VNB.t2 VNB.t4 1196.12
R221 VNB.t5 VNB.t2 1196.12
R222 VNB.t6 VNB.t5 1196.12
R223 VNB.t12 VNB.t9 1196.12
R224 VNB.t10 VNB.t12 1196.12
R225 VNB.t13 VNB.t10 1196.12
R226 VNB.t11 VNB.t13 1196.12
R227 VNB.t14 VNB.t11 1196.12
R228 VNB.t8 VNB.t14 1196.12
R229 VNB.t15 VNB.t8 1196.12
R230 VNB VNB.t16 911.327
R231 TE_B.n0 TE_B.t5 310.087
R232 TE_B.n7 TE_B.t8 220.391
R233 TE_B.n6 TE_B.t4 199.227
R234 TE_B.n0 TE_B.t6 175.127
R235 TE_B.n1 TE_B.t7 175.127
R236 TE_B.n2 TE_B.t0 175.127
R237 TE_B.n3 TE_B.t1 175.127
R238 TE_B.n4 TE_B.t2 175.127
R239 TE_B.n5 TE_B.t3 175.127
R240 TE_B.n8 TE_B.t9 158.064
R241 TE_B TE_B.n8 155.685
R242 TE_B.n7 TE_B.n6 151.028
R243 TE_B.n1 TE_B.n0 134.96
R244 TE_B.n2 TE_B.n1 134.96
R245 TE_B.n3 TE_B.n2 134.96
R246 TE_B.n4 TE_B.n3 134.96
R247 TE_B.n5 TE_B.n4 134.96
R248 TE_B.n6 TE_B.n5 110.861
R249 TE_B.n8 TE_B.n7 9.97291
R250 VPWR.n6 VPWR.t2 342.474
R251 VPWR.n14 VPWR.n3 309.726
R252 VPWR.n5 VPWR.n4 309.726
R253 VPWR.n8 VPWR.n7 309.726
R254 VPWR.n16 VPWR.n1 309.724
R255 VPWR.n1 VPWR.t3 39.8196
R256 VPWR.n9 VPWR.n5 30.8711
R257 VPWR.n3 VPWR.t5 28.2931
R258 VPWR.n3 VPWR.t4 28.2931
R259 VPWR.n4 VPWR.t7 28.2931
R260 VPWR.n4 VPWR.t6 28.2931
R261 VPWR.n7 VPWR.t1 28.2931
R262 VPWR.n7 VPWR.t0 28.2931
R263 VPWR.n1 VPWR.t8 26.4528
R264 VPWR.n14 VPWR.n13 24.8476
R265 VPWR.n16 VPWR.n15 22.9652
R266 VPWR.n15 VPWR.n14 19.577
R267 VPWR.n13 VPWR.n5 13.5534
R268 VPWR.n10 VPWR.n9 9.3005
R269 VPWR.n11 VPWR.n5 9.3005
R270 VPWR.n13 VPWR.n12 9.3005
R271 VPWR.n14 VPWR.n2 9.3005
R272 VPWR.n15 VPWR.n0 9.3005
R273 VPWR.n8 VPWR.n6 8.81261
R274 VPWR.n9 VPWR.n8 7.52991
R275 VPWR.n17 VPWR.n16 7.12063
R276 VPWR.n10 VPWR.n6 1.13618
R277 VPWR.n17 VPWR.n0 0.148519
R278 VPWR.n11 VPWR.n10 0.120292
R279 VPWR.n12 VPWR.n11 0.120292
R280 VPWR.n12 VPWR.n2 0.120292
R281 VPWR.n2 VPWR.n0 0.120292
R282 VPWR VPWR.n17 0.11354
C0 VPB TE_B 0.314762f
C1 Z VGND 0.045018f
C2 VPB A 0.252814f
C3 VPB VPWR 0.151265f
C4 TE_B A 0.005873f
C5 TE_B VPWR 0.175367f
C6 VPB Z 0.016173f
C7 TE_B Z 9.66e-19
C8 A VPWR 0.064359f
C9 A Z 0.69974f
C10 VPWR Z 0.040461f
C11 VPB VGND 0.009343f
C12 TE_B VGND 0.031971f
C13 A VGND 0.070001f
C14 VPWR VGND 0.15867f
C15 VGND VNB 0.882253f
C16 Z VNB 0.060563f
C17 VPWR VNB 0.7361f
C18 A VNB 0.747622f
C19 TE_B VNB 0.444885f
C20 VPB VNB 1.66792f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_4 VNB VPB VGND VPWR X D C B A
X0 VPWR.t5 a_27_47.t5 X.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t5 a_27_47.t6 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_188_47.t0 B.t0 a_109_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.079625 ps=0.895 w=0.65 l=0.15
X3 VPWR.t3 a_27_47.t7 X.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t0 D.t0 a_285_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.141375 ps=1.085 w=0.65 l=0.15
X5 VPWR.t6 D.t1 a_27_47.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.215 ps=1.43 w=1 l=0.15
X6 X.t3 a_27_47.t8 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X7 VGND.t4 a_27_47.t9 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t7 B.t1 a_27_47.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t1 a_27_47.t10 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X10 X.t7 a_27_47.t11 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_47.t0 C.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.155 ps=1.31 w=1 l=0.15
X12 VGND.t1 a_27_47.t12 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_47.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 a_285_47.t1 C.t1 a_188_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.085 as=0.108875 ps=0.985 w=0.65 l=0.15
X15 a_109_47.t1 A.t1 a_27_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.079625 pd=0.895 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n1 a_27_47.t3 336.387
R1 a_27_47.n12 a_27_47.n11 323.716
R2 a_27_47.n1 a_27_47.n0 315.574
R3 a_27_47.n3 a_27_47.t5 212.081
R4 a_27_47.n5 a_27_47.t6 212.081
R5 a_27_47.n7 a_27_47.t7 212.081
R6 a_27_47.n8 a_27_47.t8 212.081
R7 a_27_47.n4 a_27_47.n2 170.923
R8 a_27_47.n10 a_27_47.n9 152
R9 a_27_47.n6 a_27_47.n2 152
R10 a_27_47.n3 a_27_47.t12 139.78
R11 a_27_47.n5 a_27_47.t11 139.78
R12 a_27_47.n7 a_27_47.t9 139.78
R13 a_27_47.n8 a_27_47.t10 139.78
R14 a_27_47.n11 a_27_47.n10 90.7455
R15 a_27_47.n11 a_27_47.n1 59.8593
R16 a_27_47.n12 a_27_47.t2 58.1155
R17 a_27_47.n9 a_27_47.n8 48.2005
R18 a_27_47.n4 a_27_47.n3 36.5157
R19 a_27_47.n7 a_27_47.n6 36.5157
R20 a_27_47.n0 a_27_47.t4 26.5955
R21 a_27_47.n0 a_27_47.t1 26.5955
R22 a_27_47.t0 a_27_47.n12 26.5955
R23 a_27_47.n5 a_27_47.n4 24.8308
R24 a_27_47.n6 a_27_47.n5 24.8308
R25 a_27_47.n10 a_27_47.n2 18.9222
R26 a_27_47.n9 a_27_47.n7 13.146
R27 X.n2 X.n1 370.786
R28 X.n2 X.n0 314.952
R29 X.n5 X.n4 264.812
R30 X.n5 X.n3 201.565
R31 X X.n5 27.6485
R32 X.n1 X.t4 26.5955
R33 X.n1 X.t3 26.5955
R34 X.n0 X.t6 26.5955
R35 X.n0 X.t5 26.5955
R36 X.n4 X.t2 24.9236
R37 X.n4 X.t1 24.9236
R38 X.n3 X.t0 24.9236
R39 X.n3 X.t7 24.9236
R40 X X.n2 17.7236
R41 VPWR.n5 VPWR.t5 343.545
R42 VPWR.n15 VPWR.t1 340.301
R43 VPWR.n7 VPWR.n6 316.245
R44 VPWR.n13 VPWR.n2 309.726
R45 VPWR.n4 VPWR.n3 309.726
R46 VPWR.n3 VPWR.t6 36.4455
R47 VPWR.n8 VPWR.n7 32.0005
R48 VPWR.n12 VPWR.n4 31.2476
R49 VPWR.n2 VPWR.t0 30.5355
R50 VPWR.n2 VPWR.t7 30.5355
R51 VPWR.n3 VPWR.t2 28.5655
R52 VPWR.n6 VPWR.t4 26.5955
R53 VPWR.n6 VPWR.t3 26.5955
R54 VPWR.n13 VPWR.n12 24.4711
R55 VPWR.n15 VPWR.n14 22.9652
R56 VPWR.n14 VPWR.n13 19.9534
R57 VPWR.n8 VPWR.n4 13.177
R58 VPWR.n9 VPWR.n8 9.3005
R59 VPWR.n10 VPWR.n4 9.3005
R60 VPWR.n12 VPWR.n11 9.3005
R61 VPWR.n13 VPWR.n1 9.3005
R62 VPWR.n14 VPWR.n0 9.3005
R63 VPWR.n16 VPWR.n15 9.3005
R64 VPWR.n7 VPWR.n5 6.18988
R65 VPWR.n9 VPWR.n5 0.755914
R66 VPWR.n10 VPWR.n9 0.120292
R67 VPWR.n11 VPWR.n10 0.120292
R68 VPWR.n11 VPWR.n1 0.120292
R69 VPWR.n1 VPWR.n0 0.120292
R70 VPWR.n16 VPWR.n0 0.120292
R71 VPWR VPWR.n16 0.0213333
R72 VPB.t0 VPB.t6 343.303
R73 VPB.t6 VPB.t2 284.113
R74 VPB.t7 VPB.t0 272.274
R75 VPB.t4 VPB.t5 248.599
R76 VPB.t3 VPB.t4 248.599
R77 VPB.t2 VPB.t3 248.599
R78 VPB.t1 VPB.t7 248.599
R79 VPB VPB.t1 189.409
R80 B.n0 B.t1 241.536
R81 B B.n0 178.501
R82 B.n0 B.t0 169.237
R83 a_109_47.t0 a_109_47.t1 45.2313
R84 a_188_47.t0 a_188_47.t1 61.8467
R85 VNB.t6 VNB.t0 1666.02
R86 VNB.t5 VNB.t6 1381.23
R87 VNB.t0 VNB.t3 1352.75
R88 VNB.t2 VNB.t1 1196.12
R89 VNB.t4 VNB.t2 1196.12
R90 VNB.t3 VNB.t4 1196.12
R91 VNB.t7 VNB.t5 1124.92
R92 VNB VNB.t7 911.327
R93 D.n0 D.t1 241.536
R94 D D.n0 177.645
R95 D.n0 D.t0 164.952
R96 a_285_47.t0 a_285_47.t1 80.3082
R97 VGND.n1 VGND.t1 287.151
R98 VGND.n6 VGND.n5 200.898
R99 VGND.n3 VGND.n2 199.934
R100 VGND.n5 VGND.t0 33.2313
R101 VGND.n5 VGND.t3 26.7697
R102 VGND.n4 VGND.n3 25.977
R103 VGND.n2 VGND.t2 24.9236
R104 VGND.n2 VGND.t4 24.9236
R105 VGND.n6 VGND.n4 14.6829
R106 VGND.n4 VGND.n0 9.3005
R107 VGND.n7 VGND.n6 7.4819
R108 VGND.n3 VGND.n1 6.18988
R109 VGND.n1 VGND.n0 0.755914
R110 VGND VGND.n7 0.474279
R111 VGND.n7 VGND.n0 0.149004
R112 C.n0 C.t0 233.869
R113 C C.n0 185.012
R114 C.n0 C.t1 161.57
R115 A.n0 A.t0 230.363
R116 A.n0 A.t1 158.064
R117 A A.n0 153.367
C0 A VGND 0.013036f
C1 C VPWR 0.021684f
C2 B VGND 0.04486f
C3 D VPWR 0.021123f
C4 C X 0.004863f
C5 D X 0.009906f
C6 C VGND 0.048255f
C7 VPWR X 0.34457f
C8 D VGND 0.036941f
C9 VPB A 0.040083f
C10 VPWR VGND 0.084805f
C11 VPB B 0.026482f
C12 X VGND 0.229133f
C13 A B 0.05441f
C14 VPB C 0.033087f
C15 VPB D 0.028488f
C16 VPB VPWR 0.091263f
C17 B C 0.135912f
C18 VPB X 0.011564f
C19 B D 1.74e-20
C20 A VPWR 0.045725f
C21 VPB VGND 0.007761f
C22 C D 0.092843f
C23 B VPWR 0.022049f
C24 VGND VNB 0.488494f
C25 X VNB 0.070035f
C26 VPWR VNB 0.439634f
C27 D VNB 0.093185f
C28 C VNB 0.102095f
C29 B VNB 0.091991f
C30 A VNB 0.166716f
C31 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VPB VNB
X0 a_297_47.t1 a_27_47.t2 a_193_413.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47.t0 B.t0 a_297_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR.t5 D.t0 a_193_413.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X.t0 a_193_413.t5 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR.t3 A_N.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND.t1 D.t1 a_469_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X.t1 a_193_413.t6 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR.t4 B.t1 a_193_413.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413.t0 C.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413.t2 a_27_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47.t1 C.t1 a_369_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND.t2 A_N.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t0 a_27_47.n1 748.431
R1 a_27_47.n0 a_27_47.t3 334.723
R2 a_27_47.n0 a_27_47.t2 302.226
R3 a_27_47.n1 a_27_47.t1 293.671
R4 a_27_47.n1 a_27_47.n0 152
R5 a_193_413.n2 a_193_413.n1 604.201
R6 a_193_413.n4 a_193_413.n3 604.201
R7 a_193_413.n2 a_193_413.t1 329.884
R8 a_193_413.n3 a_193_413.n0 243.323
R9 a_193_413.n0 a_193_413.t6 241.536
R10 a_193_413.n0 a_193_413.t5 169.237
R11 a_193_413.n1 a_193_413.t2 126.644
R12 a_193_413.n3 a_193_413.n2 97.1299
R13 a_193_413.n1 a_193_413.t4 93.81
R14 a_193_413.t0 a_193_413.n4 84.4291
R15 a_193_413.n4 a_193_413.t3 63.3219
R16 a_297_47.t0 a_297_47.t1 60.0005
R17 VNB.t5 VNB.t2 2677.02
R18 VNB.t4 VNB.t1 1423.95
R19 VNB.t0 VNB.t3 1423.95
R20 VNB.t3 VNB.t4 1253.07
R21 VNB.t2 VNB.t0 1025.24
R22 VNB VNB.t5 925.567
R23 B.n0 B.t1 295.432
R24 B.n0 B.t0 237.591
R25 B.n1 B.n0 152
R26 B B.n1 8.0005
R27 B.n1 B 7.54336
R28 a_369_47.t0 a_369_47.t1 100.001
R29 D.n0 D.t0 334.723
R30 D.n0 D.t1 206.19
R31 D.n1 D.n0 152
R32 D.n1 D 10.7299
R33 D D.n1 2.07109
R34 VPWR.n7 VPWR.n3 606.444
R35 VPWR.n11 VPWR.n1 599.74
R36 VPWR.n4 VPWR.n2 585
R37 VPWR.n6 VPWR.n5 585
R38 VPWR.n5 VPWR.n4 159.476
R39 VPWR.n3 VPWR.t5 77.3934
R40 VPWR.n5 VPWR.t1 63.3219
R41 VPWR.n4 VPWR.t4 63.3219
R42 VPWR.n1 VPWR.t2 63.3219
R43 VPWR.n1 VPWR.t3 63.3219
R44 VPWR.n3 VPWR.t0 41.0422
R45 VPWR.n10 VPWR.n9 31.7084
R46 VPWR.n11 VPWR.n10 22.9652
R47 VPWR.n9 VPWR.n8 9.3005
R48 VPWR.n10 VPWR.n0 9.3005
R49 VPWR.n6 VPWR.n2 7.50395
R50 VPWR.n12 VPWR.n11 7.12063
R51 VPWR.n7 VPWR.n6 7.08138
R52 VPWR.n9 VPWR.n2 2.42809
R53 VPWR.n8 VPWR.n7 0.541003
R54 VPWR.n12 VPWR.n0 0.148519
R55 VPWR.n8 VPWR.n0 0.120292
R56 VPWR VPWR.n12 0.114842
R57 VPB.t4 VPB.t1 449.844
R58 VPB.t2 VPB.t4 366.978
R59 VPB.t5 VPB.t0 281.154
R60 VPB.t1 VPB.t5 275.235
R61 VPB.t3 VPB.t2 248.599
R62 VPB VPB.t3 192.369
R63 VGND.n1 VGND.t2 244.058
R64 VGND.n1 VGND.n0 205.976
R65 VGND.n0 VGND.t0 48.2862
R66 VGND.n0 VGND.t1 38.5719
R67 VGND VGND.n1 0.150529
R68 X.n1 X.t1 831.25
R69 X X.t1 735.458
R70 X.n0 X.t0 129.381
R71 X.n1 X.n0 68.6033
R72 X X.n1 6.15435
R73 X.n0 X 5.55208
R74 A_N.n0 A_N.t0 323.342
R75 A_N.n0 A_N.t1 194.809
R76 A_N.n1 A_N.n0 152
R77 A_N.n1 A_N 9.99502
R78 A_N A_N.n1 1.92927
R79 a_469_47.t0 a_469_47.t1 82.8576
R80 C.n0 C.t0 334.723
R81 C.n0 C.t1 206.19
R82 C.n1 C.n0 152
R83 C.n1 C 13.5116
R84 C C.n1 2.60791
C0 A_N VGND 0.020461f
C1 C VPWR 0.018191f
C2 D VPWR 0.018629f
C3 B VGND 0.036983f
C4 C X 0.004788f
C5 C VGND 0.039547f
C6 D X 0.016779f
C7 VPWR X 0.058561f
C8 D VGND 0.037199f
C9 VPB A_N 0.083174f
C10 VPWR VGND 0.072666f
C11 VPB B 0.088954f
C12 X VGND 0.05878f
C13 VPB C 0.07419f
C14 VPB D 0.076273f
C15 VPB VPWR 0.081835f
C16 B C 0.164206f
C17 A_N VPWR 0.020016f
C18 VPB X 0.010757f
C19 B VPWR 0.01856f
C20 C D 0.182698f
C21 VPB VGND 0.012312f
C22 VGND VNB 0.45592f
C23 X VNB 0.093393f
C24 VPWR VNB 0.367773f
C25 D VNB 0.123324f
C26 C VNB 0.107609f
C27 B VNB 0.120082f
C28 A_N VNB 0.198396f
C29 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND VNB VPB A_N B C D X
X0 VPWR.t3 a_193_413.t5 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47.t0 a_27_413.t2 a_193_413.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_369_47.t0 B.t0 a_297_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X.t1 a_193_413.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X4 VPWR.t6 D.t0 a_193_413.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X5 VPWR.t1 A_N.t0 a_27_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND.t3 D.t1 a_469_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X7 VGND.t1 a_193_413.t7 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X8 VPWR.t5 B.t1 a_193_413.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X9 a_193_413.t0 C.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X10 X.t2 a_193_413.t8 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X11 a_193_413.t2 a_27_413.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_469_47.t1 C.t1 a_369_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13 a_27_413.t1 A_N.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_193_413.n5 a_193_413.n4 607.588
R1 a_193_413.n1 a_193_413.n0 604.816
R2 a_193_413.n1 a_193_413.t1 328.62
R3 a_193_413.n4 a_193_413.n3 246.508
R4 a_193_413.n2 a_193_413.t5 212.081
R5 a_193_413.n3 a_193_413.t8 212.081
R6 a_193_413.n0 a_193_413.t3 157.131
R7 a_193_413.n2 a_193_413.t7 139.78
R8 a_193_413.n3 a_193_413.t6 139.78
R9 a_193_413.n4 a_193_413.n1 84.7064
R10 a_193_413.t0 a_193_413.n5 84.4291
R11 a_193_413.n3 a_193_413.n2 66.4581
R12 a_193_413.n0 a_193_413.t2 63.3219
R13 a_193_413.n5 a_193_413.t4 63.3219
R14 X X.n0 595.928
R15 X.n4 X.n0 585
R16 X X.n1 185.534
R17 X.n0 X.t2 33.4905
R18 X.n1 X.t1 31.3851
R19 X.n0 X.t3 26.5955
R20 X.n1 X.t0 24.9236
R21 X X.n3 20.7838
R22 X X.n2 11.8945
R23 X.n4 X 10.9273
R24 X X.n4 10.3029
R25 X.n3 X 4.87669
R26 X.n2 X 2.13383
R27 X.n3 X 1.82907
R28 X.n2 X 1.55202
R29 VPWR.n16 VPWR.n1 599.74
R30 VPWR.n6 VPWR.n5 599.74
R31 VPWR.n8 VPWR.n2 585
R32 VPWR.n10 VPWR.n9 585
R33 VPWR.n4 VPWR.t3 343.332
R34 VPWR.n9 VPWR.n8 159.476
R35 VPWR.n5 VPWR.t6 91.4648
R36 VPWR.n9 VPWR.t0 63.3219
R37 VPWR.n8 VPWR.t5 63.3219
R38 VPWR.n1 VPWR.t4 63.3219
R39 VPWR.n1 VPWR.t1 63.3219
R40 VPWR.n15 VPWR.n14 31.7746
R41 VPWR.n5 VPWR.t2 27.9557
R42 VPWR.n11 VPWR.n7 26.5725
R43 VPWR.n7 VPWR.n6 23.3417
R44 VPWR.n16 VPWR.n15 22.9652
R45 VPWR.n7 VPWR.n3 9.3005
R46 VPWR.n12 VPWR.n11 9.3005
R47 VPWR.n14 VPWR.n13 9.3005
R48 VPWR.n15 VPWR.n0 9.3005
R49 VPWR.n10 VPWR.n2 7.91323
R50 VPWR.n17 VPWR.n16 7.12063
R51 VPWR.n6 VPWR.n4 6.40813
R52 VPWR.n14 VPWR.n2 2.5605
R53 VPWR.n4 VPWR.n3 0.71136
R54 VPWR.n11 VPWR.n10 0.233227
R55 VPWR.n17 VPWR.n0 0.148519
R56 VPWR.n12 VPWR.n3 0.120292
R57 VPWR.n13 VPWR.n12 0.120292
R58 VPWR.n13 VPWR.n0 0.120292
R59 VPWR VPWR.n17 0.11354
R60 VPB.t5 VPB.t0 449.844
R61 VPB.t4 VPB.t5 366.978
R62 VPB.t6 VPB.t2 284.113
R63 VPB.t0 VPB.t6 275.235
R64 VPB.t2 VPB.t3 269.315
R65 VPB.t1 VPB.t4 248.599
R66 VPB VPB.t1 189.409
R67 a_27_413.t0 a_27_413.n1 749.78
R68 a_27_413.n0 a_27_413.t3 334.723
R69 a_27_413.n0 a_27_413.t2 305.803
R70 a_27_413.n1 a_27_413.t1 270.712
R71 a_27_413.n1 a_27_413.n0 152
R72 a_297_47.t0 a_297_47.t1 60.0005
R73 VNB.t1 VNB.t0 2677.02
R74 VNB.t5 VNB.t3 1423.95
R75 VNB.t4 VNB.t6 1423.95
R76 VNB.t3 VNB.t2 1295.79
R77 VNB.t6 VNB.t5 1267.31
R78 VNB.t0 VNB.t4 1025.24
R79 VNB VNB.t1 911.327
R80 B.n1 B.t0 255.46
R81 B.n0 B.t1 191.802
R82 B B.n0 159.856
R83 B.n2 B.n1 152
R84 B.n1 B.n0 44.2924
R85 B B.n2 11.9278
R86 B.n2 B 7.85505
R87 a_369_47.t0 a_369_47.t1 100.001
R88 VGND.n3 VGND.t1 289.204
R89 VGND.n13 VGND.t0 238.311
R90 VGND.n5 VGND.n4 199.739
R91 VGND.n4 VGND.t2 47.7807
R92 VGND.n4 VGND.t3 38.5719
R93 VGND.n7 VGND.n6 34.6358
R94 VGND.n7 VGND.n1 34.6358
R95 VGND.n11 VGND.n1 34.6358
R96 VGND.n12 VGND.n11 34.6358
R97 VGND.n13 VGND.n12 19.9534
R98 VGND.n6 VGND.n5 17.3181
R99 VGND.n14 VGND.n13 9.3005
R100 VGND.n6 VGND.n2 9.3005
R101 VGND.n8 VGND.n7 9.3005
R102 VGND.n9 VGND.n1 9.3005
R103 VGND.n11 VGND.n10 9.3005
R104 VGND.n12 VGND.n0 9.3005
R105 VGND.n5 VGND.n3 6.80788
R106 VGND.n3 VGND.n2 0.629752
R107 VGND.n8 VGND.n2 0.120292
R108 VGND.n9 VGND.n8 0.120292
R109 VGND.n10 VGND.n9 0.120292
R110 VGND.n10 VGND.n0 0.120292
R111 VGND.n14 VGND.n0 0.120292
R112 VGND VGND.n14 0.0213333
R113 D.n0 D.t0 334.723
R114 D.n0 D.t1 206.19
R115 D D.n0 163.055
R116 A_N.n0 A_N.t0 323.55
R117 A_N.n0 A_N.t1 195.017
R118 A_N.n1 A_N.n0 152
R119 A_N.n1 A_N 18.2405
R120 A_N A_N.n1 3.5205
R121 a_469_47.t0 a_469_47.t1 84.2862
R122 C.n0 C.t0 332.692
R123 C.n0 C.t1 204.157
R124 C C.n0 168.052
C0 VPB B 0.090475f
C1 X VGND 0.129318f
C2 VPB C 0.073665f
C3 VPB D 0.078106f
C4 B C 0.177533f
C5 VPB VPWR 0.093168f
C6 A_N VPWR 0.018806f
C7 VPB X 0.008732f
C8 B D 1.04e-19
C9 C D 0.184579f
C10 VPB VGND 0.013296f
C11 B VPWR 0.018993f
C12 A_N VGND 0.037344f
C13 C VPWR 0.018708f
C14 B VGND 0.033927f
C15 D VPWR 0.019096f
C16 C X 0.004267f
C17 D X 0.01879f
C18 C VGND 0.044472f
C19 VPWR X 0.148268f
C20 D VGND 0.036311f
C21 VPB A_N 0.080669f
C22 VPWR VGND 0.082543f
C23 VGND VNB 0.516815f
C24 X VNB 0.06398f
C25 VPWR VNB 0.421195f
C26 D VNB 0.121638f
C27 C VNB 0.109763f
C28 B VNB 0.121022f
C29 A_N VNB 0.207062f
C30 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4b_4 VNB VPB VGND VPWR A_N X D C B
X0 VPWR.t8 a_174_21.t5 X.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t1 a_174_21.t6 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_815_47.t0 B.t0 a_701_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR.t6 a_174_21.t7 X.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t4 C.t0 a_174_21.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X5 a_174_21.t2 a_27_47.t2 a_815_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.143 ps=1.09 w=0.65 l=0.15
X6 X.t7 a_174_21.t8 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR.t0 A_N.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_701_47.t1 C.t1 a_617_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_174_21.t0 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3275 ps=1.655 w=1 l=0.15
X10 a_174_21.t1 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.21 ps=1.42 w=1 l=0.15
X11 VPWR.t3 a_27_47.t3 a_174_21.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.22 ps=1.44 w=1 l=0.15
X12 X.t6 a_174_21.t9 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13 X.t5 a_174_21.t10 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_617_47.t1 D.t1 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.212875 ps=1.305 w=0.65 l=0.15
X15 VGND.t3 a_174_21.t11 X.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t2 a_174_21.t12 X.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.212875 pd=1.305 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t0 A_N.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_174_21.n10 a_174_21.n0 672.341
R1 a_174_21.n11 a_174_21.n10 585
R2 a_174_21.n9 a_174_21.t2 319.707
R3 a_174_21.n7 a_174_21.t5 212.081
R4 a_174_21.n5 a_174_21.t6 212.081
R5 a_174_21.n3 a_174_21.t7 212.081
R6 a_174_21.n2 a_174_21.t8 212.081
R7 a_174_21.n4 a_174_21.n1 177.601
R8 a_174_21.n8 a_174_21.n7 163.685
R9 a_174_21.n6 a_174_21.n1 152
R10 a_174_21.n7 a_174_21.t12 139.78
R11 a_174_21.n5 a_174_21.t10 139.78
R12 a_174_21.n3 a_174_21.t11 139.78
R13 a_174_21.n2 a_174_21.t9 139.78
R14 a_174_21.n10 a_174_21.n9 79.4358
R15 a_174_21.n3 a_174_21.n2 61.346
R16 a_174_21.n0 a_174_21.t1 60.0855
R17 a_174_21.n7 a_174_21.n6 37.9763
R18 a_174_21.n4 a_174_21.n3 35.055
R19 a_174_21.n0 a_174_21.t3 26.5955
R20 a_174_21.n11 a_174_21.t4 26.5955
R21 a_174_21.t0 a_174_21.n11 26.5955
R22 a_174_21.n5 a_174_21.n4 26.2914
R23 a_174_21.n8 a_174_21.n1 25.6005
R24 a_174_21.n6 a_174_21.n5 23.3702
R25 a_174_21.n9 a_174_21.n8 13.5534
R26 X.n2 X.n0 640.341
R27 X.n2 X.n1 585
R28 X.n5 X.n3 257.659
R29 X.n5 X.n4 206.203
R30 X.n1 X.t0 26.5955
R31 X.n1 X.t7 26.5955
R32 X.n0 X.t2 26.5955
R33 X.n0 X.t1 26.5955
R34 X.n3 X.t4 24.9236
R35 X.n3 X.t5 24.9236
R36 X.n4 X.t3 24.9236
R37 X.n4 X.t6 24.9236
R38 X X.n2 8.45764
R39 X X.n5 1.37193
R40 VPWR.n8 VPWR.t3 875.422
R41 VPWR.n18 VPWR.n1 599.74
R42 VPWR.n16 VPWR.n3 599.74
R43 VPWR.n5 VPWR.n4 599.74
R44 VPWR.n9 VPWR.n7 599.74
R45 VPWR.n4 VPWR.t1 102.441
R46 VPWR.n1 VPWR.t0 63.3219
R47 VPWR.n7 VPWR.t2 56.1455
R48 VPWR.n1 VPWR.t5 55.1136
R49 VPWR.n11 VPWR.n10 34.6358
R50 VPWR.n11 VPWR.n5 30.8711
R51 VPWR.n3 VPWR.t7 26.5955
R52 VPWR.n3 VPWR.t6 26.5955
R53 VPWR.n4 VPWR.t8 26.5955
R54 VPWR.n7 VPWR.t4 26.5955
R55 VPWR.n16 VPWR.n15 24.8476
R56 VPWR.n18 VPWR.n17 22.9652
R57 VPWR.n17 VPWR.n16 19.577
R58 VPWR.n9 VPWR.n8 15.081
R59 VPWR.n15 VPWR.n5 13.5534
R60 VPWR.n10 VPWR.n6 9.3005
R61 VPWR.n12 VPWR.n11 9.3005
R62 VPWR.n13 VPWR.n5 9.3005
R63 VPWR.n15 VPWR.n14 9.3005
R64 VPWR.n16 VPWR.n2 9.3005
R65 VPWR.n17 VPWR.n0 9.3005
R66 VPWR.n19 VPWR.n18 7.12063
R67 VPWR.n10 VPWR.n9 1.88285
R68 VPWR.n8 VPWR.n6 0.554787
R69 VPWR.n19 VPWR.n0 0.148519
R70 VPWR.n12 VPWR.n6 0.120292
R71 VPWR.n13 VPWR.n12 0.120292
R72 VPWR.n14 VPWR.n13 0.120292
R73 VPWR.n14 VPWR.n2 0.120292
R74 VPWR.n2 VPWR.n0 0.120292
R75 VPWR VPWR.n19 0.11354
R76 VPB.t8 VPB.t1 476.481
R77 VPB.t2 VPB.t3 349.221
R78 VPB.t4 VPB.t2 337.384
R79 VPB.t0 VPB.t5 281.154
R80 VPB.t1 VPB.t4 248.599
R81 VPB.t7 VPB.t8 248.599
R82 VPB.t6 VPB.t7 248.599
R83 VPB.t5 VPB.t6 248.599
R84 VPB VPB.t0 189.409
R85 B.n0 B.t1 241.536
R86 B.n0 B.t0 169.237
R87 B B.n0 154.133
R88 a_701_47.t0 a_701_47.t1 77.539
R89 a_815_47.t0 a_815_47.t1 81.2313
R90 VNB.t5 VNB.t0 2292.56
R91 VNB.t1 VNB.t4 1680.26
R92 VNB.t2 VNB.t1 1623.3
R93 VNB.t3 VNB.t8 1352.75
R94 VNB.t0 VNB.t2 1196.12
R95 VNB.t7 VNB.t5 1196.12
R96 VNB.t6 VNB.t7 1196.12
R97 VNB.t8 VNB.t6 1196.12
R98 VNB VNB.t3 911.327
R99 C.n0 C.t0 241.536
R100 C.n0 C.t1 169.237
R101 C C.n0 155.352
R102 a_27_47.t0 a_27_47.n1 663.091
R103 a_27_47.n1 a_27_47.n0 545.413
R104 a_27_47.n1 a_27_47.t1 333.159
R105 a_27_47.n0 a_27_47.t3 230.363
R106 a_27_47.n0 a_27_47.t2 158.064
R107 A_N.n0 A_N.t0 334.723
R108 A_N.n0 A_N.t1 206.19
R109 A_N.n1 A_N.n0 152
R110 A_N.n1 A_N 10.4234
R111 A_N A_N.n1 2.01193
R112 a_617_47.t0 a_617_47.t1 49.8467
R113 D.n0 D.t0 241.536
R114 D.n0 D.t1 169.237
R115 D D.n0 155.201
R116 VGND.n2 VGND.n1 204.256
R117 VGND.n4 VGND.n3 199.934
R118 VGND.n7 VGND.n6 199.739
R119 VGND.n1 VGND.t1 89.539
R120 VGND.n6 VGND.t0 54.2862
R121 VGND.n1 VGND.t2 31.3851
R122 VGND.n6 VGND.t5 25.9346
R123 VGND.n3 VGND.t4 24.9236
R124 VGND.n3 VGND.t3 24.9236
R125 VGND.n5 VGND.n4 19.577
R126 VGND.n7 VGND.n5 18.824
R127 VGND.n5 VGND.n0 9.3005
R128 VGND.n8 VGND.n7 7.32436
R129 VGND.n4 VGND.n2 6.68071
R130 VGND.n2 VGND.n0 0.628824
R131 VGND.n8 VGND.n0 0.145929
R132 VGND VGND.n8 0.116164
C0 VPB D 0.029682f
C1 X VGND 0.182187f
C2 VPB C 0.027405f
C3 VPB B 0.030373f
C4 A_N C 2.66e-20
C5 VPB VPWR 0.103284f
C6 D C 0.080037f
C7 A_N B 3.49e-20
C8 D B 4.65e-20
C9 VPB X 0.00496f
C10 A_N VPWR 0.020042f
C11 D VPWR 0.011777f
C12 C B 0.072661f
C13 VPB VGND 0.008857f
C14 A_N X 0.072262f
C15 A_N VGND 0.041506f
C16 C VPWR 0.012506f
C17 D VGND 0.009398f
C18 B VPWR 0.014791f
C19 C VGND 0.009666f
C20 B VGND 0.01114f
C21 VPWR X 0.02985f
C22 VPB A_N 0.090699f
C23 VPWR VGND 0.103639f
C24 VGND VNB 0.56902f
C25 X VNB 0.01178f
C26 VPWR VNB 0.486711f
C27 B VNB 0.106329f
C28 C VNB 0.094442f
C29 D VNB 0.094593f
C30 A_N VNB 0.16501f
C31 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4bb_1 VNB VPB VGND VPWR A_N B_N C D X
X0 VPWR.t2 D.t0 a_343_93.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47.t1 B_N.t0 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93.t0 a_223_47.t2 a_429_93.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47.t0 B_N.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR.t6 A_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND.t2 A_N.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X.t0 a_343_93.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93.t0 a_27_47.t2 a_343_93.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND.t1 D.t1 a_615_93.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93.t1 C.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93.t3 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93.t0 C.t1 a_515_93.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X.t1 a_343_93.t6 VGND.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR.t4 a_223_47.t3 a_343_93.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 D.n0 D.t0 334.723
R1 D.n1 D.n0 152
R2 D.n0 D.t1 132.282
R3 D.n1 D 16.1598
R4 D D.n1 2.76128
R5 a_343_93.n3 a_343_93.n1 601.188
R6 a_343_93.n4 a_343_93.n0 601.188
R7 a_343_93.t0 a_343_93.n4 317.348
R8 a_343_93.n3 a_343_93.n2 265.695
R9 a_343_93.n2 a_343_93.t5 224.805
R10 a_343_93.n2 a_343_93.t6 152.506
R11 a_343_93.n1 a_343_93.t2 93.81
R12 a_343_93.n1 a_343_93.t1 79.7386
R13 a_343_93.n4 a_343_93.n3 71.9064
R14 a_343_93.n0 a_343_93.t3 68.0124
R15 a_343_93.n0 a_343_93.t4 63.3219
R16 VPWR.n2 VPWR.t3 677.133
R17 VPWR.n6 VPWR.n5 605.394
R18 VPWR.n14 VPWR.n1 599.74
R19 VPWR.n7 VPWR.n4 599.74
R20 VPWR.n5 VPWR.t2 152.44
R21 VPWR.n4 VPWR.t1 89.1195
R22 VPWR.n4 VPWR.t4 75.0481
R23 VPWR.n1 VPWR.t5 68.0124
R24 VPWR.n1 VPWR.t6 63.3219
R25 VPWR.n13 VPWR.n12 34.6358
R26 VPWR.n9 VPWR.n8 34.6358
R27 VPWR.n5 VPWR.t0 27.9557
R28 VPWR.n7 VPWR.n6 14.0546
R29 VPWR.n14 VPWR.n13 12.424
R30 VPWR.n8 VPWR.n3 9.3005
R31 VPWR.n10 VPWR.n9 9.3005
R32 VPWR.n12 VPWR.n11 9.3005
R33 VPWR.n13 VPWR.n0 9.3005
R34 VPWR.n15 VPWR.n14 7.57378
R35 VPWR.n9 VPWR.n2 5.64756
R36 VPWR.n12 VPWR.n2 4.14168
R37 VPWR.n8 VPWR.n7 3.01226
R38 VPWR.n6 VPWR.n3 0.453385
R39 VPWR.n15 VPWR.n0 0.142757
R40 VPWR VPWR.n15 0.120679
R41 VPWR.n10 VPWR.n3 0.120292
R42 VPWR.n11 VPWR.n10 0.120292
R43 VPWR.n11 VPWR.n0 0.120292
R44 VPB.t5 VPB.t3 609.658
R45 VPB.t2 VPB.t0 361.06
R46 VPB.t1 VPB.t2 307.788
R47 VPB.t4 VPB.t1 295.95
R48 VPB VPB.t6 275.235
R49 VPB.t3 VPB.t4 254.518
R50 VPB.t6 VPB.t5 254.518
R51 B_N.n0 B_N.t1 376.399
R52 B_N B_N.n0 186.6
R53 B_N.n0 B_N.t0 164.319
R54 VGND.n2 VGND.n0 208.91
R55 VGND.n2 VGND.n1 205.202
R56 VGND.n0 VGND.t1 94.2862
R57 VGND.n1 VGND.t3 41.4291
R58 VGND.n1 VGND.t2 38.5719
R59 VGND.n0 VGND.t0 24.0005
R60 VGND VGND.n2 0.167403
R61 a_223_47.t0 a_223_47.n1 847.066
R62 a_223_47.n0 a_223_47.t3 334.723
R63 a_223_47.n1 a_223_47.n0 284.82
R64 a_223_47.n1 a_223_47.t1 243.571
R65 a_223_47.n0 a_223_47.t2 132.282
R66 VNB.t6 VNB.t0 2933.33
R67 VNB.t4 VNB.t3 1737.22
R68 VNB.t2 VNB.t4 1480.91
R69 VNB.t1 VNB.t2 1423.95
R70 VNB VNB.t5 1324.27
R71 VNB.t0 VNB.t1 1224.6
R72 VNB.t5 VNB.t6 1224.6
R73 a_429_93.t0 a_429_93.t1 80.0005
R74 a_515_93.t0 a_515_93.t1 100.001
R75 A_N.n0 A_N.t1 392.466
R76 A_N A_N.n0 153.647
R77 A_N.n0 A_N.t0 148.252
R78 a_27_47.t0 a_27_47.n1 773.312
R79 a_27_47.n1 a_27_47.t1 324.401
R80 a_27_47.n1 a_27_47.n0 305.635
R81 a_27_47.n0 a_27_47.t2 188.114
R82 a_27_47.n0 a_27_47.t3 166.692
R83 X X.n0 593.615
R84 X.n1 X.n0 585
R85 X X.t1 226.966
R86 X.n0 X.t0 26.5955
R87 X.n1 X 8.61589
R88 X X.n1 8.12358
R89 a_615_93.t0 a_615_93.t1 105.715
R90 C.n0 C.t0 334.723
R91 C.n1 C.n0 152
R92 C.n0 C.t1 132.282
R93 C.n1 C 17.4858
R94 C C.n1 3.06137
C0 VPB D 0.081017f
C1 VPB VPWR 0.1059f
C2 B_N C 9.56e-20
C3 VPB X 0.010318f
C4 A_N VPWR 0.031836f
C5 B_N D 6.67e-20
C6 VPB VGND 0.01669f
C7 C D 0.16344f
C8 B_N VPWR 0.016829f
C9 B_N X 4.64e-20
C10 A_N VGND 0.014613f
C11 C VPWR 0.012039f
C12 D VPWR 0.014287f
C13 B_N VGND 0.04274f
C14 C VGND 0.024978f
C15 D X 0.019253f
C16 VPWR X 0.058176f
C17 D VGND 0.041448f
C18 VPB A_N 0.084844f
C19 VPWR VGND 0.090642f
C20 VPB B_N 0.064623f
C21 X VGND 0.060874f
C22 A_N B_N 0.117058f
C23 VPB C 0.068601f
C24 VGND VNB 0.553085f
C25 X VNB 0.090815f
C26 VPWR VNB 0.453229f
C27 D VNB 0.124261f
C28 C VNB 0.106642f
C29 B_N VNB 0.134007f
C30 A_N VNB 0.143769f
C31 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4bb_2 VNB VPB VGND VPWR A_N X C D B_N
X0 a_174_21.t1 C.t0 VPWR.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21.t2 a_27_47.t2 VPWR.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X2 a_476_47.t1 a_27_47.t3 a_174_21.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VPWR.t1 a_174_21.t5 X.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X4 X.t2 a_174_21.t6 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X5 a_548_47.t1 a_505_280.t2 a_476_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR.t6 A_N.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 X.t0 a_174_21.t7 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR.t0 D.t0 a_174_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND.t0 D.t1 a_639_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR.t7 a_505_280.t3 a_174_21.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280.t0 B_N.t0 VPWR.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND.t3 a_174_21.t8 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_505_280.t1 B_N.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47.t0 C.t1 a_548_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X15 VGND.t2 A_N.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 C.n0 C.t0 405.416
R1 C.n1 C.n0 152
R2 C.n0 C.t1 135.496
R3 C.n1 C 8.45333
R4 C C.n1 7.97031
R5 VPWR.n6 VPWR.n5 605.337
R6 VPWR.n15 VPWR.n1 599.74
R7 VPWR.n8 VPWR.n7 599.307
R8 VPWR.n3 VPWR.n2 310.861
R9 VPWR.n5 VPWR.t0 143.06
R10 VPWR.n2 VPWR.t1 90.683
R11 VPWR.n7 VPWR.t4 68.0124
R12 VPWR.n1 VPWR.t6 63.3219
R13 VPWR.n7 VPWR.t7 63.3219
R14 VPWR.n5 VPWR.t3 63.3219
R15 VPWR.n1 VPWR.t2 55.1136
R16 VPWR.n2 VPWR.t5 35.1791
R17 VPWR.n10 VPWR.n9 29.9539
R18 VPWR.n14 VPWR.n13 28.3932
R19 VPWR.n15 VPWR.n14 22.9652
R20 VPWR.n9 VPWR.n8 15.4358
R21 VPWR.n9 VPWR.n4 9.3005
R22 VPWR.n11 VPWR.n10 9.3005
R23 VPWR.n13 VPWR.n12 9.3005
R24 VPWR.n14 VPWR.n0 9.3005
R25 VPWR.n16 VPWR.n15 7.12063
R26 VPWR.n8 VPWR.n6 6.98891
R27 VPWR.n10 VPWR.n3 5.67624
R28 VPWR.n13 VPWR.n3 4.97806
R29 VPWR.n6 VPWR.n4 0.500932
R30 VPWR.n16 VPWR.n0 0.148519
R31 VPWR.n11 VPWR.n4 0.120292
R32 VPWR.n12 VPWR.n11 0.120292
R33 VPWR.n12 VPWR.n0 0.120292
R34 VPWR VPWR.n16 0.11354
R35 a_174_21.n5 a_174_21.n4 665.188
R36 a_174_21.n4 a_174_21.n0 601.188
R37 a_174_21.n3 a_174_21.n2 243.249
R38 a_174_21.n3 a_174_21.t3 239.761
R39 a_174_21.n2 a_174_21.t5 212.081
R40 a_174_21.n1 a_174_21.t6 212.081
R41 a_174_21.n2 a_174_21.t8 139.78
R42 a_174_21.n1 a_174_21.t7 139.78
R43 a_174_21.n4 a_174_21.n3 112.566
R44 a_174_21.n0 a_174_21.t2 86.7743
R45 a_174_21.n0 a_174_21.t4 63.3219
R46 a_174_21.t0 a_174_21.n5 63.3219
R47 a_174_21.n5 a_174_21.t1 63.3219
R48 a_174_21.n2 a_174_21.n1 61.346
R49 VPB.t6 VPB.t3 506.075
R50 VPB.t0 VPB.t1 349.221
R51 VPB.t4 VPB.t5 281.154
R52 VPB.t3 VPB.t7 278.193
R53 VPB.t7 VPB.t2 254.518
R54 VPB.t2 VPB.t0 248.599
R55 VPB.t5 VPB.t6 248.599
R56 VPB VPB.t4 189.409
R57 a_27_47.n1 a_27_47.t1 691.24
R58 a_27_47.t0 a_27_47.n1 345.548
R59 a_27_47.n0 a_27_47.t2 326.762
R60 a_27_47.n1 a_27_47.n0 295.473
R61 a_27_47.n0 a_27_47.t3 149.409
R62 a_476_47.t0 a_476_47.t1 60.0005
R63 VNB.t5 VNB.t7 2677.02
R64 VNB.t0 VNB.t2 1680.26
R65 VNB.t1 VNB.t6 1352.75
R66 VNB.t4 VNB.t3 1295.79
R67 VNB.t3 VNB.t0 1196.12
R68 VNB.t6 VNB.t5 1196.12
R69 VNB.t7 VNB.t4 1025.24
R70 VNB VNB.t1 911.327
R71 X X.n0 595.524
R72 X X.n1 204.627
R73 X.n0 X.t3 26.5955
R74 X.n0 X.t2 26.5955
R75 X.n1 X.t1 24.9236
R76 X.n1 X.t0 24.9236
R77 a_505_280.t0 a_505_280.n1 663.091
R78 a_505_280.n0 a_505_280.t2 336.329
R79 a_505_280.n1 a_505_280.t1 336.021
R80 a_505_280.n1 a_505_280.n0 285.647
R81 a_505_280.n0 a_505_280.t3 204.583
R82 a_548_47.t0 a_548_47.t1 87.1434
R83 A_N.n0 A_N.t0 323.342
R84 A_N.n0 A_N.t1 194.809
R85 A_N.n1 A_N.n0 152
R86 A_N.n1 A_N 20.2672
R87 A_N A_N.n1 3.91161
R88 VGND.n3 VGND.t3 282.817
R89 VGND.n2 VGND.n1 213.007
R90 VGND.n6 VGND.n5 199.739
R91 VGND.n1 VGND.t0 87.1434
R92 VGND.n5 VGND.t4 41.6488
R93 VGND.n1 VGND.t1 38.5719
R94 VGND.n5 VGND.t2 38.5719
R95 VGND.n6 VGND.n4 22.9652
R96 VGND.n4 VGND.n3 19.577
R97 VGND.n4 VGND.n0 9.3005
R98 VGND.n3 VGND.n2 7.20206
R99 VGND.n7 VGND.n6 7.12063
R100 VGND.n2 VGND.n0 0.155249
R101 VGND.n7 VGND.n0 0.148519
R102 VGND VGND.n7 0.11354
R103 D.n0 D.t0 309.017
R104 D.n0 D.t1 231.897
R105 D D.n0 186.203
R106 a_639_47.t0 a_639_47.t1 77.1434
R107 B_N.n0 B_N.t0 408.63
R108 B_N B_N.n0 158.281
R109 B_N.n0 B_N.t1 132.282
C0 D VPWR 0.014752f
C1 A_N VGND 0.017266f
C2 B_N VPWR 0.015634f
C3 C VGND 0.032807f
C4 D VGND 0.051255f
C5 B_N VGND 0.045001f
C6 VPWR X 0.014124f
C7 VPB A_N 0.096861f
C8 VPWR VGND 0.093314f
C9 VPB C 0.054148f
C10 X VGND 0.074636f
C11 VPB D 0.065568f
C12 VPB B_N 0.074525f
C13 VPB VPWR 0.097965f
C14 C D 0.177344f
C15 VPB X 0.003174f
C16 A_N VPWR 0.016669f
C17 VPB VGND 0.01423f
C18 C VPWR 0.015059f
C19 D B_N 0.116523f
C20 A_N X 0.002416f
C21 VGND VNB 0.548354f
C22 X VNB 0.005428f
C23 VPWR VNB 0.445614f
C24 B_N VNB 0.162373f
C25 D VNB 0.110151f
C26 C VNB 0.108512f
C27 A_N VNB 0.199185f
C28 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4bb_4 VNB VPB VGND VPWR A_N C D X B_N
X0 VPWR.t9 a_174_21.t5 X.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_174_21.t0 a_832_21.t2 a_766_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X.t6 a_174_21.t6 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_832_21.t1 A_N.t0 VGND.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1764 ps=1.68 w=0.42 l=0.15
X4 a_766_47.t0 a_27_47.t2 a_652_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1365 ps=1.07 w=0.65 l=0.15
X5 VPWR.t7 a_174_21.t7 X.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X.t4 a_174_21.t8 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR.t1 B_N.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_652_47.t0 C.t0 a_556_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 a_832_21.t0 A_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.31165 ps=2.125 w=0.42 l=0.15
X10 X.t3 a_174_21.t9 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11 X.t2 a_174_21.t10 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_556_47.t0 D.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.11375 ps=1 w=0.65 l=0.15
X13 a_174_21.t4 D.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X14 VPWR.t4 C.t1 a_174_21.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X15 VGND.t3 a_174_21.t11 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t2 a_174_21.t12 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t2 a_832_21.t3 a_174_21.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.31165 pd=2.125 as=0.165 ps=1.33 w=1 l=0.15
X18 a_174_21.t2 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X19 VGND.t0 B_N.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_174_21.n11 a_174_21.n10 661.048
R1 a_174_21.n10 a_174_21.n9 585
R2 a_174_21.n8 a_174_21.t0 306.065
R3 a_174_21.n6 a_174_21.t5 196.013
R4 a_174_21.n4 a_174_21.t6 196.013
R5 a_174_21.n2 a_174_21.t7 196.013
R6 a_174_21.n1 a_174_21.t8 196.013
R7 a_174_21.n3 a_174_21.n0 177.601
R8 a_174_21.n7 a_174_21.n6 158.887
R9 a_174_21.n5 a_174_21.n0 152
R10 a_174_21.n6 a_174_21.t12 149.421
R11 a_174_21.n4 a_174_21.t10 149.421
R12 a_174_21.n2 a_174_21.t11 149.421
R13 a_174_21.n1 a_174_21.t9 149.421
R14 a_174_21.n10 a_174_21.n8 64.7534
R15 a_174_21.n2 a_174_21.n1 57.8405
R16 a_174_21.n6 a_174_21.n5 39.9376
R17 a_174_21.n9 a_174_21.t4 38.4155
R18 a_174_21.t1 a_174_21.n11 34.4755
R19 a_174_21.n11 a_174_21.t2 30.5355
R20 a_174_21.n4 a_174_21.n3 28.9205
R21 a_174_21.n3 a_174_21.n2 28.9205
R22 a_174_21.n9 a_174_21.t3 26.5955
R23 a_174_21.n7 a_174_21.n0 25.6005
R24 a_174_21.n5 a_174_21.n4 17.9034
R25 a_174_21.n8 a_174_21.n7 12.0476
R26 X.n2 X.n0 641.847
R27 X.n2 X.n1 585
R28 X.n5 X.n3 259.166
R29 X.n5 X.n4 206.203
R30 X.n1 X.t5 26.5955
R31 X.n1 X.t4 26.5955
R32 X.n0 X.t7 26.5955
R33 X.n0 X.t6 26.5955
R34 X.n3 X.t0 24.9236
R35 X.n3 X.t2 24.9236
R36 X.n4 X.t1 24.9236
R37 X.n4 X.t3 24.9236
R38 X X.n2 8.45764
R39 X X.n5 1.37193
R40 VPWR.n28 VPWR.n1 599.74
R41 VPWR.n26 VPWR.n3 599.74
R42 VPWR.n5 VPWR.n4 599.74
R43 VPWR.n20 VPWR.n7 599.74
R44 VPWR.n14 VPWR.n13 585
R45 VPWR.n12 VPWR.n10 585
R46 VPWR.n11 VPWR.n9 585
R47 VPWR.n12 VPWR.n11 159.476
R48 VPWR.n13 VPWR.n12 159.476
R49 VPWR.n11 VPWR.t0 107.882
R50 VPWR.n13 VPWR.t2 65.4795
R51 VPWR.n1 VPWR.t1 63.3219
R52 VPWR.n1 VPWR.t6 55.1136
R53 VPWR.n7 VPWR.t4 46.2955
R54 VPWR.n4 VPWR.t5 42.3555
R55 VPWR.n7 VPWR.t3 36.4455
R56 VPWR.n19 VPWR.n8 34.1156
R57 VPWR.n21 VPWR.n5 30.8711
R58 VPWR.n3 VPWR.t8 26.5955
R59 VPWR.n3 VPWR.t7 26.5955
R60 VPWR.n4 VPWR.t9 26.5955
R61 VPWR.n21 VPWR.n20 25.6005
R62 VPWR.n26 VPWR.n25 24.8476
R63 VPWR.n28 VPWR.n27 22.9652
R64 VPWR.n27 VPWR.n26 19.577
R65 VPWR.n20 VPWR.n19 18.824
R66 VPWR.n25 VPWR.n5 13.5534
R67 VPWR.n16 VPWR.n9 9.64031
R68 VPWR.n16 VPWR.n15 9.3005
R69 VPWR.n17 VPWR.n8 9.3005
R70 VPWR.n19 VPWR.n18 9.3005
R71 VPWR.n20 VPWR.n6 9.3005
R72 VPWR.n22 VPWR.n21 9.3005
R73 VPWR.n23 VPWR.n5 9.3005
R74 VPWR.n25 VPWR.n24 9.3005
R75 VPWR.n26 VPWR.n2 9.3005
R76 VPWR.n27 VPWR.n0 9.3005
R77 VPWR.n10 VPWR.n9 7.91323
R78 VPWR.n29 VPWR.n28 7.12063
R79 VPWR.n15 VPWR.n14 7.09868
R80 VPWR.n14 VPWR.n8 3.60777
R81 VPWR.n15 VPWR.n10 0.815045
R82 VPWR.n29 VPWR.n0 0.148519
R83 VPWR.n17 VPWR.n16 0.120292
R84 VPWR.n18 VPWR.n17 0.120292
R85 VPWR.n18 VPWR.n6 0.120292
R86 VPWR.n22 VPWR.n6 0.120292
R87 VPWR.n23 VPWR.n22 0.120292
R88 VPWR.n24 VPWR.n23 0.120292
R89 VPWR.n24 VPWR.n2 0.120292
R90 VPWR.n2 VPWR.n0 0.120292
R91 VPWR VPWR.n29 0.11354
R92 VPB.t2 VPB.t0 754.673
R93 VPB.t4 VPB.t3 337.384
R94 VPB.t9 VPB.t5 295.95
R95 VPB.t3 VPB.t2 284.113
R96 VPB.t5 VPB.t4 284.113
R97 VPB.t1 VPB.t6 281.154
R98 VPB.t8 VPB.t9 248.599
R99 VPB.t7 VPB.t8 248.599
R100 VPB.t6 VPB.t7 248.599
R101 VPB VPB.t1 189.409
R102 a_832_21.t0 a_832_21.n1 772.933
R103 a_832_21.n1 a_832_21.t1 318.067
R104 a_832_21.n1 a_832_21.n0 268.849
R105 a_832_21.n0 a_832_21.t3 212.081
R106 a_832_21.n0 a_832_21.t2 139.78
R107 a_766_47.t0 a_766_47.t1 60.9236
R108 VNB.t9 VNB.t4 3631.07
R109 VNB.t1 VNB.t3 1623.3
R110 VNB.t5 VNB.t2 1423.95
R111 VNB.t3 VNB.t9 1366.99
R112 VNB.t2 VNB.t1 1366.99
R113 VNB.t0 VNB.t8 1352.75
R114 VNB.t7 VNB.t5 1196.12
R115 VNB.t6 VNB.t7 1196.12
R116 VNB.t8 VNB.t6 1196.12
R117 VNB VNB.t0 911.327
R118 A_N.n0 A_N.t1 334.723
R119 A_N.n0 A_N.t0 206.19
R120 A_N.n1 A_N.n0 152
R121 A_N.n1 A_N 10.1338
R122 A_N A_N.n1 1.95606
R123 VGND.n5 VGND.t6 290.055
R124 VGND.n8 VGND.n2 199.934
R125 VGND.n11 VGND.n10 199.739
R126 VGND.n4 VGND.n3 198.964
R127 VGND.n10 VGND.t0 54.2862
R128 VGND.n3 VGND.t1 36.0005
R129 VGND.n3 VGND.t2 28.6159
R130 VGND.n10 VGND.t5 25.9346
R131 VGND.n2 VGND.t4 24.9236
R132 VGND.n2 VGND.t3 24.9236
R133 VGND.n8 VGND.n1 24.8476
R134 VGND.n9 VGND.n8 19.577
R135 VGND.n11 VGND.n9 18.824
R136 VGND.n4 VGND.n1 15.0593
R137 VGND.n6 VGND.n1 9.3005
R138 VGND.n8 VGND.n7 9.3005
R139 VGND.n9 VGND.n0 9.3005
R140 VGND.n5 VGND.n4 7.40753
R141 VGND.n12 VGND.n11 7.32436
R142 VGND.n6 VGND.n5 0.150738
R143 VGND.n12 VGND.n0 0.145929
R144 VGND.n7 VGND.n6 0.120292
R145 VGND.n7 VGND.n0 0.120292
R146 VGND VGND.n12 0.116164
R147 a_27_47.t0 a_27_47.n1 663.091
R148 a_27_47.n1 a_27_47.n0 546.542
R149 a_27_47.n1 a_27_47.t1 333.159
R150 a_27_47.n0 a_27_47.t3 241.536
R151 a_27_47.n0 a_27_47.t2 169.237
R152 a_652_47.t0 a_652_47.t1 77.539
R153 B_N.n0 B_N.t0 334.723
R154 B_N.n0 B_N.t1 206.19
R155 B_N.n1 B_N.n0 152
R156 B_N.n1 B_N 10.4234
R157 B_N B_N.n1 2.01193
R158 C.n0 C.t1 234.173
R159 C.n0 C.t0 161.873
R160 C C.n0 154.387
R161 a_556_47.t0 a_556_47.t1 60.9236
R162 D.n0 D.t1 241.536
R163 D.n0 D.t0 169.237
R164 D D.n0 157.625
C0 C VPWR 0.017924f
C1 D X 4.06e-19
C2 B_N VGND 0.040939f
C3 A_N VPWR 0.018476f
C4 D VGND 0.015807f
C5 A_N X 2.34e-19
C6 C VGND 0.013613f
C7 A_N VGND 0.018493f
C8 VPWR X 0.029711f
C9 VPB B_N 0.090754f
C10 VPWR VGND 0.124793f
C11 VPB D 0.028164f
C12 X VGND 0.183126f
C13 VPB C 0.033047f
C14 B_N C 3.88e-20
C15 VPB A_N 0.101357f
C16 VPB VPWR 0.12201f
C17 D C 0.083393f
C18 B_N A_N 0.002674f
C19 B_N VPWR 0.01984f
C20 VPB X 0.003626f
C21 D VPWR 0.016448f
C22 C A_N 7.38e-20
C23 VPB VGND 0.014132f
C24 B_N X 0.07454f
C25 VGND VNB 0.677453f
C26 X VNB 0.012672f
C27 VPWR VNB 0.560869f
C28 A_N VNB 0.18985f
C29 C VNB 0.103017f
C30 D VNB 0.091161f
C31 B_N VNB 0.162377f
C32 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR.t1 A.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X.t1 a_27_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X.t0 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
R0 A.n0 A.t0 260.322
R1 A.n0 A.t1 175.169
R2 A A.n0 156.325
R3 a_27_47.t0 a_27_47.n1 405.735
R4 a_27_47.n1 a_27_47.t1 294.611
R5 a_27_47.n0 a_27_47.t3 254.389
R6 a_27_47.n0 a_27_47.t2 211.01
R7 a_27_47.n1 a_27_47.n0 152
R8 VPWR VPWR.n0 327.954
R9 VPWR.n0 VPWR.t0 36.1587
R10 VPWR.n0 VPWR.t1 36.1587
R11 VPB.t1 VPB.t0 260.437
R12 VPB VPB.t1 192.369
R13 VGND VGND.n0 214.889
R14 VGND.n0 VGND.t0 33.462
R15 VGND.n0 VGND.t1 33.462
R16 X.n1 X.t0 368.521
R17 X.n0 X.t1 216.155
R18 X X.n0 78.8791
R19 X.n1 X 10.5563
R20 X X.n1 5.48477
R21 X.n0 X 5.16973
R22 VNB.t1 VNB.t0 1253.07
R23 VNB VNB.t1 897.087
C0 VPB A 0.052393f
C1 VPB VPWR 0.035491f
C2 A VPWR 0.021545f
C3 VPB X 0.012762f
C4 A X 8.48e-19
C5 VPB VGND 0.00505f
C6 A VGND 0.018425f
C7 VPWR X 0.089678f
C8 VPWR VGND 0.028968f
C9 X VGND 0.054627f
C10 VGND VNB 0.207322f
C11 X VNB 0.094114f
C12 VPWR VNB 0.175402f
C13 A VNB 0.164055f
C14 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR.t1 a_27_47.t2 X.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t2 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR.t2 A.t0 a_27_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X.t0 a_27_47.t4 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND.t1 a_27_47.t5 X.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t0 A.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.t1 a_27_47.n2 447.445
R1 a_27_47.n2 a_27_47.t0 301.502
R2 a_27_47.n0 a_27_47.t2 212.081
R3 a_27_47.n1 a_27_47.t3 212.081
R4 a_27_47.n2 a_27_47.n1 160.034
R5 a_27_47.n0 a_27_47.t5 139.78
R6 a_27_47.n1 a_27_47.t4 139.78
R7 a_27_47.n1 a_27_47.n0 61.346
R8 X.n0 X 589.769
R9 X.n1 X.n0 585
R10 X.n3 X.n2 185
R11 X X.n3 81.3181
R12 X.n0 X.t3 26.5955
R13 X.n0 X.t2 26.5955
R14 X.n2 X.t1 24.9236
R15 X.n2 X.t0 24.9236
R16 X.n1 X 15.5613
R17 X.n3 X 5.27109
R18 X X.n1 1.50638
R19 VPWR.n1 VPWR.n0 315.904
R20 VPWR.n1 VPWR.t1 257.788
R21 VPWR.n0 VPWR.t2 55.4067
R22 VPWR.n0 VPWR.t0 34.0906
R23 VPWR VPWR.n1 12.4075
R24 VPB.t2 VPB.t0 281.154
R25 VPB.t0 VPB.t1 248.599
R26 VPB VPB.t2 192.369
R27 A.n0 A.t0 276.464
R28 A.n0 A.t1 196.131
R29 A A.n0 156.325
R30 VGND.n1 VGND.n0 203.591
R31 VGND.n1 VGND.t1 162.987
R32 VGND.n0 VGND.t0 51.4291
R33 VGND.n0 VGND.t2 28.7917
R34 VGND VGND.n1 12.4075
R35 VNB.t0 VNB.t2 1352.75
R36 VNB.t2 VNB.t1 1196.12
R37 VNB VNB.t0 925.567
C0 A VGND 0.019887f
C1 VPWR X 0.168994f
C2 VPWR VGND 0.051753f
C3 X VGND 0.111264f
C4 VPB A 0.069727f
C5 VPB VPWR 0.05279f
C6 A VPWR 0.022108f
C7 VPB X 0.004428f
C8 A X 0.003062f
C9 VPB VGND 0.006417f
C10 VGND VNB 0.284185f
C11 X VNB 0.021498f
C12 VPWR VNB 0.249629f
C13 A VNB 0.187471f
C14 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR.t4 a_27_47.t2 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t2 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t2 a_27_47.t4 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X.t0 a_27_47.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X.t7 a_27_47.t6 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X.t6 a_27_47.t7 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND.t2 a_27_47.t8 X.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t1 a_27_47.t9 X.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.t0 a_27_47.n5 271.759
R1 a_27_47.n5 a_27_47.t1 270.911
R2 a_27_47.n0 a_27_47.t2 221.72
R3 a_27_47.n1 a_27_47.t3 221.72
R4 a_27_47.n2 a_27_47.t4 221.72
R5 a_27_47.n3 a_27_47.t5 221.72
R6 a_27_47.n5 a_27_47.n4 170.825
R7 a_27_47.n0 a_27_47.t9 149.421
R8 a_27_47.n1 a_27_47.t7 149.421
R9 a_27_47.n2 a_27_47.t8 149.421
R10 a_27_47.n3 a_27_47.t6 149.421
R11 a_27_47.n1 a_27_47.n0 74.9783
R12 a_27_47.n2 a_27_47.n1 74.9783
R13 a_27_47.n4 a_27_47.n2 59.8042
R14 a_27_47.n4 a_27_47.n3 15.1746
R15 X.n3 X.n1 344.096
R16 X.n3 X.n2 313.916
R17 X.n4 X.n0 230.554
R18 X X.n5 198.952
R19 X.n1 X.t1 26.5955
R20 X.n1 X.t0 26.5955
R21 X.n2 X.t3 26.5955
R22 X.n2 X.t2 26.5955
R23 X.n0 X.t5 24.9236
R24 X.n0 X.t7 24.9236
R25 X.n5 X.t4 24.9236
R26 X.n5 X.t6 24.9236
R27 X.n4 X 7.3702
R28 X X.n3 2.19848
R29 X X.n4 1.42272
R30 VPWR.n1 VPWR.n0 317.231
R31 VPWR.n4 VPWR.n3 310.502
R32 VPWR.n2 VPWR.t4 249.126
R33 VPWR.n0 VPWR.t1 26.5955
R34 VPWR.n0 VPWR.t0 26.5955
R35 VPWR.n3 VPWR.t3 26.5955
R36 VPWR.n3 VPWR.t2 26.5955
R37 VPWR.n5 VPWR.n1 23.7181
R38 VPWR.n5 VPWR.n4 15.4358
R39 VPWR VPWR.n7 11.6277
R40 VPWR.n6 VPWR.n5 9.3005
R41 VPWR.n4 VPWR.n2 6.67472
R42 VPWR.n7 VPWR.n1 5.5329
R43 VPWR.n7 VPWR.n6 2.0169
R44 VPWR.n6 VPWR.n2 0.811095
R45 VPB.t3 VPB.t4 248.599
R46 VPB.t2 VPB.t3 248.599
R47 VPB.t1 VPB.t2 248.599
R48 VPB.t0 VPB.t1 248.599
R49 VPB VPB.t0 189.409
R50 VGND.n1 VGND.n0 206.333
R51 VGND.n4 VGND.n3 200.516
R52 VGND.n2 VGND.t1 155.376
R53 VGND.n5 VGND.n1 28.9887
R54 VGND.n0 VGND.t4 24.9236
R55 VGND.n0 VGND.t0 24.9236
R56 VGND.n3 VGND.t3 24.9236
R57 VGND.n3 VGND.t2 24.9236
R58 VGND.n5 VGND.n4 15.4358
R59 VGND VGND.n7 11.1362
R60 VGND.n6 VGND.n5 9.3005
R61 VGND.n4 VGND.n2 6.67472
R62 VGND.n7 VGND.n1 5.0477
R63 VGND.n7 VGND.n6 2.26105
R64 VGND.n6 VGND.n2 0.811095
R65 VNB.t3 VNB.t1 1196.12
R66 VNB.t2 VNB.t3 1196.12
R67 VNB.t4 VNB.t2 1196.12
R68 VNB.t0 VNB.t4 1196.12
R69 VNB VNB.t0 911.327
R70 A.n0 A.t0 235.763
R71 A.n0 A.t1 163.464
R72 A A.n0 160.268
C0 VPB A 0.03609f
C1 VPB VPWR 0.071068f
C2 A VPWR 0.016006f
C3 VPB X 0.008994f
C4 A X 4.66e-19
C5 VPB VGND 0.007955f
C6 A VGND 0.019369f
C7 VPWR X 0.332544f
C8 VPWR VGND 0.072027f
C9 X VGND 0.229885f
C10 VGND VNB 0.37777f
C11 X VNB 0.039034f
C12 VPWR VNB 0.325078f
C13 A VNB 0.139971f
C14 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VPB VNB
X0 VPWR.t5 a_161_47.t4 X.t11 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47.t0 A.t0 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X.t10 a_161_47.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t3 a_161_47.t6 X.t9 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t6 A.t1 a_161_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X.t8 a_161_47.t7 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t5 a_161_47.t8 X.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t4 a_161_47.t9 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t1 a_161_47.t10 X.t7 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t6 a_161_47.t11 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X.t3 a_161_47.t12 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X.t2 a_161_47.t13 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t1 a_161_47.t14 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR.t6 A.t2 a_161_47.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t0 a_161_47.t15 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_161_47.t3 A.t3 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R0 a_161_47.n9 a_161_47.n8 247.799
R1 a_161_47.n1 a_161_47.t4 221.72
R2 a_161_47.n2 a_161_47.t5 221.72
R3 a_161_47.n3 a_161_47.t6 221.72
R4 a_161_47.n4 a_161_47.t7 221.72
R5 a_161_47.n5 a_161_47.t10 221.72
R6 a_161_47.n6 a_161_47.t11 221.72
R7 a_161_47.n8 a_161_47.n7 168.565
R8 a_161_47.n1 a_161_47.t15 149.421
R9 a_161_47.n2 a_161_47.t14 149.421
R10 a_161_47.n3 a_161_47.t9 149.421
R11 a_161_47.n4 a_161_47.t13 149.421
R12 a_161_47.n5 a_161_47.t8 149.421
R13 a_161_47.n6 a_161_47.t12 149.421
R14 a_161_47.n8 a_161_47.n0 137.588
R15 a_161_47.n2 a_161_47.n1 74.9783
R16 a_161_47.n3 a_161_47.n2 74.9783
R17 a_161_47.n4 a_161_47.n3 74.9783
R18 a_161_47.n5 a_161_47.n4 74.9783
R19 a_161_47.n7 a_161_47.n5 58.9116
R20 a_161_47.t2 a_161_47.n9 26.5955
R21 a_161_47.n9 a_161_47.t3 26.5955
R22 a_161_47.n0 a_161_47.t1 24.9236
R23 a_161_47.n0 a_161_47.t0 24.9236
R24 a_161_47.n7 a_161_47.n6 16.0672
R25 X X.n0 344.096
R26 X.n6 X.n4 311.717
R27 X.n7 X.n2 311.717
R28 X X.n1 230.554
R29 X.n6 X.n5 198.177
R30 X.n7 X.n3 198.177
R31 X.n0 X.t7 26.5955
R32 X.n0 X.t6 26.5955
R33 X.n4 X.t11 26.5955
R34 X.n4 X.t10 26.5955
R35 X.n2 X.t9 26.5955
R36 X.n2 X.t8 26.5955
R37 X.n1 X.t5 24.9236
R38 X.n1 X.t3 24.9236
R39 X.n5 X.t0 24.9236
R40 X.n5 X.t1 24.9236
R41 X.n3 X.t4 24.9236
R42 X.n3 X.t2 24.9236
R43 X.n7 X.n6 12.2187
R44 X X.n7 5.96414
R45 VPWR.n13 VPWR.n12 317.233
R46 VPWR.n6 VPWR.n5 310.502
R47 VPWR.n3 VPWR.n2 310.502
R48 VPWR.n0 VPWR.t7 257.474
R49 VPWR.n4 VPWR.t5 249.96
R50 VPWR.n15 VPWR.n14 34.6358
R51 VPWR.n11 VPWR.n3 32.0005
R52 VPWR.n2 VPWR.t2 26.5955
R53 VPWR.n2 VPWR.t1 26.5955
R54 VPWR.n5 VPWR.t4 26.5955
R55 VPWR.n5 VPWR.t3 26.5955
R56 VPWR.n12 VPWR.t0 26.5955
R57 VPWR.n12 VPWR.t6 26.5955
R58 VPWR.n7 VPWR.n6 25.977
R59 VPWR.n17 VPWR.n0 21.8358
R60 VPWR.n15 VPWR.n0 12.8005
R61 VPWR.n7 VPWR.n3 12.424
R62 VPWR.n17 VPWR.n16 9.42029
R63 VPWR.n14 VPWR.n13 9.41227
R64 VPWR.n8 VPWR.n7 9.3005
R65 VPWR.n9 VPWR.n3 9.3005
R66 VPWR.n11 VPWR.n10 9.3005
R67 VPWR.n14 VPWR.n1 9.3005
R68 VPWR.n16 VPWR.n15 9.3005
R69 VPWR.n13 VPWR.n11 7.15344
R70 VPWR.n6 VPWR.n4 6.18988
R71 VPWR VPWR.n17 6.02403
R72 VPWR.n8 VPWR.n4 0.755914
R73 VPWR.n9 VPWR.n8 0.120292
R74 VPWR.n10 VPWR.n9 0.120292
R75 VPWR.n10 VPWR.n1 0.120292
R76 VPWR.n16 VPWR.n1 0.120292
R77 VPB VPB.t7 343.303
R78 VPB.t4 VPB.t5 248.599
R79 VPB.t3 VPB.t4 248.599
R80 VPB.t2 VPB.t3 248.599
R81 VPB.t1 VPB.t2 248.599
R82 VPB.t0 VPB.t1 248.599
R83 VPB.t6 VPB.t0 248.599
R84 VPB.t7 VPB.t6 248.599
R85 A.n0 A.t2 221.72
R86 A.n2 A.t3 221.72
R87 A.n3 A.n2 185.026
R88 A.n1 A 158.934
R89 A.n0 A.t1 149.421
R90 A.n2 A.t0 149.421
R91 A.n2 A.n1 51.7709
R92 A.n1 A.n0 23.2079
R93 A.n3 A 18.4005
R94 A A.n3 8.26717
R95 VGND.n0 VGND.t7 282.565
R96 VGND.n13 VGND.n2 208.719
R97 VGND.n7 VGND.n6 200.516
R98 VGND.n4 VGND.n3 200.516
R99 VGND.n5 VGND.t0 156.209
R100 VGND.n15 VGND.n14 34.6358
R101 VGND.n12 VGND.n4 32.0005
R102 VGND.n8 VGND.n7 25.977
R103 VGND.n3 VGND.t2 24.9236
R104 VGND.n3 VGND.t5 24.9236
R105 VGND.n6 VGND.t1 24.9236
R106 VGND.n6 VGND.t4 24.9236
R107 VGND.n2 VGND.t3 24.9236
R108 VGND.n2 VGND.t6 24.9236
R109 VGND.n17 VGND.n0 21.8358
R110 VGND.n13 VGND.n12 18.824
R111 VGND.n14 VGND.n13 15.8123
R112 VGND.n15 VGND.n0 12.8005
R113 VGND.n8 VGND.n4 12.424
R114 VGND.n17 VGND.n16 9.42029
R115 VGND.n9 VGND.n8 9.3005
R116 VGND.n10 VGND.n4 9.3005
R117 VGND.n16 VGND.n15 9.3005
R118 VGND.n14 VGND.n1 9.3005
R119 VGND.n12 VGND.n11 9.3005
R120 VGND.n7 VGND.n5 6.18988
R121 VGND VGND.n17 6.02403
R122 VGND.n9 VGND.n5 0.755914
R123 VGND.n10 VGND.n9 0.120292
R124 VGND.n11 VGND.n10 0.120292
R125 VGND.n11 VGND.n1 0.120292
R126 VGND.n16 VGND.n1 0.120292
R127 VNB VNB.t7 1651.78
R128 VNB.t1 VNB.t0 1196.12
R129 VNB.t4 VNB.t1 1196.12
R130 VNB.t2 VNB.t4 1196.12
R131 VNB.t5 VNB.t2 1196.12
R132 VNB.t3 VNB.t5 1196.12
R133 VNB.t6 VNB.t3 1196.12
R134 VNB.t7 VNB.t6 1196.12
C0 A X 3.93e-19
C1 VPB VGND 0.010018f
C2 A VGND 0.041682f
C3 VPWR X 0.507648f
C4 VPWR VGND 0.101848f
C5 X VGND 0.363808f
C6 VPB A 0.075647f
C7 VPB VPWR 0.101686f
C8 A VPWR 0.050548f
C9 VPB X 0.012957f
C10 VGND VNB 0.532636f
C11 X VNB 0.050616f
C12 VPWR VNB 0.479991f
C13 A VNB 0.239842f
C14 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_8 VPB VNB VGND VPWR A X
X0 X.t7 a_27_47.t6 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X.t6 a_27_47.t7 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X.t5 a_27_47.t8 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t9 a_27_47.t9 X.t15 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X.t14 a_27_47.t10 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t5 a_27_47.t11 X.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t7 a_27_47.t12 X.t13 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47.t1 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t12 a_27_47.t13 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X.t3 a_27_47.t14 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t5 a_27_47.t15 X.t11 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X.t10 a_27_47.t16 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t9 A.t3 a_27_47.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t3 a_27_47.t17 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t3 a_27_47.t18 X.t9 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t2 a_27_47.t19 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t1 a_27_47.t20 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X.t8 a_27_47.t21 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t10 A.t4 a_27_47.t4 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND.t10 A.t5 a_27_47.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n22 a_27_47.t5 286.348
R1 a_27_47.n24 a_27_47.t4 271.051
R2 a_27_47.n4 a_27_47.t12 221.72
R3 a_27_47.n5 a_27_47.t13 221.72
R4 a_27_47.n3 a_27_47.t15 221.72
R5 a_27_47.n9 a_27_47.t16 221.72
R6 a_27_47.n11 a_27_47.t18 221.72
R7 a_27_47.n1 a_27_47.t21 221.72
R8 a_27_47.n17 a_27_47.t9 221.72
R9 a_27_47.n18 a_27_47.t10 221.72
R10 a_27_47.n25 a_27_47.n24 206.055
R11 a_27_47.n22 a_27_47.n21 198.177
R12 a_27_47.n7 a_27_47.n6 177.601
R13 a_27_47.n20 a_27_47.n19 152
R14 a_27_47.n16 a_27_47.n0 152
R15 a_27_47.n15 a_27_47.n14 152
R16 a_27_47.n13 a_27_47.n12 152
R17 a_27_47.n10 a_27_47.n2 152
R18 a_27_47.n8 a_27_47.n7 152
R19 a_27_47.n4 a_27_47.t11 149.421
R20 a_27_47.n5 a_27_47.t8 149.421
R21 a_27_47.n3 a_27_47.t20 149.421
R22 a_27_47.n9 a_27_47.t7 149.421
R23 a_27_47.n11 a_27_47.t19 149.421
R24 a_27_47.n1 a_27_47.t6 149.421
R25 a_27_47.n17 a_27_47.t17 149.421
R26 a_27_47.n18 a_27_47.t14 149.421
R27 a_27_47.n5 a_27_47.n4 74.9783
R28 a_27_47.n6 a_27_47.n5 66.0523
R29 a_27_47.n16 a_27_47.n15 60.6968
R30 a_27_47.n19 a_27_47.n17 55.3412
R31 a_27_47.n8 a_27_47.n3 51.7709
R32 a_27_47.n12 a_27_47.n1 51.7709
R33 a_27_47.n23 a_27_47.n22 48.9632
R34 a_27_47.n24 a_27_47.n23 38.7339
R35 a_27_47.n10 a_27_47.n9 37.4894
R36 a_27_47.n11 a_27_47.n10 37.4894
R37 a_27_47.t0 a_27_47.n25 26.5955
R38 a_27_47.n25 a_27_47.t1 26.5955
R39 a_27_47.n7 a_27_47.n2 25.6005
R40 a_27_47.n13 a_27_47.n2 25.6005
R41 a_27_47.n14 a_27_47.n13 25.6005
R42 a_27_47.n14 a_27_47.n0 25.6005
R43 a_27_47.n20 a_27_47.n0 25.6005
R44 a_27_47.n21 a_27_47.t3 24.9236
R45 a_27_47.n21 a_27_47.t2 24.9236
R46 a_27_47.n9 a_27_47.n8 23.2079
R47 a_27_47.n12 a_27_47.n11 23.2079
R48 a_27_47.n19 a_27_47.n18 19.6375
R49 a_27_47.n23 a_27_47.n20 18.4476
R50 a_27_47.n6 a_27_47.n3 8.92643
R51 a_27_47.n15 a_27_47.n1 8.92643
R52 a_27_47.n17 a_27_47.n16 5.35606
R53 VGND.n5 VGND.n4 200.516
R54 VGND.n10 VGND.n9 200.516
R55 VGND.n13 VGND.n12 200.516
R56 VGND.n18 VGND.n2 200.516
R57 VGND.n21 VGND.n20 200.516
R58 VGND.n6 VGND.t5 155.156
R59 VGND.n14 VGND.n11 34.6358
R60 VGND.n8 VGND.n5 32.0005
R61 VGND.n18 VGND.n1 28.9887
R62 VGND.n4 VGND.t6 24.9236
R63 VGND.n4 VGND.t1 24.9236
R64 VGND.n9 VGND.t7 24.9236
R65 VGND.n9 VGND.t2 24.9236
R66 VGND.n12 VGND.t8 24.9236
R67 VGND.n12 VGND.t3 24.9236
R68 VGND.n2 VGND.t4 24.9236
R69 VGND.n2 VGND.t9 24.9236
R70 VGND.n20 VGND.t0 24.9236
R71 VGND.n20 VGND.t10 24.9236
R72 VGND.n21 VGND.n19 22.9652
R73 VGND.n19 VGND.n18 15.4358
R74 VGND.n13 VGND.n1 9.41227
R75 VGND.n19 VGND.n0 9.3005
R76 VGND.n18 VGND.n17 9.3005
R77 VGND.n16 VGND.n1 9.3005
R78 VGND.n15 VGND.n14 9.3005
R79 VGND.n11 VGND.n3 9.3005
R80 VGND.n8 VGND.n7 9.3005
R81 VGND.n22 VGND.n21 7.12063
R82 VGND.n10 VGND.n8 6.4005
R83 VGND.n6 VGND.n5 5.79315
R84 VGND.n11 VGND.n10 3.38874
R85 VGND.n7 VGND.n6 0.656787
R86 VGND.n14 VGND.n13 0.376971
R87 VGND.n22 VGND.n0 0.148519
R88 VGND.n7 VGND.n3 0.120292
R89 VGND.n15 VGND.n3 0.120292
R90 VGND.n16 VGND.n15 0.120292
R91 VGND.n17 VGND.n16 0.120292
R92 VGND.n17 VGND.n0 0.120292
R93 VGND VGND.n22 0.11354
R94 X.n8 X.n7 374.966
R95 X.n11 X.n10 315.985
R96 X.n9 X.n5 311.717
R97 X.n8 X.n6 311.717
R98 X.n3 X.n2 261.425
R99 X X.n13 199.683
R100 X.n3 X.n1 198.177
R101 X.n4 X.n0 198.177
R102 X.n4 X.n3 63.2476
R103 X.n9 X.n8 63.2476
R104 X.n12 X.n4 50.4476
R105 X.n11 X.n9 50.4476
R106 X.n5 X.t11 26.5955
R107 X.n5 X.t10 26.5955
R108 X.n6 X.t9 26.5955
R109 X.n6 X.t8 26.5955
R110 X.n7 X.t15 26.5955
R111 X.n7 X.t14 26.5955
R112 X.n10 X.t13 26.5955
R113 X.n10 X.t12 26.5955
R114 X.n2 X.t2 24.9236
R115 X.n2 X.t3 24.9236
R116 X.n1 X.t1 24.9236
R117 X.n1 X.t7 24.9236
R118 X.n0 X.t0 24.9236
R119 X.n0 X.t6 24.9236
R120 X.n13 X.t4 24.9236
R121 X.n13 X.t5 24.9236
R122 X.n12 X 14.3064
R123 X X.n11 4.26717
R124 X X.n12 2.76128
R125 VNB.t6 VNB.t5 1196.12
R126 VNB.t1 VNB.t6 1196.12
R127 VNB.t7 VNB.t1 1196.12
R128 VNB.t2 VNB.t7 1196.12
R129 VNB.t8 VNB.t2 1196.12
R130 VNB.t3 VNB.t8 1196.12
R131 VNB.t4 VNB.t3 1196.12
R132 VNB.t9 VNB.t4 1196.12
R133 VNB.t0 VNB.t9 1196.12
R134 VNB.t10 VNB.t0 1196.12
R135 VNB VNB.t10 911.327
R136 VPWR.n3 VPWR.n2 320.976
R137 VPWR.n24 VPWR.n1 320.976
R138 VPWR.n17 VPWR.n5 310.502
R139 VPWR.n11 VPWR.n10 310.502
R140 VPWR.n9 VPWR.n8 310.502
R141 VPWR.n7 VPWR.t7 248.906
R142 VPWR.n25 VPWR.n24 43.1829
R143 VPWR.n19 VPWR.n18 34.6358
R144 VPWR.n23 VPWR.n22 34.6358
R145 VPWR.n16 VPWR.n6 34.6358
R146 VPWR.n12 VPWR.n9 32.0005
R147 VPWR.n22 VPWR.n3 27.8593
R148 VPWR.n1 VPWR.t1 26.5955
R149 VPWR.n1 VPWR.t10 26.5955
R150 VPWR.n2 VPWR.t8 26.5955
R151 VPWR.n2 VPWR.t0 26.5955
R152 VPWR.n5 VPWR.t2 26.5955
R153 VPWR.n5 VPWR.t9 26.5955
R154 VPWR.n10 VPWR.t4 26.5955
R155 VPWR.n10 VPWR.t3 26.5955
R156 VPWR.n8 VPWR.t6 26.5955
R157 VPWR.n8 VPWR.t5 26.5955
R158 VPWR.n18 VPWR.n17 9.41227
R159 VPWR.n13 VPWR.n12 9.3005
R160 VPWR.n14 VPWR.n6 9.3005
R161 VPWR.n16 VPWR.n15 9.3005
R162 VPWR.n18 VPWR.n4 9.3005
R163 VPWR.n20 VPWR.n19 9.3005
R164 VPWR.n22 VPWR.n21 9.3005
R165 VPWR.n23 VPWR.n0 9.3005
R166 VPWR.n19 VPWR.n3 6.77697
R167 VPWR.n12 VPWR.n11 6.4005
R168 VPWR.n9 VPWR.n7 5.7932
R169 VPWR.n11 VPWR.n6 3.38874
R170 VPWR.n24 VPWR.n23 0.753441
R171 VPWR.n13 VPWR.n7 0.656729
R172 VPWR.n17 VPWR.n16 0.376971
R173 VPWR.n14 VPWR.n13 0.120292
R174 VPWR.n15 VPWR.n14 0.120292
R175 VPWR.n15 VPWR.n4 0.120292
R176 VPWR.n20 VPWR.n4 0.120292
R177 VPWR.n21 VPWR.n20 0.120292
R178 VPWR.n21 VPWR.n0 0.120292
R179 VPWR.n25 VPWR.n0 0.120292
R180 VPWR VPWR.n25 0.0213333
R181 VPB.t6 VPB.t7 248.599
R182 VPB.t5 VPB.t6 248.599
R183 VPB.t4 VPB.t5 248.599
R184 VPB.t3 VPB.t4 248.599
R185 VPB.t2 VPB.t3 248.599
R186 VPB.t9 VPB.t2 248.599
R187 VPB.t8 VPB.t9 248.599
R188 VPB.t0 VPB.t8 248.599
R189 VPB.t1 VPB.t0 248.599
R190 VPB.t10 VPB.t1 248.599
R191 VPB VPB.t10 189.409
R192 A.n6 A.t4 235.763
R193 A.n1 A.t0 221.72
R194 A.n0 A.t1 221.72
R195 A.n6 A.t5 163.464
R196 A.n3 A.n2 152
R197 A.n5 A.n4 152
R198 A.n7 A.n6 152
R199 A.n1 A.t3 149.421
R200 A.n0 A.t2 149.421
R201 A.n2 A.n1 58.019
R202 A.n5 A.n0 43.7375
R203 A.n4 A.n3 21.7605
R204 A.n7 A 19.5205
R205 A.n6 A.n5 17.8524
R206 A.n2 A.n0 16.9598
R207 A A.n7 9.9205
R208 A.n3 A 5.4405
R209 A.n4 A 2.2405
C0 A X 6.16e-19
C1 VPB VGND 0.014158f
C2 A VGND 0.05431f
C3 VPWR X 0.664309f
C4 VPWR VGND 0.130194f
C5 X VGND 0.485646f
C6 VPB A 0.099483f
C7 VPB VPWR 0.129764f
C8 A VPWR 0.049241f
C9 VPB X 0.01638f
C10 VGND VNB 0.654069f
C11 X VNB 0.059666f
C12 VPWR VNB 0.555848f
C13 A VNB 0.321526f
C14 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_12 VPB VNB VGND VPWR A X
X0 VGND.t11 a_109_47.t8 X.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X.t23 a_109_47.t9 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t10 a_109_47.t10 X.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t9 a_109_47.t11 X.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND.t8 a_109_47.t12 X.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X.t22 a_109_47.t13 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t13 A.t0 a_109_47.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t7 a_109_47.t14 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X.t6 a_109_47.t15 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X.t5 a_109_47.t16 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_109_47.t6 A.t1 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR.t9 a_109_47.t17 X.t21 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X.t20 a_109_47.t18 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR.t15 A.t2 a_109_47.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t7 a_109_47.t19 X.t19 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t13 A.t3 a_109_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t14 A.t4 a_109_47.t2 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t4 a_109_47.t20 X.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 X.t18 a_109_47.t21 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t5 a_109_47.t22 X.t17 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_109_47.t3 A.t5 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 X.t3 a_109_47.t23 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 X.t16 a_109_47.t24 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t3 a_109_47.t25 X.t15 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.135 ps=1.27 w=1 l=0.15
X24 X.t2 a_109_47.t26 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 X.t1 a_109_47.t27 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t2 a_109_47.t28 X.t14 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 X.t13 a_109_47.t29 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_109_47.t4 A.t6 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 VPWR.t0 a_109_47.t30 X.t12 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_109_47.t0 A.t7 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND.t0 a_109_47.t31 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_109_47.n27 a_109_47.n26 261.425
R1 a_109_47.n31 a_109_47.n30 244.457
R2 a_109_47.n4 a_109_47.t25 221.72
R3 a_109_47.n5 a_109_47.t29 221.72
R4 a_109_47.n6 a_109_47.t30 221.72
R5 a_109_47.n7 a_109_47.t9 221.72
R6 a_109_47.n8 a_109_47.t17 221.72
R7 a_109_47.n9 a_109_47.t18 221.72
R8 a_109_47.n3 a_109_47.t19 221.72
R9 a_109_47.n13 a_109_47.t21 221.72
R10 a_109_47.n15 a_109_47.t22 221.72
R11 a_109_47.n1 a_109_47.t24 221.72
R12 a_109_47.n21 a_109_47.t28 221.72
R13 a_109_47.n22 a_109_47.t13 221.72
R14 a_109_47.n30 a_109_47.n29 206.056
R15 a_109_47.n27 a_109_47.n25 198.177
R16 a_109_47.n11 a_109_47.n10 177.601
R17 a_109_47.n24 a_109_47.n23 152
R18 a_109_47.n20 a_109_47.n0 152
R19 a_109_47.n19 a_109_47.n18 152
R20 a_109_47.n17 a_109_47.n16 152
R21 a_109_47.n14 a_109_47.n2 152
R22 a_109_47.n12 a_109_47.n11 152
R23 a_109_47.n4 a_109_47.t20 149.421
R24 a_109_47.n5 a_109_47.t15 149.421
R25 a_109_47.n6 a_109_47.t11 149.421
R26 a_109_47.n7 a_109_47.t14 149.421
R27 a_109_47.n8 a_109_47.t31 149.421
R28 a_109_47.n9 a_109_47.t16 149.421
R29 a_109_47.n3 a_109_47.t12 149.421
R30 a_109_47.n13 a_109_47.t27 149.421
R31 a_109_47.n15 a_109_47.t10 149.421
R32 a_109_47.n1 a_109_47.t26 149.421
R33 a_109_47.n21 a_109_47.t8 149.421
R34 a_109_47.n22 a_109_47.t23 149.421
R35 a_109_47.n5 a_109_47.n4 74.9783
R36 a_109_47.n6 a_109_47.n5 74.9783
R37 a_109_47.n7 a_109_47.n6 74.9783
R38 a_109_47.n8 a_109_47.n7 74.9783
R39 a_109_47.n9 a_109_47.n8 74.9783
R40 a_109_47.n10 a_109_47.n9 66.0523
R41 a_109_47.n20 a_109_47.n19 60.6968
R42 a_109_47.n23 a_109_47.n21 55.3412
R43 a_109_47.n12 a_109_47.n3 51.7709
R44 a_109_47.n16 a_109_47.n1 51.7709
R45 a_109_47.n28 a_109_47.n27 48.9632
R46 a_109_47.n30 a_109_47.n28 38.7339
R47 a_109_47.n14 a_109_47.n13 37.4894
R48 a_109_47.n15 a_109_47.n14 37.4894
R49 a_109_47.n29 a_109_47.t5 26.5955
R50 a_109_47.n29 a_109_47.t6 26.5955
R51 a_109_47.n31 a_109_47.t7 26.5955
R52 a_109_47.t4 a_109_47.n31 26.5955
R53 a_109_47.n11 a_109_47.n2 25.6005
R54 a_109_47.n17 a_109_47.n2 25.6005
R55 a_109_47.n18 a_109_47.n17 25.6005
R56 a_109_47.n18 a_109_47.n0 25.6005
R57 a_109_47.n24 a_109_47.n0 25.6005
R58 a_109_47.n26 a_109_47.t1 24.9236
R59 a_109_47.n26 a_109_47.t0 24.9236
R60 a_109_47.n25 a_109_47.t2 24.9236
R61 a_109_47.n25 a_109_47.t3 24.9236
R62 a_109_47.n13 a_109_47.n12 23.2079
R63 a_109_47.n16 a_109_47.n15 23.2079
R64 a_109_47.n23 a_109_47.n22 19.6375
R65 a_109_47.n28 a_109_47.n24 18.4476
R66 a_109_47.n10 a_109_47.n3 8.92643
R67 a_109_47.n19 a_109_47.n1 8.92643
R68 a_109_47.n21 a_109_47.n20 5.35606
R69 X.n3 X.n2 374.966
R70 X.n4 X.n0 311.717
R71 X.n3 X.n1 311.717
R72 X.n16 X.n14 311.717
R73 X.n17 X.n12 311.717
R74 X.n18 X.n10 311.717
R75 X.n8 X.n7 261.425
R76 X.n8 X.n6 198.177
R77 X.n9 X.n5 198.177
R78 X.n16 X.n15 198.177
R79 X.n17 X.n13 198.177
R80 X.n18 X.n11 198.177
R81 X.n4 X.n3 63.2476
R82 X.n9 X.n8 63.2476
R83 X X.n4 50.4476
R84 X X.n9 50.4476
R85 X.n0 X.t19 26.5955
R86 X.n0 X.t18 26.5955
R87 X.n1 X.t17 26.5955
R88 X.n1 X.t16 26.5955
R89 X.n2 X.t14 26.5955
R90 X.n2 X.t22 26.5955
R91 X.n14 X.t15 26.5955
R92 X.n14 X.t13 26.5955
R93 X.n12 X.t12 26.5955
R94 X.n12 X.t23 26.5955
R95 X.n10 X.t21 26.5955
R96 X.n10 X.t20 26.5955
R97 X.n7 X.t11 24.9236
R98 X.n7 X.t3 24.9236
R99 X.n6 X.t10 24.9236
R100 X.n6 X.t2 24.9236
R101 X.n5 X.t8 24.9236
R102 X.n5 X.t1 24.9236
R103 X.n15 X.t4 24.9236
R104 X.n15 X.t6 24.9236
R105 X.n13 X.t9 24.9236
R106 X.n13 X.t7 24.9236
R107 X.n11 X.t0 24.9236
R108 X.n11 X.t5 24.9236
R109 X.n17 X.n16 12.2187
R110 X.n18 X.n17 12.2187
R111 X X.n18 2.47323
R112 VGND.n35 VGND.t12 274.361
R113 VGND.n10 VGND.n9 200.516
R114 VGND.n7 VGND.n6 200.516
R115 VGND.n17 VGND.n16 200.516
R116 VGND.n19 VGND.n18 200.516
R117 VGND.n26 VGND.n25 200.516
R118 VGND.n29 VGND.n28 200.516
R119 VGND.n33 VGND.n2 200.516
R120 VGND.n8 VGND.t4 143.024
R121 VGND.n24 VGND.n4 34.6358
R122 VGND.n29 VGND.n27 32.0005
R123 VGND.n20 VGND.n17 28.9887
R124 VGND.n33 VGND.n1 25.977
R125 VGND.n9 VGND.t6 24.9236
R126 VGND.n9 VGND.t9 24.9236
R127 VGND.n6 VGND.t7 24.9236
R128 VGND.n6 VGND.t0 24.9236
R129 VGND.n16 VGND.t5 24.9236
R130 VGND.n16 VGND.t8 24.9236
R131 VGND.n18 VGND.t1 24.9236
R132 VGND.n18 VGND.t10 24.9236
R133 VGND.n25 VGND.t2 24.9236
R134 VGND.n25 VGND.t11 24.9236
R135 VGND.n28 VGND.t3 24.9236
R136 VGND.n28 VGND.t14 24.9236
R137 VGND.n2 VGND.t15 24.9236
R138 VGND.n2 VGND.t13 24.9236
R139 VGND.n15 VGND.n7 22.9652
R140 VGND.n11 VGND.n7 21.4593
R141 VGND.n35 VGND.n34 19.9534
R142 VGND.n34 VGND.n33 18.4476
R143 VGND.n11 VGND.n10 16.9417
R144 VGND.n17 VGND.n15 15.4358
R145 VGND.n29 VGND.n1 12.424
R146 VGND.n20 VGND.n19 9.41227
R147 VGND VGND.n35 9.38904
R148 VGND.n34 VGND.n0 9.3005
R149 VGND.n33 VGND.n32 9.3005
R150 VGND.n31 VGND.n1 9.3005
R151 VGND.n30 VGND.n29 9.3005
R152 VGND.n27 VGND.n3 9.3005
R153 VGND.n24 VGND.n23 9.3005
R154 VGND.n22 VGND.n4 9.3005
R155 VGND.n21 VGND.n20 9.3005
R156 VGND.n17 VGND.n5 9.3005
R157 VGND.n15 VGND.n14 9.3005
R158 VGND.n13 VGND.n7 9.3005
R159 VGND.n12 VGND.n11 9.3005
R160 VGND.n10 VGND.n8 6.64192
R161 VGND.n27 VGND.n26 6.4005
R162 VGND.n26 VGND.n24 3.38874
R163 VGND.n12 VGND.n8 0.78172
R164 VGND.n19 VGND.n4 0.376971
R165 VGND.n13 VGND.n12 0.120292
R166 VGND.n14 VGND.n13 0.120292
R167 VGND.n14 VGND.n5 0.120292
R168 VGND.n21 VGND.n5 0.120292
R169 VGND.n22 VGND.n21 0.120292
R170 VGND.n23 VGND.n22 0.120292
R171 VGND.n23 VGND.n3 0.120292
R172 VGND.n30 VGND.n3 0.120292
R173 VGND.n31 VGND.n30 0.120292
R174 VGND.n32 VGND.n31 0.120292
R175 VGND.n32 VGND.n0 0.120292
R176 VGND VGND.n0 0.03175
R177 VNB.t6 VNB.t4 1196.12
R178 VNB.t9 VNB.t6 1196.12
R179 VNB.t7 VNB.t9 1196.12
R180 VNB.t0 VNB.t7 1196.12
R181 VNB.t5 VNB.t0 1196.12
R182 VNB.t8 VNB.t5 1196.12
R183 VNB.t1 VNB.t8 1196.12
R184 VNB.t10 VNB.t1 1196.12
R185 VNB.t2 VNB.t10 1196.12
R186 VNB.t11 VNB.t2 1196.12
R187 VNB.t3 VNB.t11 1196.12
R188 VNB.t14 VNB.t3 1196.12
R189 VNB.t15 VNB.t14 1196.12
R190 VNB.t13 VNB.t15 1196.12
R191 VNB VNB.t13 911.327
R192 VNB VNB.t12 284.791
R193 VPWR.n37 VPWR.t12 347.57
R194 VPWR.n35 VPWR.n1 320.976
R195 VPWR.n29 VPWR.n28 320.976
R196 VPWR.n26 VPWR.n4 310.502
R197 VPWR.n20 VPWR.n19 310.502
R198 VPWR.n18 VPWR.n7 310.502
R199 VPWR.n9 VPWR.n8 310.502
R200 VPWR.n12 VPWR.n11 310.502
R201 VPWR.n10 VPWR.t3 249.179
R202 VPWR.n30 VPWR.n27 34.6358
R203 VPWR.n34 VPWR.n2 34.6358
R204 VPWR.n25 VPWR.n5 34.6358
R205 VPWR.n37 VPWR.n36 32.377
R206 VPWR.n36 VPWR.n35 30.8711
R207 VPWR.n21 VPWR.n18 28.9887
R208 VPWR.n1 VPWR.t14 26.5955
R209 VPWR.n1 VPWR.t15 26.5955
R210 VPWR.n28 VPWR.t10 26.5955
R211 VPWR.n28 VPWR.t13 26.5955
R212 VPWR.n4 VPWR.t4 26.5955
R213 VPWR.n4 VPWR.t2 26.5955
R214 VPWR.n19 VPWR.t6 26.5955
R215 VPWR.n19 VPWR.t5 26.5955
R216 VPWR.n7 VPWR.t8 26.5955
R217 VPWR.n7 VPWR.t7 26.5955
R218 VPWR.n8 VPWR.t11 26.5955
R219 VPWR.n8 VPWR.t9 26.5955
R220 VPWR.n11 VPWR.t1 26.5955
R221 VPWR.n11 VPWR.t0 26.5955
R222 VPWR.n29 VPWR.n2 24.8476
R223 VPWR.n17 VPWR.n9 22.9652
R224 VPWR.n13 VPWR.n9 21.4593
R225 VPWR.n13 VPWR.n12 16.9417
R226 VPWR.n18 VPWR.n17 15.4358
R227 VPWR VPWR.n37 11.6479
R228 VPWR.n30 VPWR.n29 9.78874
R229 VPWR.n21 VPWR.n20 9.41227
R230 VPWR.n14 VPWR.n13 9.3005
R231 VPWR.n15 VPWR.n9 9.3005
R232 VPWR.n17 VPWR.n16 9.3005
R233 VPWR.n18 VPWR.n6 9.3005
R234 VPWR.n22 VPWR.n21 9.3005
R235 VPWR.n23 VPWR.n5 9.3005
R236 VPWR.n25 VPWR.n24 9.3005
R237 VPWR.n27 VPWR.n3 9.3005
R238 VPWR.n31 VPWR.n30 9.3005
R239 VPWR.n32 VPWR.n2 9.3005
R240 VPWR.n34 VPWR.n33 9.3005
R241 VPWR.n36 VPWR.n0 9.3005
R242 VPWR.n12 VPWR.n10 6.64192
R243 VPWR.n27 VPWR.n26 6.4005
R244 VPWR.n35 VPWR.n34 3.76521
R245 VPWR.n26 VPWR.n25 3.38874
R246 VPWR.n14 VPWR.n10 0.78172
R247 VPWR.n20 VPWR.n5 0.376971
R248 VPWR.n15 VPWR.n14 0.120292
R249 VPWR.n16 VPWR.n15 0.120292
R250 VPWR.n16 VPWR.n6 0.120292
R251 VPWR.n22 VPWR.n6 0.120292
R252 VPWR.n23 VPWR.n22 0.120292
R253 VPWR.n24 VPWR.n23 0.120292
R254 VPWR.n24 VPWR.n3 0.120292
R255 VPWR.n31 VPWR.n3 0.120292
R256 VPWR.n32 VPWR.n31 0.120292
R257 VPWR.n33 VPWR.n32 0.120292
R258 VPWR.n33 VPWR.n0 0.120292
R259 VPWR VPWR.n0 0.03175
R260 VPB.t1 VPB.t3 248.599
R261 VPB.t0 VPB.t1 248.599
R262 VPB.t11 VPB.t0 248.599
R263 VPB.t9 VPB.t11 248.599
R264 VPB.t8 VPB.t9 248.599
R265 VPB.t7 VPB.t8 248.599
R266 VPB.t6 VPB.t7 248.599
R267 VPB.t5 VPB.t6 248.599
R268 VPB.t4 VPB.t5 248.599
R269 VPB.t2 VPB.t4 248.599
R270 VPB.t10 VPB.t2 248.599
R271 VPB.t13 VPB.t10 248.599
R272 VPB.t14 VPB.t13 248.599
R273 VPB.t15 VPB.t14 248.599
R274 VPB VPB.t15 189.409
R275 VPB VPB.t12 59.1905
R276 A.n9 A.t6 235.554
R277 A.n2 A.t0 221.72
R278 A.n4 A.t1 221.72
R279 A.n0 A.t2 221.72
R280 A.n9 A.t7 163.254
R281 A.n3 A.n1 152
R282 A.n6 A.n5 152
R283 A.n8 A.n7 152
R284 A.n10 A.n9 152
R285 A.n2 A.t4 149.421
R286 A.n4 A.t5 149.421
R287 A.n0 A.t3 149.421
R288 A.n3 A.n2 58.019
R289 A.n5 A.n4 43.7375
R290 A.n9 A.n8 32.1338
R291 A.n5 A.n0 31.2412
R292 A.n8 A.n0 29.4561
R293 A.n6 A.n1 21.7605
R294 A.n7 A 19.5205
R295 A.n4 A.n3 16.9598
R296 A.n10 A 11.8405
R297 A.n7 A 9.9205
R298 A A.n10 9.9205
R299 A.n1 A 5.4405
R300 A A.n6 2.2405
C0 VPB A 0.132061f
C1 VPB VPWR 0.148372f
C2 A VPWR 0.080969f
C3 VPB X 0.024481f
C4 A X 6.16e-19
C5 VPB VGND 0.01077f
C6 A VGND 0.091246f
C7 VPWR X 1.01279f
C8 VPWR VGND 0.168922f
C9 X VGND 0.751669f
C10 VGND VNB 0.835647f
C11 X VNB 0.082954f
C12 VPWR VNB 0.727686f
C13 A VNB 0.415834f
C14 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_16 VNB VPB VGND VPWR A X
X0 VGND.t5 A.t0 a_109_47.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X.t15 a_109_47.t12 VPWR.t21 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t21 a_109_47.t13 X.t31 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t20 a_109_47.t14 X.t30 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X.t14 a_109_47.t15 VPWR.t20 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t19 a_109_47.t16 X.t29 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t19 a_109_47.t17 X.t13 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_47.t11 A.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 X.t12 a_109_47.t18 VPWR.t18 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR.t4 A.t2 a_109_47.t10 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X.t28 a_109_47.t19 VGND.t18 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X.t27 a_109_47.t20 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t26 a_109_47.t21 VGND.t16 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 X.t25 a_109_47.t22 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_47.t9 A.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t17 a_109_47.t23 X.t11 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X.t24 a_109_47.t24 VGND.t14 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 X.t10 a_109_47.t25 VPWR.t16 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR.t2 A.t4 a_109_47.t8 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t15 a_109_47.t26 X.t9 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t4 A.t5 a_109_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t3 A.t6 a_109_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND.t13 a_109_47.t27 X.t23 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 X.t8 a_109_47.t28 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND.t12 a_109_47.t29 X.t22 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VPWR.t13 a_109_47.t30 X.t7 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND.t11 a_109_47.t31 X.t21 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR.t12 a_109_47.t32 X.t6 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X.t5 a_109_47.t33 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND.t10 a_109_47.t34 X.t20 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_109_47.t2 A.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_109_47.t1 A.t8 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 X.t4 a_109_47.t35 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR.t9 a_109_47.t36 X.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X.t19 a_109_47.t37 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 X.t18 a_109_47.t38 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 VPWR.t1 A.t9 a_109_47.t7 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X.t2 a_109_47.t39 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 X.t17 a_109_47.t40 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_109_47.t6 A.t10 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR.t7 a_109_47.t41 X.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR.t6 a_109_47.t42 X.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_109_47.t0 A.t11 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND.t6 a_109_47.t43 X.t16 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A.n3 A.t9 221.72
R1 A.n2 A.t1 221.72
R2 A.n7 A.t2 221.72
R3 A.n9 A.t3 221.72
R4 A.n12 A.t4 221.72
R5 A.n10 A.t10 221.72
R6 A.n11 A.n1 173.761
R7 A A.n4 171.84
R8 A.n6 A.n5 152
R9 A.n8 A.n0 152
R10 A.n15 A.n14 152
R11 A.n13 A.n1 152
R12 A.n3 A.t0 149.421
R13 A.n2 A.t8 149.421
R14 A.n7 A.t6 149.421
R15 A.n9 A.t7 149.421
R16 A.n12 A.t5 149.421
R17 A.n10 A.t11 149.421
R18 A.n14 A.n13 60.6968
R19 A.n9 A.n8 55.3412
R20 A.n12 A.n11 51.7709
R21 A.n4 A.n3 48.2005
R22 A.n7 A.n6 41.0598
R23 A.n6 A.n2 33.919
R24 A.n4 A.n2 26.7783
R25 A.n11 A.n10 23.2079
R26 A.n5 A.n0 21.7605
R27 A.n15 A.n1 21.7605
R28 A.n8 A.n7 19.6375
R29 A A.n15 16.0005
R30 A.n13 A.n12 8.92643
R31 A A.n0 5.7605
R32 A.n14 A.n9 5.35606
R33 A.n5 A 1.9205
R34 a_109_47.n61 a_109_47.n60 244.457
R35 a_109_47.n15 a_109_47.t42 221.72
R36 a_109_47.n17 a_109_47.t15 221.72
R37 a_109_47.n14 a_109_47.t17 221.72
R38 a_109_47.n22 a_109_47.t18 221.72
R39 a_109_47.n24 a_109_47.t30 221.72
R40 a_109_47.n25 a_109_47.t33 221.72
R41 a_109_47.n31 a_109_47.t36 221.72
R42 a_109_47.n33 a_109_47.t39 221.72
R43 a_109_47.n10 a_109_47.t41 221.72
R44 a_109_47.n38 a_109_47.t12 221.72
R45 a_109_47.n8 a_109_47.t23 221.72
R46 a_109_47.n44 a_109_47.t25 221.72
R47 a_109_47.n46 a_109_47.t26 221.72
R48 a_109_47.n6 a_109_47.t28 221.72
R49 a_109_47.n52 a_109_47.t32 221.72
R50 a_109_47.n53 a_109_47.t35 221.72
R51 a_109_47.n58 a_109_47.n57 206.056
R52 a_109_47.n60 a_109_47.n59 206.056
R53 a_109_47.n55 a_109_47.n54 152
R54 a_109_47.n51 a_109_47.n5 152
R55 a_109_47.n50 a_109_47.n49 152
R56 a_109_47.n48 a_109_47.n47 152
R57 a_109_47.n45 a_109_47.n7 152
R58 a_109_47.n43 a_109_47.n42 152
R59 a_109_47.n41 a_109_47.n40 152
R60 a_109_47.n39 a_109_47.n9 152
R61 a_109_47.n37 a_109_47.n36 152
R62 a_109_47.n35 a_109_47.n34 152
R63 a_109_47.n32 a_109_47.n11 152
R64 a_109_47.n30 a_109_47.n29 152
R65 a_109_47.n28 a_109_47.n12 152
R66 a_109_47.n27 a_109_47.n26 152
R67 a_109_47.n23 a_109_47.n13 152
R68 a_109_47.n21 a_109_47.n20 152
R69 a_109_47.n19 a_109_47.n18 152
R70 a_109_47.n15 a_109_47.t34 149.421
R71 a_109_47.n17 a_109_47.t40 149.421
R72 a_109_47.n14 a_109_47.t31 149.421
R73 a_109_47.n22 a_109_47.t24 149.421
R74 a_109_47.n24 a_109_47.t29 149.421
R75 a_109_47.n25 a_109_47.t22 149.421
R76 a_109_47.n31 a_109_47.t27 149.421
R77 a_109_47.n33 a_109_47.t20 149.421
R78 a_109_47.n10 a_109_47.t14 149.421
R79 a_109_47.n38 a_109_47.t19 149.421
R80 a_109_47.n8 a_109_47.t43 149.421
R81 a_109_47.n44 a_109_47.t21 149.421
R82 a_109_47.n46 a_109_47.t16 149.421
R83 a_109_47.n6 a_109_47.t38 149.421
R84 a_109_47.n52 a_109_47.t13 149.421
R85 a_109_47.n53 a_109_47.t37 149.421
R86 a_109_47.n2 a_109_47.n0 137.189
R87 a_109_47.n2 a_109_47.n1 98.788
R88 a_109_47.n4 a_109_47.n3 98.788
R89 a_109_47.n19 a_109_47.n16 90.1038
R90 a_109_47.n30 a_109_47.n12 60.6968
R91 a_109_47.n40 a_109_47.n39 60.6968
R92 a_109_47.n51 a_109_47.n50 60.6968
R93 a_109_47.n18 a_109_47.n17 58.9116
R94 a_109_47.n26 a_109_47.n25 58.9116
R95 a_109_47.n38 a_109_47.n37 55.3412
R96 a_109_47.n54 a_109_47.n52 55.3412
R97 a_109_47.n43 a_109_47.n8 51.7709
R98 a_109_47.n47 a_109_47.n6 51.7709
R99 a_109_47.n32 a_109_47.n31 48.2005
R100 a_109_47.n21 a_109_47.n14 44.6301
R101 a_109_47.n24 a_109_47.n23 44.6301
R102 a_109_47.n34 a_109_47.n10 41.0598
R103 a_109_47.n16 a_109_47.n15 39.7878
R104 a_109_47.n4 a_109_47.n2 38.4005
R105 a_109_47.n60 a_109_47.n58 38.4005
R106 a_109_47.n45 a_109_47.n44 37.4894
R107 a_109_47.n46 a_109_47.n45 37.4894
R108 a_109_47.n34 a_109_47.n33 33.919
R109 a_109_47.n56 a_109_47.n4 31.0755
R110 a_109_47.n58 a_109_47.n56 31.0755
R111 a_109_47.n22 a_109_47.n21 30.3486
R112 a_109_47.n23 a_109_47.n22 30.3486
R113 a_109_47.n33 a_109_47.n32 26.7783
R114 a_109_47.n57 a_109_47.t7 26.5955
R115 a_109_47.n57 a_109_47.t11 26.5955
R116 a_109_47.n59 a_109_47.t10 26.5955
R117 a_109_47.n59 a_109_47.t9 26.5955
R118 a_109_47.n61 a_109_47.t8 26.5955
R119 a_109_47.t6 a_109_47.n61 26.5955
R120 a_109_47.n17 a_109_47.n16 25.6591
R121 a_109_47.n0 a_109_47.t4 24.9236
R122 a_109_47.n0 a_109_47.t0 24.9236
R123 a_109_47.n1 a_109_47.t3 24.9236
R124 a_109_47.n1 a_109_47.t2 24.9236
R125 a_109_47.n3 a_109_47.t5 24.9236
R126 a_109_47.n3 a_109_47.t1 24.9236
R127 a_109_47.n44 a_109_47.n43 23.2079
R128 a_109_47.n47 a_109_47.n46 23.2079
R129 a_109_47.n20 a_109_47.n19 21.7605
R130 a_109_47.n20 a_109_47.n13 21.7605
R131 a_109_47.n27 a_109_47.n13 21.7605
R132 a_109_47.n28 a_109_47.n27 21.7605
R133 a_109_47.n29 a_109_47.n28 21.7605
R134 a_109_47.n29 a_109_47.n11 21.7605
R135 a_109_47.n35 a_109_47.n11 21.7605
R136 a_109_47.n36 a_109_47.n35 21.7605
R137 a_109_47.n36 a_109_47.n9 21.7605
R138 a_109_47.n41 a_109_47.n9 21.7605
R139 a_109_47.n42 a_109_47.n41 21.7605
R140 a_109_47.n42 a_109_47.n7 21.7605
R141 a_109_47.n48 a_109_47.n7 21.7605
R142 a_109_47.n49 a_109_47.n48 21.7605
R143 a_109_47.n49 a_109_47.n5 21.7605
R144 a_109_47.n55 a_109_47.n5 21.7605
R145 a_109_47.n56 a_109_47.n55 20.8005
R146 a_109_47.n37 a_109_47.n10 19.6375
R147 a_109_47.n54 a_109_47.n53 19.6375
R148 a_109_47.n18 a_109_47.n14 16.0672
R149 a_109_47.n26 a_109_47.n24 16.0672
R150 a_109_47.n31 a_109_47.n30 12.4968
R151 a_109_47.n40 a_109_47.n8 8.92643
R152 a_109_47.n50 a_109_47.n6 8.92643
R153 a_109_47.n39 a_109_47.n38 5.35606
R154 a_109_47.n52 a_109_47.n51 5.35606
R155 a_109_47.n25 a_109_47.n12 1.78569
R156 VGND.n18 VGND.t10 291.125
R157 VGND.n17 VGND.n16 208.719
R158 VGND.n22 VGND.n14 208.719
R159 VGND.n12 VGND.n11 208.719
R160 VGND.n29 VGND.n10 208.719
R161 VGND.n31 VGND.n30 208.719
R162 VGND.n37 VGND.n7 208.719
R163 VGND.n40 VGND.n39 208.719
R164 VGND.n46 VGND.n4 208.719
R165 VGND.n49 VGND.n48 208.719
R166 VGND.n55 VGND.n1 208.719
R167 VGND.n57 VGND.t0 161.302
R168 VGND.n21 VGND.n15 34.6358
R169 VGND.n24 VGND.n23 34.6358
R170 VGND.n28 VGND.n27 34.6358
R171 VGND.n36 VGND.n8 34.6358
R172 VGND.n41 VGND.n38 34.6358
R173 VGND.n45 VGND.n5 34.6358
R174 VGND.n50 VGND.n47 34.6358
R175 VGND.n54 VGND.n2 34.6358
R176 VGND.n32 VGND.n31 33.8829
R177 VGND.n57 VGND.n56 32.377
R178 VGND.n56 VGND.n55 30.8711
R179 VGND.n18 VGND.n17 29.7335
R180 VGND.n32 VGND.n29 29.3652
R181 VGND.n37 VGND.n36 27.8593
R182 VGND.n16 VGND.t7 24.9236
R183 VGND.n16 VGND.t11 24.9236
R184 VGND.n14 VGND.t14 24.9236
R185 VGND.n14 VGND.t12 24.9236
R186 VGND.n11 VGND.t15 24.9236
R187 VGND.n11 VGND.t13 24.9236
R188 VGND.n10 VGND.t17 24.9236
R189 VGND.n10 VGND.t20 24.9236
R190 VGND.n30 VGND.t18 24.9236
R191 VGND.n30 VGND.t6 24.9236
R192 VGND.n7 VGND.t16 24.9236
R193 VGND.n7 VGND.t19 24.9236
R194 VGND.n39 VGND.t8 24.9236
R195 VGND.n39 VGND.t21 24.9236
R196 VGND.n4 VGND.t9 24.9236
R197 VGND.n4 VGND.t5 24.9236
R198 VGND.n48 VGND.t1 24.9236
R199 VGND.n48 VGND.t3 24.9236
R200 VGND.n1 VGND.t2 24.9236
R201 VGND.n1 VGND.t4 24.9236
R202 VGND.n49 VGND.n2 24.8476
R203 VGND.n27 VGND.n12 23.3417
R204 VGND.n41 VGND.n40 21.8358
R205 VGND.n47 VGND.n46 18.824
R206 VGND.n22 VGND.n21 17.3181
R207 VGND.n23 VGND.n22 17.3181
R208 VGND.n46 VGND.n45 15.8123
R209 VGND.n40 VGND.n5 12.8005
R210 VGND.n58 VGND.n57 11.5593
R211 VGND.n17 VGND.n15 11.2946
R212 VGND.n24 VGND.n12 11.2946
R213 VGND.n50 VGND.n49 9.78874
R214 VGND.n19 VGND.n15 9.3005
R215 VGND.n21 VGND.n20 9.3005
R216 VGND.n23 VGND.n13 9.3005
R217 VGND.n25 VGND.n24 9.3005
R218 VGND.n27 VGND.n26 9.3005
R219 VGND.n28 VGND.n9 9.3005
R220 VGND.n33 VGND.n32 9.3005
R221 VGND.n34 VGND.n8 9.3005
R222 VGND.n36 VGND.n35 9.3005
R223 VGND.n38 VGND.n6 9.3005
R224 VGND.n42 VGND.n41 9.3005
R225 VGND.n43 VGND.n5 9.3005
R226 VGND.n45 VGND.n44 9.3005
R227 VGND.n47 VGND.n3 9.3005
R228 VGND.n51 VGND.n50 9.3005
R229 VGND.n52 VGND.n2 9.3005
R230 VGND.n54 VGND.n53 9.3005
R231 VGND.n56 VGND.n0 9.3005
R232 VGND.n38 VGND.n37 6.77697
R233 VGND.n29 VGND.n28 5.27109
R234 VGND.n55 VGND.n54 3.76521
R235 VGND.n19 VGND.n18 1.35766
R236 VGND.n31 VGND.n8 0.753441
R237 VGND.n20 VGND.n19 0.120292
R238 VGND.n20 VGND.n13 0.120292
R239 VGND.n25 VGND.n13 0.120292
R240 VGND.n26 VGND.n25 0.120292
R241 VGND.n26 VGND.n9 0.120292
R242 VGND.n33 VGND.n9 0.120292
R243 VGND.n34 VGND.n33 0.120292
R244 VGND.n35 VGND.n34 0.120292
R245 VGND.n35 VGND.n6 0.120292
R246 VGND.n42 VGND.n6 0.120292
R247 VGND.n43 VGND.n42 0.120292
R248 VGND.n44 VGND.n43 0.120292
R249 VGND.n44 VGND.n3 0.120292
R250 VGND.n51 VGND.n3 0.120292
R251 VGND.n52 VGND.n51 0.120292
R252 VGND.n53 VGND.n52 0.120292
R253 VGND.n53 VGND.n0 0.120292
R254 VGND.n58 VGND.n0 0.120292
R255 VGND VGND.n58 0.0213333
R256 VNB.t7 VNB.t10 1196.12
R257 VNB.t11 VNB.t7 1196.12
R258 VNB.t14 VNB.t11 1196.12
R259 VNB.t12 VNB.t14 1196.12
R260 VNB.t15 VNB.t12 1196.12
R261 VNB.t13 VNB.t15 1196.12
R262 VNB.t17 VNB.t13 1196.12
R263 VNB.t20 VNB.t17 1196.12
R264 VNB.t18 VNB.t20 1196.12
R265 VNB.t6 VNB.t18 1196.12
R266 VNB.t16 VNB.t6 1196.12
R267 VNB.t19 VNB.t16 1196.12
R268 VNB.t8 VNB.t19 1196.12
R269 VNB.t21 VNB.t8 1196.12
R270 VNB.t9 VNB.t21 1196.12
R271 VNB.t5 VNB.t9 1196.12
R272 VNB.t1 VNB.t5 1196.12
R273 VNB.t3 VNB.t1 1196.12
R274 VNB.t2 VNB.t3 1196.12
R275 VNB.t4 VNB.t2 1196.12
R276 VNB.t0 VNB.t4 1196.12
R277 VNB VNB.t0 911.327
R278 VPWR.n18 VPWR.t6 356.132
R279 VPWR.n55 VPWR.n1 320.976
R280 VPWR.n49 VPWR.n48 320.976
R281 VPWR.n46 VPWR.n4 320.976
R282 VPWR.n40 VPWR.n39 320.976
R283 VPWR.n37 VPWR.n7 320.976
R284 VPWR.n31 VPWR.n30 320.976
R285 VPWR.n29 VPWR.n10 320.976
R286 VPWR.n12 VPWR.n11 320.976
R287 VPWR.n22 VPWR.n14 320.976
R288 VPWR.n17 VPWR.n16 320.976
R289 VPWR.n57 VPWR.t0 257.474
R290 VPWR.n21 VPWR.n15 34.6358
R291 VPWR.n24 VPWR.n23 34.6358
R292 VPWR.n28 VPWR.n27 34.6358
R293 VPWR.n36 VPWR.n8 34.6358
R294 VPWR.n41 VPWR.n38 34.6358
R295 VPWR.n45 VPWR.n5 34.6358
R296 VPWR.n50 VPWR.n47 34.6358
R297 VPWR.n54 VPWR.n2 34.6358
R298 VPWR.n32 VPWR.n31 33.8829
R299 VPWR.n57 VPWR.n56 32.377
R300 VPWR.n56 VPWR.n55 30.8711
R301 VPWR.n18 VPWR.n17 29.7335
R302 VPWR.n32 VPWR.n29 29.3652
R303 VPWR.n37 VPWR.n36 27.8593
R304 VPWR.n1 VPWR.t3 26.5955
R305 VPWR.n1 VPWR.t2 26.5955
R306 VPWR.n48 VPWR.t5 26.5955
R307 VPWR.n48 VPWR.t4 26.5955
R308 VPWR.n4 VPWR.t10 26.5955
R309 VPWR.n4 VPWR.t1 26.5955
R310 VPWR.n39 VPWR.t14 26.5955
R311 VPWR.n39 VPWR.t12 26.5955
R312 VPWR.n7 VPWR.t16 26.5955
R313 VPWR.n7 VPWR.t15 26.5955
R314 VPWR.n30 VPWR.t21 26.5955
R315 VPWR.n30 VPWR.t17 26.5955
R316 VPWR.n10 VPWR.t8 26.5955
R317 VPWR.n10 VPWR.t7 26.5955
R318 VPWR.n11 VPWR.t11 26.5955
R319 VPWR.n11 VPWR.t9 26.5955
R320 VPWR.n14 VPWR.t18 26.5955
R321 VPWR.n14 VPWR.t13 26.5955
R322 VPWR.n16 VPWR.t20 26.5955
R323 VPWR.n16 VPWR.t19 26.5955
R324 VPWR.n49 VPWR.n2 24.8476
R325 VPWR.n27 VPWR.n12 23.3417
R326 VPWR.n41 VPWR.n40 21.8358
R327 VPWR.n47 VPWR.n46 18.824
R328 VPWR.n22 VPWR.n21 17.3181
R329 VPWR.n23 VPWR.n22 17.3181
R330 VPWR.n46 VPWR.n45 15.8123
R331 VPWR.n40 VPWR.n5 12.8005
R332 VPWR.n58 VPWR.n57 11.5593
R333 VPWR.n17 VPWR.n15 11.2946
R334 VPWR.n24 VPWR.n12 11.2946
R335 VPWR.n50 VPWR.n49 9.78874
R336 VPWR.n19 VPWR.n15 9.3005
R337 VPWR.n21 VPWR.n20 9.3005
R338 VPWR.n23 VPWR.n13 9.3005
R339 VPWR.n25 VPWR.n24 9.3005
R340 VPWR.n27 VPWR.n26 9.3005
R341 VPWR.n28 VPWR.n9 9.3005
R342 VPWR.n33 VPWR.n32 9.3005
R343 VPWR.n34 VPWR.n8 9.3005
R344 VPWR.n36 VPWR.n35 9.3005
R345 VPWR.n38 VPWR.n6 9.3005
R346 VPWR.n42 VPWR.n41 9.3005
R347 VPWR.n43 VPWR.n5 9.3005
R348 VPWR.n45 VPWR.n44 9.3005
R349 VPWR.n47 VPWR.n3 9.3005
R350 VPWR.n51 VPWR.n50 9.3005
R351 VPWR.n52 VPWR.n2 9.3005
R352 VPWR.n54 VPWR.n53 9.3005
R353 VPWR.n56 VPWR.n0 9.3005
R354 VPWR.n38 VPWR.n37 6.77697
R355 VPWR.n29 VPWR.n28 5.27109
R356 VPWR.n55 VPWR.n54 3.76521
R357 VPWR.n19 VPWR.n18 1.35766
R358 VPWR.n31 VPWR.n8 0.753441
R359 VPWR.n20 VPWR.n19 0.120292
R360 VPWR.n20 VPWR.n13 0.120292
R361 VPWR.n25 VPWR.n13 0.120292
R362 VPWR.n26 VPWR.n25 0.120292
R363 VPWR.n26 VPWR.n9 0.120292
R364 VPWR.n33 VPWR.n9 0.120292
R365 VPWR.n34 VPWR.n33 0.120292
R366 VPWR.n35 VPWR.n34 0.120292
R367 VPWR.n35 VPWR.n6 0.120292
R368 VPWR.n42 VPWR.n6 0.120292
R369 VPWR.n43 VPWR.n42 0.120292
R370 VPWR.n44 VPWR.n43 0.120292
R371 VPWR.n44 VPWR.n3 0.120292
R372 VPWR.n51 VPWR.n3 0.120292
R373 VPWR.n52 VPWR.n51 0.120292
R374 VPWR.n53 VPWR.n52 0.120292
R375 VPWR.n53 VPWR.n0 0.120292
R376 VPWR.n58 VPWR.n0 0.120292
R377 VPWR VPWR.n58 0.0213333
R378 X.n2 X.n0 244.457
R379 X.n2 X.n1 206.056
R380 X.n4 X.n3 206.056
R381 X.n6 X.n5 206.056
R382 X.n8 X.n7 206.056
R383 X.n10 X.n9 206.056
R384 X.n12 X.n11 206.056
R385 X.n14 X.n13 206.056
R386 X.n17 X.n15 137.189
R387 X.n17 X.n16 98.788
R388 X.n19 X.n18 98.788
R389 X.n21 X.n20 98.788
R390 X.n23 X.n22 98.788
R391 X.n25 X.n24 98.788
R392 X.n27 X.n26 98.788
R393 X.n29 X.n28 98.788
R394 X X.n29 40.4711
R395 X.n19 X.n17 38.4005
R396 X.n21 X.n19 38.4005
R397 X.n23 X.n21 38.4005
R398 X.n25 X.n23 38.4005
R399 X.n27 X.n25 38.4005
R400 X.n29 X.n27 38.4005
R401 X.n4 X.n2 38.4005
R402 X.n6 X.n4 38.4005
R403 X.n8 X.n6 38.4005
R404 X.n10 X.n8 38.4005
R405 X.n12 X.n10 38.4005
R406 X.n14 X.n12 38.4005
R407 X X.n14 33.7342
R408 X.n0 X.t6 26.5955
R409 X.n0 X.t4 26.5955
R410 X.n1 X.t9 26.5955
R411 X.n1 X.t8 26.5955
R412 X.n3 X.t11 26.5955
R413 X.n3 X.t10 26.5955
R414 X.n5 X.t1 26.5955
R415 X.n5 X.t15 26.5955
R416 X.n7 X.t3 26.5955
R417 X.n7 X.t2 26.5955
R418 X.n9 X.t7 26.5955
R419 X.n9 X.t5 26.5955
R420 X.n11 X.t13 26.5955
R421 X.n11 X.t12 26.5955
R422 X.n13 X.t0 26.5955
R423 X.n13 X.t14 26.5955
R424 X.n15 X.t31 24.9236
R425 X.n15 X.t19 24.9236
R426 X.n16 X.t29 24.9236
R427 X.n16 X.t18 24.9236
R428 X.n18 X.t16 24.9236
R429 X.n18 X.t26 24.9236
R430 X.n20 X.t30 24.9236
R431 X.n20 X.t28 24.9236
R432 X.n22 X.t23 24.9236
R433 X.n22 X.t27 24.9236
R434 X.n24 X.t22 24.9236
R435 X.n24 X.t25 24.9236
R436 X.n26 X.t21 24.9236
R437 X.n26 X.t24 24.9236
R438 X.n28 X.t20 24.9236
R439 X.n28 X.t17 24.9236
R440 VPB.t20 VPB.t6 248.599
R441 VPB.t19 VPB.t20 248.599
R442 VPB.t18 VPB.t19 248.599
R443 VPB.t13 VPB.t18 248.599
R444 VPB.t11 VPB.t13 248.599
R445 VPB.t9 VPB.t11 248.599
R446 VPB.t8 VPB.t9 248.599
R447 VPB.t7 VPB.t8 248.599
R448 VPB.t21 VPB.t7 248.599
R449 VPB.t17 VPB.t21 248.599
R450 VPB.t16 VPB.t17 248.599
R451 VPB.t15 VPB.t16 248.599
R452 VPB.t14 VPB.t15 248.599
R453 VPB.t12 VPB.t14 248.599
R454 VPB.t10 VPB.t12 248.599
R455 VPB.t1 VPB.t10 248.599
R456 VPB.t5 VPB.t1 248.599
R457 VPB.t4 VPB.t5 248.599
R458 VPB.t3 VPB.t4 248.599
R459 VPB.t2 VPB.t3 248.599
R460 VPB.t0 VPB.t2 248.599
R461 VPB VPB.t0 189.409
C0 VPB A 0.18511f
C1 VPB VPWR 0.200549f
C2 A VPWR 0.115105f
C3 VPB X 0.054017f
C4 A X 0.001696f
C5 VPB VGND 0.013036f
C6 A VGND 0.109982f
C7 VPWR X 1.52599f
C8 VPWR VGND 0.207673f
C9 X VGND 1.10184f
C10 VGND VNB 1.12477f
C11 X VNB 0.122283f
C12 VPWR VNB 0.962735f
C13 A VNB 0.577934f
C14 VPB VNB 2.0223f
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufbuf_8 VNB VPB VGND VPWR A X
X0 a_318_47.t5 a_206_47.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t6 a_318_47.t6 X.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 a_206_47.t3 a_318_47.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 X.t15 a_318_47.t7 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X.t6 a_318_47.t8 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t8 a_318_47.t9 X.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X.t4 a_318_47.t10 VPWR.t9 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t2 a_206_47.t4 a_318_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR.t10 a_318_47.t11 X.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t2 a_318_47.t12 VPWR.t11 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_318_47.t1 a_206_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X.t14 a_318_47.t13 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_206_47.t0 a_27_47.t2 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13 X.t13 a_318_47.t14 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_206_47.t1 a_27_47.t3 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X15 VPWR.t3 a_318_47.t15 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t0 a_206_47.t6 a_318_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t8 a_318_47.t16 X.t12 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t7 a_318_47.t17 X.t11 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VGND.t6 a_318_47.t18 X.t10 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 X.t0 a_318_47.t19 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND.t5 a_318_47.t20 X.t9 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t0 a_206_47.t7 a_318_47.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t5 A.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X24 VGND.t3 A.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 X.t8 a_318_47.t21 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_206_47.t1 a_206_47.n6 251.038
R1 a_206_47.n0 a_206_47.t7 221.72
R2 a_206_47.n2 a_206_47.t2 221.72
R3 a_206_47.n3 a_206_47.t3 221.72
R4 a_206_47.n5 a_206_47.n1 173.761
R5 a_206_47.n6 a_206_47.t0 156.28
R6 a_206_47.n5 a_206_47.n4 152
R7 a_206_47.n0 a_206_47.t6 149.421
R8 a_206_47.n2 a_206_47.t5 149.421
R9 a_206_47.n3 a_206_47.t4 149.421
R10 a_206_47.n6 a_206_47.n5 53.7605
R11 a_206_47.n1 a_206_47.n0 51.7709
R12 a_206_47.n4 a_206_47.n2 37.4894
R13 a_206_47.n4 a_206_47.n3 37.4894
R14 a_206_47.n2 a_206_47.n1 23.2079
R15 VPWR.n34 VPWR.n1 636.577
R16 VPWR.n12 VPWR.t6 358.002
R17 VPWR.n27 VPWR.n4 320.976
R18 VPWR.n25 VPWR.n5 320.976
R19 VPWR.n19 VPWR.n18 320.976
R20 VPWR.n16 VPWR.n8 320.976
R21 VPWR.n11 VPWR.n10 320.976
R22 VPWR.n1 VPWR.t12 50.6025
R23 VPWR.n35 VPWR.n34 43.1829
R24 VPWR.n1 VPWR.t5 41.5552
R25 VPWR.n15 VPWR.n9 34.6358
R26 VPWR.n20 VPWR.n17 34.6358
R27 VPWR.n24 VPWR.n6 34.6358
R28 VPWR.n28 VPWR.n2 34.6358
R29 VPWR.n32 VPWR.n2 34.6358
R30 VPWR.n33 VPWR.n32 34.6358
R31 VPWR.n26 VPWR.n25 33.5064
R32 VPWR.n27 VPWR.n26 29.7417
R33 VPWR.n19 VPWR.n6 27.4829
R34 VPWR.n4 VPWR.t2 26.5955
R35 VPWR.n4 VPWR.t1 26.5955
R36 VPWR.n5 VPWR.t4 26.5955
R37 VPWR.n5 VPWR.t0 26.5955
R38 VPWR.n18 VPWR.t11 26.5955
R39 VPWR.n18 VPWR.t3 26.5955
R40 VPWR.n8 VPWR.t9 26.5955
R41 VPWR.n8 VPWR.t10 26.5955
R42 VPWR.n10 VPWR.t7 26.5955
R43 VPWR.n10 VPWR.t8 26.5955
R44 VPWR.n12 VPWR.n11 25.7221
R45 VPWR.n17 VPWR.n16 21.4593
R46 VPWR.n11 VPWR.n9 15.4358
R47 VPWR.n16 VPWR.n15 13.177
R48 VPWR.n13 VPWR.n9 9.3005
R49 VPWR.n15 VPWR.n14 9.3005
R50 VPWR.n17 VPWR.n7 9.3005
R51 VPWR.n21 VPWR.n20 9.3005
R52 VPWR.n22 VPWR.n6 9.3005
R53 VPWR.n24 VPWR.n23 9.3005
R54 VPWR.n26 VPWR.n3 9.3005
R55 VPWR.n29 VPWR.n28 9.3005
R56 VPWR.n30 VPWR.n2 9.3005
R57 VPWR.n32 VPWR.n31 9.3005
R58 VPWR.n33 VPWR.n0 9.3005
R59 VPWR.n20 VPWR.n19 7.15344
R60 VPWR.n28 VPWR.n27 4.89462
R61 VPWR.n13 VPWR.n12 1.2279
R62 VPWR.n25 VPWR.n24 1.12991
R63 VPWR.n34 VPWR.n33 0.753441
R64 VPWR.n14 VPWR.n13 0.120292
R65 VPWR.n14 VPWR.n7 0.120292
R66 VPWR.n21 VPWR.n7 0.120292
R67 VPWR.n22 VPWR.n21 0.120292
R68 VPWR.n23 VPWR.n22 0.120292
R69 VPWR.n23 VPWR.n3 0.120292
R70 VPWR.n29 VPWR.n3 0.120292
R71 VPWR.n30 VPWR.n29 0.120292
R72 VPWR.n31 VPWR.n30 0.120292
R73 VPWR.n31 VPWR.n0 0.120292
R74 VPWR.n35 VPWR.n0 0.120292
R75 VPWR VPWR.n35 0.0213333
R76 a_318_47.n22 a_318_47.t4 271.051
R77 a_318_47.n5 a_318_47.t6 221.72
R78 a_318_47.n6 a_318_47.t8 221.72
R79 a_318_47.n7 a_318_47.t9 221.72
R80 a_318_47.n9 a_318_47.t10 221.72
R81 a_318_47.n11 a_318_47.t11 221.72
R82 a_318_47.n3 a_318_47.t12 221.72
R83 a_318_47.n17 a_318_47.t15 221.72
R84 a_318_47.n18 a_318_47.t19 221.72
R85 a_318_47.n23 a_318_47.n22 206.055
R86 a_318_47.n1 a_318_47.t2 176.525
R87 a_318_47.n8 a_318_47.n4 173.761
R88 a_318_47.n20 a_318_47.n19 152
R89 a_318_47.n16 a_318_47.n2 152
R90 a_318_47.n15 a_318_47.n14 152
R91 a_318_47.n13 a_318_47.n12 152
R92 a_318_47.n10 a_318_47.n4 152
R93 a_318_47.n5 a_318_47.t18 149.421
R94 a_318_47.n6 a_318_47.t21 149.421
R95 a_318_47.n7 a_318_47.t16 149.421
R96 a_318_47.n9 a_318_47.t7 149.421
R97 a_318_47.n11 a_318_47.t20 149.421
R98 a_318_47.n3 a_318_47.t14 149.421
R99 a_318_47.n17 a_318_47.t17 149.421
R100 a_318_47.n18 a_318_47.t13 149.421
R101 a_318_47.n1 a_318_47.n0 98.788
R102 a_318_47.n6 a_318_47.n5 74.9783
R103 a_318_47.n7 a_318_47.n6 74.9783
R104 a_318_47.n16 a_318_47.n15 60.6968
R105 a_318_47.n12 a_318_47.n3 55.3412
R106 a_318_47.n19 a_318_47.n17 51.7709
R107 a_318_47.n8 a_318_47.n7 48.2005
R108 a_318_47.n11 a_318_47.n10 41.0598
R109 a_318_47.n10 a_318_47.n9 33.919
R110 a_318_47.n21 a_318_47.n1 32.0005
R111 a_318_47.n22 a_318_47.n21 32.0005
R112 a_318_47.n9 a_318_47.n8 26.7783
R113 a_318_47.n23 a_318_47.t3 26.5955
R114 a_318_47.t5 a_318_47.n23 26.5955
R115 a_318_47.n0 a_318_47.t0 24.9236
R116 a_318_47.n0 a_318_47.t1 24.9236
R117 a_318_47.n19 a_318_47.n18 23.2079
R118 a_318_47.n13 a_318_47.n4 21.7605
R119 a_318_47.n14 a_318_47.n13 21.7605
R120 a_318_47.n14 a_318_47.n2 21.7605
R121 a_318_47.n20 a_318_47.n2 21.7605
R122 a_318_47.n21 a_318_47.n20 21.7605
R123 a_318_47.n12 a_318_47.n11 19.6375
R124 a_318_47.n17 a_318_47.n16 8.92643
R125 a_318_47.n15 a_318_47.n3 5.35606
R126 VPB.t12 VPB.t1 574.144
R127 VPB.t11 VPB.t12 287.072
R128 VPB.t9 VPB.t10 248.599
R129 VPB.t8 VPB.t9 248.599
R130 VPB.t7 VPB.t8 248.599
R131 VPB.t6 VPB.t7 248.599
R132 VPB.t5 VPB.t6 248.599
R133 VPB.t4 VPB.t5 248.599
R134 VPB.t3 VPB.t4 248.599
R135 VPB.t0 VPB.t3 248.599
R136 VPB.t2 VPB.t0 248.599
R137 VPB.t1 VPB.t2 248.599
R138 VPB VPB.t11 189.409
R139 X.n2 X.n0 244.457
R140 X.n2 X.n1 206.056
R141 X.n4 X.n3 206.056
R142 X.n6 X.n5 206.056
R143 X.n9 X.n7 137.189
R144 X.n9 X.n8 98.788
R145 X.n11 X.n10 98.788
R146 X.n13 X.n12 98.788
R147 X.n11 X.n9 38.4005
R148 X.n13 X.n11 38.4005
R149 X.n4 X.n2 38.4005
R150 X.n6 X.n4 38.4005
R151 X X.n13 36.3299
R152 X X.n6 29.5931
R153 X.n0 X.t1 26.5955
R154 X.n0 X.t0 26.5955
R155 X.n1 X.t3 26.5955
R156 X.n1 X.t2 26.5955
R157 X.n3 X.t5 26.5955
R158 X.n3 X.t4 26.5955
R159 X.n5 X.t7 26.5955
R160 X.n5 X.t6 26.5955
R161 X.n7 X.t11 24.9236
R162 X.n7 X.t14 24.9236
R163 X.n8 X.t9 24.9236
R164 X.n8 X.t13 24.9236
R165 X.n10 X.t12 24.9236
R166 X.n10 X.t15 24.9236
R167 X.n12 X.t10 24.9236
R168 X.n12 X.t8 24.9236
R169 VGND.n12 VGND.t6 292.995
R170 VGND.n11 VGND.n10 208.719
R171 VGND.n16 VGND.n8 208.719
R172 VGND.n19 VGND.n18 208.719
R173 VGND.n25 VGND.n5 208.719
R174 VGND.n27 VGND.n4 208.719
R175 VGND.n34 VGND.n1 208.719
R176 VGND.n1 VGND.t12 44.0005
R177 VGND.n35 VGND.n34 43.1829
R178 VGND.n1 VGND.t3 38.5719
R179 VGND.n15 VGND.n9 34.6358
R180 VGND.n20 VGND.n17 34.6358
R181 VGND.n24 VGND.n6 34.6358
R182 VGND.n28 VGND.n2 34.6358
R183 VGND.n32 VGND.n2 34.6358
R184 VGND.n33 VGND.n32 34.6358
R185 VGND.n26 VGND.n25 33.5064
R186 VGND.n27 VGND.n26 29.7417
R187 VGND.n19 VGND.n6 27.4829
R188 VGND.n12 VGND.n11 25.7221
R189 VGND.n10 VGND.t4 24.9236
R190 VGND.n10 VGND.t8 24.9236
R191 VGND.n8 VGND.t11 24.9236
R192 VGND.n8 VGND.t5 24.9236
R193 VGND.n18 VGND.t9 24.9236
R194 VGND.n18 VGND.t7 24.9236
R195 VGND.n5 VGND.t10 24.9236
R196 VGND.n5 VGND.t0 24.9236
R197 VGND.n4 VGND.t1 24.9236
R198 VGND.n4 VGND.t2 24.9236
R199 VGND.n17 VGND.n16 21.4593
R200 VGND.n11 VGND.n9 15.4358
R201 VGND.n16 VGND.n15 13.177
R202 VGND.n13 VGND.n9 9.3005
R203 VGND.n15 VGND.n14 9.3005
R204 VGND.n17 VGND.n7 9.3005
R205 VGND.n21 VGND.n20 9.3005
R206 VGND.n22 VGND.n6 9.3005
R207 VGND.n24 VGND.n23 9.3005
R208 VGND.n26 VGND.n3 9.3005
R209 VGND.n29 VGND.n28 9.3005
R210 VGND.n30 VGND.n2 9.3005
R211 VGND.n32 VGND.n31 9.3005
R212 VGND.n33 VGND.n0 9.3005
R213 VGND.n20 VGND.n19 7.15344
R214 VGND.n28 VGND.n27 4.89462
R215 VGND.n13 VGND.n12 1.2279
R216 VGND.n25 VGND.n24 1.12991
R217 VGND.n34 VGND.n33 0.753441
R218 VGND.n14 VGND.n13 0.120292
R219 VGND.n14 VGND.n7 0.120292
R220 VGND.n21 VGND.n7 0.120292
R221 VGND.n22 VGND.n21 0.120292
R222 VGND.n23 VGND.n22 0.120292
R223 VGND.n23 VGND.n3 0.120292
R224 VGND.n29 VGND.n3 0.120292
R225 VGND.n30 VGND.n29 0.120292
R226 VGND.n31 VGND.n30 0.120292
R227 VGND.n31 VGND.n0 0.120292
R228 VGND.n35 VGND.n0 0.120292
R229 VGND VGND.n35 0.0213333
R230 VNB.t12 VNB.t2 2762.46
R231 VNB.t3 VNB.t12 1381.23
R232 VNB.t4 VNB.t6 1196.12
R233 VNB.t8 VNB.t4 1196.12
R234 VNB.t11 VNB.t8 1196.12
R235 VNB.t5 VNB.t11 1196.12
R236 VNB.t9 VNB.t5 1196.12
R237 VNB.t7 VNB.t9 1196.12
R238 VNB.t10 VNB.t7 1196.12
R239 VNB.t0 VNB.t10 1196.12
R240 VNB.t1 VNB.t0 1196.12
R241 VNB.t2 VNB.t1 1196.12
R242 VNB VNB.t3 911.327
R243 a_27_47.t1 a_27_47.n1 398.351
R244 a_27_47.n1 a_27_47.t0 269.166
R245 a_27_47.n0 a_27_47.t3 239.986
R246 a_27_47.n0 a_27_47.t2 167.685
R247 a_27_47.n1 a_27_47.n0 152
R248 A.n0 A.t1 195.017
R249 A.n0 A.t0 172.524
R250 A A.n0 160
C0 X VGND 0.538027f
C1 VPB A 0.044244f
C2 VPB VPWR 0.15858f
C3 A VPWR 0.010259f
C4 VPB X 0.031607f
C5 VPB VGND 0.013151f
C6 A X 4.27e-19
C7 VPWR X 0.736898f
C8 A VGND 0.014854f
C9 VPWR VGND 0.140018f
C10 VGND VNB 0.786457f
C11 X VNB 0.076386f
C12 VPWR VNB 0.676923f
C13 A VNB 0.168818f
C14 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s15_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s15_2 VNB VPB VPWR VGND X A
X0 VPWR.t1 A.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.20085 pd=1.435 as=0.27 ps=2.54 w=1 l=0.15
X1 VGND.t4 a_362_333.t2 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.2058 pd=1.82 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VPWR.t3 a_228_47.t2 a_362_333.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.3136 pd=1.71 as=0.2173 ps=2.17 w=0.82 l=0.15
X3 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.128725 pd=1.085 as=0.1134 ps=1.38 w=0.42 l=0.15
X4 X.t2 a_362_333.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3136 ps=1.71 w=1 l=0.15
X5 X.t0 a_362_333.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.179575 ps=1.36 w=0.42 l=0.15
X6 VPWR.t0 a_362_333.t5 X.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.49 pd=2.98 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND.t2 a_228_47.t3 a_362_333.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.179575 pd=1.36 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_228_47.t1 a_27_47.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3116 pd=2.4 as=0.20085 ps=1.435 w=0.82 l=0.15
X9 a_228_47.t0 a_27_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.26325 pd=2.11 as=0.128725 ps=1.085 w=0.65 l=0.15
R0 A.n0 A.t0 241.144
R1 A.n0 A.t1 205.798
R2 A.n1 A.n0 152
R3 A.n1 A 7.7622
R4 A A.n1 1.49837
R5 a_27_47.t0 a_27_47.n1 408.616
R6 a_27_47.n1 a_27_47.t1 296.027
R7 a_27_47.n0 a_27_47.t2 270.358
R8 a_27_47.n0 a_27_47.t3 169.138
R9 a_27_47.n1 a_27_47.n0 165.554
R10 VPWR.n12 VPWR.n1 601.292
R11 VPWR.n5 VPWR.n4 601.292
R12 VPWR.n3 VPWR.t0 391.373
R13 VPWR.n4 VPWR.t3 117.721
R14 VPWR.n1 VPWR.t2 54.0554
R15 VPWR.n4 VPWR.t4 49.6583
R16 VPWR.n1 VPWR.t1 47.2559
R17 VPWR.n6 VPWR.n2 34.6358
R18 VPWR.n10 VPWR.n2 34.6358
R19 VPWR.n11 VPWR.n10 34.6358
R20 VPWR.n12 VPWR.n11 16.5652
R21 VPWR.n5 VPWR.n3 15.4623
R22 VPWR.n7 VPWR.n6 9.3005
R23 VPWR.n8 VPWR.n2 9.3005
R24 VPWR.n10 VPWR.n9 9.3005
R25 VPWR.n11 VPWR.n0 9.3005
R26 VPWR.n13 VPWR.n12 7.42022
R27 VPWR.n6 VPWR.n5 1.50638
R28 VPWR.n7 VPWR.n3 0.550633
R29 VPWR.n13 VPWR.n0 0.14471
R30 VPWR.n8 VPWR.n7 0.120292
R31 VPWR.n9 VPWR.n8 0.120292
R32 VPWR.n9 VPWR.n0 0.120292
R33 VPWR VPWR.n13 0.117399
R34 VPB.t2 VPB.t3 642.212
R35 VPB.t3 VPB.t4 509.034
R36 VPB.t1 VPB.t2 346.262
R37 VPB.t4 VPB.t0 254.518
R38 VPB VPB.t1 195.327
R39 a_362_333.t1 a_362_333.n3 427.473
R40 a_362_333.n3 a_362_333.t0 335.214
R41 a_362_333.n0 a_362_333.t5 221.72
R42 a_362_333.n1 a_362_333.t3 221.72
R43 a_362_333.n0 a_362_333.t2 186.374
R44 a_362_333.n1 a_362_333.t4 186.374
R45 a_362_333.n3 a_362_333.n2 167.435
R46 a_362_333.n2 a_362_333.n0 74.9783
R47 a_362_333.n2 a_362_333.n1 1.78569
R48 X X.n0 589.668
R49 X.n3 X.n0 585
R50 X X.n1 189.655
R51 X.n1 X.t3 40.0005
R52 X.n1 X.t0 40.0005
R53 X.n0 X.t1 27.5805
R54 X.n0 X.t2 27.5805
R55 X X.n2 8.0005
R56 X X.n3 7.2005
R57 X.n2 X 2.62614
R58 X.n3 X 1.86717
R59 X.n2 X 1.06717
R60 VGND.n2 VGND.t4 312.063
R61 VGND.n12 VGND.n11 201.292
R62 VGND.n4 VGND.n3 200.516
R63 VGND.n3 VGND.t2 126.858
R64 VGND.n3 VGND.t3 62.8576
R65 VGND.n11 VGND.t0 55.7148
R66 VGND.n11 VGND.t1 51.8906
R67 VGND.n5 VGND.n1 34.6358
R68 VGND.n9 VGND.n1 34.6358
R69 VGND.n10 VGND.n9 34.6358
R70 VGND.n12 VGND.n10 17.6946
R71 VGND.n4 VGND.n2 15.4623
R72 VGND.n6 VGND.n5 9.3005
R73 VGND.n7 VGND.n1 9.3005
R74 VGND.n9 VGND.n8 9.3005
R75 VGND.n10 VGND.n0 9.3005
R76 VGND.n13 VGND.n12 7.37348
R77 VGND.n5 VGND.n4 1.50638
R78 VGND.n6 VGND.n2 0.550633
R79 VGND.n13 VGND.n0 0.145304
R80 VGND.n7 VGND.n6 0.120292
R81 VGND.n8 VGND.n7 0.120292
R82 VGND.n8 VGND.n0 0.120292
R83 VGND VGND.n13 0.116797
R84 VNB.t1 VNB.t2 3089.97
R85 VNB.t2 VNB.t3 2449.19
R86 VNB.t0 VNB.t1 1666.02
R87 VNB.t3 VNB.t4 1224.6
R88 VNB VNB.t0 939.807
R89 a_228_47.t1 a_228_47.n1 384.07
R90 a_228_47.n1 a_228_47.t0 265.829
R91 a_228_47.n0 a_228_47.t2 250.641
R92 a_228_47.n0 a_228_47.t3 149.421
R93 a_228_47.n1 a_228_47.n0 104.15
C0 VPWR VGND 0.09873f
C1 X VGND 0.127998f
C2 VPB A 0.039653f
C3 VPB VPWR 0.100822f
C4 VPB X 0.006105f
C5 A VPWR 0.018453f
C6 VPB VGND 0.010683f
C7 A VGND 0.018096f
C8 VPWR X 0.183274f
C9 VGND VNB 0.517666f
C10 X VNB 0.039216f
C11 VPWR VNB 0.446224f
C12 A VNB 0.177772f
C13 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s15_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s15_1 VGND VPWR X A VPB VNB
X0 VPWR.t0 A.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.346 pd=1.71 as=0.265 ps=2.53 w=1 l=0.15
X1 a_282_47.t1 a_27_47.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.222125 ps=1.36 w=0.65 l=0.15
X2 X.t1 a_394_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.2181 ps=1.36 w=0.42 l=0.15
X3 VGND.t3 a_282_47.t2 a_394_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.2181 pd=1.36 as=0.17225 ps=1.83 w=0.65 l=0.15
X4 X.t0 a_394_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.3406 ps=1.71 w=1 l=0.15
X5 a_282_47.t0 a_27_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2173 pd=2.17 as=0.346 ps=1.71 w=0.82 l=0.15
X6 VGND.t0 A.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.222125 pd=1.36 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 VPWR.t1 a_282_47.t3 a_394_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.3406 pd=1.71 as=0.2173 ps=2.17 w=0.82 l=0.15
R0 A.n0 A.t0 236.18
R1 A.n0 A.t1 206.093
R2 A A.n0 163.852
R3 a_27_47.t1 a_27_47.n1 371.791
R4 a_27_47.n1 a_27_47.t0 273.277
R5 a_27_47.n0 a_27_47.t3 250.641
R6 a_27_47.n1 a_27_47.n0 216.268
R7 a_27_47.n0 a_27_47.t2 139.78
R8 VPWR.n2 VPWR.n1 322.675
R9 VPWR.n2 VPWR.n0 316.846
R10 VPWR.n0 VPWR.t1 112.889
R11 VPWR.n1 VPWR.t2 110.654
R12 VPWR.n0 VPWR.t3 33.5289
R13 VPWR.n1 VPWR.t0 29.5213
R14 VPWR VPWR.n2 0.162202
R15 VPB.t2 VPB.t1 577.104
R16 VPB.t1 VPB.t3 509.034
R17 VPB.t0 VPB.t2 509.034
R18 VPB VPB.t0 195.327
R19 VGND.n2 VGND.n1 206.156
R20 VGND.n2 VGND.n0 205.825
R21 VGND.n1 VGND.t2 95.0774
R22 VGND.n0 VGND.t3 90.462
R23 VGND.n0 VGND.t1 51.7368
R24 VGND.n1 VGND.t0 43.5829
R25 VGND VGND.n2 0.16023
R26 a_282_47.t0 a_282_47.n1 378.688
R27 a_282_47.n0 a_282_47.t3 239.393
R28 a_282_47.n1 a_282_47.t1 154.595
R29 a_282_47.n0 a_282_47.t2 141.387
R30 a_282_47.n1 a_282_47.n0 125.847
R31 VNB.t2 VNB.t3 2776.7
R32 VNB.t3 VNB.t1 2449.19
R33 VNB.t0 VNB.t2 2449.19
R34 VNB VNB.t0 939.807
R35 a_394_47.t0 a_394_47.n1 388.079
R36 a_394_47.n1 a_394_47.t1 341.154
R37 a_394_47.n0 a_394_47.t3 235.304
R38 a_394_47.n0 a_394_47.t2 201.71
R39 a_394_47.n1 a_394_47.n0 152
R40 X X.n0 592.149
R41 X.n2 X.n0 585
R42 X X.t1 226.496
R43 X.n0 X.t0 27.5805
R44 X X.n1 12.244
R45 X.n2 X 7.14855
R46 X.n1 X 6.67876
R47 X X.n2 4.15634
R48 X.n1 X 3.99011
C0 A VPWR 0.019211f
C1 X VGND 0.071815f
C2 X VPB 0.012922f
C3 VGND VPB 0.007419f
C4 VGND A 0.016578f
C5 X VPWR 0.11463f
C6 VPB A 0.038069f
C7 VGND VPWR 0.080247f
C8 VPB VPWR 0.082105f
C9 VGND VNB 0.441721f
C10 X VNB 0.09455f
C11 VPWR VNB 0.363409f
C12 A VNB 0.165238f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR.t15 A.t0 a_110_47.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR.t11 a_110_47.t8 X.t23 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X.t22 a_110_47.t9 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X.t21 a_110_47.t10 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_47.t6 A.t1 VPWR.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 a_110_47.t3 A.t2 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 X.t11 a_110_47.t11 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 a_110_47.t5 A.t3 VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND.t14 A.t4 a_110_47.t2 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND.t10 a_110_47.t12 X.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VPWR.t8 a_110_47.t13 X.t20 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 X.t19 a_110_47.t14 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND.t13 A.t5 a_110_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR.t6 a_110_47.t15 X.t18 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X14 VGND.t9 a_110_47.t16 X.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X.t17 a_110_47.t17 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X16 a_110_47.t0 A.t6 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X17 VPWR.t12 A.t7 a_110_47.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 X.t16 a_110_47.t18 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND.t8 a_110_47.t19 X.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 VGND.t7 a_110_47.t20 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 X.t6 a_110_47.t21 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 X.t15 a_110_47.t22 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 X.t14 a_110_47.t23 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 X.t5 a_110_47.t24 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X25 VPWR.t1 a_110_47.t25 X.t13 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 X.t12 a_110_47.t26 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 X.t4 a_110_47.t27 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 X.t3 a_110_47.t28 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X.t2 a_110_47.t29 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X.t1 a_110_47.t30 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X31 X.t0 a_110_47.t31 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
R0 A.n0 A.t7 184.768
R1 A.n1 A.t3 184.768
R2 A.n2 A.t0 184.768
R3 A.n3 A.t1 184.768
R4 A A.n3 173.609
R5 A.n0 A.t4 146.208
R6 A.n1 A.t2 146.208
R7 A.n2 A.t5 146.208
R8 A.n3 A.t6 146.208
R9 A.n1 A.n0 40.6397
R10 A.n2 A.n1 40.6397
R11 A.n3 A.n2 40.6397
R12 a_110_47.n56 a_110_47.n55 330.308
R13 a_110_47.n58 a_110_47.n57 327.252
R14 a_110_47.n57 a_110_47.n2 217.256
R15 a_110_47.n56 a_110_47.n54 217.256
R16 a_110_47.n18 a_110_47.n16 212.081
R17 a_110_47.n19 a_110_47.t26 212.081
R18 a_110_47.n20 a_110_47.n14 212.081
R19 a_110_47.n22 a_110_47.t14 212.081
R20 a_110_47.n24 a_110_47.n12 212.081
R21 a_110_47.n1 a_110_47.t22 212.081
R22 a_110_47.n29 a_110_47.n9 212.081
R23 a_110_47.n7 a_110_47.t17 212.081
R24 a_110_47.n34 a_110_47.t15 212.081
R25 a_110_47.n0 a_110_47.t10 212.081
R26 a_110_47.n39 a_110_47.t25 212.081
R27 a_110_47.n41 a_110_47.t18 212.081
R28 a_110_47.n42 a_110_47.t13 212.081
R29 a_110_47.n48 a_110_47.t9 212.081
R30 a_110_47.n50 a_110_47.t8 212.081
R31 a_110_47.n51 a_110_47.t23 212.081
R32 a_110_47.n21 a_110_47.n11 169.409
R33 a_110_47.n18 a_110_47.n17 162.274
R34 a_110_47.n19 a_110_47.t21 162.274
R35 a_110_47.n20 a_110_47.n15 162.274
R36 a_110_47.n22 a_110_47.t27 162.274
R37 a_110_47.n24 a_110_47.n13 162.274
R38 a_110_47.n1 a_110_47.t29 162.274
R39 a_110_47.n29 a_110_47.n10 162.274
R40 a_110_47.n7 a_110_47.t31 162.274
R41 a_110_47.n34 a_110_47.t12 162.274
R42 a_110_47.n0 a_110_47.t11 162.274
R43 a_110_47.n39 a_110_47.t16 162.274
R44 a_110_47.n41 a_110_47.t24 162.274
R45 a_110_47.n42 a_110_47.t19 162.274
R46 a_110_47.n48 a_110_47.t28 162.274
R47 a_110_47.n50 a_110_47.t20 162.274
R48 a_110_47.n51 a_110_47.t30 162.274
R49 a_110_47.n53 a_110_47.n52 152
R50 a_110_47.n49 a_110_47.n3 152
R51 a_110_47.n47 a_110_47.n46 152
R52 a_110_47.n45 a_110_47.n4 152
R53 a_110_47.n44 a_110_47.n43 152
R54 a_110_47.n40 a_110_47.n5 152
R55 a_110_47.n38 a_110_47.n37 152
R56 a_110_47.n36 a_110_47.n0 152
R57 a_110_47.n35 a_110_47.n6 152
R58 a_110_47.n33 a_110_47.n32 152
R59 a_110_47.n31 a_110_47.n30 152
R60 a_110_47.n28 a_110_47.n8 152
R61 a_110_47.n1 a_110_47.n27 152
R62 a_110_47.n26 a_110_47.n25 152
R63 a_110_47.n23 a_110_47.n11 152
R64 a_110_47.n19 a_110_47.n18 55.2698
R65 a_110_47.n20 a_110_47.n19 55.2698
R66 a_110_47.n57 a_110_47.n56 44.0325
R67 a_110_47.n25 a_110_47.n1 43.7018
R68 a_110_47.n28 a_110_47.n1 43.7018
R69 a_110_47.n0 a_110_47.n35 43.7018
R70 a_110_47.n47 a_110_47.n4 43.7018
R71 a_110_47.n38 a_110_47.n0 43.7018
R72 a_110_47.n57 a_110_47.n53 43.5205
R73 a_110_47.n2 a_110_47.t2 40.0005
R74 a_110_47.n2 a_110_47.t3 40.0005
R75 a_110_47.n54 a_110_47.t1 40.0005
R76 a_110_47.n54 a_110_47.t0 40.0005
R77 a_110_47.n49 a_110_47.n48 39.8458
R78 a_110_47.n43 a_110_47.n42 35.9898
R79 a_110_47.n21 a_110_47.n20 35.3472
R80 a_110_47.n34 a_110_47.n33 33.4192
R81 a_110_47.n30 a_110_47.n29 32.7765
R82 a_110_47.n24 a_110_47.n23 31.4912
R83 a_110_47.n40 a_110_47.n39 30.8485
R84 a_110_47.n52 a_110_47.n50 28.2778
R85 a_110_47.n55 a_110_47.t7 27.5805
R86 a_110_47.n55 a_110_47.t6 27.5805
R87 a_110_47.t4 a_110_47.n58 27.5805
R88 a_110_47.n58 a_110_47.t5 27.5805
R89 a_110_47.n52 a_110_47.n51 26.9925
R90 a_110_47.n41 a_110_47.n40 24.4218
R91 a_110_47.n23 a_110_47.n22 23.7792
R92 a_110_47.n30 a_110_47.n7 22.4938
R93 a_110_47.n33 a_110_47.n7 21.2085
R94 a_110_47.n22 a_110_47.n21 19.9232
R95 a_110_47.n43 a_110_47.n41 19.2805
R96 a_110_47.n26 a_110_47.n11 17.4085
R97 a_110_47.n27 a_110_47.n26 17.4085
R98 a_110_47.n27 a_110_47.n8 17.4085
R99 a_110_47.n31 a_110_47.n8 17.4085
R100 a_110_47.n32 a_110_47.n31 17.4085
R101 a_110_47.n32 a_110_47.n6 17.4085
R102 a_110_47.n36 a_110_47.n6 17.4085
R103 a_110_47.n37 a_110_47.n36 17.4085
R104 a_110_47.n37 a_110_47.n5 17.4085
R105 a_110_47.n44 a_110_47.n5 17.4085
R106 a_110_47.n45 a_110_47.n44 17.4085
R107 a_110_47.n46 a_110_47.n45 17.4085
R108 a_110_47.n46 a_110_47.n3 17.4085
R109 a_110_47.n53 a_110_47.n3 17.4085
R110 a_110_47.n50 a_110_47.n49 15.4245
R111 a_110_47.n39 a_110_47.n38 12.8538
R112 a_110_47.n25 a_110_47.n24 12.2112
R113 a_110_47.n29 a_110_47.n28 10.9258
R114 a_110_47.n35 a_110_47.n34 10.2832
R115 a_110_47.n42 a_110_47.n4 7.7125
R116 a_110_47.n48 a_110_47.n47 3.8565
R117 VPWR.n14 VPWR.t0 780.891
R118 VPWR.n17 VPWR.t3 776.202
R119 VPWR.n13 VPWR.t7 776.202
R120 VPWR.n11 VPWR.n10 610.861
R121 VPWR.n30 VPWR.n5 609.37
R122 VPWR.n7 VPWR.n6 609.37
R123 VPWR.n23 VPWR.n9 609.37
R124 VPWR.n40 VPWR.t14 340.211
R125 VPWR.n38 VPWR.n2 315.334
R126 VPWR.n32 VPWR.n31 315.089
R127 VPWR.n29 VPWR.n28 33.6462
R128 VPWR.n25 VPWR.n24 33.6462
R129 VPWR.n22 VPWR.n11 33.6462
R130 VPWR.n33 VPWR.n32 30.7205
R131 VPWR.n18 VPWR.n17 29.2576
R132 VPWR.n2 VPWR.t13 27.5805
R133 VPWR.n2 VPWR.t15 27.5805
R134 VPWR.n31 VPWR.t2 27.5805
R135 VPWR.n31 VPWR.t12 27.5805
R136 VPWR.n5 VPWR.t10 27.5805
R137 VPWR.n5 VPWR.t11 27.5805
R138 VPWR.n6 VPWR.t4 27.5805
R139 VPWR.n6 VPWR.t8 27.5805
R140 VPWR.n9 VPWR.t9 27.5805
R141 VPWR.n9 VPWR.t1 27.5805
R142 VPWR.n10 VPWR.t6 27.5805
R143 VPWR.n38 VPWR.n37 27.1064
R144 VPWR.n10 VPWR.t5 26.5955
R145 VPWR.n16 VPWR.n13 24.8691
R146 VPWR.n39 VPWR.n38 22.5887
R147 VPWR.n40 VPWR.n39 22.5887
R148 VPWR.n17 VPWR.n16 20.1148
R149 VPWR.n37 VPWR.n3 18.0711
R150 VPWR.n18 VPWR.n11 15.7262
R151 VPWR.n33 VPWR.n30 13.1662
R152 VPWR.n23 VPWR.n22 10.2405
R153 VPWR.n20 VPWR.n11 9.56172
R154 VPWR.n17 VPWR.n12 9.56172
R155 VPWR.n16 VPWR.n15 9.3005
R156 VPWR.n19 VPWR.n18 9.3005
R157 VPWR.n22 VPWR.n21 9.3005
R158 VPWR.n24 VPWR.n8 9.3005
R159 VPWR.n26 VPWR.n25 9.3005
R160 VPWR.n28 VPWR.n27 9.3005
R161 VPWR.n29 VPWR.n4 9.3005
R162 VPWR.n34 VPWR.n33 9.3005
R163 VPWR.n35 VPWR.n3 9.3005
R164 VPWR.n37 VPWR.n36 9.3005
R165 VPWR.n38 VPWR.n1 9.3005
R166 VPWR.n39 VPWR.n0 9.3005
R167 VPWR.n41 VPWR.n40 9.3005
R168 VPWR.n28 VPWR.n7 8.77764
R169 VPWR.n14 VPWR.n13 6.86786
R170 VPWR.n25 VPWR.n7 5.85193
R171 VPWR.n24 VPWR.n23 4.38907
R172 VPWR.n30 VPWR.n29 1.46336
R173 VPWR.n15 VPWR.n14 0.595283
R174 VPWR.n32 VPWR.n3 0.246654
R175 VPWR.n15 VPWR.n12 0.120292
R176 VPWR.n19 VPWR.n12 0.120292
R177 VPWR.n20 VPWR.n19 0.120292
R178 VPWR.n21 VPWR.n20 0.120292
R179 VPWR.n21 VPWR.n8 0.120292
R180 VPWR.n26 VPWR.n8 0.120292
R181 VPWR.n27 VPWR.n26 0.120292
R182 VPWR.n27 VPWR.n4 0.120292
R183 VPWR.n34 VPWR.n4 0.120292
R184 VPWR.n35 VPWR.n34 0.120292
R185 VPWR.n36 VPWR.n35 0.120292
R186 VPWR.n36 VPWR.n1 0.120292
R187 VPWR.n1 VPWR.n0 0.120292
R188 VPWR.n41 VPWR.n0 0.120292
R189 VPWR VPWR.n41 0.0226354
R190 VPB.t7 VPB.t0 509.034
R191 VPB.t3 VPB.t7 509.034
R192 VPB.t5 VPB.t3 509.034
R193 VPB.t9 VPB.t6 254.518
R194 VPB.t1 VPB.t9 254.518
R195 VPB.t4 VPB.t1 254.518
R196 VPB.t8 VPB.t4 254.518
R197 VPB.t10 VPB.t8 254.518
R198 VPB.t11 VPB.t10 254.518
R199 VPB.t2 VPB.t11 254.518
R200 VPB.t12 VPB.t2 254.518
R201 VPB.t13 VPB.t12 254.518
R202 VPB.t15 VPB.t13 254.518
R203 VPB.t14 VPB.t15 254.518
R204 VPB.t6 VPB.t5 251.559
R205 VPB VPB.t14 145.017
R206 X.n12 X.n10 333.392
R207 X.n19 X.t19 328.971
R208 X.n17 X.t17 328.971
R209 X.n18 X.t15 328.971
R210 X.n20 X.t12 325.442
R211 X.n12 X.n11 301.392
R212 X.n14 X.n13 301.392
R213 X.n16 X.n15 301.392
R214 X.n2 X.n0 248.638
R215 X.n7 X.t0 243.463
R216 X.n8 X.t2 243.463
R217 X.n9 X.t4 243.463
R218 X X.t6 239.607
R219 X.n2 X.n1 203.463
R220 X.n4 X.n3 203.463
R221 X.n6 X.n5 202.456
R222 X.n4 X.n2 45.177
R223 X.n8 X.n7 45.177
R224 X.n9 X.n8 45.177
R225 X.n6 X.n4 44.0476
R226 X.n7 X.n6 44.0476
R227 X.n0 X.t7 40.0005
R228 X.n0 X.t1 40.0005
R229 X.n1 X.t8 40.0005
R230 X.n1 X.t3 40.0005
R231 X.n3 X.t9 40.0005
R232 X.n3 X.t5 40.0005
R233 X.n5 X.t10 40.0005
R234 X.n5 X.t11 40.0005
R235 X.n14 X.n12 32.0005
R236 X.n16 X.n14 32.0005
R237 X.n18 X.n17 32.0005
R238 X.n19 X.n18 32.0005
R239 X.n17 X.n16 31.2005
R240 X.n10 X.t23 27.5805
R241 X.n10 X.t14 27.5805
R242 X.n11 X.t20 27.5805
R243 X.n11 X.t22 27.5805
R244 X.n13 X.t13 27.5805
R245 X.n13 X.t16 27.5805
R246 X.n15 X.t18 27.5805
R247 X.n15 X.t21 27.5805
R248 X.n21 X.n9 13.177
R249 X.n20 X.n19 10.4484
R250 X.n21 X 3.13183
R251 X X.n20 1.75844
R252 X X.n21 0.604792
R253 VGND.n10 VGND.t6 250.282
R254 VGND.n9 VGND.t4 245.481
R255 VGND.n13 VGND.t2 245.481
R256 VGND.n39 VGND.t12 240.948
R257 VGND.n33 VGND.n32 206.909
R258 VGND.n37 VGND.n2 206.909
R259 VGND.n7 VGND.n6 205.899
R260 VGND.n20 VGND.n19 205.899
R261 VGND.n23 VGND.n22 204.692
R262 VGND.n30 VGND.n29 204.692
R263 VGND.n6 VGND.t10 40.0005
R264 VGND.n19 VGND.t11 40.0005
R265 VGND.n19 VGND.t9 40.0005
R266 VGND.n22 VGND.t5 40.0005
R267 VGND.n22 VGND.t8 40.0005
R268 VGND.n29 VGND.t3 40.0005
R269 VGND.n29 VGND.t7 40.0005
R270 VGND.n32 VGND.t1 40.0005
R271 VGND.n32 VGND.t14 40.0005
R272 VGND.n2 VGND.t15 40.0005
R273 VGND.n2 VGND.t13 40.0005
R274 VGND.n6 VGND.t0 38.5719
R275 VGND.n18 VGND.n7 34.6358
R276 VGND.n24 VGND.n21 34.6358
R277 VGND.n28 VGND.n4 34.6358
R278 VGND.n33 VGND.n31 31.624
R279 VGND.n14 VGND.n13 29.7417
R280 VGND.n37 VGND.n1 27.1064
R281 VGND.n12 VGND.n9 25.224
R282 VGND.n38 VGND.n37 22.5887
R283 VGND.n39 VGND.n38 22.5887
R284 VGND.n13 VGND.n12 20.7064
R285 VGND.n33 VGND.n1 18.0711
R286 VGND.n14 VGND.n7 16.1887
R287 VGND.n31 VGND.n30 13.5534
R288 VGND.n20 VGND.n18 11.6711
R289 VGND.n40 VGND.n39 9.3005
R290 VGND.n12 VGND.n11 9.3005
R291 VGND.n13 VGND.n8 9.3005
R292 VGND.n15 VGND.n14 9.3005
R293 VGND.n16 VGND.n7 9.3005
R294 VGND.n18 VGND.n17 9.3005
R295 VGND.n21 VGND.n5 9.3005
R296 VGND.n25 VGND.n24 9.3005
R297 VGND.n26 VGND.n4 9.3005
R298 VGND.n28 VGND.n27 9.3005
R299 VGND.n31 VGND.n3 9.3005
R300 VGND.n34 VGND.n33 9.3005
R301 VGND.n35 VGND.n1 9.3005
R302 VGND.n37 VGND.n36 9.3005
R303 VGND.n38 VGND.n0 9.3005
R304 VGND.n23 VGND.n4 9.03579
R305 VGND.n10 VGND.n9 6.78128
R306 VGND.n24 VGND.n23 6.02403
R307 VGND.n21 VGND.n20 4.51815
R308 VGND.n30 VGND.n28 1.50638
R309 VGND.n11 VGND.n10 0.56336
R310 VGND.n11 VGND.n8 0.120292
R311 VGND.n15 VGND.n8 0.120292
R312 VGND.n16 VGND.n15 0.120292
R313 VGND.n17 VGND.n16 0.120292
R314 VGND.n17 VGND.n5 0.120292
R315 VGND.n25 VGND.n5 0.120292
R316 VGND.n26 VGND.n25 0.120292
R317 VGND.n27 VGND.n26 0.120292
R318 VGND.n27 VGND.n3 0.120292
R319 VGND.n34 VGND.n3 0.120292
R320 VGND.n35 VGND.n34 0.120292
R321 VGND.n36 VGND.n35 0.120292
R322 VGND.n36 VGND.n0 0.120292
R323 VGND.n40 VGND.n0 0.120292
R324 VGND VGND.n40 0.0226354
R325 VNB.t4 VNB.t6 2449.19
R326 VNB.t2 VNB.t4 2449.19
R327 VNB.t0 VNB.t2 2449.19
R328 VNB.t11 VNB.t10 1224.6
R329 VNB.t9 VNB.t11 1224.6
R330 VNB.t5 VNB.t9 1224.6
R331 VNB.t8 VNB.t5 1224.6
R332 VNB.t3 VNB.t8 1224.6
R333 VNB.t7 VNB.t3 1224.6
R334 VNB.t1 VNB.t7 1224.6
R335 VNB.t14 VNB.t1 1224.6
R336 VNB.t15 VNB.t14 1224.6
R337 VNB.t13 VNB.t15 1224.6
R338 VNB.t12 VNB.t13 1224.6
R339 VNB.t10 VNB.t0 1210.36
R340 VNB VNB.t12 697.736
C0 A VGND 0.115353f
C1 VPWR X 1.36494f
C2 VPWR VGND 0.187357f
C3 X VGND 0.976879f
C4 VPB A 0.133397f
C5 VPB VPWR 0.183858f
C6 A VPWR 0.111641f
C7 VPB X 0.03148f
C8 VPB VGND 0.011388f
C9 A X 0.002918f
C10 VGND VNB 1.01442f
C11 X VNB 0.110579f
C12 VPWR VNB 0.834786f
C13 A VNB 0.494734f
C14 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_8 X A VPB VNB VGND VPWR
X0 VPWR.t1 A.t0 a_110_47.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR.t9 a_110_47.t4 X.t15 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X.t14 a_110_47.t5 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47.t2 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X.t4 a_110_47.t6 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X.t13 a_110_47.t7 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND.t8 a_110_47.t8 X.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR.t6 a_110_47.t9 X.t12 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND.t1 A.t2 a_110_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND.t7 a_110_47.t10 X.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47.t1 A.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR.t5 a_110_47.t11 X.t11 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X.t10 a_110_47.t12 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND.t6 a_110_47.t13 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND.t5 a_110_47.t14 X.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X.t9 a_110_47.t15 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X.t7 a_110_47.t16 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR.t2 a_110_47.t17 X.t8 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X.t6 a_110_47.t18 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X.t5 a_110_47.t19 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A.n0 A.t0 184.768
R1 A.n1 A.t1 184.768
R2 A A.n1 173.609
R3 A.n0 A.t2 146.208
R4 A.n1 A.t3 146.208
R5 A.n1 A.n0 40.6397
R6 a_110_47.n21 a_110_47.n20 316.591
R7 a_110_47.n20 a_110_47.n0 217.256
R8 a_110_47.n3 a_110_47.t17 212.081
R9 a_110_47.n4 a_110_47.t12 212.081
R10 a_110_47.n5 a_110_47.t9 212.081
R11 a_110_47.n7 a_110_47.t5 212.081
R12 a_110_47.n8 a_110_47.t4 212.081
R13 a_110_47.n14 a_110_47.t15 212.081
R14 a_110_47.n16 a_110_47.t11 212.081
R15 a_110_47.n17 a_110_47.t7 212.081
R16 a_110_47.n10 a_110_47.n6 169.409
R17 a_110_47.n3 a_110_47.t10 162.274
R18 a_110_47.n4 a_110_47.t16 162.274
R19 a_110_47.n5 a_110_47.t13 162.274
R20 a_110_47.n7 a_110_47.t18 162.274
R21 a_110_47.n8 a_110_47.t14 162.274
R22 a_110_47.n14 a_110_47.t19 162.274
R23 a_110_47.n16 a_110_47.t8 162.274
R24 a_110_47.n17 a_110_47.t6 162.274
R25 a_110_47.n19 a_110_47.n18 152
R26 a_110_47.n15 a_110_47.n1 152
R27 a_110_47.n13 a_110_47.n12 152
R28 a_110_47.n11 a_110_47.n2 152
R29 a_110_47.n10 a_110_47.n9 152
R30 a_110_47.n4 a_110_47.n3 55.2698
R31 a_110_47.n5 a_110_47.n4 55.2698
R32 a_110_47.n13 a_110_47.n2 43.7018
R33 a_110_47.n20 a_110_47.n19 43.5205
R34 a_110_47.n0 a_110_47.t0 40.0005
R35 a_110_47.n0 a_110_47.t1 40.0005
R36 a_110_47.n15 a_110_47.n14 39.8458
R37 a_110_47.n9 a_110_47.n8 35.9898
R38 a_110_47.n6 a_110_47.n5 30.8485
R39 a_110_47.n18 a_110_47.n16 28.2778
R40 a_110_47.n21 a_110_47.t3 27.5805
R41 a_110_47.t2 a_110_47.n21 27.5805
R42 a_110_47.n18 a_110_47.n17 26.9925
R43 a_110_47.n7 a_110_47.n6 24.4218
R44 a_110_47.n9 a_110_47.n7 19.2805
R45 a_110_47.n11 a_110_47.n10 17.4085
R46 a_110_47.n12 a_110_47.n11 17.4085
R47 a_110_47.n12 a_110_47.n1 17.4085
R48 a_110_47.n19 a_110_47.n1 17.4085
R49 a_110_47.n16 a_110_47.n15 15.4245
R50 a_110_47.n8 a_110_47.n2 7.7125
R51 a_110_47.n14 a_110_47.n13 3.8565
R52 VPWR.n9 VPWR.t2 787.674
R53 VPWR.n4 VPWR.n3 609.615
R54 VPWR.n13 VPWR.n6 609.615
R55 VPWR.n8 VPWR.n7 609.615
R56 VPWR.n21 VPWR.t0 350.705
R57 VPWR.n19 VPWR.n2 327.238
R58 VPWR.n12 VPWR.n11 34.6358
R59 VPWR.n14 VPWR.n4 31.624
R60 VPWR.n2 VPWR.t7 27.5805
R61 VPWR.n2 VPWR.t1 27.5805
R62 VPWR.n3 VPWR.t3 27.5805
R63 VPWR.n3 VPWR.t5 27.5805
R64 VPWR.n6 VPWR.t8 27.5805
R65 VPWR.n6 VPWR.t9 27.5805
R66 VPWR.n7 VPWR.t4 27.5805
R67 VPWR.n7 VPWR.t6 27.5805
R68 VPWR.n19 VPWR.n18 27.1064
R69 VPWR.n20 VPWR.n19 22.5887
R70 VPWR.n21 VPWR.n20 22.5887
R71 VPWR.n18 VPWR.n4 18.0711
R72 VPWR.n14 VPWR.n13 13.5534
R73 VPWR.n9 VPWR.n8 12.6411
R74 VPWR.n11 VPWR.n10 9.3005
R75 VPWR.n12 VPWR.n5 9.3005
R76 VPWR.n15 VPWR.n14 9.3005
R77 VPWR.n16 VPWR.n4 9.3005
R78 VPWR.n18 VPWR.n17 9.3005
R79 VPWR.n19 VPWR.n1 9.3005
R80 VPWR.n20 VPWR.n0 9.3005
R81 VPWR.n22 VPWR.n21 9.3005
R82 VPWR.n11 VPWR.n8 9.03579
R83 VPWR.n13 VPWR.n12 1.50638
R84 VPWR.n10 VPWR.n9 1.09422
R85 VPWR.n10 VPWR.n5 0.120292
R86 VPWR.n15 VPWR.n5 0.120292
R87 VPWR.n16 VPWR.n15 0.120292
R88 VPWR.n17 VPWR.n16 0.120292
R89 VPWR.n17 VPWR.n1 0.120292
R90 VPWR.n1 VPWR.n0 0.120292
R91 VPWR.n22 VPWR.n0 0.120292
R92 VPWR VPWR.n22 0.0226354
R93 VPB.t4 VPB.t2 254.518
R94 VPB.t6 VPB.t4 254.518
R95 VPB.t8 VPB.t6 254.518
R96 VPB.t9 VPB.t8 254.518
R97 VPB.t3 VPB.t9 254.518
R98 VPB.t5 VPB.t3 254.518
R99 VPB.t7 VPB.t5 254.518
R100 VPB.t1 VPB.t7 254.518
R101 VPB.t0 VPB.t1 254.518
R102 VPB VPB.t0 195.327
R103 X.n7 X.n5 333.392
R104 X.n7 X.n6 301.392
R105 X.n9 X.n8 301.392
R106 X.n11 X.n10 298.296
R107 X.n2 X.n0 248.638
R108 X.n2 X.n1 203.463
R109 X.n4 X.n3 203.463
R110 X X.n13 199.673
R111 X.n4 X.n2 45.177
R112 X.n0 X.t3 40.0005
R113 X.n0 X.t4 40.0005
R114 X.n1 X.t0 40.0005
R115 X.n1 X.t5 40.0005
R116 X.n3 X.t1 40.0005
R117 X.n3 X.t6 40.0005
R118 X.n13 X.t2 40.0005
R119 X.n13 X.t7 40.0005
R120 X.n9 X.n7 32.0005
R121 X.n5 X.t11 27.5805
R122 X.n5 X.t13 27.5805
R123 X.n6 X.t15 27.5805
R124 X.n6 X.t9 27.5805
R125 X.n8 X.t12 27.5805
R126 X.n8 X.t14 27.5805
R127 X.n10 X.t8 27.5805
R128 X.n10 X.t10 27.5805
R129 X.n12 X.n4 27.1064
R130 X.n11 X.n9 19.2005
R131 X.n12 X 3.76132
R132 X X.n11 2.2438
R133 X X.n12 0.726273
R134 VGND.n7 VGND.t7 249.72
R135 VGND.n21 VGND.t0 244.853
R136 VGND.n19 VGND.n2 206.909
R137 VGND.n6 VGND.n5 204.692
R138 VGND.n12 VGND.n11 204.692
R139 VGND.n15 VGND.n14 204.692
R140 VGND.n5 VGND.t4 40.0005
R141 VGND.n5 VGND.t6 40.0005
R142 VGND.n11 VGND.t3 40.0005
R143 VGND.n11 VGND.t5 40.0005
R144 VGND.n14 VGND.t2 40.0005
R145 VGND.n14 VGND.t8 40.0005
R146 VGND.n2 VGND.t9 40.0005
R147 VGND.n2 VGND.t1 40.0005
R148 VGND.n10 VGND.n4 34.6358
R149 VGND.n15 VGND.n13 31.624
R150 VGND.n19 VGND.n1 27.1064
R151 VGND.n20 VGND.n19 22.5887
R152 VGND.n21 VGND.n20 22.5887
R153 VGND.n15 VGND.n1 18.0711
R154 VGND.n13 VGND.n12 13.5534
R155 VGND.n7 VGND.n6 12.6486
R156 VGND.n22 VGND.n21 9.3005
R157 VGND.n8 VGND.n4 9.3005
R158 VGND.n10 VGND.n9 9.3005
R159 VGND.n13 VGND.n3 9.3005
R160 VGND.n16 VGND.n15 9.3005
R161 VGND.n17 VGND.n1 9.3005
R162 VGND.n19 VGND.n18 9.3005
R163 VGND.n20 VGND.n0 9.3005
R164 VGND.n6 VGND.n4 9.03579
R165 VGND.n12 VGND.n10 1.50638
R166 VGND.n8 VGND.n7 1.08558
R167 VGND.n9 VGND.n8 0.120292
R168 VGND.n9 VGND.n3 0.120292
R169 VGND.n16 VGND.n3 0.120292
R170 VGND.n17 VGND.n16 0.120292
R171 VGND.n18 VGND.n17 0.120292
R172 VGND.n18 VGND.n0 0.120292
R173 VGND.n22 VGND.n0 0.120292
R174 VGND VGND.n22 0.0226354
R175 VNB.t4 VNB.t7 1224.6
R176 VNB.t6 VNB.t4 1224.6
R177 VNB.t3 VNB.t6 1224.6
R178 VNB.t5 VNB.t3 1224.6
R179 VNB.t2 VNB.t5 1224.6
R180 VNB.t8 VNB.t2 1224.6
R181 VNB.t9 VNB.t8 1224.6
R182 VNB.t1 VNB.t9 1224.6
R183 VNB.t0 VNB.t1 1224.6
R184 VNB VNB.t0 939.807
C0 VPWR VGND 0.106233f
C1 X VGND 0.492094f
C2 VPB A 0.070741f
C3 VPB VPWR 0.11643f
C4 A VPWR 0.081114f
C5 VPB X 0.022318f
C6 VPB VGND 0.00944f
C7 A X 0.001679f
C8 A VGND 0.069477f
C9 VPWR X 0.71159f
C10 VGND VNB 0.607928f
C11 X VNB 0.081251f
C12 VPWR VNB 0.526748f
C13 A VNB 0.28981f
C14 VPB VNB 1.04774f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR.t4 A.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND.t3 a_27_47.t2 X.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND.t2 a_27_47.t3 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X.t7 a_27_47.t4 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X.t2 a_27_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND.t4 A.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR.t1 a_27_47.t6 X.t6 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X.t3 a_27_47.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X.t5 a_27_47.t8 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR.t3 a_27_47.t9 X.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n0 A.t0 238.59
R1 A.n0 A.t1 203.244
R2 A A.n0 154.012
R3 a_27_47.t0 a_27_47.n9 416.464
R4 a_27_47.n9 a_27_47.t1 304.067
R5 a_27_47.n6 a_27_47.t8 223.19
R6 a_27_47.n3 a_27_47.t6 221.72
R7 a_27_47.n0 a_27_47.t4 221.72
R8 a_27_47.n1 a_27_47.t9 221.72
R9 a_27_47.n3 a_27_47.t2 185.38
R10 a_27_47.n6 a_27_47.t7 184.768
R11 a_27_47.n1 a_27_47.t3 184.768
R12 a_27_47.n0 a_27_47.t5 184.768
R13 a_27_47.n4 a_27_47.n2 177.601
R14 a_27_47.n8 a_27_47.n7 152
R15 a_27_47.n5 a_27_47.n2 152
R16 a_27_47.n9 a_27_47.n8 82.4476
R17 a_27_47.n4 a_27_47.n3 56.9641
R18 a_27_47.n7 a_27_47.n6 49.0769
R19 a_27_47.n5 a_27_47.n0 41.1896
R20 a_27_47.n1 a_27_47.n5 33.3023
R21 a_27_47.n7 a_27_47.n1 26.2914
R22 a_27_47.n8 a_27_47.n2 25.6005
R23 a_27_47.n0 a_27_47.n4 18.4041
R24 VPWR.n4 VPWR.n3 604.076
R25 VPWR.n2 VPWR.t1 350.644
R26 VPWR.n6 VPWR.n1 311.659
R27 VPWR.n1 VPWR.t0 37.4305
R28 VPWR.n1 VPWR.t4 27.5805
R29 VPWR.n3 VPWR.t2 27.5805
R30 VPWR.n3 VPWR.t3 27.5805
R31 VPWR.n5 VPWR.n4 24.4711
R32 VPWR.n6 VPWR.n5 20.7064
R33 VPWR.n5 VPWR.n0 9.3005
R34 VPWR.n7 VPWR.n6 7.30743
R35 VPWR.n4 VPWR.n2 6.71867
R36 VPWR.n2 VPWR.n0 0.647964
R37 VPWR.n7 VPWR.n0 0.146144
R38 VPWR VPWR.n7 0.117248
R39 VPB.t4 VPB.t1 284.113
R40 VPB.t3 VPB.t2 254.518
R41 VPB.t0 VPB.t3 254.518
R42 VPB.t1 VPB.t0 254.518
R43 VPB VPB.t4 195.327
R44 X.n5 X.n3 647.148
R45 X.n2 X.n0 243.627
R46 X.n2 X.n1 200.262
R47 X.n5 X.n4 194.441
R48 X.n0 X.t1 40.0005
R49 X.n0 X.t3 40.0005
R50 X.n1 X.t0 40.0005
R51 X.n1 X.t2 40.0005
R52 X.n4 X.t6 27.5805
R53 X.n4 X.t7 27.5805
R54 X.n3 X.t4 27.5805
R55 X.n3 X.t5 27.5805
R56 X X.n6 19.2609
R57 X.n6 X.n5 15.5262
R58 X.n7 X 9.00791
R59 X.n7 X.n2 6.77697
R60 X.n6 X 2.70819
R61 X X.n7 1.73877
R62 VGND.n1 VGND.t3 249.87
R63 VGND.n3 VGND.n2 205.078
R64 VGND.n6 VGND.n5 203.619
R65 VGND.n5 VGND.t0 55.7148
R66 VGND.n2 VGND.t1 40.0005
R67 VGND.n2 VGND.t2 40.0005
R68 VGND.n5 VGND.t4 40.0005
R69 VGND.n4 VGND.n3 24.4711
R70 VGND.n6 VGND.n4 24.0946
R71 VGND.n4 VGND.n0 9.3005
R72 VGND.n7 VGND.n6 7.27268
R73 VGND.n3 VGND.n1 6.71867
R74 VGND.n1 VGND.n0 0.647964
R75 VGND.n7 VGND.n0 0.146586
R76 VGND VGND.n7 0.116801
R77 VNB.t4 VNB.t0 1381.23
R78 VNB.t1 VNB.t3 1224.6
R79 VNB.t2 VNB.t1 1224.6
R80 VNB.t0 VNB.t2 1224.6
R81 VNB VNB.t4 939.807
C0 VPB A 0.032139f
C1 VPB VPWR 0.063172f
C2 A VPWR 0.021953f
C3 VPB X 0.012159f
C4 VPB VGND 0.005825f
C5 A X 0.013951f
C6 A VGND 0.043094f
C7 VPWR X 0.316967f
C8 VPWR VGND 0.057043f
C9 X VGND 0.21559f
C10 VGND VNB 0.357713f
C11 X VNB 0.067008f
C12 VPWR VNB 0.307647f
C13 A VNB 0.147639f
C14 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR.t2 a_27_47.t2 X.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X.t1 a_27_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X.t0 a_27_47.t4 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND.t1 a_27_47.t5 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 A.n0 A.t0 224.984
R1 A.n0 A.t1 187.714
R2 A A.n0 153.957
R3 a_27_47.t0 a_27_47.n3 403.579
R4 a_27_47.n3 a_27_47.t1 305.671
R5 a_27_47.n3 a_27_47.n2 219.434
R6 a_27_47.n0 a_27_47.t3 189.588
R7 a_27_47.n0 a_27_47.t2 189.588
R8 a_27_47.n1 a_27_47.t5 96.4005
R9 a_27_47.n1 a_27_47.t4 96.4005
R10 a_27_47.n2 a_27_47.n1 35.0935
R11 a_27_47.n2 a_27_47.n0 19.8724
R12 VPWR.n1 VPWR.t2 842.768
R13 VPWR.n1 VPWR.n0 318.115
R14 VPWR.n0 VPWR.t1 36.4455
R15 VPWR.n0 VPWR.t0 27.5805
R16 VPWR VPWR.n1 0.565825
R17 VPB.t0 VPB.t1 281.154
R18 VPB.t1 VPB.t2 248.599
R19 VPB VPB.t0 195.327
R20 X X.n0 623.909
R21 X X.n1 216.464
R22 X.n1 X.t3 38.5719
R23 X.n1 X.t0 38.5719
R24 X.n0 X.t2 26.5955
R25 X.n0 X.t1 26.5955
R26 VGND.n1 VGND.t1 245.523
R27 VGND.n1 VGND.n0 209.065
R28 VGND.n0 VGND.t2 52.8576
R29 VGND.n0 VGND.t0 40.0005
R30 VGND VGND.n1 0.549826
R31 VNB.t0 VNB.t2 1352.75
R32 VNB.t2 VNB.t1 1196.12
R33 VNB VNB.t0 939.807
C0 VPB A 0.033457f
C1 VPB VPWR 0.043784f
C2 A VPWR 0.021971f
C3 VPB X 0.008368f
C4 VPB VGND 0.00461f
C5 A X 0.012264f
C6 A VGND 0.045291f
C7 VPWR X 0.139126f
C8 VPWR VGND 0.038085f
C9 X VGND 0.11464f
C10 VGND VNB 0.262974f
C11 X VNB 0.07314f
C12 VPWR VNB 0.220607f
C13 A VNB 0.147598f
C14 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR.t1 a_75_212.t2 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212.t1 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND.t1 a_75_212.t3 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
R0 a_75_212.t0 a_75_212.n1 407.228
R1 a_75_212.n1 a_75_212.t1 294.341
R2 a_75_212.n0 a_75_212.t2 254.389
R3 a_75_212.n0 a_75_212.t3 211.01
R4 a_75_212.n1 a_75_212.n0 152
R5 X.n1 X.t1 368.521
R6 X.n0 X.t0 216.155
R7 X X.n0 82.2255
R8 X.n1 X 10.5563
R9 X X.n1 5.48477
R10 X.n0 X 5.16973
R11 VPWR VPWR.n0 317.971
R12 VPWR.n0 VPWR.t0 36.1587
R13 VPWR.n0 VPWR.t1 36.1587
R14 VPB.t0 VPB.t1 260.437
R15 VPB VPB.t0 91.745
R16 A.n0 A.t1 260.322
R17 A.n0 A.t0 175.169
R18 A A.n0 154.133
R19 VGND VGND.n0 205.657
R20 VGND.n0 VGND.t0 33.462
R21 VGND.n0 VGND.t1 33.462
R22 VNB.t0 VNB.t1 1253.07
R23 VNB VNB.t0 441.425
C0 A VPWR 0.021742f
C1 X VPWR 0.089604f
C2 VPB VGND 0.005071f
C3 A VGND 0.018424f
C4 X VGND 0.054484f
C5 VPWR VGND 0.028869f
C6 VPB A 0.052491f
C7 VPB X 0.012788f
C8 A X 8.48e-19
C9 VPB VPWR 0.035518f
C10 VGND VNB 0.20733f
C11 VPWR VNB 0.175531f
C12 X VNB 0.094159f
C13 A VNB 0.164205f
C14 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufinv_16 VNB VPB VGND VPWR A Y
X0 a_361_47.t7 a_27_47.t6 VGND.t21 VNB.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR.t18 a_361_47.t12 Y.t15 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_361_47.t6 a_27_47.t7 VGND.t20 VNB.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y.t31 a_361_47.t13 VGND.t22 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t17 a_361_47.t14 Y.t14 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t30 a_361_47.t15 VGND.t23 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t13 a_361_47.t16 VPWR.t16 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t24 a_27_47.t8 a_361_47.t11 VPB.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t15 a_361_47.t17 Y.t12 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR.t14 a_361_47.t18 Y.t11 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t24 a_361_47.t19 Y.t29 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_361_47.t10 a_27_47.t9 VPWR.t23 VPB.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t0 a_361_47.t20 Y.t28 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t1 a_361_47.t21 Y.t27 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t2 a_361_47.t22 Y.t26 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t3 a_361_47.t23 Y.t25 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y.t10 a_361_47.t24 VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND.t4 a_361_47.t25 Y.t24 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR.t12 a_361_47.t26 Y.t9 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_27_47.t1 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 Y.t8 a_361_47.t27 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_27_47.t2 A.t2 VGND.t13 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_361_47.t5 a_27_47.t10 VGND.t19 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 Y.t7 a_361_47.t28 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t23 a_361_47.t29 VGND.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t22 a_27_47.t11 a_361_47.t9 VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t22 a_361_47.t30 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y.t6 a_361_47.t31 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y.t21 a_361_47.t32 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_361_47.t8 a_27_47.t12 VPWR.t21 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VPWR.t8 a_361_47.t33 Y.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 Y.t20 a_361_47.t34 VGND.t8 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t14 A.t3 a_27_47.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 VGND.t18 a_27_47.t13 a_361_47.t4 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 VPWR.t20 a_27_47.t14 a_361_47.t1 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y.t4 a_361_47.t35 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VGND.t17 a_27_47.t15 a_361_47.t3 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 VGND.t16 a_27_47.t16 a_361_47.t2 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_361_47.t0 a_27_47.t17 VPWR.t19 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X40 VPWR.t6 a_361_47.t36 Y.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR.t5 a_361_47.t37 Y.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X42 VGND.t9 a_361_47.t38 Y.t19 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 VGND.t10 a_361_47.t39 Y.t18 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X44 VPWR.t2 A.t4 a_27_47.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X45 Y.t1 a_361_47.t40 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 Y.t17 a_361_47.t41 VGND.t11 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 Y.t0 a_361_47.t42 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 VGND.t15 A.t5 a_27_47.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X49 Y.t16 a_361_47.t43 VGND.t12 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_27_47.n20 a_27_47.t4 271.051
R1 a_27_47.n5 a_27_47.t11 221.72
R2 a_27_47.n7 a_27_47.t12 221.72
R3 a_27_47.n9 a_27_47.t14 221.72
R4 a_27_47.n3 a_27_47.t17 221.72
R5 a_27_47.n15 a_27_47.t8 221.72
R6 a_27_47.n16 a_27_47.t9 221.72
R7 a_27_47.n21 a_27_47.n20 206.055
R8 a_27_47.n1 a_27_47.t5 176.525
R9 a_27_47.n6 a_27_47.n4 173.761
R10 a_27_47.n18 a_27_47.n17 152
R11 a_27_47.n14 a_27_47.n2 152
R12 a_27_47.n13 a_27_47.n12 152
R13 a_27_47.n11 a_27_47.n10 152
R14 a_27_47.n8 a_27_47.n4 152
R15 a_27_47.n5 a_27_47.t16 149.421
R16 a_27_47.n7 a_27_47.t7 149.421
R17 a_27_47.n9 a_27_47.t15 149.421
R18 a_27_47.n3 a_27_47.t6 149.421
R19 a_27_47.n15 a_27_47.t13 149.421
R20 a_27_47.n16 a_27_47.t10 149.421
R21 a_27_47.n1 a_27_47.n0 98.788
R22 a_27_47.n14 a_27_47.n13 60.6968
R23 a_27_47.n10 a_27_47.n3 55.3412
R24 a_27_47.n17 a_27_47.n15 51.7709
R25 a_27_47.n6 a_27_47.n5 48.2005
R26 a_27_47.n9 a_27_47.n8 41.0598
R27 a_27_47.n8 a_27_47.n7 33.919
R28 a_27_47.n19 a_27_47.n1 32.0005
R29 a_27_47.n20 a_27_47.n19 32.0005
R30 a_27_47.n7 a_27_47.n6 26.7783
R31 a_27_47.t0 a_27_47.n21 26.5955
R32 a_27_47.n21 a_27_47.t1 26.5955
R33 a_27_47.n0 a_27_47.t3 24.9236
R34 a_27_47.n0 a_27_47.t2 24.9236
R35 a_27_47.n17 a_27_47.n16 23.2079
R36 a_27_47.n11 a_27_47.n4 21.7605
R37 a_27_47.n12 a_27_47.n11 21.7605
R38 a_27_47.n12 a_27_47.n2 21.7605
R39 a_27_47.n18 a_27_47.n2 21.7605
R40 a_27_47.n19 a_27_47.n18 21.7605
R41 a_27_47.n10 a_27_47.n9 19.6375
R42 a_27_47.n15 a_27_47.n14 8.92643
R43 a_27_47.n13 a_27_47.n3 5.35606
R44 VGND.n22 VGND.t24 290.193
R45 VGND.n21 VGND.n20 208.719
R46 VGND.n26 VGND.n18 208.719
R47 VGND.n29 VGND.n28 208.719
R48 VGND.n35 VGND.n15 208.719
R49 VGND.n13 VGND.n12 208.719
R50 VGND.n42 VGND.n11 208.719
R51 VGND.n44 VGND.n43 208.719
R52 VGND.n50 VGND.n8 208.719
R53 VGND.n53 VGND.n52 208.719
R54 VGND.n59 VGND.n5 208.719
R55 VGND.n3 VGND.n2 208.719
R56 VGND.n66 VGND.n1 208.719
R57 VGND.n67 VGND.n66 43.1829
R58 VGND.n22 VGND.n21 37.7583
R59 VGND.n25 VGND.n19 34.6358
R60 VGND.n30 VGND.n27 34.6358
R61 VGND.n34 VGND.n16 34.6358
R62 VGND.n37 VGND.n36 34.6358
R63 VGND.n41 VGND.n40 34.6358
R64 VGND.n49 VGND.n9 34.6358
R65 VGND.n54 VGND.n51 34.6358
R66 VGND.n58 VGND.n6 34.6358
R67 VGND.n61 VGND.n60 34.6358
R68 VGND.n65 VGND.n64 34.6358
R69 VGND.n45 VGND.n42 32.377
R70 VGND.n45 VGND.n44 30.8711
R71 VGND.n64 VGND.n3 27.8593
R72 VGND.n26 VGND.n25 26.3534
R73 VGND.n40 VGND.n13 26.3534
R74 VGND.n20 VGND.t11 24.9236
R75 VGND.n20 VGND.t10 24.9236
R76 VGND.n18 VGND.t8 24.9236
R77 VGND.n18 VGND.t9 24.9236
R78 VGND.n28 VGND.t7 24.9236
R79 VGND.n28 VGND.t4 24.9236
R80 VGND.n15 VGND.t6 24.9236
R81 VGND.n15 VGND.t3 24.9236
R82 VGND.n12 VGND.t5 24.9236
R83 VGND.n12 VGND.t1 24.9236
R84 VGND.n11 VGND.t22 24.9236
R85 VGND.n11 VGND.t0 24.9236
R86 VGND.n43 VGND.t12 24.9236
R87 VGND.n43 VGND.t2 24.9236
R88 VGND.n8 VGND.t23 24.9236
R89 VGND.n8 VGND.t16 24.9236
R90 VGND.n52 VGND.t20 24.9236
R91 VGND.n52 VGND.t17 24.9236
R92 VGND.n5 VGND.t21 24.9236
R93 VGND.n5 VGND.t18 24.9236
R94 VGND.n2 VGND.t19 24.9236
R95 VGND.n2 VGND.t14 24.9236
R96 VGND.n1 VGND.t13 24.9236
R97 VGND.n1 VGND.t15 24.9236
R98 VGND.n50 VGND.n49 24.8476
R99 VGND.n60 VGND.n59 21.8358
R100 VGND.n30 VGND.n29 20.3299
R101 VGND.n36 VGND.n35 20.3299
R102 VGND.n54 VGND.n53 18.824
R103 VGND.n53 VGND.n6 15.8123
R104 VGND.n29 VGND.n16 14.3064
R105 VGND.n35 VGND.n34 14.3064
R106 VGND.n59 VGND.n58 12.8005
R107 VGND.n51 VGND.n50 9.78874
R108 VGND.n23 VGND.n19 9.3005
R109 VGND.n25 VGND.n24 9.3005
R110 VGND.n27 VGND.n17 9.3005
R111 VGND.n31 VGND.n30 9.3005
R112 VGND.n32 VGND.n16 9.3005
R113 VGND.n34 VGND.n33 9.3005
R114 VGND.n36 VGND.n14 9.3005
R115 VGND.n38 VGND.n37 9.3005
R116 VGND.n40 VGND.n39 9.3005
R117 VGND.n41 VGND.n10 9.3005
R118 VGND.n46 VGND.n45 9.3005
R119 VGND.n47 VGND.n9 9.3005
R120 VGND.n49 VGND.n48 9.3005
R121 VGND.n51 VGND.n7 9.3005
R122 VGND.n55 VGND.n54 9.3005
R123 VGND.n56 VGND.n6 9.3005
R124 VGND.n58 VGND.n57 9.3005
R125 VGND.n60 VGND.n4 9.3005
R126 VGND.n62 VGND.n61 9.3005
R127 VGND.n64 VGND.n63 9.3005
R128 VGND.n65 VGND.n0 9.3005
R129 VGND.n27 VGND.n26 8.28285
R130 VGND.n37 VGND.n13 8.28285
R131 VGND.n61 VGND.n3 6.77697
R132 VGND.n44 VGND.n9 3.76521
R133 VGND.n23 VGND.n22 2.4189
R134 VGND.n21 VGND.n19 2.25932
R135 VGND.n42 VGND.n41 2.25932
R136 VGND.n66 VGND.n65 0.753441
R137 VGND.n24 VGND.n23 0.120292
R138 VGND.n24 VGND.n17 0.120292
R139 VGND.n31 VGND.n17 0.120292
R140 VGND.n32 VGND.n31 0.120292
R141 VGND.n33 VGND.n32 0.120292
R142 VGND.n33 VGND.n14 0.120292
R143 VGND.n38 VGND.n14 0.120292
R144 VGND.n39 VGND.n38 0.120292
R145 VGND.n39 VGND.n10 0.120292
R146 VGND.n46 VGND.n10 0.120292
R147 VGND.n47 VGND.n46 0.120292
R148 VGND.n48 VGND.n47 0.120292
R149 VGND.n48 VGND.n7 0.120292
R150 VGND.n55 VGND.n7 0.120292
R151 VGND.n56 VGND.n55 0.120292
R152 VGND.n57 VGND.n56 0.120292
R153 VGND.n57 VGND.n4 0.120292
R154 VGND.n62 VGND.n4 0.120292
R155 VGND.n63 VGND.n62 0.120292
R156 VGND.n63 VGND.n0 0.120292
R157 VGND.n67 VGND.n0 0.120292
R158 VGND VGND.n67 0.0213333
R159 a_361_47.n3 a_361_47.n1 244.457
R160 a_361_47.n16 a_361_47.t17 221.72
R161 a_361_47.n18 a_361_47.t28 221.72
R162 a_361_47.n15 a_361_47.t37 221.72
R163 a_361_47.n23 a_361_47.t42 221.72
R164 a_361_47.n25 a_361_47.t14 221.72
R165 a_361_47.n26 a_361_47.t16 221.72
R166 a_361_47.n32 a_361_47.t18 221.72
R167 a_361_47.n34 a_361_47.t31 221.72
R168 a_361_47.n11 a_361_47.t33 221.72
R169 a_361_47.n39 a_361_47.t35 221.72
R170 a_361_47.n9 a_361_47.t36 221.72
R171 a_361_47.n45 a_361_47.t40 221.72
R172 a_361_47.n47 a_361_47.t12 221.72
R173 a_361_47.n7 a_361_47.t24 221.72
R174 a_361_47.n53 a_361_47.t26 221.72
R175 a_361_47.n54 a_361_47.t27 221.72
R176 a_361_47.n3 a_361_47.n2 206.056
R177 a_361_47.n5 a_361_47.n4 206.056
R178 a_361_47.n20 a_361_47.n17 173.761
R179 a_361_47.n56 a_361_47.n55 152
R180 a_361_47.n52 a_361_47.n6 152
R181 a_361_47.n51 a_361_47.n50 152
R182 a_361_47.n49 a_361_47.n48 152
R183 a_361_47.n46 a_361_47.n8 152
R184 a_361_47.n44 a_361_47.n43 152
R185 a_361_47.n42 a_361_47.n41 152
R186 a_361_47.n40 a_361_47.n10 152
R187 a_361_47.n38 a_361_47.n37 152
R188 a_361_47.n36 a_361_47.n35 152
R189 a_361_47.n33 a_361_47.n12 152
R190 a_361_47.n31 a_361_47.n30 152
R191 a_361_47.n29 a_361_47.n13 152
R192 a_361_47.n28 a_361_47.n27 152
R193 a_361_47.n24 a_361_47.n14 152
R194 a_361_47.n22 a_361_47.n21 152
R195 a_361_47.n20 a_361_47.n19 152
R196 a_361_47.n16 a_361_47.t19 149.421
R197 a_361_47.n18 a_361_47.t41 149.421
R198 a_361_47.n15 a_361_47.t39 149.421
R199 a_361_47.n23 a_361_47.t34 149.421
R200 a_361_47.n25 a_361_47.t38 149.421
R201 a_361_47.n26 a_361_47.t32 149.421
R202 a_361_47.n32 a_361_47.t25 149.421
R203 a_361_47.n34 a_361_47.t30 149.421
R204 a_361_47.n11 a_361_47.t23 149.421
R205 a_361_47.n39 a_361_47.t29 149.421
R206 a_361_47.n9 a_361_47.t21 149.421
R207 a_361_47.n45 a_361_47.t13 149.421
R208 a_361_47.n47 a_361_47.t20 149.421
R209 a_361_47.n7 a_361_47.t43 149.421
R210 a_361_47.n53 a_361_47.t22 149.421
R211 a_361_47.n54 a_361_47.t15 149.421
R212 a_361_47.n60 a_361_47.n0 137.189
R213 a_361_47.n59 a_361_47.n58 98.788
R214 a_361_47.n61 a_361_47.n60 98.788
R215 a_361_47.n17 a_361_47.n16 73.1931
R216 a_361_47.n31 a_361_47.n13 60.6968
R217 a_361_47.n41 a_361_47.n40 60.6968
R218 a_361_47.n52 a_361_47.n51 60.6968
R219 a_361_47.n19 a_361_47.n18 58.9116
R220 a_361_47.n27 a_361_47.n26 58.9116
R221 a_361_47.n39 a_361_47.n38 55.3412
R222 a_361_47.n55 a_361_47.n53 55.3412
R223 a_361_47.n44 a_361_47.n9 51.7709
R224 a_361_47.n48 a_361_47.n7 51.7709
R225 a_361_47.n33 a_361_47.n32 48.2005
R226 a_361_47.n22 a_361_47.n15 44.6301
R227 a_361_47.n25 a_361_47.n24 44.6301
R228 a_361_47.n35 a_361_47.n11 41.0598
R229 a_361_47.n5 a_361_47.n3 38.4005
R230 a_361_47.n60 a_361_47.n59 38.4005
R231 a_361_47.n46 a_361_47.n45 37.4894
R232 a_361_47.n47 a_361_47.n46 37.4894
R233 a_361_47.n35 a_361_47.n34 33.919
R234 a_361_47.n57 a_361_47.n5 31.0755
R235 a_361_47.n59 a_361_47.n57 31.0755
R236 a_361_47.n23 a_361_47.n22 30.3486
R237 a_361_47.n24 a_361_47.n23 30.3486
R238 a_361_47.n34 a_361_47.n33 26.7783
R239 a_361_47.n1 a_361_47.t11 26.5955
R240 a_361_47.n1 a_361_47.t10 26.5955
R241 a_361_47.n2 a_361_47.t1 26.5955
R242 a_361_47.n2 a_361_47.t0 26.5955
R243 a_361_47.n4 a_361_47.t9 26.5955
R244 a_361_47.n4 a_361_47.t8 26.5955
R245 a_361_47.n58 a_361_47.t2 24.9236
R246 a_361_47.n58 a_361_47.t6 24.9236
R247 a_361_47.n0 a_361_47.t4 24.9236
R248 a_361_47.n0 a_361_47.t5 24.9236
R249 a_361_47.n61 a_361_47.t3 24.9236
R250 a_361_47.t7 a_361_47.n61 24.9236
R251 a_361_47.n45 a_361_47.n44 23.2079
R252 a_361_47.n48 a_361_47.n47 23.2079
R253 a_361_47.n21 a_361_47.n20 21.7605
R254 a_361_47.n21 a_361_47.n14 21.7605
R255 a_361_47.n28 a_361_47.n14 21.7605
R256 a_361_47.n29 a_361_47.n28 21.7605
R257 a_361_47.n30 a_361_47.n29 21.7605
R258 a_361_47.n30 a_361_47.n12 21.7605
R259 a_361_47.n36 a_361_47.n12 21.7605
R260 a_361_47.n37 a_361_47.n36 21.7605
R261 a_361_47.n37 a_361_47.n10 21.7605
R262 a_361_47.n42 a_361_47.n10 21.7605
R263 a_361_47.n43 a_361_47.n42 21.7605
R264 a_361_47.n43 a_361_47.n8 21.7605
R265 a_361_47.n49 a_361_47.n8 21.7605
R266 a_361_47.n50 a_361_47.n49 21.7605
R267 a_361_47.n50 a_361_47.n6 21.7605
R268 a_361_47.n56 a_361_47.n6 21.7605
R269 a_361_47.n57 a_361_47.n56 20.8005
R270 a_361_47.n38 a_361_47.n11 19.6375
R271 a_361_47.n55 a_361_47.n54 19.6375
R272 a_361_47.n19 a_361_47.n15 16.0672
R273 a_361_47.n27 a_361_47.n25 16.0672
R274 a_361_47.n32 a_361_47.n31 12.4968
R275 a_361_47.n41 a_361_47.n9 8.92643
R276 a_361_47.n51 a_361_47.n7 8.92643
R277 a_361_47.n40 a_361_47.n39 5.35606
R278 a_361_47.n53 a_361_47.n52 5.35606
R279 a_361_47.n18 a_361_47.n17 1.78569
R280 a_361_47.n26 a_361_47.n13 1.78569
R281 VNB.t4 VNB.t16 1196.12
R282 VNB.t5 VNB.t4 1196.12
R283 VNB.t7 VNB.t5 1196.12
R284 VNB.t6 VNB.t7 1196.12
R285 VNB.t8 VNB.t6 1196.12
R286 VNB.t11 VNB.t8 1196.12
R287 VNB.t9 VNB.t11 1196.12
R288 VNB.t12 VNB.t9 1196.12
R289 VNB.t10 VNB.t12 1196.12
R290 VNB.t14 VNB.t10 1196.12
R291 VNB.t18 VNB.t14 1196.12
R292 VNB.t15 VNB.t18 1196.12
R293 VNB.t3 VNB.t15 1196.12
R294 VNB.t13 VNB.t3 1196.12
R295 VNB.t17 VNB.t13 1196.12
R296 VNB.t19 VNB.t17 1196.12
R297 VNB.t23 VNB.t19 1196.12
R298 VNB.t20 VNB.t23 1196.12
R299 VNB.t24 VNB.t20 1196.12
R300 VNB.t21 VNB.t24 1196.12
R301 VNB.t22 VNB.t21 1196.12
R302 VNB.t1 VNB.t22 1196.12
R303 VNB.t0 VNB.t1 1196.12
R304 VNB.t2 VNB.t0 1196.12
R305 VNB VNB.t2 911.327
R306 Y.n2 Y.n0 244.457
R307 Y.n2 Y.n1 206.056
R308 Y.n4 Y.n3 206.056
R309 Y.n6 Y.n5 206.056
R310 Y.n8 Y.n7 206.056
R311 Y.n10 Y.n9 206.056
R312 Y.n12 Y.n11 206.056
R313 Y.n14 Y.n13 206.056
R314 Y.n17 Y.n15 137.189
R315 Y.n17 Y.n16 98.788
R316 Y.n19 Y.n18 98.788
R317 Y.n21 Y.n20 98.788
R318 Y.n23 Y.n22 98.788
R319 Y.n25 Y.n24 98.788
R320 Y.n27 Y.n26 98.788
R321 Y.n29 Y.n28 98.788
R322 Y.n19 Y.n17 38.4005
R323 Y.n21 Y.n19 38.4005
R324 Y.n23 Y.n21 38.4005
R325 Y.n25 Y.n23 38.4005
R326 Y.n27 Y.n25 38.4005
R327 Y.n29 Y.n27 38.4005
R328 Y.n4 Y.n2 38.4005
R329 Y.n6 Y.n4 38.4005
R330 Y.n8 Y.n6 38.4005
R331 Y.n10 Y.n8 38.4005
R332 Y.n12 Y.n10 38.4005
R333 Y.n14 Y.n12 38.4005
R334 Y.n0 Y.t9 26.5955
R335 Y.n0 Y.t8 26.5955
R336 Y.n1 Y.t15 26.5955
R337 Y.n1 Y.t10 26.5955
R338 Y.n3 Y.t3 26.5955
R339 Y.n3 Y.t1 26.5955
R340 Y.n5 Y.t5 26.5955
R341 Y.n5 Y.t4 26.5955
R342 Y.n7 Y.t11 26.5955
R343 Y.n7 Y.t6 26.5955
R344 Y.n9 Y.t14 26.5955
R345 Y.n9 Y.t13 26.5955
R346 Y.n11 Y.t2 26.5955
R347 Y.n11 Y.t0 26.5955
R348 Y.n13 Y.t12 26.5955
R349 Y.n13 Y.t7 26.5955
R350 Y Y.n29 26.4424
R351 Y.n15 Y.t26 24.9236
R352 Y.n15 Y.t30 24.9236
R353 Y.n16 Y.t28 24.9236
R354 Y.n16 Y.t16 24.9236
R355 Y.n18 Y.t27 24.9236
R356 Y.n18 Y.t31 24.9236
R357 Y.n20 Y.t25 24.9236
R358 Y.n20 Y.t23 24.9236
R359 Y.n22 Y.t24 24.9236
R360 Y.n22 Y.t22 24.9236
R361 Y.n24 Y.t19 24.9236
R362 Y.n24 Y.t21 24.9236
R363 Y.n26 Y.t18 24.9236
R364 Y.n26 Y.t20 24.9236
R365 Y.n28 Y.t29 24.9236
R366 Y.n28 Y.t17 24.9236
R367 Y Y.n14 17.1333
R368 VPWR.n22 VPWR.t15 355.2
R369 VPWR.n3 VPWR.n2 320.976
R370 VPWR.n59 VPWR.n5 320.976
R371 VPWR.n53 VPWR.n52 320.976
R372 VPWR.n50 VPWR.n8 320.976
R373 VPWR.n44 VPWR.n43 320.976
R374 VPWR.n42 VPWR.n11 320.976
R375 VPWR.n13 VPWR.n12 320.976
R376 VPWR.n35 VPWR.n15 320.976
R377 VPWR.n29 VPWR.n28 320.976
R378 VPWR.n26 VPWR.n18 320.976
R379 VPWR.n21 VPWR.n20 320.976
R380 VPWR.n66 VPWR.n1 320.976
R381 VPWR.n67 VPWR.n66 43.1829
R382 VPWR.n22 VPWR.n21 37.7583
R383 VPWR.n25 VPWR.n19 34.6358
R384 VPWR.n30 VPWR.n27 34.6358
R385 VPWR.n34 VPWR.n16 34.6358
R386 VPWR.n37 VPWR.n36 34.6358
R387 VPWR.n41 VPWR.n40 34.6358
R388 VPWR.n49 VPWR.n9 34.6358
R389 VPWR.n54 VPWR.n51 34.6358
R390 VPWR.n58 VPWR.n6 34.6358
R391 VPWR.n61 VPWR.n60 34.6358
R392 VPWR.n65 VPWR.n64 34.6358
R393 VPWR.n45 VPWR.n42 32.377
R394 VPWR.n45 VPWR.n44 30.8711
R395 VPWR.n64 VPWR.n3 27.8593
R396 VPWR.n1 VPWR.t1 26.5955
R397 VPWR.n1 VPWR.t2 26.5955
R398 VPWR.n2 VPWR.t23 26.5955
R399 VPWR.n2 VPWR.t0 26.5955
R400 VPWR.n5 VPWR.t19 26.5955
R401 VPWR.n5 VPWR.t24 26.5955
R402 VPWR.n52 VPWR.t21 26.5955
R403 VPWR.n52 VPWR.t20 26.5955
R404 VPWR.n8 VPWR.t11 26.5955
R405 VPWR.n8 VPWR.t22 26.5955
R406 VPWR.n43 VPWR.t13 26.5955
R407 VPWR.n43 VPWR.t12 26.5955
R408 VPWR.n11 VPWR.t4 26.5955
R409 VPWR.n11 VPWR.t18 26.5955
R410 VPWR.n12 VPWR.t7 26.5955
R411 VPWR.n12 VPWR.t6 26.5955
R412 VPWR.n15 VPWR.t9 26.5955
R413 VPWR.n15 VPWR.t8 26.5955
R414 VPWR.n28 VPWR.t16 26.5955
R415 VPWR.n28 VPWR.t14 26.5955
R416 VPWR.n18 VPWR.t3 26.5955
R417 VPWR.n18 VPWR.t17 26.5955
R418 VPWR.n20 VPWR.t10 26.5955
R419 VPWR.n20 VPWR.t5 26.5955
R420 VPWR.n26 VPWR.n25 26.3534
R421 VPWR.n40 VPWR.n13 26.3534
R422 VPWR.n50 VPWR.n49 24.8476
R423 VPWR.n60 VPWR.n59 21.8358
R424 VPWR.n30 VPWR.n29 20.3299
R425 VPWR.n36 VPWR.n35 20.3299
R426 VPWR.n54 VPWR.n53 18.824
R427 VPWR.n53 VPWR.n6 15.8123
R428 VPWR.n29 VPWR.n16 14.3064
R429 VPWR.n35 VPWR.n34 14.3064
R430 VPWR.n59 VPWR.n58 12.8005
R431 VPWR.n51 VPWR.n50 9.78874
R432 VPWR.n23 VPWR.n19 9.3005
R433 VPWR.n25 VPWR.n24 9.3005
R434 VPWR.n27 VPWR.n17 9.3005
R435 VPWR.n31 VPWR.n30 9.3005
R436 VPWR.n32 VPWR.n16 9.3005
R437 VPWR.n34 VPWR.n33 9.3005
R438 VPWR.n36 VPWR.n14 9.3005
R439 VPWR.n38 VPWR.n37 9.3005
R440 VPWR.n40 VPWR.n39 9.3005
R441 VPWR.n41 VPWR.n10 9.3005
R442 VPWR.n46 VPWR.n45 9.3005
R443 VPWR.n47 VPWR.n9 9.3005
R444 VPWR.n49 VPWR.n48 9.3005
R445 VPWR.n51 VPWR.n7 9.3005
R446 VPWR.n55 VPWR.n54 9.3005
R447 VPWR.n56 VPWR.n6 9.3005
R448 VPWR.n58 VPWR.n57 9.3005
R449 VPWR.n60 VPWR.n4 9.3005
R450 VPWR.n62 VPWR.n61 9.3005
R451 VPWR.n64 VPWR.n63 9.3005
R452 VPWR.n65 VPWR.n0 9.3005
R453 VPWR.n27 VPWR.n26 8.28285
R454 VPWR.n37 VPWR.n13 8.28285
R455 VPWR.n61 VPWR.n3 6.77697
R456 VPWR.n44 VPWR.n9 3.76521
R457 VPWR.n23 VPWR.n22 2.4189
R458 VPWR.n21 VPWR.n19 2.25932
R459 VPWR.n42 VPWR.n41 2.25932
R460 VPWR.n66 VPWR.n65 0.753441
R461 VPWR.n24 VPWR.n23 0.120292
R462 VPWR.n24 VPWR.n17 0.120292
R463 VPWR.n31 VPWR.n17 0.120292
R464 VPWR.n32 VPWR.n31 0.120292
R465 VPWR.n33 VPWR.n32 0.120292
R466 VPWR.n33 VPWR.n14 0.120292
R467 VPWR.n38 VPWR.n14 0.120292
R468 VPWR.n39 VPWR.n38 0.120292
R469 VPWR.n39 VPWR.n10 0.120292
R470 VPWR.n46 VPWR.n10 0.120292
R471 VPWR.n47 VPWR.n46 0.120292
R472 VPWR.n48 VPWR.n47 0.120292
R473 VPWR.n48 VPWR.n7 0.120292
R474 VPWR.n55 VPWR.n7 0.120292
R475 VPWR.n56 VPWR.n55 0.120292
R476 VPWR.n57 VPWR.n56 0.120292
R477 VPWR.n57 VPWR.n4 0.120292
R478 VPWR.n62 VPWR.n4 0.120292
R479 VPWR.n63 VPWR.n62 0.120292
R480 VPWR.n63 VPWR.n0 0.120292
R481 VPWR.n67 VPWR.n0 0.120292
R482 VPWR VPWR.n67 0.0213333
R483 VPB.t10 VPB.t15 248.599
R484 VPB.t5 VPB.t10 248.599
R485 VPB.t3 VPB.t5 248.599
R486 VPB.t17 VPB.t3 248.599
R487 VPB.t16 VPB.t17 248.599
R488 VPB.t14 VPB.t16 248.599
R489 VPB.t9 VPB.t14 248.599
R490 VPB.t8 VPB.t9 248.599
R491 VPB.t7 VPB.t8 248.599
R492 VPB.t6 VPB.t7 248.599
R493 VPB.t4 VPB.t6 248.599
R494 VPB.t18 VPB.t4 248.599
R495 VPB.t13 VPB.t18 248.599
R496 VPB.t12 VPB.t13 248.599
R497 VPB.t11 VPB.t12 248.599
R498 VPB.t22 VPB.t11 248.599
R499 VPB.t21 VPB.t22 248.599
R500 VPB.t20 VPB.t21 248.599
R501 VPB.t19 VPB.t20 248.599
R502 VPB.t24 VPB.t19 248.599
R503 VPB.t23 VPB.t24 248.599
R504 VPB.t0 VPB.t23 248.599
R505 VPB.t1 VPB.t0 248.599
R506 VPB.t2 VPB.t1 248.599
R507 VPB VPB.t2 189.409
R508 A.n0 A.t0 221.72
R509 A.n2 A.t1 221.72
R510 A.n3 A.t4 221.72
R511 A.n5 A.n1 173.761
R512 A.n5 A.n4 152
R513 A.n0 A.t3 149.421
R514 A.n2 A.t2 149.421
R515 A.n3 A.t5 149.421
R516 A.n1 A.n0 51.7709
R517 A.n4 A.n2 37.4894
R518 A.n4 A.n3 37.4894
R519 A A.n5 33.9205
R520 A.n2 A.n1 23.2079
C0 VPB A 0.08817f
C1 VPB VPWR 0.208345f
C2 VPB Y 0.034848f
C3 A VPWR 0.049802f
C4 VPB VGND 0.012723f
C5 A VGND 0.04463f
C6 VPWR Y 1.45006f
C7 VPWR VGND 0.2259f
C8 Y VGND 1.053f
C9 VGND VNB 1.19187f
C10 Y VNB 0.077469f
C11 VPWR VNB 1.01898f
C12 A VNB 0.299674f
C13 VPB VNB 2.19949f
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufinv_8 VNB VPB VGND VPWR A Y
X0 VPWR.t11 a_215_47.t6 Y.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t3 a_109_47.t2 a_215_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 VGND.t2 a_109_47.t3 a_215_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t11 a_215_47.t7 Y.t15 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t6 a_215_47.t8 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t10 a_215_47.t9 Y.t14 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t13 a_215_47.t10 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y.t12 a_215_47.t11 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t11 a_215_47.t12 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y.t10 a_215_47.t13 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR.t9 a_215_47.t14 Y.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y.t4 a_215_47.t15 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t5 a_215_47.t16 Y.t9 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t4 a_215_47.t17 Y.t8 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t2 a_109_47.t4 a_215_47.t4 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_215_47.t0 a_109_47.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR.t7 a_215_47.t18 Y.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_215_47.t3 a_109_47.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR.t3 a_109_47.t7 a_215_47.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y.t2 a_215_47.t19 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t5 a_215_47.t20 Y.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_109_47.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 Y.t0 a_215_47.t21 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_109_47.t1 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_215_47.n28 a_215_47.t5 271.051
R1 a_215_47.n7 a_215_47.t18 221.72
R2 a_215_47.n9 a_215_47.t19 221.72
R3 a_215_47.n5 a_215_47.t20 221.72
R4 a_215_47.n15 a_215_47.t21 221.72
R5 a_215_47.n17 a_215_47.t6 221.72
R6 a_215_47.n3 a_215_47.t8 221.72
R7 a_215_47.n23 a_215_47.t14 221.72
R8 a_215_47.n24 a_215_47.t15 221.72
R9 a_215_47.n29 a_215_47.n28 206.055
R10 a_215_47.n1 a_215_47.t2 176.525
R11 a_215_47.n8 a_215_47.n6 173.761
R12 a_215_47.n26 a_215_47.n25 152
R13 a_215_47.n22 a_215_47.n2 152
R14 a_215_47.n21 a_215_47.n20 152
R15 a_215_47.n19 a_215_47.n18 152
R16 a_215_47.n16 a_215_47.n4 152
R17 a_215_47.n14 a_215_47.n13 152
R18 a_215_47.n12 a_215_47.n11 152
R19 a_215_47.n10 a_215_47.n6 152
R20 a_215_47.n7 a_215_47.t16 149.421
R21 a_215_47.n9 a_215_47.t11 149.421
R22 a_215_47.n5 a_215_47.t17 149.421
R23 a_215_47.n15 a_215_47.t13 149.421
R24 a_215_47.n17 a_215_47.t9 149.421
R25 a_215_47.n3 a_215_47.t12 149.421
R26 a_215_47.n23 a_215_47.t7 149.421
R27 a_215_47.n24 a_215_47.t10 149.421
R28 a_215_47.n1 a_215_47.n0 98.788
R29 a_215_47.n11 a_215_47.n10 60.6968
R30 a_215_47.n22 a_215_47.n21 60.6968
R31 a_215_47.n9 a_215_47.n8 58.9116
R32 a_215_47.n18 a_215_47.n3 55.3412
R33 a_215_47.n25 a_215_47.n23 51.7709
R34 a_215_47.n14 a_215_47.n5 48.2005
R35 a_215_47.n17 a_215_47.n16 41.0598
R36 a_215_47.n16 a_215_47.n15 33.919
R37 a_215_47.n27 a_215_47.n1 32.0005
R38 a_215_47.n28 a_215_47.n27 32.0005
R39 a_215_47.n15 a_215_47.n14 26.7783
R40 a_215_47.n29 a_215_47.t4 26.5955
R41 a_215_47.t0 a_215_47.n29 26.5955
R42 a_215_47.n0 a_215_47.t1 24.9236
R43 a_215_47.n0 a_215_47.t3 24.9236
R44 a_215_47.n25 a_215_47.n24 23.2079
R45 a_215_47.n12 a_215_47.n6 21.7605
R46 a_215_47.n13 a_215_47.n12 21.7605
R47 a_215_47.n13 a_215_47.n4 21.7605
R48 a_215_47.n19 a_215_47.n4 21.7605
R49 a_215_47.n20 a_215_47.n19 21.7605
R50 a_215_47.n20 a_215_47.n2 21.7605
R51 a_215_47.n26 a_215_47.n2 21.7605
R52 a_215_47.n27 a_215_47.n26 21.7605
R53 a_215_47.n18 a_215_47.n17 19.6375
R54 a_215_47.n8 a_215_47.n7 16.0672
R55 a_215_47.n11 a_215_47.n5 12.4968
R56 a_215_47.n23 a_215_47.n22 8.92643
R57 a_215_47.n21 a_215_47.n3 5.35606
R58 a_215_47.n10 a_215_47.n9 1.78569
R59 Y.n2 Y.n0 244.457
R60 Y.n2 Y.n1 206.056
R61 Y.n4 Y.n3 206.056
R62 Y.n6 Y.n5 206.056
R63 Y.n9 Y.n7 137.189
R64 Y.n9 Y.n8 98.788
R65 Y.n11 Y.n10 98.788
R66 Y.n13 Y.n12 98.788
R67 Y Y.n13 39.9699
R68 Y.n11 Y.n9 38.4005
R69 Y.n13 Y.n11 38.4005
R70 Y.n4 Y.n2 38.4005
R71 Y.n6 Y.n4 38.4005
R72 Y Y.n6 33.3206
R73 Y.n0 Y.t5 26.5955
R74 Y.n0 Y.t4 26.5955
R75 Y.n1 Y.t7 26.5955
R76 Y.n1 Y.t6 26.5955
R77 Y.n3 Y.t1 26.5955
R78 Y.n3 Y.t0 26.5955
R79 Y.n5 Y.t3 26.5955
R80 Y.n5 Y.t2 26.5955
R81 Y.n7 Y.t15 24.9236
R82 Y.n7 Y.t13 24.9236
R83 Y.n8 Y.t14 24.9236
R84 Y.n8 Y.t11 24.9236
R85 Y.n10 Y.t8 24.9236
R86 Y.n10 Y.t10 24.9236
R87 Y.n12 Y.t9 24.9236
R88 Y.n12 Y.t12 24.9236
R89 VPWR.n11 VPWR.t7 356.132
R90 VPWR.n24 VPWR.n23 320.976
R91 VPWR.n22 VPWR.n3 320.976
R92 VPWR.n5 VPWR.n4 320.976
R93 VPWR.n15 VPWR.n7 320.976
R94 VPWR.n10 VPWR.n9 320.976
R95 VPWR.n31 VPWR.t0 257.474
R96 VPWR.n14 VPWR.n8 34.6358
R97 VPWR.n17 VPWR.n16 34.6358
R98 VPWR.n21 VPWR.n20 34.6358
R99 VPWR.n29 VPWR.n1 34.6358
R100 VPWR.n30 VPWR.n29 34.6358
R101 VPWR.n25 VPWR.n24 33.8829
R102 VPWR.n31 VPWR.n30 32.377
R103 VPWR.n11 VPWR.n10 29.7335
R104 VPWR.n25 VPWR.n22 29.3652
R105 VPWR.n23 VPWR.t1 26.5955
R106 VPWR.n23 VPWR.t3 26.5955
R107 VPWR.n3 VPWR.t8 26.5955
R108 VPWR.n3 VPWR.t2 26.5955
R109 VPWR.n4 VPWR.t10 26.5955
R110 VPWR.n4 VPWR.t9 26.5955
R111 VPWR.n7 VPWR.t4 26.5955
R112 VPWR.n7 VPWR.t11 26.5955
R113 VPWR.n9 VPWR.t6 26.5955
R114 VPWR.n9 VPWR.t5 26.5955
R115 VPWR.n20 VPWR.n5 23.3417
R116 VPWR.n15 VPWR.n14 17.3181
R117 VPWR.n16 VPWR.n15 17.3181
R118 VPWR.n32 VPWR.n31 11.5593
R119 VPWR.n10 VPWR.n8 11.2946
R120 VPWR.n17 VPWR.n5 11.2946
R121 VPWR.n12 VPWR.n8 9.3005
R122 VPWR.n14 VPWR.n13 9.3005
R123 VPWR.n16 VPWR.n6 9.3005
R124 VPWR.n18 VPWR.n17 9.3005
R125 VPWR.n20 VPWR.n19 9.3005
R126 VPWR.n21 VPWR.n2 9.3005
R127 VPWR.n26 VPWR.n25 9.3005
R128 VPWR.n27 VPWR.n1 9.3005
R129 VPWR.n29 VPWR.n28 9.3005
R130 VPWR.n30 VPWR.n0 9.3005
R131 VPWR.n22 VPWR.n21 5.27109
R132 VPWR.n12 VPWR.n11 1.35766
R133 VPWR.n24 VPWR.n1 0.753441
R134 VPWR.n13 VPWR.n12 0.120292
R135 VPWR.n13 VPWR.n6 0.120292
R136 VPWR.n18 VPWR.n6 0.120292
R137 VPWR.n19 VPWR.n18 0.120292
R138 VPWR.n19 VPWR.n2 0.120292
R139 VPWR.n26 VPWR.n2 0.120292
R140 VPWR.n27 VPWR.n26 0.120292
R141 VPWR.n28 VPWR.n27 0.120292
R142 VPWR.n28 VPWR.n0 0.120292
R143 VPWR.n32 VPWR.n0 0.120292
R144 VPWR VPWR.n32 0.0213333
R145 VPB.t0 VPB.t3 556.386
R146 VPB.t6 VPB.t7 248.599
R147 VPB.t5 VPB.t6 248.599
R148 VPB.t4 VPB.t5 248.599
R149 VPB.t11 VPB.t4 248.599
R150 VPB.t10 VPB.t11 248.599
R151 VPB.t9 VPB.t10 248.599
R152 VPB.t8 VPB.t9 248.599
R153 VPB.t2 VPB.t8 248.599
R154 VPB.t1 VPB.t2 248.599
R155 VPB.t3 VPB.t1 248.599
R156 VPB VPB.t0 189.409
R157 a_109_47.t0 a_109_47.n6 252.399
R158 a_109_47.n0 a_109_47.t4 221.72
R159 a_109_47.n2 a_109_47.t5 221.72
R160 a_109_47.n3 a_109_47.t7 221.72
R161 a_109_47.n5 a_109_47.n1 173.761
R162 a_109_47.n6 a_109_47.t1 154.221
R163 a_109_47.n5 a_109_47.n4 152
R164 a_109_47.n0 a_109_47.t3 149.421
R165 a_109_47.n2 a_109_47.t6 149.421
R166 a_109_47.n3 a_109_47.t2 149.421
R167 a_109_47.n6 a_109_47.n5 55.0405
R168 a_109_47.n1 a_109_47.n0 51.7709
R169 a_109_47.n4 a_109_47.n2 37.4894
R170 a_109_47.n4 a_109_47.n3 37.4894
R171 a_109_47.n2 a_109_47.n1 23.2079
R172 VGND.n11 VGND.t5 291.125
R173 VGND.n10 VGND.n9 208.719
R174 VGND.n15 VGND.n7 208.719
R175 VGND.n5 VGND.n4 208.719
R176 VGND.n22 VGND.n3 208.719
R177 VGND.n24 VGND.n23 208.719
R178 VGND.n31 VGND.t0 161.302
R179 VGND.n14 VGND.n8 34.6358
R180 VGND.n17 VGND.n16 34.6358
R181 VGND.n21 VGND.n20 34.6358
R182 VGND.n29 VGND.n1 34.6358
R183 VGND.n30 VGND.n29 34.6358
R184 VGND.n25 VGND.n24 33.8829
R185 VGND.n31 VGND.n30 32.377
R186 VGND.n11 VGND.n10 29.7335
R187 VGND.n25 VGND.n22 29.3652
R188 VGND.n9 VGND.t8 24.9236
R189 VGND.n9 VGND.t4 24.9236
R190 VGND.n7 VGND.t6 24.9236
R191 VGND.n7 VGND.t10 24.9236
R192 VGND.n4 VGND.t7 24.9236
R193 VGND.n4 VGND.t11 24.9236
R194 VGND.n3 VGND.t9 24.9236
R195 VGND.n3 VGND.t2 24.9236
R196 VGND.n23 VGND.t1 24.9236
R197 VGND.n23 VGND.t3 24.9236
R198 VGND.n20 VGND.n5 23.3417
R199 VGND.n15 VGND.n14 17.3181
R200 VGND.n16 VGND.n15 17.3181
R201 VGND.n32 VGND.n31 11.5593
R202 VGND.n10 VGND.n8 11.2946
R203 VGND.n17 VGND.n5 11.2946
R204 VGND.n12 VGND.n8 9.3005
R205 VGND.n14 VGND.n13 9.3005
R206 VGND.n16 VGND.n6 9.3005
R207 VGND.n18 VGND.n17 9.3005
R208 VGND.n20 VGND.n19 9.3005
R209 VGND.n21 VGND.n2 9.3005
R210 VGND.n26 VGND.n25 9.3005
R211 VGND.n27 VGND.n1 9.3005
R212 VGND.n29 VGND.n28 9.3005
R213 VGND.n30 VGND.n0 9.3005
R214 VGND.n22 VGND.n21 5.27109
R215 VGND.n12 VGND.n11 1.35766
R216 VGND.n24 VGND.n1 0.753441
R217 VGND.n13 VGND.n12 0.120292
R218 VGND.n13 VGND.n6 0.120292
R219 VGND.n18 VGND.n6 0.120292
R220 VGND.n19 VGND.n18 0.120292
R221 VGND.n19 VGND.n2 0.120292
R222 VGND.n26 VGND.n2 0.120292
R223 VGND.n27 VGND.n26 0.120292
R224 VGND.n28 VGND.n27 0.120292
R225 VGND.n28 VGND.n0 0.120292
R226 VGND.n32 VGND.n0 0.120292
R227 VGND VGND.n32 0.0213333
R228 VNB.t0 VNB.t3 2677.02
R229 VNB.t8 VNB.t5 1196.12
R230 VNB.t4 VNB.t8 1196.12
R231 VNB.t6 VNB.t4 1196.12
R232 VNB.t10 VNB.t6 1196.12
R233 VNB.t7 VNB.t10 1196.12
R234 VNB.t11 VNB.t7 1196.12
R235 VNB.t9 VNB.t11 1196.12
R236 VNB.t2 VNB.t9 1196.12
R237 VNB.t1 VNB.t2 1196.12
R238 VNB.t3 VNB.t1 1196.12
R239 VNB VNB.t0 911.327
R240 A.n0 A.t0 230.155
R241 A A.n0 160
R242 A.n0 A.t1 157.856
C0 VPB A 0.044154f
C1 VPB VPWR 0.149338f
C2 A VPWR 0.043015f
C3 VPB Y 0.031887f
C4 VPB VGND 0.012762f
C5 A VGND 0.042931f
C6 VPWR Y 0.738422f
C7 VPWR VGND 0.131565f
C8 Y VGND 0.540408f
C9 VGND VNB 0.770145f
C10 Y VNB 0.076047f
C11 VPWR VNB 0.669033f
C12 A VNB 0.152757f
C13 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufbuf_16 VNB VPB VGND VPWR A X
X0 X.t15 a_549_47.t12 VPWR.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t31 a_549_47.t13 VGND.t15 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t24 a_215_47.t6 a_549_47.t8 VPB.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t22 a_109_47.t2 a_215_47.t2 VNB.t22 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 X.t14 a_549_47.t14 VPWR.t15 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t23 a_109_47.t3 a_215_47.t3 VNB.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND.t24 a_215_47.t7 a_549_47.t9 VNB.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_549_47.t10 a_215_47.t8 VPWR.t25 VPB.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t14 a_549_47.t15 X.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t25 a_215_47.t9 a_549_47.t11 VNB.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t14 a_549_47.t16 X.t30 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t13 a_549_47.t17 X.t29 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t12 a_549_47.t18 VPWR.t13 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X.t28 a_549_47.t19 VGND.t12 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_549_47.t0 a_215_47.t10 VGND.t18 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR.t12 a_549_47.t20 X.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X.t27 a_549_47.t21 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t11 a_549_47.t22 X.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 X.t9 a_549_47.t23 VPWR.t10 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_549_47.t1 a_215_47.t11 VGND.t19 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_549_47.t2 a_215_47.t12 VGND.t20 VNB.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 X.t26 a_549_47.t24 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 X.t8 a_549_47.t25 VPWR.t9 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR.t17 a_215_47.t13 a_549_47.t3 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t8 a_549_47.t26 X.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND.t9 a_549_47.t27 X.t25 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t7 a_549_47.t28 X.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_549_47.t4 a_215_47.t14 VPWR.t18 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X.t5 a_549_47.t29 VPWR.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND.t8 a_549_47.t30 X.t24 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VGND.t7 a_549_47.t31 X.t23 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 X.t4 a_549_47.t32 VPWR.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VGND.t21 a_215_47.t15 a_549_47.t5 VNB.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t6 a_549_47.t33 X.t22 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 VGND.t5 a_549_47.t34 X.t21 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 VPWR.t22 a_109_47.t4 a_215_47.t4 VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND.t4 a_549_47.t35 X.t20 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 a_215_47.t5 a_109_47.t5 VPWR.t23 VPB.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 VPWR.t4 a_549_47.t36 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 X.t19 a_549_47.t37 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 a_215_47.t0 a_109_47.t6 VGND.t16 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 VPWR.t16 a_109_47.t7 a_215_47.t1 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X42 X.t2 a_549_47.t38 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X43 VPWR.t19 a_215_47.t16 a_549_47.t6 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 X.t18 a_549_47.t39 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X45 X.t17 a_549_47.t40 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 a_109_47.t1 A.t0 VPWR.t21 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X47 VPWR.t2 a_549_47.t41 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 a_549_47.t7 a_215_47.t17 VPWR.t20 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X49 VPWR.t1 a_549_47.t42 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X50 a_109_47.t0 A.t1 VGND.t17 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X51 X.t16 a_549_47.t43 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 a_549_47.n61 a_549_47.n60 244.457
R1 a_549_47.n15 a_549_47.t26 221.72
R2 a_549_47.n17 a_549_47.t29 221.72
R3 a_549_47.n14 a_549_47.t41 221.72
R4 a_549_47.n22 a_549_47.t12 221.72
R5 a_549_47.n24 a_549_47.t22 221.72
R6 a_549_47.n25 a_549_47.t25 221.72
R7 a_549_47.n31 a_549_47.t28 221.72
R8 a_549_47.n33 a_549_47.t32 221.72
R9 a_549_47.n10 a_549_47.t42 221.72
R10 a_549_47.n38 a_549_47.t14 221.72
R11 a_549_47.n8 a_549_47.t15 221.72
R12 a_549_47.n44 a_549_47.t18 221.72
R13 a_549_47.n46 a_549_47.t20 221.72
R14 a_549_47.n6 a_549_47.t23 221.72
R15 a_549_47.n52 a_549_47.t36 221.72
R16 a_549_47.n53 a_549_47.t38 221.72
R17 a_549_47.n58 a_549_47.n57 206.056
R18 a_549_47.n60 a_549_47.n59 206.056
R19 a_549_47.n19 a_549_47.n16 173.761
R20 a_549_47.n55 a_549_47.n54 152
R21 a_549_47.n51 a_549_47.n5 152
R22 a_549_47.n50 a_549_47.n49 152
R23 a_549_47.n48 a_549_47.n47 152
R24 a_549_47.n45 a_549_47.n7 152
R25 a_549_47.n43 a_549_47.n42 152
R26 a_549_47.n41 a_549_47.n40 152
R27 a_549_47.n39 a_549_47.n9 152
R28 a_549_47.n37 a_549_47.n36 152
R29 a_549_47.n35 a_549_47.n34 152
R30 a_549_47.n32 a_549_47.n11 152
R31 a_549_47.n30 a_549_47.n29 152
R32 a_549_47.n28 a_549_47.n12 152
R33 a_549_47.n27 a_549_47.n26 152
R34 a_549_47.n23 a_549_47.n13 152
R35 a_549_47.n21 a_549_47.n20 152
R36 a_549_47.n19 a_549_47.n18 152
R37 a_549_47.n15 a_549_47.t31 149.421
R38 a_549_47.n17 a_549_47.t37 149.421
R39 a_549_47.n14 a_549_47.t27 149.421
R40 a_549_47.n22 a_549_47.t19 149.421
R41 a_549_47.n24 a_549_47.t17 149.421
R42 a_549_47.n25 a_549_47.t13 149.421
R43 a_549_47.n31 a_549_47.t16 149.421
R44 a_549_47.n33 a_549_47.t43 149.421
R45 a_549_47.n10 a_549_47.t35 149.421
R46 a_549_47.n38 a_549_47.t40 149.421
R47 a_549_47.n8 a_549_47.t34 149.421
R48 a_549_47.n44 a_549_47.t39 149.421
R49 a_549_47.n46 a_549_47.t33 149.421
R50 a_549_47.n6 a_549_47.t24 149.421
R51 a_549_47.n52 a_549_47.t30 149.421
R52 a_549_47.n53 a_549_47.t21 149.421
R53 a_549_47.n2 a_549_47.n0 137.189
R54 a_549_47.n2 a_549_47.n1 98.788
R55 a_549_47.n4 a_549_47.n3 98.788
R56 a_549_47.n16 a_549_47.n15 73.1931
R57 a_549_47.n30 a_549_47.n12 60.6968
R58 a_549_47.n40 a_549_47.n39 60.6968
R59 a_549_47.n51 a_549_47.n50 60.6968
R60 a_549_47.n18 a_549_47.n17 58.9116
R61 a_549_47.n26 a_549_47.n25 58.9116
R62 a_549_47.n38 a_549_47.n37 55.3412
R63 a_549_47.n54 a_549_47.n52 55.3412
R64 a_549_47.n43 a_549_47.n8 51.7709
R65 a_549_47.n47 a_549_47.n6 51.7709
R66 a_549_47.n32 a_549_47.n31 48.2005
R67 a_549_47.n21 a_549_47.n14 44.6301
R68 a_549_47.n24 a_549_47.n23 44.6301
R69 a_549_47.n34 a_549_47.n10 41.0598
R70 a_549_47.n4 a_549_47.n2 38.4005
R71 a_549_47.n60 a_549_47.n58 38.4005
R72 a_549_47.n45 a_549_47.n44 37.4894
R73 a_549_47.n46 a_549_47.n45 37.4894
R74 a_549_47.n34 a_549_47.n33 33.919
R75 a_549_47.n56 a_549_47.n4 31.0755
R76 a_549_47.n58 a_549_47.n56 31.0755
R77 a_549_47.n22 a_549_47.n21 30.3486
R78 a_549_47.n23 a_549_47.n22 30.3486
R79 a_549_47.n33 a_549_47.n32 26.7783
R80 a_549_47.n57 a_549_47.t6 26.5955
R81 a_549_47.n57 a_549_47.t7 26.5955
R82 a_549_47.n59 a_549_47.t8 26.5955
R83 a_549_47.n59 a_549_47.t10 26.5955
R84 a_549_47.t3 a_549_47.n61 26.5955
R85 a_549_47.n61 a_549_47.t4 26.5955
R86 a_549_47.n0 a_549_47.t9 24.9236
R87 a_549_47.n0 a_549_47.t0 24.9236
R88 a_549_47.n1 a_549_47.t11 24.9236
R89 a_549_47.n1 a_549_47.t1 24.9236
R90 a_549_47.n3 a_549_47.t5 24.9236
R91 a_549_47.n3 a_549_47.t2 24.9236
R92 a_549_47.n44 a_549_47.n43 23.2079
R93 a_549_47.n47 a_549_47.n46 23.2079
R94 a_549_47.n20 a_549_47.n19 21.7605
R95 a_549_47.n20 a_549_47.n13 21.7605
R96 a_549_47.n27 a_549_47.n13 21.7605
R97 a_549_47.n28 a_549_47.n27 21.7605
R98 a_549_47.n29 a_549_47.n28 21.7605
R99 a_549_47.n29 a_549_47.n11 21.7605
R100 a_549_47.n35 a_549_47.n11 21.7605
R101 a_549_47.n36 a_549_47.n35 21.7605
R102 a_549_47.n36 a_549_47.n9 21.7605
R103 a_549_47.n41 a_549_47.n9 21.7605
R104 a_549_47.n42 a_549_47.n41 21.7605
R105 a_549_47.n42 a_549_47.n7 21.7605
R106 a_549_47.n48 a_549_47.n7 21.7605
R107 a_549_47.n49 a_549_47.n48 21.7605
R108 a_549_47.n49 a_549_47.n5 21.7605
R109 a_549_47.n55 a_549_47.n5 21.7605
R110 a_549_47.n56 a_549_47.n55 20.8005
R111 a_549_47.n37 a_549_47.n10 19.6375
R112 a_549_47.n54 a_549_47.n53 19.6375
R113 a_549_47.n18 a_549_47.n14 16.0672
R114 a_549_47.n26 a_549_47.n24 16.0672
R115 a_549_47.n31 a_549_47.n30 12.4968
R116 a_549_47.n40 a_549_47.n8 8.92643
R117 a_549_47.n50 a_549_47.n6 8.92643
R118 a_549_47.n39 a_549_47.n38 5.35606
R119 a_549_47.n52 a_549_47.n51 5.35606
R120 a_549_47.n17 a_549_47.n16 1.78569
R121 a_549_47.n25 a_549_47.n12 1.78569
R122 VPWR.n21 VPWR.t8 354.659
R123 VPWR.n64 VPWR.n63 320.976
R124 VPWR.n62 VPWR.n3 320.976
R125 VPWR.n5 VPWR.n4 320.976
R126 VPWR.n55 VPWR.n7 320.976
R127 VPWR.n49 VPWR.n48 320.976
R128 VPWR.n46 VPWR.n10 320.976
R129 VPWR.n12 VPWR.n11 320.976
R130 VPWR.n40 VPWR.n14 320.976
R131 VPWR.n34 VPWR.n33 320.976
R132 VPWR.n31 VPWR.n17 320.976
R133 VPWR.n25 VPWR.n24 320.976
R134 VPWR.n22 VPWR.n20 320.976
R135 VPWR.n71 VPWR.t21 257.474
R136 VPWR.n22 VPWR.n21 36.5149
R137 VPWR.n26 VPWR.n23 34.6358
R138 VPWR.n30 VPWR.n18 34.6358
R139 VPWR.n35 VPWR.n32 34.6358
R140 VPWR.n39 VPWR.n15 34.6358
R141 VPWR.n42 VPWR.n41 34.6358
R142 VPWR.n50 VPWR.n47 34.6358
R143 VPWR.n54 VPWR.n8 34.6358
R144 VPWR.n57 VPWR.n56 34.6358
R145 VPWR.n61 VPWR.n60 34.6358
R146 VPWR.n69 VPWR.n1 34.6358
R147 VPWR.n70 VPWR.n69 34.6358
R148 VPWR.n45 VPWR.n12 33.8829
R149 VPWR.n65 VPWR.n64 33.8829
R150 VPWR.n71 VPWR.n70 32.377
R151 VPWR.n46 VPWR.n45 29.3652
R152 VPWR.n65 VPWR.n62 29.3652
R153 VPWR.n41 VPWR.n40 27.8593
R154 VPWR.n63 VPWR.t23 26.5955
R155 VPWR.n63 VPWR.t16 26.5955
R156 VPWR.n3 VPWR.t18 26.5955
R157 VPWR.n3 VPWR.t22 26.5955
R158 VPWR.n4 VPWR.t25 26.5955
R159 VPWR.n4 VPWR.t17 26.5955
R160 VPWR.n7 VPWR.t20 26.5955
R161 VPWR.n7 VPWR.t24 26.5955
R162 VPWR.n48 VPWR.t3 26.5955
R163 VPWR.n48 VPWR.t19 26.5955
R164 VPWR.n10 VPWR.t10 26.5955
R165 VPWR.n10 VPWR.t4 26.5955
R166 VPWR.n11 VPWR.t13 26.5955
R167 VPWR.n11 VPWR.t12 26.5955
R168 VPWR.n14 VPWR.t15 26.5955
R169 VPWR.n14 VPWR.t14 26.5955
R170 VPWR.n33 VPWR.t5 26.5955
R171 VPWR.n33 VPWR.t1 26.5955
R172 VPWR.n17 VPWR.t9 26.5955
R173 VPWR.n17 VPWR.t7 26.5955
R174 VPWR.n24 VPWR.t0 26.5955
R175 VPWR.n24 VPWR.t11 26.5955
R176 VPWR.n20 VPWR.t6 26.5955
R177 VPWR.n20 VPWR.t2 26.5955
R178 VPWR.n26 VPWR.n25 24.8476
R179 VPWR.n50 VPWR.n49 23.3417
R180 VPWR.n60 VPWR.n5 23.3417
R181 VPWR.n34 VPWR.n15 21.8358
R182 VPWR.n31 VPWR.n30 18.824
R183 VPWR.n55 VPWR.n54 17.3181
R184 VPWR.n56 VPWR.n55 17.3181
R185 VPWR.n32 VPWR.n31 15.8123
R186 VPWR.n35 VPWR.n34 12.8005
R187 VPWR.n72 VPWR.n71 11.5593
R188 VPWR.n49 VPWR.n8 11.2946
R189 VPWR.n57 VPWR.n5 11.2946
R190 VPWR.n25 VPWR.n18 9.78874
R191 VPWR.n23 VPWR.n19 9.3005
R192 VPWR.n27 VPWR.n26 9.3005
R193 VPWR.n28 VPWR.n18 9.3005
R194 VPWR.n30 VPWR.n29 9.3005
R195 VPWR.n32 VPWR.n16 9.3005
R196 VPWR.n36 VPWR.n35 9.3005
R197 VPWR.n37 VPWR.n15 9.3005
R198 VPWR.n39 VPWR.n38 9.3005
R199 VPWR.n41 VPWR.n13 9.3005
R200 VPWR.n43 VPWR.n42 9.3005
R201 VPWR.n45 VPWR.n44 9.3005
R202 VPWR.n47 VPWR.n9 9.3005
R203 VPWR.n51 VPWR.n50 9.3005
R204 VPWR.n52 VPWR.n8 9.3005
R205 VPWR.n54 VPWR.n53 9.3005
R206 VPWR.n56 VPWR.n6 9.3005
R207 VPWR.n58 VPWR.n57 9.3005
R208 VPWR.n60 VPWR.n59 9.3005
R209 VPWR.n61 VPWR.n2 9.3005
R210 VPWR.n66 VPWR.n65 9.3005
R211 VPWR.n67 VPWR.n1 9.3005
R212 VPWR.n69 VPWR.n68 9.3005
R213 VPWR.n70 VPWR.n0 9.3005
R214 VPWR.n40 VPWR.n39 6.77697
R215 VPWR.n47 VPWR.n46 5.27109
R216 VPWR.n62 VPWR.n61 5.27109
R217 VPWR.n23 VPWR.n22 3.76521
R218 VPWR.n21 VPWR.n19 2.15642
R219 VPWR.n42 VPWR.n12 0.753441
R220 VPWR.n64 VPWR.n1 0.753441
R221 VPWR.n27 VPWR.n19 0.120292
R222 VPWR.n28 VPWR.n27 0.120292
R223 VPWR.n29 VPWR.n28 0.120292
R224 VPWR.n29 VPWR.n16 0.120292
R225 VPWR.n36 VPWR.n16 0.120292
R226 VPWR.n37 VPWR.n36 0.120292
R227 VPWR.n38 VPWR.n37 0.120292
R228 VPWR.n38 VPWR.n13 0.120292
R229 VPWR.n43 VPWR.n13 0.120292
R230 VPWR.n44 VPWR.n43 0.120292
R231 VPWR.n44 VPWR.n9 0.120292
R232 VPWR.n51 VPWR.n9 0.120292
R233 VPWR.n52 VPWR.n51 0.120292
R234 VPWR.n53 VPWR.n52 0.120292
R235 VPWR.n53 VPWR.n6 0.120292
R236 VPWR.n58 VPWR.n6 0.120292
R237 VPWR.n59 VPWR.n58 0.120292
R238 VPWR.n59 VPWR.n2 0.120292
R239 VPWR.n66 VPWR.n2 0.120292
R240 VPWR.n67 VPWR.n66 0.120292
R241 VPWR.n68 VPWR.n67 0.120292
R242 VPWR.n68 VPWR.n0 0.120292
R243 VPWR.n72 VPWR.n0 0.120292
R244 VPWR VPWR.n72 0.0213333
R245 X.n2 X.n0 244.457
R246 X.n2 X.n1 206.056
R247 X.n4 X.n3 206.056
R248 X.n6 X.n5 206.056
R249 X.n8 X.n7 206.056
R250 X.n10 X.n9 206.056
R251 X.n12 X.n11 206.056
R252 X.n14 X.n13 206.056
R253 X.n17 X.n15 137.189
R254 X.n17 X.n16 98.788
R255 X.n19 X.n18 98.788
R256 X.n21 X.n20 98.788
R257 X.n23 X.n22 98.788
R258 X.n25 X.n24 98.788
R259 X.n27 X.n26 98.788
R260 X.n29 X.n28 98.788
R261 X.n19 X.n17 38.4005
R262 X.n21 X.n19 38.4005
R263 X.n23 X.n21 38.4005
R264 X.n25 X.n23 38.4005
R265 X.n27 X.n25 38.4005
R266 X.n29 X.n27 38.4005
R267 X.n4 X.n2 38.4005
R268 X.n6 X.n4 38.4005
R269 X.n8 X.n6 38.4005
R270 X.n10 X.n8 38.4005
R271 X.n12 X.n10 38.4005
R272 X.n14 X.n12 38.4005
R273 X X.n29 27.4829
R274 X.n0 X.t3 26.5955
R275 X.n0 X.t2 26.5955
R276 X.n1 X.t11 26.5955
R277 X.n1 X.t9 26.5955
R278 X.n3 X.t13 26.5955
R279 X.n3 X.t12 26.5955
R280 X.n5 X.t0 26.5955
R281 X.n5 X.t14 26.5955
R282 X.n7 X.t6 26.5955
R283 X.n7 X.t4 26.5955
R284 X.n9 X.t10 26.5955
R285 X.n9 X.t8 26.5955
R286 X.n11 X.t1 26.5955
R287 X.n11 X.t15 26.5955
R288 X.n13 X.t7 26.5955
R289 X.n13 X.t5 26.5955
R290 X.n15 X.t24 24.9236
R291 X.n15 X.t27 24.9236
R292 X.n16 X.t22 24.9236
R293 X.n16 X.t26 24.9236
R294 X.n18 X.t21 24.9236
R295 X.n18 X.t18 24.9236
R296 X.n20 X.t20 24.9236
R297 X.n20 X.t17 24.9236
R298 X.n22 X.t30 24.9236
R299 X.n22 X.t16 24.9236
R300 X.n24 X.t29 24.9236
R301 X.n24 X.t31 24.9236
R302 X.n26 X.t25 24.9236
R303 X.n26 X.t28 24.9236
R304 X.n28 X.t23 24.9236
R305 X.n28 X.t19 24.9236
R306 X X.n14 17.4436
R307 VPB.t21 VPB.t16 556.386
R308 VPB.t5 VPB.t7 248.599
R309 VPB.t1 VPB.t5 248.599
R310 VPB.t15 VPB.t1 248.599
R311 VPB.t10 VPB.t15 248.599
R312 VPB.t8 VPB.t10 248.599
R313 VPB.t6 VPB.t8 248.599
R314 VPB.t4 VPB.t6 248.599
R315 VPB.t0 VPB.t4 248.599
R316 VPB.t14 VPB.t0 248.599
R317 VPB.t13 VPB.t14 248.599
R318 VPB.t12 VPB.t13 248.599
R319 VPB.t11 VPB.t12 248.599
R320 VPB.t9 VPB.t11 248.599
R321 VPB.t3 VPB.t9 248.599
R322 VPB.t2 VPB.t3 248.599
R323 VPB.t19 VPB.t2 248.599
R324 VPB.t20 VPB.t19 248.599
R325 VPB.t24 VPB.t20 248.599
R326 VPB.t25 VPB.t24 248.599
R327 VPB.t17 VPB.t25 248.599
R328 VPB.t18 VPB.t17 248.599
R329 VPB.t22 VPB.t18 248.599
R330 VPB.t23 VPB.t22 248.599
R331 VPB.t16 VPB.t23 248.599
R332 VPB VPB.t21 189.409
R333 VGND.n21 VGND.t7 289.651
R334 VGND.n22 VGND.n20 208.719
R335 VGND.n25 VGND.n24 208.719
R336 VGND.n31 VGND.n17 208.719
R337 VGND.n34 VGND.n33 208.719
R338 VGND.n40 VGND.n14 208.719
R339 VGND.n12 VGND.n11 208.719
R340 VGND.n46 VGND.n10 208.719
R341 VGND.n49 VGND.n48 208.719
R342 VGND.n55 VGND.n7 208.719
R343 VGND.n5 VGND.n4 208.719
R344 VGND.n62 VGND.n3 208.719
R345 VGND.n64 VGND.n63 208.719
R346 VGND.n71 VGND.t17 161.302
R347 VGND.n22 VGND.n21 36.5149
R348 VGND.n26 VGND.n23 34.6358
R349 VGND.n30 VGND.n18 34.6358
R350 VGND.n35 VGND.n32 34.6358
R351 VGND.n39 VGND.n15 34.6358
R352 VGND.n42 VGND.n41 34.6358
R353 VGND.n50 VGND.n47 34.6358
R354 VGND.n54 VGND.n8 34.6358
R355 VGND.n57 VGND.n56 34.6358
R356 VGND.n61 VGND.n60 34.6358
R357 VGND.n69 VGND.n1 34.6358
R358 VGND.n70 VGND.n69 34.6358
R359 VGND.n45 VGND.n12 33.8829
R360 VGND.n65 VGND.n64 33.8829
R361 VGND.n71 VGND.n70 32.377
R362 VGND.n46 VGND.n45 29.3652
R363 VGND.n65 VGND.n62 29.3652
R364 VGND.n41 VGND.n40 27.8593
R365 VGND.n20 VGND.t3 24.9236
R366 VGND.n20 VGND.t9 24.9236
R367 VGND.n24 VGND.t12 24.9236
R368 VGND.n24 VGND.t13 24.9236
R369 VGND.n17 VGND.t15 24.9236
R370 VGND.n17 VGND.t14 24.9236
R371 VGND.n33 VGND.t0 24.9236
R372 VGND.n33 VGND.t4 24.9236
R373 VGND.n14 VGND.t1 24.9236
R374 VGND.n14 VGND.t5 24.9236
R375 VGND.n11 VGND.t2 24.9236
R376 VGND.n11 VGND.t6 24.9236
R377 VGND.n10 VGND.t10 24.9236
R378 VGND.n10 VGND.t8 24.9236
R379 VGND.n48 VGND.t11 24.9236
R380 VGND.n48 VGND.t21 24.9236
R381 VGND.n7 VGND.t20 24.9236
R382 VGND.n7 VGND.t25 24.9236
R383 VGND.n4 VGND.t19 24.9236
R384 VGND.n4 VGND.t24 24.9236
R385 VGND.n3 VGND.t18 24.9236
R386 VGND.n3 VGND.t23 24.9236
R387 VGND.n63 VGND.t16 24.9236
R388 VGND.n63 VGND.t22 24.9236
R389 VGND.n26 VGND.n25 24.8476
R390 VGND.n50 VGND.n49 23.3417
R391 VGND.n60 VGND.n5 23.3417
R392 VGND.n34 VGND.n15 21.8358
R393 VGND.n31 VGND.n30 18.824
R394 VGND.n55 VGND.n54 17.3181
R395 VGND.n56 VGND.n55 17.3181
R396 VGND.n32 VGND.n31 15.8123
R397 VGND.n35 VGND.n34 12.8005
R398 VGND.n72 VGND.n71 11.5593
R399 VGND.n49 VGND.n8 11.2946
R400 VGND.n57 VGND.n5 11.2946
R401 VGND.n25 VGND.n18 9.78874
R402 VGND.n23 VGND.n19 9.3005
R403 VGND.n27 VGND.n26 9.3005
R404 VGND.n28 VGND.n18 9.3005
R405 VGND.n30 VGND.n29 9.3005
R406 VGND.n32 VGND.n16 9.3005
R407 VGND.n36 VGND.n35 9.3005
R408 VGND.n37 VGND.n15 9.3005
R409 VGND.n39 VGND.n38 9.3005
R410 VGND.n41 VGND.n13 9.3005
R411 VGND.n43 VGND.n42 9.3005
R412 VGND.n45 VGND.n44 9.3005
R413 VGND.n47 VGND.n9 9.3005
R414 VGND.n51 VGND.n50 9.3005
R415 VGND.n52 VGND.n8 9.3005
R416 VGND.n54 VGND.n53 9.3005
R417 VGND.n56 VGND.n6 9.3005
R418 VGND.n58 VGND.n57 9.3005
R419 VGND.n60 VGND.n59 9.3005
R420 VGND.n61 VGND.n2 9.3005
R421 VGND.n66 VGND.n65 9.3005
R422 VGND.n67 VGND.n1 9.3005
R423 VGND.n69 VGND.n68 9.3005
R424 VGND.n70 VGND.n0 9.3005
R425 VGND.n40 VGND.n39 6.77697
R426 VGND.n47 VGND.n46 5.27109
R427 VGND.n62 VGND.n61 5.27109
R428 VGND.n23 VGND.n22 3.76521
R429 VGND.n21 VGND.n19 2.15642
R430 VGND.n42 VGND.n12 0.753441
R431 VGND.n64 VGND.n1 0.753441
R432 VGND.n27 VGND.n19 0.120292
R433 VGND.n28 VGND.n27 0.120292
R434 VGND.n29 VGND.n28 0.120292
R435 VGND.n29 VGND.n16 0.120292
R436 VGND.n36 VGND.n16 0.120292
R437 VGND.n37 VGND.n36 0.120292
R438 VGND.n38 VGND.n37 0.120292
R439 VGND.n38 VGND.n13 0.120292
R440 VGND.n43 VGND.n13 0.120292
R441 VGND.n44 VGND.n43 0.120292
R442 VGND.n44 VGND.n9 0.120292
R443 VGND.n51 VGND.n9 0.120292
R444 VGND.n52 VGND.n51 0.120292
R445 VGND.n53 VGND.n52 0.120292
R446 VGND.n53 VGND.n6 0.120292
R447 VGND.n58 VGND.n6 0.120292
R448 VGND.n59 VGND.n58 0.120292
R449 VGND.n59 VGND.n2 0.120292
R450 VGND.n66 VGND.n2 0.120292
R451 VGND.n67 VGND.n66 0.120292
R452 VGND.n68 VGND.n67 0.120292
R453 VGND.n68 VGND.n0 0.120292
R454 VGND.n72 VGND.n0 0.120292
R455 VGND VGND.n72 0.0213333
R456 VNB.t17 VNB.t22 2677.02
R457 VNB.t3 VNB.t7 1196.12
R458 VNB.t9 VNB.t3 1196.12
R459 VNB.t12 VNB.t9 1196.12
R460 VNB.t13 VNB.t12 1196.12
R461 VNB.t15 VNB.t13 1196.12
R462 VNB.t14 VNB.t15 1196.12
R463 VNB.t0 VNB.t14 1196.12
R464 VNB.t4 VNB.t0 1196.12
R465 VNB.t1 VNB.t4 1196.12
R466 VNB.t5 VNB.t1 1196.12
R467 VNB.t2 VNB.t5 1196.12
R468 VNB.t6 VNB.t2 1196.12
R469 VNB.t10 VNB.t6 1196.12
R470 VNB.t8 VNB.t10 1196.12
R471 VNB.t11 VNB.t8 1196.12
R472 VNB.t21 VNB.t11 1196.12
R473 VNB.t20 VNB.t21 1196.12
R474 VNB.t25 VNB.t20 1196.12
R475 VNB.t19 VNB.t25 1196.12
R476 VNB.t24 VNB.t19 1196.12
R477 VNB.t18 VNB.t24 1196.12
R478 VNB.t23 VNB.t18 1196.12
R479 VNB.t16 VNB.t23 1196.12
R480 VNB.t22 VNB.t16 1196.12
R481 VNB VNB.t17 911.327
R482 a_215_47.t1 a_215_47.n21 271.051
R483 a_215_47.n5 a_215_47.t16 221.72
R484 a_215_47.n7 a_215_47.t17 221.72
R485 a_215_47.n9 a_215_47.t6 221.72
R486 a_215_47.n3 a_215_47.t8 221.72
R487 a_215_47.n15 a_215_47.t13 221.72
R488 a_215_47.n16 a_215_47.t14 221.72
R489 a_215_47.n21 a_215_47.n20 206.056
R490 a_215_47.n1 a_215_47.t2 176.525
R491 a_215_47.n6 a_215_47.n4 173.761
R492 a_215_47.n18 a_215_47.n17 152
R493 a_215_47.n14 a_215_47.n2 152
R494 a_215_47.n13 a_215_47.n12 152
R495 a_215_47.n11 a_215_47.n10 152
R496 a_215_47.n8 a_215_47.n4 152
R497 a_215_47.n5 a_215_47.t15 149.421
R498 a_215_47.n7 a_215_47.t12 149.421
R499 a_215_47.n9 a_215_47.t9 149.421
R500 a_215_47.n3 a_215_47.t11 149.421
R501 a_215_47.n15 a_215_47.t7 149.421
R502 a_215_47.n16 a_215_47.t10 149.421
R503 a_215_47.n1 a_215_47.n0 98.788
R504 a_215_47.n14 a_215_47.n13 60.6968
R505 a_215_47.n10 a_215_47.n3 55.3412
R506 a_215_47.n17 a_215_47.n15 51.7709
R507 a_215_47.n6 a_215_47.n5 48.2005
R508 a_215_47.n9 a_215_47.n8 41.0598
R509 a_215_47.n8 a_215_47.n7 33.919
R510 a_215_47.n19 a_215_47.n1 32.0005
R511 a_215_47.n21 a_215_47.n19 32.0005
R512 a_215_47.n7 a_215_47.n6 26.7783
R513 a_215_47.n20 a_215_47.t4 26.5955
R514 a_215_47.n20 a_215_47.t5 26.5955
R515 a_215_47.n0 a_215_47.t3 24.9236
R516 a_215_47.n0 a_215_47.t0 24.9236
R517 a_215_47.n17 a_215_47.n16 23.2079
R518 a_215_47.n11 a_215_47.n4 21.7605
R519 a_215_47.n12 a_215_47.n11 21.7605
R520 a_215_47.n12 a_215_47.n2 21.7605
R521 a_215_47.n18 a_215_47.n2 21.7605
R522 a_215_47.n19 a_215_47.n18 21.7605
R523 a_215_47.n10 a_215_47.n9 19.6375
R524 a_215_47.n15 a_215_47.n14 8.92643
R525 a_215_47.n13 a_215_47.n3 5.35606
R526 a_109_47.t1 a_109_47.n6 250.655
R527 a_109_47.n0 a_109_47.t4 221.72
R528 a_109_47.n2 a_109_47.t5 221.72
R529 a_109_47.n3 a_109_47.t7 221.72
R530 a_109_47.n5 a_109_47.n1 173.761
R531 a_109_47.n6 a_109_47.t0 156.129
R532 a_109_47.n5 a_109_47.n4 152
R533 a_109_47.n0 a_109_47.t3 149.421
R534 a_109_47.n2 a_109_47.t6 149.421
R535 a_109_47.n3 a_109_47.t2 149.421
R536 a_109_47.n1 a_109_47.n0 51.7709
R537 a_109_47.n6 a_109_47.n5 49.6005
R538 a_109_47.n4 a_109_47.n2 37.4894
R539 a_109_47.n4 a_109_47.n3 37.4894
R540 a_109_47.n2 a_109_47.n1 23.2079
R541 A.n0 A.t0 230.363
R542 A A.n0 160
R543 A.n0 A.t1 158.064
C0 VPB A 0.043416f
C1 VGND VPB 0.015325f
C2 VPB VPWR 0.237419f
C3 VGND A 0.041236f
C4 A VPWR 0.041524f
C5 VPB X 0.034218f
C6 VGND VPWR 0.245724f
C7 VGND X 1.05198f
C8 VPWR X 1.44943f
C9 VGND VNB 1.31889f
C10 X VNB 0.076881f
C11 VPWR VNB 1.13547f
C12 A VNB 0.151434f
C13 VPB VNB 2.37668f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s18_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s18_1 VPWR VGND X A VPB VNB
X0 VPWR.t1 A.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.3184 pd=1.68 as=0.265 ps=2.53 w=1 l=0.15
X1 X.t0 a_394_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.20835 ps=1.33 w=0.42 l=0.15
X2 VGND.t2 a_282_47.t2 a_394_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.20835 pd=1.33 as=0.17225 ps=1.83 w=0.65 l=0.18
X3 X.t1 a_394_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.3229 ps=1.68 w=1 l=0.15
X4 a_282_47.t1 a_27_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2173 pd=2.17 as=0.3184 ps=1.68 w=0.82 l=0.18
X5 VGND.t0 A.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.20835 pd=1.33 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 a_282_47.t0 a_27_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.20835 ps=1.33 w=0.65 l=0.18
X7 VPWR.t2 a_282_47.t3 a_394_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.3229 pd=1.68 as=0.2173 ps=2.17 w=0.82 l=0.18
R0 A.n0 A.t0 227.417
R1 A.n0 A.t1 206.093
R2 A A.n0 163.379
R3 a_27_47.t1 a_27_47.n1 371.348
R4 a_27_47.n1 a_27_47.t0 272.812
R5 a_27_47.n1 a_27_47.n0 206.398
R6 a_27_47.n0 a_27_47.t2 187.445
R7 a_27_47.n0 a_27_47.t3 124.517
R8 VPWR.n2 VPWR.n0 318.279
R9 VPWR.n2 VPWR.n1 316.774
R10 VPWR.n1 VPWR.t3 112.269
R11 VPWR.n0 VPWR.t2 108.627
R12 VPWR.n1 VPWR.t1 36.8562
R13 VPWR.n0 VPWR.t0 36.264
R14 VPWR VPWR.n2 0.161481
R15 VPB.t3 VPB.t2 594.861
R16 VPB.t2 VPB.t0 500.156
R17 VPB.t1 VPB.t3 500.156
R18 VPB VPB.t1 195.327
R19 a_394_47.t0 a_394_47.n1 405.026
R20 a_394_47.n1 a_394_47.t1 341.154
R21 a_394_47.n0 a_394_47.t3 227.417
R22 a_394_47.n0 a_394_47.t2 205.215
R23 a_394_47.n1 a_394_47.n0 152
R24 VGND.n2 VGND.n1 206.156
R25 VGND.n2 VGND.n0 205.825
R26 VGND.n1 VGND.t3 89.539
R27 VGND.n0 VGND.t2 84.9236
R28 VGND.n0 VGND.t1 51.7368
R29 VGND.n1 VGND.t0 47.1214
R30 VGND VGND.n2 0.16023
R31 X X.n0 591.227
R32 X.n2 X.n0 585
R33 X X.t0 226.517
R34 X.n0 X.t1 27.5805
R35 X X.n1 12.5161
R36 X.n1 X 6.82717
R37 X.n2 X 6.22753
R38 X X.n2 5.53564
R39 X.n1 X 4.04261
R40 VNB.t3 VNB.t2 2862.14
R41 VNB.t2 VNB.t1 2406.47
R42 VNB.t0 VNB.t3 2406.47
R43 VNB VNB.t0 939.807
R44 a_282_47.t1 a_282_47.n1 377.663
R45 a_282_47.n0 a_282_47.t3 201.838
R46 a_282_47.n1 a_282_47.t0 154.595
R47 a_282_47.n0 a_282_47.t2 132.55
R48 a_282_47.n1 a_282_47.n0 114.349
C0 VPB VGND 0.007099f
C1 A VGND 0.016568f
C2 VPWR X 0.110863f
C3 VPWR VGND 0.079827f
C4 X VGND 0.076926f
C5 VPB A 0.036819f
C6 VPB VPWR 0.081668f
C7 A VPWR 0.019256f
C8 VPB X 0.012748f
C9 VGND VNB 0.440506f
C10 X VNB 0.095068f
C11 VPWR VNB 0.364774f
C12 A VNB 0.165494f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s18_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s18_2 VNB VPB VGND VPWR A X
X0 a_227_47.t0 a_27_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.11735 ps=1.05 w=0.65 l=0.18
X1 VGND.t3 a_334_47.t2 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.59 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND.t2 a_227_47.t2 a_334_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1446 pd=1.125 as=0.17225 ps=1.83 w=0.65 l=0.18
X3 VPWR.t2 a_227_47.t3 a_334_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.21725 pd=1.475 as=0.2173 ps=2.17 w=0.82 l=0.18
X4 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1865 pd=1.4 as=0.27 ps=2.54 w=1 l=0.15
X5 X.t1 a_334_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1446 ps=1.125 w=0.42 l=0.15
X6 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.11735 pd=1.05 as=0.1134 ps=1.38 w=0.42 l=0.15
X7 X.t0 a_334_47.t4 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.21725 ps=1.475 w=1 l=0.15
X8 a_227_47.t1 a_27_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2173 pd=2.17 as=0.1865 ps=1.4 w=0.82 l=0.18
X9 VPWR.t3 a_334_47.t5 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.375 pd=2.75 as=0.14 ps=1.28 w=1 l=0.15
R0 a_27_47.t0 a_27_47.n1 376.536
R1 a_27_47.n1 a_27_47.t1 277.043
R2 a_27_47.n0 a_27_47.t3 228.585
R3 a_27_47.n1 a_27_47.n0 152
R4 a_27_47.n0 a_27_47.t2 144.236
R5 VGND.n4 VGND.t3 279.418
R6 VGND.n10 VGND.n9 200.516
R7 VGND.n3 VGND.n2 198.839
R8 VGND.n2 VGND.t4 71.4291
R9 VGND.n9 VGND.t1 55.7148
R10 VGND.n2 VGND.t2 44.5719
R11 VGND.n9 VGND.t0 43.9126
R12 VGND.n7 VGND.n1 34.6358
R13 VGND.n8 VGND.n7 34.6358
R14 VGND.n10 VGND.n8 17.6946
R15 VGND.n5 VGND.n1 9.3005
R16 VGND.n7 VGND.n6 9.3005
R17 VGND.n8 VGND.n0 9.3005
R18 VGND.n11 VGND.n10 7.37348
R19 VGND.n4 VGND.n3 7.21628
R20 VGND.n3 VGND.n1 7.15344
R21 VGND.n5 VGND.n4 0.509445
R22 VGND.n11 VGND.n0 0.145304
R23 VGND.n6 VGND.n5 0.120292
R24 VGND.n6 VGND.n0 0.120292
R25 VGND VGND.n11 0.116797
R26 a_227_47.t1 a_227_47.n1 376.832
R27 a_227_47.n1 a_227_47.t0 254.155
R28 a_227_47.n0 a_227_47.t3 208.868
R29 a_227_47.n0 a_227_47.t2 124.517
R30 a_227_47.n1 a_227_47.n0 121.129
R31 VNB.t0 VNB.t2 2790.94
R32 VNB.t2 VNB.t4 1822.65
R33 VNB.t1 VNB.t0 1609.06
R34 VNB.t4 VNB.t3 1224.6
R35 VNB VNB.t1 939.807
R36 a_334_47.t1 a_334_47.n2 399.522
R37 a_334_47.n2 a_334_47.t0 276.228
R38 a_334_47.n1 a_334_47.t5 221.72
R39 a_334_47.n0 a_334_47.t4 221.72
R40 a_334_47.n1 a_334_47.t2 186.374
R41 a_334_47.n0 a_334_47.t3 186.374
R42 a_334_47.n2 a_334_47.n0 168.189
R43 a_334_47.n0 a_334_47.n1 76.7635
R44 X.n0 X 590.298
R45 X.n1 X.n0 585
R46 X.n3 X.n2 185
R47 X X.n3 88.9364
R48 X.n2 X.t2 40.0005
R49 X.n2 X.t1 40.0005
R50 X.n0 X.t3 27.5805
R51 X.n0 X.t0 27.5805
R52 X X.n1 5.29705
R53 X.n1 X 4.70855
R54 X.n3 X 0.28814
R55 VPWR.n5 VPWR.t3 369.036
R56 VPWR.n10 VPWR.n1 311.858
R57 VPWR.n4 VPWR.n3 307.899
R58 VPWR.n3 VPWR.t2 56.4578
R59 VPWR.n3 VPWR.t4 54.4632
R60 VPWR.n1 VPWR.t0 47.2559
R61 VPWR.n1 VPWR.t1 45.6468
R62 VPWR.n8 VPWR.n2 34.6358
R63 VPWR.n9 VPWR.n8 34.6358
R64 VPWR.n10 VPWR.n9 16.5652
R65 VPWR.n6 VPWR.n2 9.3005
R66 VPWR.n8 VPWR.n7 9.3005
R67 VPWR.n9 VPWR.n0 9.3005
R68 VPWR.n11 VPWR.n10 7.42022
R69 VPWR.n5 VPWR.n4 7.18504
R70 VPWR.n4 VPWR.n2 4.51815
R71 VPWR.n6 VPWR.n5 0.515269
R72 VPWR.n11 VPWR.n0 0.14471
R73 VPWR.n7 VPWR.n6 0.120292
R74 VPWR.n7 VPWR.n0 0.120292
R75 VPWR VPWR.n11 0.117399
R76 VPB.t1 VPB.t2 580.062
R77 VPB.t2 VPB.t4 378.817
R78 VPB.t0 VPB.t1 334.425
R79 VPB.t4 VPB.t3 254.518
R80 VPB VPB.t0 195.327
R81 A.n0 A.t0 240.012
R82 A.n0 A.t1 204.666
R83 A A.n0 166.587
C0 A VPWR 0.019195f
C1 VPB X 0.006377f
C2 VPB VGND 0.009395f
C3 A VGND 0.017169f
C4 VPWR X 0.193393f
C5 VPWR VGND 0.086461f
C6 X VGND 0.116813f
C7 VPB A 0.034491f
C8 VPB VPWR 0.08852f
C9 VGND VNB 0.46727f
C10 X VNB 0.042103f
C11 VPWR VNB 0.400673f
C12 A VNB 0.161118f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s25_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 VNB VPB VPWR VGND A X
X0 a_244_47.t1 a_27_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2173 pd=2.17 as=0.19265 ps=1.415 w=0.82 l=0.25
X1 VPWR.t1 a_244_47.t2 a_355_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2726 pd=1.61 as=0.2173 ps=2.17 w=0.82 l=0.25
X2 X.t1 a_355_47.t2 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.495 pd=2.99 as=0.2726 ps=1.61 w=1 l=0.15
X3 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.19265 pd=1.415 as=0.27 ps=2.54 w=1 l=0.15
X4 VGND.t2 A.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1228 pd=1.065 as=0.1134 ps=1.38 w=0.42 l=0.15
X5 VGND.t1 a_244_47.t3 a_355_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1856 pd=1.26 as=0.17225 ps=1.83 w=0.65 l=0.25
X6 X.t0 a_355_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.2079 pd=1.83 as=0.1856 ps=1.26 w=0.42 l=0.15
X7 a_244_47.t0 a_27_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1228 ps=1.065 w=0.65 l=0.25
R0 a_27_47.t0 a_27_47.n1 370.902
R1 a_27_47.n1 a_27_47.t1 271.635
R2 a_27_47.n0 a_27_47.t2 165.006
R3 a_27_47.n1 a_27_47.n0 152
R4 a_27_47.n0 a_27_47.t3 104.275
R5 VPWR.n2 VPWR.n1 316.625
R6 VPWR.n2 VPWR.n0 307.483
R7 VPWR.n0 VPWR.t1 93.6956
R8 VPWR.n1 VPWR.t3 50.4517
R9 VPWR.n0 VPWR.t2 49.6583
R10 VPWR.n1 VPWR.t0 46.0547
R11 VPWR VPWR.n2 0.173195
R12 a_244_47.t1 a_244_47.n1 373.861
R13 a_244_47.n1 a_244_47.t0 285.937
R14 a_244_47.n0 a_244_47.t2 150.385
R15 a_244_47.n1 a_244_47.n0 123.716
R16 a_244_47.n0 a_244_47.t3 89.6525
R17 VPB.t3 VPB.t2 633.333
R18 VPB.t2 VPB.t1 479.44
R19 VPB.t0 VPB.t3 364.019
R20 VPB VPB.t0 195.327
R21 a_355_47.t1 a_355_47.n1 413.627
R22 a_355_47.n1 a_355_47.t0 288.815
R23 a_355_47.n0 a_355_47.t2 241.536
R24 a_355_47.n0 a_355_47.t3 206.19
R25 a_355_47.n1 a_355_47.n0 152
R26 X.n0 X 589
R27 X.n1 X.n0 585
R28 X X.t0 225.553
R29 X.n0 X.t1 27.5805
R30 X.n2 X 5.02907
R31 X X.n2 4.20872
R32 X X.n1 4.0005
R33 X.n1 X 3.77193
R34 X.n2 X 2.74336
R35 A.n0 A.t0 235.98
R36 A.n0 A.t1 200.633
R37 A A.n0 160.882
R38 VGND.n2 VGND.n0 206.192
R39 VGND.n2 VGND.n1 192.191
R40 VGND.n1 VGND.t1 72.0005
R41 VGND.n0 VGND.t2 54.2862
R42 VGND.n1 VGND.t0 51.7368
R43 VGND.n0 VGND.t3 48.6159
R44 VGND VGND.n2 0.166916
R45 VNB.t3 VNB.t1 3047.25
R46 VNB.t1 VNB.t0 2306.8
R47 VNB.t2 VNB.t3 1751.46
R48 VNB VNB.t2 939.807
C0 VPB A 0.038194f
C1 VPB VPWR 0.079396f
C2 A VPWR 0.019203f
C3 VPB X 0.01394f
C4 VPB VGND 0.007517f
C5 A VGND 0.017771f
C6 VPWR X 0.131051f
C7 VPWR VGND 0.075125f
C8 X VGND 0.106391f
C9 VGND VNB 0.439033f
C10 X VNB 0.101906f
C11 VPWR VNB 0.364864f
C12 A VNB 0.167891f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s25_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s25_2 VNB VPB VPWR VGND A X
X0 X.t3 a_331_47.t2 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.097 ps=0.975 w=0.42 l=0.15
X1 VPWR.t4 A.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND.t0 a_225_47.t2 a_331_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.25
X3 VPWR.t3 a_331_47.t3 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.175 ps=1.35 w=1 l=0.15
X4 VGND.t3 A.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 VPWR.t1 a_225_47.t3 a_331_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.325 as=0.2132 ps=2.16 w=0.82 l=0.25
X6 a_225_47.t0 a_27_47.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.25
X7 X.t0 a_331_47.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.15575 ps=1.325 w=1 l=0.15
X8 a_225_47.t1 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=2.16 as=0.15575 ps=1.325 w=0.82 l=0.25
X9 VGND.t1 a_331_47.t5 X.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1407 pd=1.51 as=0.0735 ps=0.77 w=0.42 l=0.15
R0 a_331_47.t1 a_331_47.n2 444.337
R1 a_331_47.n2 a_331_47.t0 317.281
R2 a_331_47.n0 a_331_47.t3 207.261
R3 a_331_47.n1 a_331_47.t4 207.261
R4 a_331_47.n0 a_331_47.t5 173.52
R5 a_331_47.n1 a_331_47.t2 173.52
R6 a_331_47.n2 a_331_47.n1 159.469
R7 a_331_47.n1 a_331_47.n0 67.8878
R8 VGND.n4 VGND.t1 266.692
R9 VGND.n10 VGND.n9 199.934
R10 VGND.n3 VGND.n2 199.739
R11 VGND.n2 VGND.t2 54.2862
R12 VGND.n9 VGND.t3 54.2862
R13 VGND.n7 VGND.n1 34.6358
R14 VGND.n8 VGND.n7 34.6358
R15 VGND.n2 VGND.t0 25.9346
R16 VGND.n9 VGND.t4 25.9346
R17 VGND.n10 VGND.n8 18.4476
R18 VGND.n4 VGND.n3 12.0788
R19 VGND.n8 VGND.n0 9.3005
R20 VGND.n7 VGND.n6 9.3005
R21 VGND.n5 VGND.n1 9.3005
R22 VGND.n11 VGND.n10 7.34101
R23 VGND.n3 VGND.n1 4.89462
R24 VGND.n5 VGND.n4 0.546561
R25 VGND.n11 VGND.n0 0.145717
R26 VGND.n6 VGND.n5 0.120292
R27 VGND.n6 VGND.n0 0.120292
R28 VGND VGND.n11 0.117681
R29 X X.n0 591.696
R30 X.n3 X.n0 585
R31 X.n2 X.n1 185
R32 X.n1 X.t3 61.4291
R33 X.n0 X.t0 42.3555
R34 X.n1 X.t2 38.5719
R35 X.n0 X.t1 26.5955
R36 X X.n2 14.8468
R37 X X.n3 13.1943
R38 X.n2 X 0.985115
R39 X.n3 X 0.197423
R40 VNB.t4 VNB.t0 2961.81
R41 VNB.t0 VNB.t2 1495.15
R42 VNB.t3 VNB.t4 1495.15
R43 VNB.t2 VNB.t1 1423.95
R44 VNB VNB.t3 939.807
R45 A.n0 A.t0 236.18
R46 A.n0 A.t1 196.452
R47 A.n1 A.n0 152
R48 A.n1 A 8.89806
R49 A A.n1 1.71757
R50 a_27_47.t0 a_27_47.n1 383.807
R51 a_27_47.n1 a_27_47.t1 288.111
R52 a_27_47.n0 a_27_47.t3 170.256
R53 a_27_47.n1 a_27_47.n0 152
R54 a_27_47.n0 a_27_47.t2 109.523
R55 VPWR.n10 VPWR.n1 599.74
R56 VPWR.n5 VPWR.t3 359.997
R57 VPWR.n4 VPWR.n3 310.502
R58 VPWR.n1 VPWR.t4 42.451
R59 VPWR.n3 VPWR.t2 42.451
R60 VPWR.n8 VPWR.n2 34.6358
R61 VPWR.n9 VPWR.n8 34.6358
R62 VPWR.n1 VPWR.t0 32.4334
R63 VPWR.n3 VPWR.t1 32.4334
R64 VPWR.n10 VPWR.n9 18.4476
R65 VPWR.n5 VPWR.n4 12.0788
R66 VPWR.n6 VPWR.n2 9.3005
R67 VPWR.n8 VPWR.n7 9.3005
R68 VPWR.n9 VPWR.n0 9.3005
R69 VPWR.n11 VPWR.n10 7.34101
R70 VPWR.n4 VPWR.n2 4.89462
R71 VPWR.n6 VPWR.n5 0.546561
R72 VPWR.n11 VPWR.n0 0.145717
R73 VPWR.n7 VPWR.n6 0.120292
R74 VPWR.n7 VPWR.n0 0.120292
R75 VPWR VPWR.n11 0.117681
R76 VPB.t0 VPB.t1 615.577
R77 VPB.t1 VPB.t2 310.748
R78 VPB.t4 VPB.t0 310.748
R79 VPB.t2 VPB.t3 295.95
R80 VPB VPB.t4 195.327
R81 a_225_47.t1 a_225_47.n1 415.272
R82 a_225_47.n1 a_225_47.t0 232.905
R83 a_225_47.n0 a_225_47.t3 144.601
R84 a_225_47.n1 a_225_47.n0 106.916
R85 a_225_47.n0 a_225_47.t2 83.8685
C0 VPB A 0.037074f
C1 VPB VPWR 0.089946f
C2 VPB X 0.007725f
C3 A VPWR 0.019486f
C4 VPB VGND 0.007938f
C5 A VGND 0.018073f
C6 VPWR X 0.182026f
C7 VPWR VGND 0.07686f
C8 X VGND 0.119053f
C9 VGND VNB 0.459855f
C10 X VNB 0.058352f
C11 VPWR VNB 0.399828f
C12 A VNB 0.176436f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s50_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 VNB VPB VGND VPWR A X
X0 a_283_47.t1 a_27_47.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2173 pd=2.17 as=0.1701 ps=1.36 w=0.82 l=0.5
X1 VPWR.t0 A.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1701 pd=1.36 as=0.27 ps=2.54 w=1 l=0.15
X2 VPWR.t3 a_283_47.t2 a_390_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.325 as=0.2173 ps=2.17 w=0.82 l=0.5
X3 VGND.t3 a_283_47.t3 a_390_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.17225 ps=1.83 w=0.65 l=0.5
X4 X.t1 a_390_47.t2 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.355 pd=2.71 as=0.15575 ps=1.325 w=1 l=0.15
X5 VGND.t0 A.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10435 pd=1.01 as=0.1134 ps=1.38 w=0.42 l=0.15
X6 a_283_47.t0 a_27_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10435 ps=1.01 w=0.65 l=0.5
X7 X.t0 a_390_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1491 pd=1.55 as=0.097 ps=0.975 w=0.42 l=0.15
R0 a_27_47.t1 a_27_47.n1 373.57
R1 a_27_47.n1 a_27_47.t0 274.204
R2 a_27_47.n1 a_27_47.n0 152
R3 a_27_47.n0 a_27_47.t2 88.2065
R4 a_27_47.n0 a_27_47.t3 57.8405
R5 VPWR.n2 VPWR.n0 317.854
R6 VPWR.n2 VPWR.n1 317.5
R7 VPWR.n1 VPWR.t0 47.2559
R8 VPWR.n0 VPWR.t2 41.2498
R9 VPWR.n1 VPWR.t1 36.0371
R10 VPWR.n0 VPWR.t3 33.6346
R11 VPWR VPWR.n2 0.161102
R12 a_283_47.t1 a_283_47.n1 357.372
R13 a_283_47.n1 a_283_47.t0 237.718
R14 a_283_47.n1 a_283_47.n0 194.657
R15 a_283_47.n0 a_283_47.t2 88.2065
R16 a_283_47.n0 a_283_47.t3 57.8405
R17 VPB.t1 VPB.t2 769.471
R18 VPB.t0 VPB.t1 405.452
R19 VPB.t2 VPB.t3 384.736
R20 VPB VPB.t0 195.327
R21 A.n0 A.t0 237.558
R22 A.n0 A.t1 203.13
R23 A A.n0 165.099
R24 a_390_47.t1 a_390_47.n1 381.88
R25 a_390_47.n1 a_390_47.t0 256.656
R26 a_390_47.n0 a_390_47.t2 241.536
R27 a_390_47.n0 a_390_47.t3 206.19
R28 a_390_47.n1 a_390_47.n0 174.498
R29 VGND.n2 VGND.n0 207.871
R30 VGND.n2 VGND.n1 207.549
R31 VGND.n1 VGND.t0 55.7148
R32 VGND.n0 VGND.t1 52.8576
R33 VGND.n1 VGND.t2 34.506
R34 VGND.n0 VGND.t3 27.3631
R35 VGND VGND.n2 0.159137
R36 VNB.t2 VNB.t3 3702.27
R37 VNB.t0 VNB.t2 1950.81
R38 VNB.t3 VNB.t1 1851.13
R39 VNB VNB.t0 939.807
R40 X.n0 X 590.532
R41 X.n1 X.n0 585
R42 X.n2 X.t0 229.286
R43 X.n0 X.t1 30.5355
R44 X X.n2 12.8795
R45 X X.n1 5.53136
R46 X.n1 X 5.21532
R47 X.n2 X 0.316549
C0 VPWR X 0.111102f
C1 A VGND 0.017183f
C2 VPWR VGND 0.074926f
C3 X VGND 0.085045f
C4 VPB A 0.034868f
C5 VPB VPWR 0.078949f
C6 A VPWR 0.019195f
C7 VPB X 0.01322f
C8 VPB VGND 0.007266f
C9 VGND VNB 0.439163f
C10 X VNB 0.097664f
C11 VPWR VNB 0.36659f
C12 A VNB 0.162604f
C13 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s50_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 VNB VPB VGND VPWR A X
X0 VPWR.t2 a_283_47.t2 a_390_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1578 pd=1.33 as=0.2132 ps=2.16 w=0.82 l=0.5
X1 a_283_47.t0 a_27_47.t2 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2173 pd=2.17 as=0.1701 ps=1.36 w=0.82 l=0.5
X2 VPWR.t3 a_390_47.t2 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.1375 ps=1.275 w=1 l=0.15
X3 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1701 pd=1.36 as=0.27 ps=2.54 w=1 l=0.15
X4 X.t2 a_390_47.t3 VPWR.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.1578 ps=1.33 w=1 l=0.15
X5 VGND.t2 a_283_47.t3 a_390_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.09805 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.5
X6 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10435 pd=1.01 as=0.1134 ps=1.38 w=0.42 l=0.15
X7 VGND.t4 a_390_47.t4 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1638 pd=1.62 as=0.05775 ps=0.695 w=0.42 l=0.15
X8 a_283_47.t1 a_27_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10435 ps=1.01 w=0.65 l=0.5
X9 X.t0 a_390_47.t5 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.09805 ps=0.98 w=0.42 l=0.15
R0 a_283_47.t0 a_283_47.n1 375.146
R1 a_283_47.n1 a_283_47.t1 240.79
R2 a_283_47.n1 a_283_47.n0 196.012
R3 a_283_47.n0 a_283_47.t2 88.2065
R4 a_283_47.n0 a_283_47.t3 57.8405
R5 a_390_47.t1 a_390_47.n2 385.106
R6 a_390_47.n1 a_390_47.t3 308.481
R7 a_390_47.n1 a_390_47.t5 273.134
R8 a_390_47.n2 a_390_47.t0 259.091
R9 a_390_47.n0 a_390_47.t2 221.72
R10 a_390_47.n0 a_390_47.t4 186.374
R11 a_390_47.n2 a_390_47.n1 171.201
R12 a_390_47.n1 a_390_47.n0 86.582
R13 VPWR.n3 VPWR.t3 376.341
R14 VPWR.n5 VPWR.n4 311.858
R15 VPWR.n12 VPWR.n1 311.858
R16 VPWR.n1 VPWR.t0 47.2559
R17 VPWR.n4 VPWR.t4 42.451
R18 VPWR.n1 VPWR.t1 36.0371
R19 VPWR.n6 VPWR.n2 34.6358
R20 VPWR.n10 VPWR.n2 34.6358
R21 VPWR.n11 VPWR.n10 34.6358
R22 VPWR.n4 VPWR.t2 33.6346
R23 VPWR.n12 VPWR.n11 16.5652
R24 VPWR.n6 VPWR.n5 11.6711
R25 VPWR.n7 VPWR.n6 9.3005
R26 VPWR.n8 VPWR.n2 9.3005
R27 VPWR.n10 VPWR.n9 9.3005
R28 VPWR.n11 VPWR.n0 9.3005
R29 VPWR.n13 VPWR.n12 7.42022
R30 VPWR.n5 VPWR.n3 7.16456
R31 VPWR.n7 VPWR.n3 0.511327
R32 VPWR.n13 VPWR.n0 0.14471
R33 VPWR.n8 VPWR.n7 0.120292
R34 VPWR.n9 VPWR.n8 0.120292
R35 VPWR.n9 VPWR.n0 0.120292
R36 VPWR VPWR.n13 0.117399
R37 VPB.t1 VPB.t2 766.511
R38 VPB.t0 VPB.t1 405.452
R39 VPB.t2 VPB.t3 387.695
R40 VPB.t3 VPB.t4 251.559
R41 VPB VPB.t0 195.327
R42 a_27_47.t0 a_27_47.n1 381.271
R43 a_27_47.n1 a_27_47.t1 281.692
R44 a_27_47.n0 a_27_47.t2 88.2065
R45 a_27_47.n1 a_27_47.n0 76.0005
R46 a_27_47.n0 a_27_47.t3 57.8405
R47 X.n0 X 590.091
R48 X.n1 X.n0 585
R49 X.n4 X.n3 185
R50 X.n3 X.t0 40.0005
R51 X.n3 X.t1 38.5719
R52 X.n0 X.t2 27.5805
R53 X.n0 X.t3 26.5955
R54 X X.n4 10.6602
R55 X.n2 X 7.41868
R56 X X.n1 5.09141
R57 X.n1 X 4.8005
R58 X X.n2 3.88621
R59 X.n2 X 2.47323
R60 X.n4 X 1.30959
R61 A.n0 A.t0 235.763
R62 A.n0 A.t1 200.417
R63 A A.n0 162.058
R64 VGND.n2 VGND.t4 290.932
R65 VGND.n12 VGND.n11 201.486
R66 VGND.n4 VGND.n3 200.516
R67 VGND.n11 VGND.t0 55.7148
R68 VGND.n3 VGND.t3 54.2862
R69 VGND.n5 VGND.n1 34.6358
R70 VGND.n9 VGND.n1 34.6358
R71 VGND.n10 VGND.n9 34.6358
R72 VGND.n11 VGND.t1 34.506
R73 VGND.n3 VGND.t2 27.3631
R74 VGND.n12 VGND.n10 17.6946
R75 VGND.n5 VGND.n4 11.6711
R76 VGND.n6 VGND.n5 9.3005
R77 VGND.n7 VGND.n1 9.3005
R78 VGND.n9 VGND.n8 9.3005
R79 VGND.n10 VGND.n0 9.3005
R80 VGND.n13 VGND.n12 7.37348
R81 VGND.n4 VGND.n2 7.16456
R82 VGND.n6 VGND.n2 0.511327
R83 VGND.n13 VGND.n0 0.145304
R84 VGND.n7 VGND.n6 0.120292
R85 VGND.n8 VGND.n7 0.120292
R86 VGND.n8 VGND.n0 0.120292
R87 VGND VGND.n13 0.116797
R88 VNB.t1 VNB.t2 3688.03
R89 VNB.t0 VNB.t1 1950.81
R90 VNB.t2 VNB.t3 1865.37
R91 VNB.t3 VNB.t4 1210.36
R92 VNB VNB.t0 939.807
C0 VPB A 0.037279f
C1 VPB VPWR 0.093567f
C2 VPB X 0.008283f
C3 A VPWR 0.019341f
C4 VPB VGND 0.009784f
C5 A VGND 0.0174f
C6 VPWR X 0.18123f
C7 VPWR VGND 0.09342f
C8 X VGND 0.116559f
C9 VGND VNB 0.508583f
C10 X VNB 0.047975f
C11 VPWR VNB 0.432988f
C12 A VNB 0.16658f
C13 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_1 VPB VNB VGND VPWR A Y
X0 Y.t2 A.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2184 ps=2.2 w=0.84 l=0.15
X1 VGND.t0 A.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR.t1 A.t2 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=2.24 as=0.1134 ps=1.11 w=0.84 l=0.15
R0 A A.n1 283.014
R1 A.n0 A.t2 231.907
R2 A.n1 A.t0 231.361
R3 A.n0 A.t1 170.308
R4 A.n1 A.n0 54.0627
R5 VPWR.n0 VPWR.t0 420.894
R6 VPWR.n0 VPWR.t1 412.313
R7 VPWR VPWR.n0 0.491159
R8 Y Y.n0 312.298
R9 Y Y.t0 236.453
R10 Y.n0 Y.t1 31.6612
R11 Y.n0 Y.t2 31.6612
R12 VPB.t1 VPB.t0 248.599
R13 VPB VPB.t1 192.369
R14 VGND VGND.t0 250.06
R15 VNB VNB.t0 2107.44
C0 Y VPB 0.013031f
C1 Y A 0.154012f
C2 VGND VPB 0.005364f
C3 VGND A 0.042592f
C4 Y VPWR 0.200797f
C5 VGND VPWR 0.031792f
C6 Y VGND 0.110165f
C7 VPB A 0.09475f
C8 VPB VPWR 0.050631f
C9 A VPWR 0.051918f
C10 VGND VNB 0.225418f
C11 Y VNB 0.067492f
C12 VPWR VNB 0.233909f
C13 A VNB 0.30727f
C14 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_2 VNB VPB VPWR VGND A Y
X0 Y.t4 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 Y.t2 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR.t1 A.t2 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND.t0 A.t3 Y.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR.t0 A.t4 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n1 A.t4 221.72
R1 A.n0 A.t1 221.72
R2 A.n7 A.t2 218.507
R3 A.n1 A.t3 189.052
R4 A.n2 A.t0 183.161
R5 A.n8 A.n7 181.087
R6 A.n4 A.n3 152
R7 A.n6 A.n5 152
R8 A.n3 A.n1 63.2789
R9 A.n6 A.n0 45.6184
R10 A.n7 A.n6 27.9589
R11 A.n5 A.n4 19.3427
R12 A.n8 A 16.2138
R13 A.n3 A.n2 10.3291
R14 A A.n8 9.95606
R15 A.n4 A 3.69828
R16 A.n5 A 3.12939
R17 A.n2 A.n0 2.58264
R18 VGND.n0 VGND.t1 249.679
R19 VGND.n0 VGND.t0 245.364
R20 VGND VGND.n0 0.591777
R21 Y.n2 Y.t1 436.959
R22 Y.n2 Y.n1 311.849
R23 Y.n3 Y.n0 222.707
R24 Y.n0 Y.t3 40.0005
R25 Y.n0 Y.t4 40.0005
R26 Y.n1 Y.t0 27.5805
R27 Y.n1 Y.t2 27.5805
R28 Y Y.n2 20.0072
R29 Y.n3 Y 13.4862
R30 Y Y.n3 2.05764
R31 VNB VNB.t1 2264.08
R32 VNB.t1 VNB.t0 1224.6
R33 VPWR.n1 VPWR.t0 351.911
R34 VPWR.n1 VPWR.n0 322.545
R35 VPWR.n0 VPWR.t2 27.5805
R36 VPWR.n0 VPWR.t1 27.5805
R37 VPWR VPWR.n1 0.564421
R38 VPB.t2 VPB.t0 254.518
R39 VPB.t1 VPB.t2 254.518
R40 VPB VPB.t1 207.166
C0 VPWR VGND 0.037876f
C1 VPB A 0.10832f
C2 VPB Y 0.019743f
C3 VPB VPWR 0.049692f
C4 A Y 0.239306f
C5 A VPWR 0.068296f
C6 VPB VGND 0.005436f
C7 A VGND 0.074863f
C8 Y VPWR 0.297003f
C9 Y VGND 0.12414f
C10 VGND VNB 0.292563f
C11 VPWR VNB 0.235802f
C12 Y VNB 0.109357f
C13 A VNB 0.373936f
C14 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_4 VNB VPB VPWR VGND A Y
X0 Y.t9 A.t0 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND.t3 A.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1659 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND.t2 A.t2 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR.t4 A.t3 Y.t8 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR.t3 A.t4 Y.t7 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y.t1 A.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y.t6 A.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y.t0 A.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1386 ps=1.5 w=0.42 l=0.15
X8 Y.t5 A.t8 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR.t0 A.t9 Y.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n2 A.t4 276.168
R1 A.n8 A.t6 247.606
R2 A.n3 A.t0 221.72
R3 A.n5 A.t9 221.72
R4 A.n13 A.t8 221.72
R5 A.n7 A.t3 221.72
R6 A.n3 A.t1 186.374
R7 A.n5 A.t5 186.374
R8 A.n13 A.t2 186.374
R9 A.n7 A.t7 186.374
R10 A.n2 A.n1 152
R11 A.n4 A.n0 152
R12 A.n15 A.n14 152
R13 A.n12 A.n11 152
R14 A.n10 A.n6 152
R15 A.n9 A.n8 152
R16 A.n12 A.n6 60.6968
R17 A.n14 A.n13 54.4486
R18 A.n8 A.n7 50.8783
R19 A.n4 A.n3 38.382
R20 A.n5 A.n4 38.382
R21 A.n3 A.n2 22.3153
R22 A.n14 A.n5 22.3153
R23 A.n1 A.n0 19.3427
R24 A.n10 A.n9 19.3427
R25 A A.n15 17.3516
R26 A.n11 A 15.6449
R27 A.n11 A 10.5249
R28 A.n7 A.n6 9.81902
R29 A.n15 A 8.81828
R30 A.n13 A.n12 6.24865
R31 A.n1 A 4.83606
R32 A A.n10 3.69828
R33 A.n9 A 3.12939
R34 A A.n0 1.99161
R35 VPWR.n5 VPWR.t3 343.014
R36 VPWR.n10 VPWR.t2 338.598
R37 VPWR.n8 VPWR.n2 317.058
R38 VPWR.n4 VPWR.n3 317.058
R39 VPWR.n2 VPWR.t1 27.5805
R40 VPWR.n2 VPWR.t4 27.5805
R41 VPWR.n3 VPWR.t5 27.5805
R42 VPWR.n3 VPWR.t0 27.5805
R43 VPWR.n9 VPWR.n8 25.6005
R44 VPWR.n8 VPWR.n7 24.0946
R45 VPWR.n7 VPWR.n4 21.0829
R46 VPWR.n10 VPWR.n9 19.577
R47 VPWR.n7 VPWR.n6 9.3005
R48 VPWR.n8 VPWR.n1 9.3005
R49 VPWR.n9 VPWR.n0 9.3005
R50 VPWR.n11 VPWR.n10 9.3005
R51 VPWR.n5 VPWR.n4 6.83453
R52 VPWR.n6 VPWR.n5 0.660185
R53 VPWR.n6 VPWR.n1 0.120292
R54 VPWR.n1 VPWR.n0 0.120292
R55 VPWR.n11 VPWR.n0 0.120292
R56 VPWR VPWR.n11 0.0226354
R57 Y.n5 Y.n4 312.226
R58 Y.n7 Y.n6 312.226
R59 Y.n9 Y.n8 311.849
R60 Y.n1 Y.n0 203.322
R61 Y.n3 Y.n2 202.97
R62 Y.n5 Y.n3 137.036
R63 Y.n10 Y.n1 51.9534
R64 Y.n7 Y.n5 45.5534
R65 Y.n3 Y.n1 45.177
R66 Y.n9 Y.n7 45.177
R67 Y.n0 Y.t3 40.0005
R68 Y.n0 Y.t1 40.0005
R69 Y.n2 Y.t2 40.0005
R70 Y.n2 Y.t0 40.0005
R71 Y.n4 Y.t8 27.5805
R72 Y.n4 Y.t6 27.5805
R73 Y.n6 Y.t4 27.5805
R74 Y.n6 Y.t5 27.5805
R75 Y.n8 Y.t7 27.5805
R76 Y.n8 Y.t9 27.5805
R77 Y Y.n9 23.4672
R78 Y.n10 Y 12.5872
R79 Y Y.n10 1.9205
R80 VPB.t5 VPB.t3 254.518
R81 VPB.t0 VPB.t5 254.518
R82 VPB.t1 VPB.t0 254.518
R83 VPB.t4 VPB.t1 254.518
R84 VPB.t2 VPB.t4 254.518
R85 VPB VPB.t2 219.004
R86 VGND.n1 VGND.t3 247.148
R87 VGND.n5 VGND.t0 241.923
R88 VGND.n3 VGND.n2 204.201
R89 VGND.n2 VGND.t1 40.0005
R90 VGND.n2 VGND.t2 40.0005
R91 VGND.n4 VGND.n3 23.3417
R92 VGND.n5 VGND.n4 21.8358
R93 VGND.n4 VGND.n0 9.3005
R94 VGND.n6 VGND.n5 7.30743
R95 VGND.n3 VGND.n1 6.81041
R96 VGND.n1 VGND.n0 0.58231
R97 VGND.n6 VGND.n0 0.146144
R98 VGND VGND.n6 0.117248
R99 VNB VNB.t0 2278.32
R100 VNB.t1 VNB.t3 1224.6
R101 VNB.t2 VNB.t1 1224.6
R102 VNB.t0 VNB.t2 1224.6
C0 A Y 0.619963f
C1 VPB VGND 0.005933f
C2 A VGND 0.085045f
C3 VPWR Y 0.577663f
C4 VPWR VGND 0.066899f
C5 Y VGND 0.318259f
C6 VPB A 0.192877f
C7 VPB VPWR 0.075396f
C8 VPB Y 0.024482f
C9 A VPWR 0.132942f
C10 VGND VNB 0.426146f
C11 Y VNB 0.144678f
C12 VPWR VNB 0.369651f
C13 A VNB 0.602468f
C14 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfbbn_1 VGND VPWR VPB VNB Q Q_N RESET_B SET_B D CLK_N
X0 a_791_47.t0 SET_B.t0 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09735 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1 a_1555_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1094 pd=1.03 as=0.07035 ps=0.755 w=0.42 l=0.15
X2 VPWR.t6 RESET_B.t0 a_941_21.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1539 pd=1.335 as=0.1696 ps=1.81 w=0.64 l=0.15
X3 a_1415_315.t1 SET_B.t1 VPWR.t11 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1323 pd=1.22 as=0.09555 ps=0.875 w=0.42 l=0.15
X4 a_791_47.t1 a_941_21.t1 a_647_21.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VGND.t0 a_1415_315.t2 a_1363_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X6 a_1340_413.t0 a_27_47.t2 a_1256_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.07875 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR.t13 CLK_N.t0 a_27_47.t0 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_381_47.t1 D.t0 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_473_413.t2 a_193_47.t2 a_381_47.t0 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X10 VPWR.t0 a_1415_315.t3 a_2136_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_1256_413.t0 a_193_47.t3 a_1112_329.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1743 ps=1.41 w=0.42 l=0.15
X12 a_581_47.t1 a_27_47.t3 a_473_413.t1 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X13 a_647_21.t2 a_473_413.t4 a_791_47.t2 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.09735 ps=0.97 w=0.64 l=0.15
X14 a_647_21.t1 SET_B.t2 VPWR.t12 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X15 VPWR.t10 a_941_21.t2 a_891_329.t1 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.2247 pd=1.375 as=0.1134 ps=1.11 w=0.84 l=0.15
X16 a_557_413.t1 a_193_47.t4 a_473_413.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_193_47.t1 a_27_47.t4 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 Q.t0 a_2136_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X19 a_473_413.t0 a_27_47.t5 a_381_47.t3 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X20 a_891_329.t0 a_473_413.t5 a_647_21.t3 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X21 Q_N.t0 a_1415_315.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1539 ps=1.335 w=1 l=0.15
X22 Q.t1 a_2136_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 VPWR.t4 a_647_21.t4 a_557_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X24 a_1112_329.t0 a_647_21.t5 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1743 pd=1.41 as=0.2247 ps=1.375 w=0.84 l=0.15
X25 VGND.t4 a_647_21.t6 a_581_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X26 VGND.t1 a_1415_315.t5 a_2136_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_193_47.t0 a_27_47.t6 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 VPWR.t9 a_941_21.t3 a_1672_329.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X29 VPWR.t2 a_1415_315.t6 a_1340_413.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.07875 ps=0.795 w=0.42 l=0.15
X30 Q_N.t1 a_1415_315.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X31 a_381_47.t2 D.t1 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_1672_329.t0 a_1256_413.t2 a_1415_315.t0 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.1323 ps=1.22 w=0.84 l=0.15
X33 VGND.t8 CLK_N.t1 a_27_47.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 SET_B.n0 SET_B.t2 389.618
R1 SET_B.n2 SET_B.t1 383.033
R2 SET_B.n3 SET_B.n2 176.9
R3 SET_B.n3 SET_B.n0 157.042
R4 SET_B.n2 SET_B.n1 148.35
R5 SET_B.n0 SET_B.t0 142.569
R6 SET_B SET_B.n3 5.0092
R7 SET_B.n3 SET_B 3.29747
R8 VGND.n20 VGND.t0 256.322
R9 VGND.n42 VGND.t6 237.274
R10 VGND.n13 VGND.t2 226.882
R11 VGND.n12 VGND.n11 207.585
R12 VGND.n4 VGND.n3 205.707
R13 VGND.n45 VGND.n44 199.739
R14 VGND.n3 VGND.t4 81.4291
R15 VGND.n11 VGND.t1 54.2862
R16 VGND.n3 VGND.t5 38.5719
R17 VGND.n44 VGND.t7 38.5719
R18 VGND.n44 VGND.t8 38.5719
R19 VGND.n14 VGND.n10 34.6358
R20 VGND.n18 VGND.n10 34.6358
R21 VGND.n19 VGND.n18 34.6358
R22 VGND.n21 VGND.n19 34.6358
R23 VGND.n25 VGND.n8 34.6358
R24 VGND.n26 VGND.n25 34.6358
R25 VGND.n27 VGND.n26 34.6358
R26 VGND.n31 VGND.n6 34.6358
R27 VGND.n32 VGND.n31 34.6358
R28 VGND.n33 VGND.n32 34.6358
R29 VGND.n37 VGND.n36 34.6358
R30 VGND.n38 VGND.n37 34.6358
R31 VGND.n38 VGND.n1 34.6358
R32 VGND.n11 VGND.t3 25.9346
R33 VGND.n45 VGND.n43 22.9652
R34 VGND.n14 VGND.n13 22.2123
R35 VGND.n42 VGND.n1 21.4593
R36 VGND.n43 VGND.n42 21.0829
R37 VGND.n33 VGND.n4 18.0711
R38 VGND.n36 VGND.n4 16.5652
R39 VGND.n15 VGND.n14 9.3005
R40 VGND.n16 VGND.n10 9.3005
R41 VGND.n18 VGND.n17 9.3005
R42 VGND.n19 VGND.n9 9.3005
R43 VGND.n22 VGND.n21 9.3005
R44 VGND.n23 VGND.n8 9.3005
R45 VGND.n25 VGND.n24 9.3005
R46 VGND.n26 VGND.n7 9.3005
R47 VGND.n28 VGND.n27 9.3005
R48 VGND.n29 VGND.n6 9.3005
R49 VGND.n31 VGND.n30 9.3005
R50 VGND.n32 VGND.n5 9.3005
R51 VGND.n34 VGND.n33 9.3005
R52 VGND.n36 VGND.n35 9.3005
R53 VGND.n37 VGND.n2 9.3005
R54 VGND.n39 VGND.n38 9.3005
R55 VGND.n40 VGND.n1 9.3005
R56 VGND.n42 VGND.n41 9.3005
R57 VGND.n43 VGND.n0 9.3005
R58 VGND.n20 VGND.n8 9.03579
R59 VGND.n27 VGND.n6 8.28285
R60 VGND.n46 VGND.n45 7.12063
R61 VGND.n13 VGND.n12 7.10028
R62 VGND.n21 VGND.n20 1.12991
R63 VGND.n15 VGND.n12 0.218617
R64 VGND.n46 VGND.n0 0.148519
R65 VGND.n16 VGND.n15 0.120292
R66 VGND.n17 VGND.n16 0.120292
R67 VGND.n17 VGND.n9 0.120292
R68 VGND.n22 VGND.n9 0.120292
R69 VGND.n23 VGND.n22 0.120292
R70 VGND.n24 VGND.n23 0.120292
R71 VGND.n24 VGND.n7 0.120292
R72 VGND.n28 VGND.n7 0.120292
R73 VGND.n29 VGND.n28 0.120292
R74 VGND.n30 VGND.n29 0.120292
R75 VGND.n30 VGND.n5 0.120292
R76 VGND.n34 VGND.n5 0.120292
R77 VGND.n35 VGND.n34 0.120292
R78 VGND.n35 VGND.n2 0.120292
R79 VGND.n39 VGND.n2 0.120292
R80 VGND.n40 VGND.n39 0.120292
R81 VGND.n41 VGND.n40 0.120292
R82 VGND.n41 VGND.n0 0.120292
R83 VGND VGND.n46 0.114842
R84 a_791_47.t1 a_791_47.n0 468.514
R85 a_791_47.n0 a_791_47.t2 42.9469
R86 a_791_47.n0 a_791_47.t0 38.5719
R87 VNB.t0 VNB.t2 8144.98
R88 VNB.t8 VNB.t0 6934.63
R89 VNB.t2 VNB.t1 2677.02
R90 VNB.t10 VNB.t7 2677.02
R91 VNB.t4 VNB.t6 1623.3
R92 VNB.t5 VNB.t9 1495.15
R93 VNB.t6 VNB.t11 1366.99
R94 VNB.t9 VNB.t4 1366.99
R95 VNB.t1 VNB.t3 1352.75
R96 VNB.t7 VNB.t5 1352.75
R97 VNB.t11 VNB.t8 1196.12
R98 VNB.t12 VNB.t10 1196.12
R99 VNB VNB.t12 683.495
R100 a_27_47.n2 a_27_47.t5 533.949
R101 a_27_47.t0 a_27_47.n6 425.406
R102 a_27_47.n1 a_27_47.t2 348.024
R103 a_27_47.n1 a_27_47.n0 285.697
R104 a_27_47.n4 a_27_47.t1 266.572
R105 a_27_47.n5 a_27_47.t6 262.945
R106 a_27_47.n5 a_27_47.t4 227.597
R107 a_27_47.n3 a_27_47.n2 164.76
R108 a_27_47.n6 a_27_47.n5 152
R109 a_27_47.n2 a_27_47.t3 141.923
R110 a_27_47.n6 a_27_47.n4 21.4266
R111 a_27_47.n3 a_27_47.n1 16.586
R112 a_27_47.n4 a_27_47.n3 11.2483
R113 a_1256_413.n2 a_1256_413.n1 928.213
R114 a_1256_413.n1 a_1256_413.t2 236.934
R115 a_1256_413.n1 a_1256_413.n0 191.946
R116 a_1256_413.n2 a_1256_413.t1 63.3219
R117 a_1256_413.t0 a_1256_413.n2 63.3219
R118 RESET_B.n1 RESET_B.n0 202.559
R119 RESET_B.n1 RESET_B.t0 173.638
R120 RESET_B RESET_B.n1 154.111
R121 a_941_21.t0 a_941_21.n3 737.593
R122 a_941_21.n3 a_941_21.n2 211.821
R123 a_941_21.n1 a_941_21.n0 211.737
R124 a_941_21.n2 a_941_21.t1 210.474
R125 a_941_21.n1 a_941_21.t3 205.31
R126 a_941_21.n2 a_941_21.t2 204.048
R127 a_941_21.n3 a_941_21.n1 161.433
R128 VPWR.n20 VPWR.t9 793.365
R129 VPWR.n14 VPWR.n13 732.75
R130 VPWR.n47 VPWR.t7 666.351
R131 VPWR.n49 VPWR.n1 604.394
R132 VPWR.n41 VPWR.n5 599.485
R133 VPWR.n27 VPWR.n26 585
R134 VPWR.n16 VPWR.n15 321.743
R135 VPWR.n35 VPWR.n8 310.502
R136 VPWR.n26 VPWR.t2 121.953
R137 VPWR.n26 VPWR.t11 91.4648
R138 VPWR.n5 VPWR.t12 91.4648
R139 VPWR.n5 VPWR.t4 86.7743
R140 VPWR.n8 VPWR.t5 86.7743
R141 VPWR.n13 VPWR.t6 63.1021
R142 VPWR.n15 VPWR.t0 58.4849
R143 VPWR.n1 VPWR.t8 41.5552
R144 VPWR.n1 VPWR.t13 41.5552
R145 VPWR.n8 VPWR.t10 38.6969
R146 VPWR.n42 VPWR.n3 34.6358
R147 VPWR.n46 VPWR.n3 34.6358
R148 VPWR.n36 VPWR.n6 34.6358
R149 VPWR.n40 VPWR.n6 34.6358
R150 VPWR.n29 VPWR.n28 34.6358
R151 VPWR.n29 VPWR.n9 34.6358
R152 VPWR.n33 VPWR.n9 34.6358
R153 VPWR.n34 VPWR.n33 34.6358
R154 VPWR.n21 VPWR.n11 34.6358
R155 VPWR.n15 VPWR.t3 31.831
R156 VPWR.n42 VPWR.n41 31.2476
R157 VPWR.n25 VPWR.n11 28.9134
R158 VPWR.n13 VPWR.t1 28.0332
R159 VPWR.n49 VPWR.n48 22.9652
R160 VPWR.n47 VPWR.n46 21.4593
R161 VPWR.n48 VPWR.n47 21.0829
R162 VPWR.n28 VPWR.n27 18.1464
R163 VPWR.n21 VPWR.n20 14.7924
R164 VPWR.n19 VPWR.n18 10.706
R165 VPWR.n18 VPWR.n14 10.1241
R166 VPWR.n41 VPWR.n40 9.41227
R167 VPWR.n18 VPWR.n17 9.3005
R168 VPWR.n19 VPWR.n12 9.3005
R169 VPWR.n22 VPWR.n21 9.3005
R170 VPWR.n23 VPWR.n11 9.3005
R171 VPWR.n25 VPWR.n24 9.3005
R172 VPWR.n28 VPWR.n10 9.3005
R173 VPWR.n30 VPWR.n29 9.3005
R174 VPWR.n31 VPWR.n9 9.3005
R175 VPWR.n33 VPWR.n32 9.3005
R176 VPWR.n34 VPWR.n7 9.3005
R177 VPWR.n37 VPWR.n36 9.3005
R178 VPWR.n38 VPWR.n6 9.3005
R179 VPWR.n40 VPWR.n39 9.3005
R180 VPWR.n41 VPWR.n4 9.3005
R181 VPWR.n43 VPWR.n42 9.3005
R182 VPWR.n44 VPWR.n3 9.3005
R183 VPWR.n46 VPWR.n45 9.3005
R184 VPWR.n47 VPWR.n2 9.3005
R185 VPWR.n48 VPWR.n0 9.3005
R186 VPWR.n16 VPWR.n14 7.84423
R187 VPWR.n50 VPWR.n49 7.12063
R188 VPWR.n35 VPWR.n34 6.4005
R189 VPWR.n36 VPWR.n35 3.38874
R190 VPWR.n20 VPWR.n19 2.67686
R191 VPWR.n27 VPWR.n25 2.44414
R192 VPWR.n17 VPWR.n16 0.210873
R193 VPWR.n50 VPWR.n0 0.148519
R194 VPWR.n17 VPWR.n12 0.120292
R195 VPWR.n22 VPWR.n12 0.120292
R196 VPWR.n23 VPWR.n22 0.120292
R197 VPWR.n24 VPWR.n23 0.120292
R198 VPWR.n24 VPWR.n10 0.120292
R199 VPWR.n30 VPWR.n10 0.120292
R200 VPWR.n31 VPWR.n30 0.120292
R201 VPWR.n32 VPWR.n31 0.120292
R202 VPWR.n32 VPWR.n7 0.120292
R203 VPWR.n37 VPWR.n7 0.120292
R204 VPWR.n38 VPWR.n37 0.120292
R205 VPWR.n39 VPWR.n38 0.120292
R206 VPWR.n39 VPWR.n4 0.120292
R207 VPWR.n43 VPWR.n4 0.120292
R208 VPWR.n44 VPWR.n43 0.120292
R209 VPWR.n45 VPWR.n44 0.120292
R210 VPWR.n45 VPWR.n2 0.120292
R211 VPWR.n2 VPWR.n0 0.120292
R212 VPWR VPWR.n50 0.114842
R213 VPB.t14 VPB.t6 559.346
R214 VPB.t1 VPB.t0 556.386
R215 VPB.t11 VPB.t8 556.386
R216 VPB.t5 VPB.t7 426.168
R217 VPB.t15 VPB.t5 405.452
R218 VPB.t2 VPB.t17 358.101
R219 VPB.t9 VPB.t4 355.14
R220 VPB.t16 VPB.t18 319.627
R221 VPB.t17 VPB.t10 313.707
R222 VPB.t4 VPB.t16 313.707
R223 VPB.t13 VPB.t2 310.748
R224 VPB.t6 VPB.t1 287.072
R225 VPB.t0 VPB.t3 281.154
R226 VPB.t8 VPB.t12 272.274
R227 VPB.t7 VPB.t13 248.599
R228 VPB.t18 VPB.t15 248.599
R229 VPB.t12 VPB.t9 248.599
R230 VPB.t19 VPB.t11 248.599
R231 VPB.t10 VPB.t14 213.084
R232 VPB VPB.t19 142.056
R233 a_1415_315.n4 a_1415_315.n3 594.413
R234 a_1415_315.n2 a_1415_315.t2 383.241
R235 a_1415_315.n3 a_1415_315.n1 348.959
R236 a_1415_315.n1 a_1415_315.t4 268.313
R237 a_1415_315.n0 a_1415_315.t3 231.945
R238 a_1415_315.n1 a_1415_315.t7 222.792
R239 a_1415_315.n3 a_1415_315.n2 204.841
R240 a_1415_315.n0 a_1415_315.t5 164.464
R241 a_1415_315.n1 a_1415_315.n0 151.742
R242 a_1415_315.n2 a_1415_315.t6 139.028
R243 a_1415_315.n4 a_1415_315.t1 91.4648
R244 a_1415_315.t0 a_1415_315.n4 57.4588
R245 a_647_21.n7 a_647_21.n0 598.178
R246 a_647_21.n8 a_647_21.n7 585
R247 a_647_21.n6 a_647_21.t6 387.961
R248 a_647_21.n3 a_647_21.t5 299.911
R249 a_647_21.n5 a_647_21.n3 215.817
R250 a_647_21.n5 a_647_21.n4 202.456
R251 a_647_21.n7 a_647_21.n6 190.656
R252 a_647_21.n3 a_647_21.n2 167.63
R253 a_647_21.n6 a_647_21.t4 143.746
R254 a_647_21.n1 a_647_21.t1 110.227
R255 a_647_21.n7 a_647_21.n5 81.1737
R256 a_647_21.t3 a_647_21.n0 63.3219
R257 a_647_21.t3 a_647_21.n8 63.3219
R258 a_647_21.n4 a_647_21.t0 25.313
R259 a_647_21.n4 a_647_21.t2 25.313
R260 a_647_21.n1 a_647_21.n0 9.38145
R261 a_647_21.n8 a_647_21.n1 9.38145
R262 a_1363_47.n0 a_1363_47.t0 11.0774
R263 a_1340_413.t0 a_1340_413.t1 175.893
R264 CLK_N.n0 CLK_N.t0 272.062
R265 CLK_N.n0 CLK_N.t1 236.716
R266 CLK_N.n1 CLK_N.n0 152
R267 CLK_N CLK_N.n1 7.6805
R268 CLK_N.n1 CLK_N 4.75479
R269 D.n0 D.t0 331.51
R270 D.n0 D.t1 209.403
R271 D.n1 D.n0 152
R272 D.n1 D 8.58587
R273 D D.n1 2.02977
R274 a_381_47.n1 a_381_47.n0 959.148
R275 a_381_47.n1 a_381_47.t3 82.0838
R276 a_381_47.n0 a_381_47.t0 63.3338
R277 a_381_47.t1 a_381_47.n1 63.3219
R278 a_381_47.n0 a_381_47.t2 29.7268
R279 a_193_47.n1 a_193_47.n0 525.917
R280 a_193_47.t0 a_193_47.n4 367.062
R281 a_193_47.n2 a_193_47.t2 314.652
R282 a_193_47.n2 a_193_47.t4 307.325
R283 a_193_47.n4 a_193_47.t1 302.7
R284 a_193_47.n3 a_193_47.n1 171.565
R285 a_193_47.n1 a_193_47.t3 148.35
R286 a_193_47.n4 a_193_47.n3 10.4313
R287 a_193_47.n3 a_193_47.n2 9.3005
R288 a_473_413.n3 a_473_413.n2 707.533
R289 a_473_413.n2 a_473_413.n0 288.925
R290 a_473_413.n1 a_473_413.t4 216.9
R291 a_473_413.n2 a_473_413.n1 216.829
R292 a_473_413.n1 a_473_413.t5 210.474
R293 a_473_413.n0 a_473_413.t1 63.3338
R294 a_473_413.n3 a_473_413.t3 63.3219
R295 a_473_413.t0 a_473_413.n3 63.3219
R296 a_473_413.n0 a_473_413.t2 61.6672
R297 a_2136_47.t0 a_2136_47.n1 384.125
R298 a_2136_47.n1 a_2136_47.t1 243.28
R299 a_2136_47.n0 a_2136_47.t2 239.04
R300 a_2136_47.n1 a_2136_47.n0 175.079
R301 a_2136_47.n0 a_2136_47.t3 166.739
R302 a_1112_329.t0 a_1112_329.t1 236.869
R303 a_581_47.t0 a_581_47.t1 93.5174
R304 a_891_329.t0 a_891_329.t1 63.3219
R305 a_557_413.t0 a_557_413.t1 211.071
R306 Q.n1 Q.t0 353.606
R307 Q.n0 Q.t1 209.923
R308 Q Q.n0 67.6928
R309 Q.n1 Q 9.10538
R310 Q Q.n1 7.47898
R311 Q.n0 Q 6.64665
R312 Q_N.n1 Q_N.t0 353.795
R313 Q_N.n0 Q_N.t1 209.923
R314 Q_N Q_N.n0 79.4391
R315 Q_N.n1 Q_N 8.2361
R316 Q_N Q_N.n1 6.90173
R317 Q_N.n0 Q_N 5.61454
R318 a_1672_329.t0 a_1672_329.t1 49.2505
C0 a_1159_47# SET_B 0.004595f
C1 a_1555_47# VPB 8.96e-20
C2 SET_B VGND 0.311388f
C3 VPB Q 0.012255f
C4 a_1159_47# VPWR 6.2e-19
C5 VPWR VGND 0.080126f
C6 SET_B RESET_B 0.002286f
C7 a_1159_47# VGND 0.010753f
C8 SET_B Q_N 3.72e-19
C9 VPWR RESET_B 0.009905f
C10 a_1555_47# SET_B 0.013084f
C11 VPWR Q_N 0.061418f
C12 SET_B Q 1.24e-19
C13 VGND RESET_B 0.028219f
C14 a_1555_47# VPWR 1.3e-19
C15 VPB CLK_N 0.070636f
C16 VGND Q_N 0.086175f
C17 VPWR Q 0.099186f
C18 VPB D 0.081727f
C19 a_1555_47# VGND 0.156913f
C20 RESET_B Q_N 0.001702f
C21 VGND Q 0.06431f
C22 a_1555_47# RESET_B 3.78e-20
C23 VPB SET_B 0.146534f
C24 RESET_B Q 6.25e-20
C25 VPB VPWR 0.255196f
C26 VPB VGND 0.015088f
C27 CLK_N VPWR 0.019577f
C28 CLK_N VGND 0.019603f
C29 D VPWR 0.015279f
C30 VPB RESET_B 0.047578f
C31 VPB Q_N 0.01022f
C32 SET_B VPWR 0.025523f
C33 D VGND 0.013433f
C34 Q VNB 0.094482f
C35 Q_N VNB 0.013515f
C36 RESET_B VNB 0.133134f
C37 VGND VNB 1.30409f
C38 VPWR VNB 1.05366f
C39 SET_B VNB 0.264325f
C40 D VNB 0.125408f
C41 CLK_N VNB 0.196714f
C42 VPB VNB 2.37668f
C43 a_1555_47# VNB 0.008712f
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
R0 VGND.n6 VGND.t2 538.312
R1 VGND.n4 VGND.t0 219.992
R2 VGND.n16 VGND.n15 214.956
R3 VGND.n17 VGND.t1 214.456
R4 VGND.n6 VGND.n5 152
R5 VGND.n8 VGND.n7 152
R6 VGND.n15 VGND.n14 152
R7 VGND.t2 VGND.n2 68.6994
R8 VGND.n7 VGND.n6 62.9556
R9 VGND.n7 VGND.n2 31.4781
R10 VGND.n15 VGND.n2 31.4781
R11 VGND.n18 VGND.n17 9.56351
R12 VGND.n1 VGND.n0 9.3005
R13 VGND.n13 VGND.n12 9.3005
R14 VGND.n11 VGND.n3 9.3005
R15 VGND.n10 VGND.n9 9.3005
R16 VGND.n5 VGND.n4 5.29077
R17 VGND.n13 VGND.n1 4.03338
R18 VGND.n9 VGND.n5 3.59502
R19 VGND.n14 VGND.n3 3.59502
R20 VGND.n17 VGND.n16 2.63064
R21 VGND.n9 VGND.n8 2.01694
R22 VGND.n8 VGND.n3 2.01694
R23 VGND.n16 VGND.n1 1.14023
R24 VGND.n14 VGND.n13 0.438856
R25 VGND.n10 VGND.n4 0.283314
R26 VGND.n11 VGND.n10 0.120292
R27 VGND.n12 VGND.n11 0.120292
R28 VGND.n12 VGND.n0 0.120292
R29 VGND.n18 VGND.n0 0.120292
R30 VGND VGND.n18 0.0226354
R31 VPWR.n15 VPWR.t2 571.745
R32 VPWR.n29 VPWR.t1 388.656
R33 VPWR.n8 VPWR.t0 388.656
R34 VPWR.n13 VPWR.n6 214.956
R35 VPWR.n15 VPWR.n3 152
R36 VPWR.n17 VPWR.n16 152
R37 VPWR.n13 VPWR.n12 152
R38 VPWR.t2 VPWR.n14 107.793
R39 VPWR.n16 VPWR.n15 62.9556
R40 VPWR.n16 VPWR.n14 32.4617
R41 VPWR.n14 VPWR.n13 30.4944
R42 VPWR.n9 VPWR.n8 9.63602
R43 VPWR.n30 VPWR.n29 9.60526
R44 VPWR.n9 VPWR.n7 9.3005
R45 VPWR.n11 VPWR.n10 9.3005
R46 VPWR.n5 VPWR.n4 9.3005
R47 VPWR.n19 VPWR.n18 9.3005
R48 VPWR.n21 VPWR.n20 9.3005
R49 VPWR.n22 VPWR.n2 9.3005
R50 VPWR.n24 VPWR.n23 9.3005
R51 VPWR.n25 VPWR.n1 9.3005
R52 VPWR.n27 VPWR.n26 9.3005
R53 VPWR.n28 VPWR.n0 9.3005
R54 VPWR.n23 VPWR.n22 4.67352
R55 VPWR.n23 VPWR.n1 4.67352
R56 VPWR.n27 VPWR.n1 4.67352
R57 VPWR.n28 VPWR.n27 4.67352
R58 VPWR.n29 VPWR.n28 4.36875
R59 VPWR.n22 VPWR.n21 4.21352
R60 VPWR.n11 VPWR.n7 3.30837
R61 VPWR.n18 VPWR.n3 3.09263
R62 VPWR.n12 VPWR.n5 2.80499
R63 VPWR.n8 VPWR.n6 2.30162
R64 VPWR.n17 VPWR.n5 1.79825
R65 VPWR.n18 VPWR.n17 1.51061
R66 VPWR.n7 VPWR.n6 0.791511
R67 VPWR.n12 VPWR.n11 0.503871
R68 VPWR.n21 VPWR.n3 0.21623
R69 VPWR.n10 VPWR.n9 0.120292
R70 VPWR.n10 VPWR.n4 0.120292
R71 VPWR.n19 VPWR.n4 0.120292
R72 VPWR.n20 VPWR.n19 0.120292
R73 VPWR.n20 VPWR.n2 0.120292
R74 VPWR.n24 VPWR.n2 0.120292
R75 VPWR.n25 VPWR.n24 0.120292
R76 VPWR.n26 VPWR.n25 0.120292
R77 VPWR.n26 VPWR.n0 0.120292
R78 VPWR.n30 VPWR.n0 0.120292
R79 VPWR VPWR.n30 0.0226354
R80 VPB VPB.t0 1547.82
R81 VNB VNB.t0 7447.25
C0 VPB VGND 0.336433f
C1 VPB VPWR 0.142266f
C2 VGND VPWR 2.00892f
C3 VPWR VNB 1.70051f
C4 VGND VNB 1.467109f
C5 VPB VNB 1.13634f
C6 VPWR.n0 VNB 0.030298f
C7 VPWR.n1 VNB 0.079533f
C8 VPWR.n2 VNB 0.030298f
C9 VPWR.n3 VNB 0.056178f
C10 VPWR.n4 VNB 0.030298f
C11 VPWR.n5 VNB 0.078161f
C12 VPWR.n6 VNB 0.062459f
C13 VPWR.n7 VNB 0.069612f
C14 VPWR.t0 VNB 0.025643f
C15 VPWR.n8 VNB 0.083476f
C16 VPWR.n9 VNB 0.061021f
C17 VPWR.n10 VNB 0.030298f
C18 VPWR.n11 VNB 0.064727f
C19 VPWR.n12 VNB 0.056178f
C20 VPWR.n13 VNB 0.055949f
C21 VPWR.n14 VNB 0.153591f
C22 VPWR.t2 VNB 0.144582f
C23 VPWR.n15 VNB 0.072439f
C24 VPWR.n16 VNB 0.032611f
C25 VPWR.n17 VNB 0.056178f
C26 VPWR.n18 VNB 0.078161f
C27 VPWR.n19 VNB 0.030298f
C28 VPWR.n20 VNB 0.030298f
C29 VPWR.n21 VNB 0.055906f
C30 VPWR.n22 VNB 0.078117f
C31 VPWR.n23 VNB 0.079533f
C32 VPWR.n24 VNB 0.030298f
C33 VPWR.n25 VNB 0.030298f
C34 VPWR.n26 VNB 0.030298f
C35 VPWR.n27 VNB 0.079533f
C36 VPWR.n28 VNB 0.07694f
C37 VPWR.t1 VNB 0.025643f
C38 VPWR.n29 VNB 0.070029f
C39 VPWR.n30 VNB 0.018763f
C40 VGND.n0 VNB 0.031105f
C41 VGND.n1 VNB 0.060675f
C42 VGND.n2 VNB 0.235961f
C43 VGND.n3 VNB 0.065817f
C44 VGND.t0 VNB 0.021017f
C45 VGND.n4 VNB 0.458709f
C46 VGND.n5 VNB 0.133885f
C47 VGND.t2 VNB 0.284279f
C48 VGND.n6 VNB 0.073843f
C49 VGND.n7 VNB 0.033134f
C50 VGND.n8 VNB 0.047306f
C51 VGND.n9 VNB 0.065817f
C52 VGND.n10 VNB 0.099589f
C53 VGND.n11 VNB 0.031105f
C54 VGND.n12 VNB 0.031105f
C55 VGND.n13 VNB 0.052448f
C56 VGND.n14 VNB 0.047306f
C57 VGND.n15 VNB 0.056808f
C58 VGND.n16 VNB 0.054026f
C59 VGND.t1 VNB 0.018097f
C60 VGND.n17 VNB 0.06601f
C61 VGND.n18 VNB 0.019276f
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
R0 VGND.n4 VGND.t0 219.518
R1 VGND.n10 VGND.t1 214.456
R2 VGND.n9 VGND.n8 200.692
R3 VGND.n3 VGND.n2 190.399
R4 VGND.n8 VGND.n7 152
R5 VGND.n2 VGND.t2 34.2973
R6 VGND.n11 VGND.n10 9.56351
R7 VGND.n1 VGND.n0 9.3005
R8 VGND.n6 VGND.n5 9.3005
R9 VGND.n4 VGND.n3 5.14426
R10 VGND.n8 VGND.n2 4.85762
R11 VGND.n6 VGND.n3 3.50735
R12 VGND.n7 VGND.n1 3.2005
R13 VGND.n10 VGND.n9 2.63064
R14 VGND.n9 VGND.n1 1.14023
R15 VGND.n7 VGND.n6 0.833377
R16 VGND.n5 VGND.n4 0.53311
R17 VGND.n5 VGND.n0 0.120292
R18 VGND.n11 VGND.n0 0.120292
R19 VGND VGND.n11 0.0226354
R20 VPWR.n18 VPWR.t1 388.656
R21 VPWR.n5 VPWR.t0 388.656
R22 VPWR.n9 VPWR.n4 202.66
R23 VPWR.n11 VPWR.n10 190.165
R24 VPWR.n9 VPWR.n8 152
R25 VPWR.n10 VPWR.t2 50.5057
R26 VPWR.n6 VPWR.n5 9.63602
R27 VPWR.n19 VPWR.n18 9.60526
R28 VPWR.n7 VPWR.n6 9.3005
R29 VPWR.n3 VPWR.n2 9.3005
R30 VPWR.n13 VPWR.n12 9.3005
R31 VPWR.n14 VPWR.n1 9.3005
R32 VPWR.n16 VPWR.n15 9.3005
R33 VPWR.n17 VPWR.n0 9.3005
R34 VPWR.n10 VPWR.n9 7.11866
R35 VPWR.n16 VPWR.n1 4.67352
R36 VPWR.n17 VPWR.n16 4.67352
R37 VPWR.n18 VPWR.n17 4.36875
R38 VPWR.n12 VPWR.n1 4.18384
R39 VPWR.n11 VPWR.n3 3.16454
R40 VPWR.n8 VPWR.n7 2.76904
R41 VPWR.n5 VPWR.n4 2.1578
R42 VPWR.n7 VPWR.n4 0.935332
R43 VPWR.n8 VPWR.n3 0.539826
R44 VPWR.n12 VPWR.n11 0.14432
R45 VPWR.n6 VPWR.n2 0.120292
R46 VPWR.n13 VPWR.n2 0.120292
R47 VPWR.n14 VPWR.n13 0.120292
R48 VPWR.n15 VPWR.n14 0.120292
R49 VPWR.n15 VPWR.n0 0.120292
R50 VPWR.n19 VPWR.n0 0.120292
R51 VPWR VPWR.n19 0.0226354
R52 VPB VPB.t0 1003.27
R53 VNB VNB.t0 4827.18
C0 VPB VGND 0.219503f
C1 VPB VPWR 0.104823f
C2 VGND VPWR 1.27274f
C3 VPWR VNB 1.14152f
C4 VGND VNB 0.991595f
C5 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
R0 VGND.n1 VGND.t0 219.12
R1 VGND.n0 VGND.t1 214.456
R2 VGND.n0 VGND.t2 121.927
R3 VGND.n1 VGND.n0 4.29166
R4 VGND VGND.n1 0.929743
R5 VPWR.n3 VPWR.t0 390.471
R6 VPWR.n8 VPWR.t1 388.656
R7 VPWR.n2 VPWR.t2 129.344
R8 VPWR.n9 VPWR.n8 9.60526
R9 VPWR.n4 VPWR.n1 9.3005
R10 VPWR.n6 VPWR.n5 9.3005
R11 VPWR.n7 VPWR.n0 9.3005
R12 VPWR.n2 VPWR.n1 4.67352
R13 VPWR.n6 VPWR.n1 4.67352
R14 VPWR.n7 VPWR.n6 4.67352
R15 VPWR.n8 VPWR.n7 4.36875
R16 VPWR.n4 VPWR.n3 3.98687
R17 VPWR.n3 VPWR.n2 1.73763
R18 VPWR.n5 VPWR.n4 0.120292
R19 VPWR.n5 VPWR.n0 0.120292
R20 VPWR.n9 VPWR.n0 0.120292
R21 VPWR VPWR.n9 0.0226354
R22 VPB VPB.t0 730.997
R23 VNB VNB.t0 3517.15
C0 VPWR VGND 0.903312f
C1 VPB VGND 0.161065f
C2 VPWR VPB 0.085759f
C3 VPWR VNB 0.867393f
C4 VGND VNB 0.761362f
C5 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
R0 VGND.n1 VGND.t2 218.308
R1 VGND.n0 VGND.t0 218.243
R2 VGND.n2 VGND.t1 214.456
R3 VGND.n3 VGND.n2 9.70901
R4 VGND.n1 VGND.n0 6.78155
R5 VGND.n2 VGND.n1 2.7239
R6 VGND.n3 VGND.n0 1.75362
R7 VGND VGND.n3 0.0226354
R8 VPWR.n6 VPWR.t1 388.656
R9 VPWR.n2 VPWR.t0 388.656
R10 VPWR.n1 VPWR.t2 210.964
R11 VPWR.n3 VPWR.n2 9.72505
R12 VPWR.n7 VPWR.n6 9.60526
R13 VPWR.n4 VPWR.n3 9.3005
R14 VPWR.n5 VPWR.n0 9.3005
R15 VPWR.n5 VPWR.n4 4.67352
R16 VPWR.n6 VPWR.n5 4.36875
R17 VPWR.n4 VPWR.n1 2.33701
R18 VPWR.n2 VPWR.n1 2.03225
R19 VPWR.n3 VPWR.n0 0.120292
R20 VPWR.n7 VPWR.n0 0.120292
R21 VPWR VPWR.n7 0.0226354
R22 VPB VPB.t0 458.724
R23 VNB VNB.t0 2207.12
C0 VPWR VGND 0.545943f
C1 VPB VGND 0.116247f
C2 VPWR VPB 0.078686f
C3 VPWR VNB 0.61942f
C4 VGND VNB 0.553666f
C5 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_3.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
R0 VGND.n1 VGND.t2 259.082
R1 VGND.n0 VGND.t0 216.798
R2 VGND.n2 VGND.t1 214.456
R3 VGND.n3 VGND.n2 9.71789
R4 VGND.n1 VGND.n0 7.01592
R5 VGND.n3 VGND.n0 3.76277
R6 VGND.n2 VGND.n1 1.18311
R7 VGND VGND.n3 0.0226354
R8 VPWR.n1 VPWR.t0 381.443
R9 VPWR.n4 VPWR.t1 381.443
R10 VPWR.n2 VPWR.t2 242.282
R11 VPWR.n1 VPWR.n0 9.72505
R12 VPWR.n5 VPWR.n4 9.60526
R13 VPWR.n3 VPWR.n0 9.3005
R14 VPWR.n4 VPWR.n3 4.36875
R15 VPWR.n3 VPWR.n2 3.50526
R16 VPWR.n2 VPWR.n1 0.863992
R17 VPWR.n5 VPWR.n0 0.120292
R18 VPWR VPWR.n5 0.0226354
R19 VPB VPB.t0 315.767
R20 VNB VNB.t0 1487.5
C0 VPWR VPB 0.062496f
C1 VGND VPB 0.079664f
C2 VGND VPWR 0.352999f
C3 VPWR VNB 0.469966f
C4 VGND VNB 0.427318f
C5 VPB VNB 0.338976f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinvlp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinvlp_4 VNB VPB VPWR VGND A Y
X0 Y.t3 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 VGND.t0 A.t1 a_268_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X2 Y.t2 A.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X3 Y.t4 A.t3 a_110_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X4 VPWR.t1 A.t4 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X5 a_110_47.t1 A.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X6 a_268_47.t0 A.t6 Y.t5 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X7 VPWR.t0 A.t7 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
R0 A.n0 A.t7 198.819
R1 A A.n6 177.44
R2 A.n6 A.t5 155.847
R3 A.n4 A.t3 155.847
R4 A.n2 A.t6 155.847
R5 A.n0 A.t1 155.847
R6 A.n1 A.t2 127.249
R7 A.n3 A.t4 127.249
R8 A.n5 A.t0 127.249
R9 A.n2 A.n1 46.7399
R10 A.n5 A.n4 45.2793
R11 A.n4 A.n3 32.1338
R12 A.n3 A.n2 30.6732
R13 A.n6 A.n5 7.30353
R14 A.n1 A.n0 5.84292
R15 VPWR.n3 VPWR.t0 250.6
R16 VPWR.n7 VPWR.t3 244.496
R17 VPWR.n2 VPWR.n1 217.226
R18 VPWR.n6 VPWR.n5 34.6358
R19 VPWR.n1 VPWR.t2 27.5805
R20 VPWR.n1 VPWR.t1 27.5805
R21 VPWR.n7 VPWR.n6 19.9534
R22 VPWR.n3 VPWR.n2 16.4308
R23 VPWR.n5 VPWR.n4 9.3005
R24 VPWR.n6 VPWR.n0 9.3005
R25 VPWR.n8 VPWR.n7 9.3005
R26 VPWR.n4 VPWR.n3 0.687989
R27 VPWR.n5 VPWR.n2 0.376971
R28 VPWR.n4 VPWR.n0 0.120292
R29 VPWR.n8 VPWR.n0 0.120292
R30 VPWR VPWR.n8 0.0226354
R31 Y Y.n0 592.644
R32 Y.n6 Y.n0 585
R33 Y.n5 Y.n0 585
R34 Y.n4 Y.n1 254.282
R35 Y.n3 Y.n2 187.862
R36 Y.n2 Y.t5 30.546
R37 Y.n2 Y.t4 30.546
R38 Y.n0 Y.t1 27.5805
R39 Y.n0 Y.t3 27.5805
R40 Y.n1 Y.t0 27.5805
R41 Y.n1 Y.t2 27.5805
R42 Y Y.n3 10.6672
R43 Y Y.n4 10.3116
R44 Y.n6 Y 7.11161
R45 Y.n5 Y 6.57828
R46 Y Y.n5 5.51161
R47 Y Y.n6 4.97828
R48 Y.n4 Y 1.77828
R49 Y.n3 Y 1.42272
R50 VPB.t2 VPB.t0 313.707
R51 VPB.t1 VPB.t2 313.707
R52 VPB.t3 VPB.t1 313.707
R53 VPB VPB.t3 224.923
R54 a_268_47.t0 a_268_47.t1 45.8187
R55 VGND.n0 VGND.t0 241.893
R56 VGND.n0 VGND.t1 239.114
R57 VGND VGND.n0 0.0966988
R58 VNB.t2 VNB.t0 1224.6
R59 VNB.t0 VNB.t3 1025.24
R60 VNB.t1 VNB.t2 1025.24
R61 VNB VNB.t1 939.807
R62 a_110_47.t0 a_110_47.t1 45.8187
C0 VPB A 0.159652f
C1 VPB VPWR 0.077158f
C2 VPB Y 0.010649f
C3 A VPWR 0.16526f
C4 VPB VGND 0.006616f
C5 A Y 0.245402f
C6 VPWR Y 0.438512f
C7 A VGND 0.10133f
C8 VPWR VGND 0.068202f
C9 Y VGND 0.17274f
C10 VGND VNB 0.399829f
C11 Y VNB 0.040509f
C12 VPWR VNB 0.367813f
C13 A VNB 0.577528f
C14 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinvlp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinvlp_2 VGND VPWR A Y VPB VNB
X0 Y.t1 A.t0 a_150_67.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.67 as=0.066 ps=0.79 w=0.55 l=0.15
X1 VPWR.t1 A.t1 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.14 ps=1.28 w=1 l=0.25
X2 a_150_67.t0 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.79 as=0.15675 ps=1.67 w=0.55 l=0.15
X3 Y.t2 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
R0 A.n0 A.t1 189.266
R1 A A.n2 159.07
R2 A.n2 A.t3 140.941
R3 A.n1 A.t2 130.166
R4 A.n0 A.t0 122.108
R5 A.n1 A.n0 77.9238
R6 A.n2 A.n1 6.07294
R7 a_150_67.t0 a_150_67.t1 52.3641
R8 Y Y.n0 313.966
R9 Y.n1 Y.t1 215.546
R10 Y.n0 Y.t0 27.5805
R11 Y.n0 Y.t2 27.5805
R12 Y Y.n1 3.87904
R13 Y.n1 Y 3.12491
R14 VNB VNB.t0 1509.39
R15 VNB.t0 VNB.t1 1110.68
R16 VPWR.n0 VPWR.t0 343.81
R17 VPWR.n0 VPWR.t1 278.623
R18 VPWR VPWR.n0 0.225632
R19 VPB.t0 VPB.t1 313.707
R20 VPB VPB.t0 301.87
R21 VGND VGND.t0 244.752
C0 VPB A 0.094415f
C1 VPB VPWR 0.05899f
C2 A VPWR 0.093831f
C3 VPB Y 0.006017f
C4 A Y 0.137056f
C5 VPWR Y 0.185535f
C6 VPB VGND 0.005971f
C7 A VGND 0.052752f
C8 VPWR VGND 0.047424f
C9 Y VGND 0.108763f
C10 VGND VNB 0.293177f
C11 Y VNB 0.062881f
C12 VPWR VNB 0.276303f
C13 A VNB 0.337243f
C14 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND.t15 A.t0 Y.t39 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 Y.t23 A.t1 VPWR.t23 VPB.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR.t22 A.t2 Y.t22 VPB.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X3 Y.t21 A.t3 VPWR.t21 VPB.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND.t14 A.t4 Y.t38 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR.t20 A.t5 Y.t20 VPB.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y.t37 A.t6 VGND.t13 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND.t12 A.t7 Y.t36 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VPWR.t19 A.t8 Y.t19 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR.t18 A.t9 Y.t18 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 Y.t35 A.t10 VGND.t11 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 Y.t17 A.t11 VPWR.t17 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VPWR.t16 A.t12 Y.t16 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2175 ps=1.435 w=1 l=0.15
X13 VGND.t10 A.t13 Y.t34 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 Y.t15 A.t14 VPWR.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.275 ps=2.55 w=1 l=0.15
X15 VPWR.t14 A.t15 Y.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y.t13 A.t16 VPWR.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 Y.t12 A.t17 VPWR.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 Y.t33 A.t18 VGND.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VGND.t8 A.t19 Y.t32 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 Y.t31 A.t20 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 VGND.t6 A.t21 Y.t30 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 Y.t11 A.t22 VPWR.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR.t10 A.t23 Y.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 Y.t9 A.t24 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.1575 ps=1.315 w=1 l=0.15
X25 Y.t8 A.t25 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 VPWR.t7 A.t26 Y.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 Y.t29 A.t27 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 Y.t6 A.t28 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR.t5 A.t29 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR.t4 A.t30 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 Y.t28 A.t31 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 VGND.t3 A.t32 Y.t27 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR.t3 A.t33 Y.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 Y.t26 A.t34 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.09135 pd=0.855 as=0.06615 ps=0.735 w=0.42 l=0.15
X35 Y.t2 A.t35 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 Y.t25 A.t36 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X37 VPWR.t1 A.t37 Y.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 Y.t0 A.t38 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND.t0 A.t39 Y.t24 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.09135 ps=0.855 w=0.42 l=0.15
R0 A.n5 A.t30 218.106
R1 A.n34 A.t14 218.106
R2 A.n6 A.t28 204.048
R3 A.n9 A.t29 204.048
R4 A.n2 A.t17 204.048
R5 A.n16 A.t5 204.048
R6 A.n17 A.t38 204.048
R7 A.n18 A.t26 204.048
R8 A.n19 A.t16 204.048
R9 A.n20 A.t15 204.048
R10 A.n21 A.t3 204.048
R11 A.n22 A.t37 204.048
R12 A.n23 A.t25 204.048
R13 A.n24 A.t12 204.048
R14 A.n25 A.t24 204.048
R15 A.n26 A.t2 204.048
R16 A.n27 A.t35 204.048
R17 A.n28 A.t23 204.048
R18 A.n29 A.t11 204.048
R19 A.n30 A.t9 204.048
R20 A.n31 A.t1 204.048
R21 A.n40 A.t33 204.048
R22 A.n38 A.t22 204.048
R23 A.n33 A.t8 204.048
R24 A.n16 A.t0 175.127
R25 A.n17 A.t10 175.127
R26 A.n18 A.t4 175.127
R27 A.n19 A.t18 175.127
R28 A.n20 A.t7 175.127
R29 A.n21 A.t20 175.127
R30 A.n22 A.t32 175.127
R31 A.n23 A.t27 175.127
R32 A.n24 A.t39 175.127
R33 A.n25 A.t34 175.127
R34 A.n26 A.t13 175.127
R35 A.n27 A.t6 175.127
R36 A.n28 A.t19 175.127
R37 A.n29 A.t31 175.127
R38 A.n30 A.t21 175.127
R39 A.n31 A.t36 175.127
R40 A.n5 A.n4 163.453
R41 A.n35 A.n34 163.453
R42 A.n15 A.n14 163.117
R43 A.n7 A.n4 152
R44 A.n11 A.n10 152
R45 A.n8 A.n3 152
R46 A.n42 A.n41 152
R47 A.n39 A.n1 152
R48 A.n37 A.n36 152
R49 A.n35 A.n32 152
R50 A.n25 A.n24 78.3255
R51 A.n26 A.n25 62.2588
R52 A.n17 A.n16 57.5727
R53 A.n18 A.n17 57.5727
R54 A.n19 A.n18 57.5727
R55 A.n20 A.n19 57.5727
R56 A.n21 A.n20 57.5727
R57 A.n22 A.n21 57.5727
R58 A.n23 A.n22 57.5727
R59 A.n24 A.n23 57.5727
R60 A.n27 A.n26 57.5727
R61 A.n28 A.n27 57.5727
R62 A.n29 A.n28 57.5727
R63 A.n30 A.n29 57.5727
R64 A.n31 A.n30 57.5727
R65 A.n10 A.n7 45.5227
R66 A.n37 A.n32 45.5227
R67 A.n6 A.n5 43.5144
R68 A.n34 A.n33 43.5144
R69 A.n9 A.n8 35.4811
R70 A.n39 A.n38 35.4811
R71 A.n16 A.n15 34.1422
R72 A.n41 A.n31 34.1422
R73 A.n15 A.n2 23.4311
R74 A.n41 A.n40 23.4311
R75 A.n8 A.n2 22.0922
R76 A.n40 A.n39 22.0922
R77 A A.n0 12.1637
R78 A.n11 A.n3 11.4531
R79 A.n42 A.n1 11.4531
R80 A.n36 A.n1 11.4531
R81 A.n36 A.n35 11.4531
R82 A.n10 A.n9 10.0422
R83 A.n38 A.n37 10.0422
R84 A.n13 A.n12 9.5505
R85 A.n1 A.n0 9.5505
R86 A.n14 A.n13 9.3005
R87 A.n12 A.n4 7.74787
R88 A.n13 A.n0 6.47061
R89 A.n12 A.n11 3.70576
R90 A.n7 A.n6 2.00883
R91 A.n33 A.n32 2.00883
R92 A A.n42 1.17945
R93 A.n14 A.n3 0.337342
R94 Y.n24 Y.n22 341.416
R95 Y.n10 Y.n8 304.63
R96 Y.n24 Y.n23 304.307
R97 Y.n3 Y.n2 303.625
R98 Y.n5 Y.n4 300.87
R99 Y.n31 Y.n29 300.798
R100 Y.n13 Y.n12 300.476
R101 Y.n28 Y.n15 300.226
R102 Y.n27 Y.n17 300.226
R103 Y.n26 Y.n19 300.226
R104 Y.n25 Y.n21 300.226
R105 Y.n3 Y.n1 244.12
R106 Y.n7 Y.n6 240.183
R107 Y.n10 Y.n9 239.965
R108 Y.n11 Y.n0 236.733
R109 Y.n28 Y.n14 234.665
R110 Y.n27 Y.n16 234.665
R111 Y.n26 Y.n18 234.665
R112 Y.n25 Y.n20 234.665
R113 Y Y.n30 221.499
R114 Y.n30 Y.t24 75.7148
R115 Y.n29 Y.t9 53.1905
R116 Y.n30 Y.t26 48.5719
R117 Y.n26 Y.n25 44.0325
R118 Y.n27 Y.n26 44.0325
R119 Y.n28 Y.n27 44.0325
R120 Y.n5 Y.n3 43.9423
R121 Y.n25 Y.n24 43.5815
R122 Y.n14 Y.t27 40.0005
R123 Y.n14 Y.t29 40.0005
R124 Y.n16 Y.t36 40.0005
R125 Y.n16 Y.t31 40.0005
R126 Y.n18 Y.t38 40.0005
R127 Y.n18 Y.t33 40.0005
R128 Y.n20 Y.t39 40.0005
R129 Y.n20 Y.t35 40.0005
R130 Y.n6 Y.t30 40.0005
R131 Y.n6 Y.t25 40.0005
R132 Y.n9 Y.t32 40.0005
R133 Y.n9 Y.t28 40.0005
R134 Y.n0 Y.t34 40.0005
R135 Y.n0 Y.t37 40.0005
R136 Y.n31 Y.n28 39.4245
R137 Y.n31 Y.n13 39.2935
R138 Y.n11 Y.n10 37.1205
R139 Y.n10 Y.n7 36.8645
R140 Y.n29 Y.t16 32.5055
R141 Y.n15 Y.t1 27.5805
R142 Y.n15 Y.t8 27.5805
R143 Y.n17 Y.t14 27.5805
R144 Y.n17 Y.t21 27.5805
R145 Y.n19 Y.t7 27.5805
R146 Y.n19 Y.t13 27.5805
R147 Y.n21 Y.t20 27.5805
R148 Y.n21 Y.t0 27.5805
R149 Y.n22 Y.t4 27.5805
R150 Y.n22 Y.t6 27.5805
R151 Y.n23 Y.t5 27.5805
R152 Y.n23 Y.t12 27.5805
R153 Y.n1 Y.t19 27.5805
R154 Y.n1 Y.t15 27.5805
R155 Y.n2 Y.t3 27.5805
R156 Y.n2 Y.t11 27.5805
R157 Y.n4 Y.t18 27.5805
R158 Y.n4 Y.t23 27.5805
R159 Y.n8 Y.t10 27.5805
R160 Y.n8 Y.t17 27.5805
R161 Y.n12 Y.t22 27.5805
R162 Y.n12 Y.t2 27.5805
R163 Y Y.n31 3.8405
R164 Y.n31 Y 3.24317
R165 Y.n7 Y.n5 0.395986
R166 Y.n13 Y.n11 0.13249
R167 VGND.n7 VGND.t15 251.076
R168 VGND.n40 VGND.t1 246.096
R169 VGND.n19 VGND.n18 210.316
R170 VGND.n9 VGND.n8 206.494
R171 VGND.n12 VGND.n11 206.494
R172 VGND.n22 VGND.n21 206.494
R173 VGND.n28 VGND.n27 206.494
R174 VGND.n31 VGND.n30 206.494
R175 VGND.n38 VGND.n37 206.494
R176 VGND.n27 VGND.t10 47.1434
R177 VGND.n27 VGND.t2 42.8576
R178 VGND.n8 VGND.t11 40.0005
R179 VGND.n8 VGND.t14 40.0005
R180 VGND.n11 VGND.t9 40.0005
R181 VGND.n11 VGND.t12 40.0005
R182 VGND.n18 VGND.t7 40.0005
R183 VGND.n18 VGND.t3 40.0005
R184 VGND.n21 VGND.t5 40.0005
R185 VGND.n21 VGND.t0 40.0005
R186 VGND.n30 VGND.t13 40.0005
R187 VGND.n30 VGND.t8 40.0005
R188 VGND.n37 VGND.t4 40.0005
R189 VGND.n37 VGND.t6 40.0005
R190 VGND.n13 VGND.n10 34.6358
R191 VGND.n17 VGND.n5 34.6358
R192 VGND.n26 VGND.n3 34.6358
R193 VGND.n32 VGND.n29 34.6358
R194 VGND.n36 VGND.n1 34.6358
R195 VGND.n22 VGND.n20 34.2593
R196 VGND.n40 VGND.n39 30.4946
R197 VGND.n9 VGND.n7 19.3233
R198 VGND.n22 VGND.n3 15.0593
R199 VGND.n39 VGND.n38 14.3064
R200 VGND.n20 VGND.n19 10.5417
R201 VGND.n31 VGND.n1 9.78874
R202 VGND.n10 VGND.n6 9.3005
R203 VGND.n14 VGND.n13 9.3005
R204 VGND.n15 VGND.n5 9.3005
R205 VGND.n17 VGND.n16 9.3005
R206 VGND.n20 VGND.n4 9.3005
R207 VGND.n23 VGND.n22 9.3005
R208 VGND.n24 VGND.n3 9.3005
R209 VGND.n26 VGND.n25 9.3005
R210 VGND.n29 VGND.n2 9.3005
R211 VGND.n33 VGND.n32 9.3005
R212 VGND.n34 VGND.n1 9.3005
R213 VGND.n36 VGND.n35 9.3005
R214 VGND.n39 VGND.n0 9.3005
R215 VGND.n13 VGND.n12 8.65932
R216 VGND.n28 VGND.n26 7.52991
R217 VGND.n19 VGND.n17 7.15344
R218 VGND.n29 VGND.n28 7.15344
R219 VGND.n41 VGND.n40 6.82589
R220 VGND.n12 VGND.n5 6.02403
R221 VGND.n32 VGND.n31 4.89462
R222 VGND.n10 VGND.n9 1.50638
R223 VGND.n7 VGND.n6 1.46762
R224 VGND VGND.n41 0.465247
R225 VGND.n38 VGND.n36 0.376971
R226 VGND.n41 VGND.n0 0.159177
R227 VGND.n14 VGND.n6 0.120292
R228 VGND.n15 VGND.n14 0.120292
R229 VGND.n16 VGND.n15 0.120292
R230 VGND.n16 VGND.n4 0.120292
R231 VGND.n23 VGND.n4 0.120292
R232 VGND.n24 VGND.n23 0.120292
R233 VGND.n25 VGND.n24 0.120292
R234 VGND.n25 VGND.n2 0.120292
R235 VGND.n33 VGND.n2 0.120292
R236 VGND.n34 VGND.n33 0.120292
R237 VGND.n35 VGND.n34 0.120292
R238 VGND.n35 VGND.n0 0.120292
R239 VNB VNB.t1 5866.67
R240 VNB.t2 VNB.t0 1666.02
R241 VNB.t10 VNB.t2 1324.27
R242 VNB.t11 VNB.t15 1224.6
R243 VNB.t14 VNB.t11 1224.6
R244 VNB.t9 VNB.t14 1224.6
R245 VNB.t12 VNB.t9 1224.6
R246 VNB.t7 VNB.t12 1224.6
R247 VNB.t3 VNB.t7 1224.6
R248 VNB.t5 VNB.t3 1224.6
R249 VNB.t0 VNB.t5 1224.6
R250 VNB.t13 VNB.t10 1224.6
R251 VNB.t8 VNB.t13 1224.6
R252 VNB.t4 VNB.t8 1224.6
R253 VNB.t6 VNB.t4 1224.6
R254 VNB.t1 VNB.t6 1224.6
R255 VPWR.n20 VPWR.t4 348.663
R256 VPWR.n4 VPWR.n3 315.781
R257 VPWR.n8 VPWR.n7 315.781
R258 VPWR.n44 VPWR.n10 315.781
R259 VPWR.n37 VPWR.n14 315.781
R260 VPWR.n31 VPWR.n30 315.781
R261 VPWR.n28 VPWR.n17 315.781
R262 VPWR.n19 VPWR.n18 315.781
R263 VPWR.n22 VPWR.n21 315.781
R264 VPWR.n39 VPWR.n13 315.361
R265 VPWR.n57 VPWR.n2 315.334
R266 VPWR.n51 VPWR.n6 315.334
R267 VPWR.n59 VPWR.t15 248.843
R268 VPWR.n50 VPWR.n49 34.6358
R269 VPWR.n46 VPWR.n45 34.6358
R270 VPWR.n43 VPWR.n11 34.6358
R271 VPWR.n39 VPWR.n38 34.6358
R272 VPWR.n36 VPWR.n15 34.6358
R273 VPWR.n32 VPWR.n29 34.6358
R274 VPWR.n27 VPWR.n19 32.0005
R275 VPWR.n10 VPWR.t22 31.5205
R276 VPWR.n52 VPWR.n4 30.8711
R277 VPWR.n10 VPWR.t9 30.5355
R278 VPWR.n13 VPWR.t8 28.5655
R279 VPWR.n2 VPWR.t11 27.5805
R280 VPWR.n2 VPWR.t19 27.5805
R281 VPWR.n3 VPWR.t23 27.5805
R282 VPWR.n3 VPWR.t3 27.5805
R283 VPWR.n6 VPWR.t17 27.5805
R284 VPWR.n6 VPWR.t18 27.5805
R285 VPWR.n7 VPWR.t2 27.5805
R286 VPWR.n7 VPWR.t10 27.5805
R287 VPWR.n14 VPWR.t21 27.5805
R288 VPWR.n14 VPWR.t1 27.5805
R289 VPWR.n30 VPWR.t13 27.5805
R290 VPWR.n30 VPWR.t14 27.5805
R291 VPWR.n17 VPWR.t0 27.5805
R292 VPWR.n17 VPWR.t7 27.5805
R293 VPWR.n18 VPWR.t12 27.5805
R294 VPWR.n18 VPWR.t20 27.5805
R295 VPWR.n21 VPWR.t6 27.5805
R296 VPWR.n21 VPWR.t5 27.5805
R297 VPWR.n23 VPWR.n22 27.4829
R298 VPWR.n13 VPWR.t16 26.5955
R299 VPWR.n57 VPWR.n56 26.3534
R300 VPWR.n58 VPWR.n57 23.3417
R301 VPWR.n59 VPWR.n58 21.4593
R302 VPWR.n56 VPWR.n4 19.2005
R303 VPWR.n23 VPWR.n19 18.0711
R304 VPWR.n39 VPWR.n11 15.0593
R305 VPWR.n52 VPWR.n51 14.3064
R306 VPWR.n28 VPWR.n27 13.5534
R307 VPWR.n38 VPWR.n37 10.9181
R308 VPWR.n49 VPWR.n8 10.1652
R309 VPWR.n24 VPWR.n23 9.3005
R310 VPWR.n25 VPWR.n19 9.3005
R311 VPWR.n27 VPWR.n26 9.3005
R312 VPWR.n29 VPWR.n16 9.3005
R313 VPWR.n33 VPWR.n32 9.3005
R314 VPWR.n34 VPWR.n15 9.3005
R315 VPWR.n36 VPWR.n35 9.3005
R316 VPWR.n38 VPWR.n12 9.3005
R317 VPWR.n40 VPWR.n39 9.3005
R318 VPWR.n41 VPWR.n11 9.3005
R319 VPWR.n43 VPWR.n42 9.3005
R320 VPWR.n45 VPWR.n9 9.3005
R321 VPWR.n47 VPWR.n46 9.3005
R322 VPWR.n49 VPWR.n48 9.3005
R323 VPWR.n50 VPWR.n5 9.3005
R324 VPWR.n53 VPWR.n52 9.3005
R325 VPWR.n54 VPWR.n4 9.3005
R326 VPWR.n56 VPWR.n55 9.3005
R327 VPWR.n57 VPWR.n1 9.3005
R328 VPWR.n58 VPWR.n0 9.3005
R329 VPWR.n60 VPWR.n59 9.3005
R330 VPWR.n32 VPWR.n31 9.03579
R331 VPWR.n44 VPWR.n43 8.28285
R332 VPWR.n45 VPWR.n44 7.15344
R333 VPWR.n22 VPWR.n20 6.56401
R334 VPWR.n31 VPWR.n15 6.4005
R335 VPWR.n46 VPWR.n8 5.27109
R336 VPWR.n37 VPWR.n36 4.51815
R337 VPWR.n29 VPWR.n28 1.88285
R338 VPWR.n51 VPWR.n50 0.753441
R339 VPWR.n24 VPWR.n20 0.652261
R340 VPWR.n25 VPWR.n24 0.120292
R341 VPWR.n26 VPWR.n25 0.120292
R342 VPWR.n26 VPWR.n16 0.120292
R343 VPWR.n33 VPWR.n16 0.120292
R344 VPWR.n34 VPWR.n33 0.120292
R345 VPWR.n35 VPWR.n34 0.120292
R346 VPWR.n35 VPWR.n12 0.120292
R347 VPWR.n40 VPWR.n12 0.120292
R348 VPWR.n41 VPWR.n40 0.120292
R349 VPWR.n42 VPWR.n41 0.120292
R350 VPWR.n42 VPWR.n9 0.120292
R351 VPWR.n47 VPWR.n9 0.120292
R352 VPWR.n48 VPWR.n47 0.120292
R353 VPWR.n48 VPWR.n5 0.120292
R354 VPWR.n53 VPWR.n5 0.120292
R355 VPWR.n54 VPWR.n53 0.120292
R356 VPWR.n55 VPWR.n54 0.120292
R357 VPWR.n55 VPWR.n1 0.120292
R358 VPWR.n1 VPWR.n0 0.120292
R359 VPWR.n60 VPWR.n0 0.120292
R360 VPWR VPWR.n60 0.0226354
R361 VPB.t9 VPB.t16 346.262
R362 VPB.t22 VPB.t9 275.235
R363 VPB.t6 VPB.t4 254.518
R364 VPB.t5 VPB.t6 254.518
R365 VPB.t12 VPB.t5 254.518
R366 VPB.t20 VPB.t12 254.518
R367 VPB.t0 VPB.t20 254.518
R368 VPB.t7 VPB.t0 254.518
R369 VPB.t13 VPB.t7 254.518
R370 VPB.t14 VPB.t13 254.518
R371 VPB.t21 VPB.t14 254.518
R372 VPB.t1 VPB.t21 254.518
R373 VPB.t8 VPB.t1 254.518
R374 VPB.t16 VPB.t8 254.518
R375 VPB.t2 VPB.t22 254.518
R376 VPB.t10 VPB.t2 254.518
R377 VPB.t17 VPB.t10 254.518
R378 VPB.t18 VPB.t17 254.518
R379 VPB.t23 VPB.t18 254.518
R380 VPB.t3 VPB.t23 254.518
R381 VPB.t11 VPB.t3 254.518
R382 VPB.t19 VPB.t11 254.518
R383 VPB.t15 VPB.t19 254.518
R384 VPB VPB.t15 201.246
C0 VPB A 0.781151f
C1 VPB VPWR 0.211998f
C2 A VPWR 0.766039f
C3 VPB Y 0.049071f
C4 A Y 1.79028f
C5 VPB VGND 0.008785f
C6 VPWR Y 2.08506f
C7 A VGND 0.797755f
C8 VPWR VGND 0.057369f
C9 Y VGND 0.805589f
C10 VGND VNB 1.29662f
C11 Y VNB 0.178563f
C12 VPWR VNB 1.039886f
C13 A VNB 2.36217f
C14 VPB VNB 2.19949f
C15 VPWR.n0 VNB 0.034337f
C16 VPWR.t15 VNB 0.043952f
C17 VPWR.n1 VNB 0.034337f
C18 VPWR.t11 VNB 0.010886f
C19 VPWR.t19 VNB 0.010886f
C20 VPWR.n2 VNB 0.023793f
C21 VPWR.t23 VNB 0.010886f
C22 VPWR.t3 VNB 0.010886f
C23 VPWR.n3 VNB 0.02379f
C24 VPWR.n4 VNB 0.045237f
C25 VPWR.n5 VNB 0.034337f
C26 VPWR.t17 VNB 0.010886f
C27 VPWR.t18 VNB 0.010886f
C28 VPWR.n6 VNB 0.023793f
C29 VPWR.t2 VNB 0.010886f
C30 VPWR.t10 VNB 0.010886f
C31 VPWR.n7 VNB 0.02379f
C32 VPWR.n8 VNB 0.039157f
C33 VPWR.n9 VNB 0.034337f
C34 VPWR.t9 VNB 0.012052f
C35 VPWR.t22 VNB 0.012441f
C36 VPWR.n10 VNB 0.026512f
C37 VPWR.n11 VNB 0.008724f
C38 VPWR.n12 VNB 0.034337f
C39 VPWR.t8 VNB 0.011274f
C40 VPWR.t16 VNB 0.010497f
C41 VPWR.n13 VNB 0.023776f
C42 VPWR.t21 VNB 0.010886f
C43 VPWR.t1 VNB 0.010886f
C44 VPWR.n14 VNB 0.02379f
C45 VPWR.n15 VNB 0.007204f
C46 VPWR.n16 VNB 0.034337f
C47 VPWR.t0 VNB 0.010886f
C48 VPWR.t7 VNB 0.010886f
C49 VPWR.n17 VNB 0.02379f
C50 VPWR.t12 VNB 0.010886f
C51 VPWR.t20 VNB 0.010886f
C52 VPWR.n18 VNB 0.02379f
C53 VPWR.n19 VNB 0.045237f
C54 VPWR.t4 VNB 0.041518f
C55 VPWR.n20 VNB 0.068181f
C56 VPWR.t6 VNB 0.010886f
C57 VPWR.t5 VNB 0.010886f
C58 VPWR.n21 VNB 0.02379f
C59 VPWR.n22 VNB 0.046695f
C60 VPWR.n23 VNB 0.007997f
C61 VPWR.n24 VNB 0.115081f
C62 VPWR.n25 VNB 0.034337f
C63 VPWR.n26 VNB 0.034337f
C64 VPWR.n27 VNB 0.007997f
C65 VPWR.n28 VNB 0.039157f
C66 VPWR.n29 VNB 0.006411f
C67 VPWR.t13 VNB 0.010886f
C68 VPWR.t14 VNB 0.010886f
C69 VPWR.n30 VNB 0.02379f
C70 VPWR.n31 VNB 0.039157f
C71 VPWR.n32 VNB 0.007667f
C72 VPWR.n33 VNB 0.034337f
C73 VPWR.n34 VNB 0.034337f
C74 VPWR.n35 VNB 0.034337f
C75 VPWR.n36 VNB 0.006874f
C76 VPWR.n37 VNB 0.039157f
C77 VPWR.n38 VNB 0.007997f
C78 VPWR.n39 VNB 0.045718f
C79 VPWR.n40 VNB 0.034337f
C80 VPWR.n41 VNB 0.034337f
C81 VPWR.n42 VNB 0.034337f
C82 VPWR.n43 VNB 0.007535f
C83 VPWR.n44 VNB 0.039157f
C84 VPWR.n45 VNB 0.007336f
C85 VPWR.n46 VNB 0.007006f
C86 VPWR.n47 VNB 0.034337f
C87 VPWR.n48 VNB 0.034337f
C88 VPWR.n49 VNB 0.007865f
C89 VPWR.n50 VNB 0.006213f
C90 VPWR.n51 VNB 0.039842f
C91 VPWR.n52 VNB 0.007931f
C92 VPWR.n53 VNB 0.034337f
C93 VPWR.n54 VNB 0.034337f
C94 VPWR.n55 VNB 0.034337f
C95 VPWR.n56 VNB 0.007997f
C96 VPWR.n57 VNB 0.045922f
C97 VPWR.n58 VNB 0.007865f
C98 VPWR.n59 VNB 0.052866f
C99 VPWR.n60 VNB 0.020341f
C100 Y.t34 VNB 0.0053f
C101 Y.t37 VNB 0.0053f
C102 Y.n0 VNB 0.016747f
C103 Y.t19 VNB 0.01262f
C104 Y.t15 VNB 0.01262f
C105 Y.n1 VNB 0.036238f
C106 Y.t3 VNB 0.01262f
C107 Y.t11 VNB 0.01262f
C108 Y.n2 VNB 0.026854f
C109 Y.n3 VNB 0.116194f
C110 Y.t18 VNB 0.01262f
C111 Y.t23 VNB 0.01262f
C112 Y.n4 VNB 0.02637f
C113 Y.n5 VNB 0.014932f
C114 Y.t30 VNB 0.0053f
C115 Y.t25 VNB 0.0053f
C116 Y.n6 VNB 0.016659f
C117 Y.n7 VNB 0.087868f
C118 Y.t10 VNB 0.01262f
C119 Y.t17 VNB 0.01262f
C120 Y.n8 VNB 0.026986f
C121 Y.t32 VNB 0.0053f
C122 Y.t28 VNB 0.0053f
C123 Y.n9 VNB 0.018103f
C124 Y.n10 VNB 0.123069f
C125 Y.n11 VNB 0.092281f
C126 Y.t22 VNB 0.01262f
C127 Y.t2 VNB 0.01262f
C128 Y.n12 VNB 0.02634f
C129 Y.n13 VNB 0.017297f
C130 Y.t27 VNB 0.0053f
C131 Y.t29 VNB 0.0053f
C132 Y.n14 VNB 0.016801f
C133 Y.t1 VNB 0.01262f
C134 Y.t8 VNB 0.01262f
C135 Y.n15 VNB 0.026342f
C136 Y.t36 VNB 0.0053f
C137 Y.t31 VNB 0.0053f
C138 Y.n16 VNB 0.016801f
C139 Y.t14 VNB 0.01262f
C140 Y.t21 VNB 0.01262f
C141 Y.n17 VNB 0.026342f
C142 Y.t38 VNB 0.0053f
C143 Y.t33 VNB 0.0053f
C144 Y.n18 VNB 0.016801f
C145 Y.t7 VNB 0.01262f
C146 Y.t13 VNB 0.01262f
C147 Y.n19 VNB 0.026342f
C148 Y.t39 VNB 0.0053f
C149 Y.t35 VNB 0.0053f
C150 Y.n20 VNB 0.016801f
C151 Y.t20 VNB 0.01262f
C152 Y.t0 VNB 0.01262f
C153 Y.n21 VNB 0.026342f
C154 Y.t4 VNB 0.01262f
C155 Y.t6 VNB 0.01262f
C156 Y.n22 VNB 0.033037f
C157 Y.t5 VNB 0.01262f
C158 Y.t12 VNB 0.01262f
C159 Y.n23 VNB 0.026849f
C160 Y.n24 VNB 0.116515f
C161 Y.n25 VNB 0.113688f
C162 Y.n26 VNB 0.117997f
C163 Y.n27 VNB 0.117997f
C164 Y.n28 VNB 0.115968f
C165 Y.t16 VNB 0.014874f
C166 Y.t9 VNB 0.024339f
C167 Y.n29 VNB 0.040991f
C168 Y.t24 VNB 0.010033f
C169 Y.t26 VNB 0.006436f
C170 Y.n30 VNB 0.023374f
C171 Y.n31 VNB 0.099286f
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_8 VNB VPB VGND VPWR A Y
X0 Y.t13 A.t0 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 VPWR.t11 A.t1 Y.t19 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y.t12 A.t2 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 Y.t11 A.t3 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y.t18 A.t4 VPWR.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t9 A.t5 Y.t17 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t8 A.t6 Y.t16 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t10 A.t7 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 Y.t15 A.t8 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t3 A.t9 Y.t9 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 Y.t14 A.t10 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1375 ps=1.275 w=1 l=0.15
X11 VPWR.t5 A.t11 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t2 A.t12 Y.t8 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR.t4 A.t13 Y.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t3 A.t14 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t1 A.t15 Y.t7 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VPWR.t2 A.t16 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y.t1 A.t17 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y.t0 A.t18 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND.t0 A.t19 Y.t6 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
R0 A.n8 A.t11 225.911
R1 A.n41 A.t18 205.375
R2 A.n7 A.t8 192.8
R3 A.n11 A.t13 192.8
R4 A.n5 A.t14 192.8
R5 A.n18 A.t16 192.8
R6 A.n23 A.t17 192.8
R7 A.n3 A.t1 192.8
R8 A.n30 A.t4 192.8
R9 A.n33 A.t6 192.8
R10 A.n1 A.t10 192.8
R11 A.n40 A.t5 192.8
R12 A.n9 A.n8 169.067
R13 A.n10 A.n9 152
R14 A.n14 A.n13 152
R15 A.n16 A.n15 152
R16 A.n20 A.n19 152
R17 A.n22 A.n21 152
R18 A.n26 A.n25 152
R19 A.n28 A.n27 152
R20 A.n31 A.n2 152
R21 A.n36 A.n35 152
R22 A.n38 A.n37 152
R23 A.n39 A.n0 152
R24 A.n42 A.n41 152
R25 A.n34 A.t0 117.287
R26 A.n32 A.t15 117.287
R27 A.n29 A.t7 117.287
R28 A.n24 A.t12 117.287
R29 A.n4 A.t3 117.287
R30 A.n17 A.t9 117.287
R31 A.n12 A.t2 117.287
R32 A.n6 A.t19 117.287
R33 A.n39 A.n38 28.5014
R34 A.n24 A.n23 24.3101
R35 A.n41 A.n40 22.6335
R36 A.n28 A.n3 21.3762
R37 A.n7 A.n6 20.957
R38 A.n13 A.n11 19.6996
R39 A.n35 A.n34 18.8614
R40 A.n19 A.n4 17.1848
R41 A.n21 A.n20 17.0672
R42 A.n36 A.n2 17.0672
R43 A.n42 A.n0 17.0672
R44 A.n27 A 16.5652
R45 A.n15 A 15.5613
R46 A.n31 A.n30 14.6701
R47 A.n14 A 13.5534
R48 A.n12 A.n5 13.4127
R49 A.n16 A.n5 12.9935
R50 A.n18 A.n17 12.5744
R51 A.n26 A 12.5495
R52 A.n37 A 11.5456
R53 A.n37 A 11.5456
R54 A.n22 A.n4 11.317
R55 A.n32 A.n31 11.317
R56 A A.n26 10.5417
R57 A.n30 A.n29 10.0596
R58 A.n17 A.n16 9.6405
R59 A A.n14 9.53776
R60 A.n33 A.n32 9.22137
R61 A.n11 A.n10 8.80224
R62 A.n34 A.n1 8.38311
R63 A.n35 A.n33 7.96398
R64 A.n15 A 7.52991
R65 A.n25 A.n3 7.12572
R66 A.n27 A 6.52599
R67 A.n19 A.n18 6.28746
R68 A.n40 A.n39 5.86833
R69 A A.n36 5.52207
R70 A A.n0 5.52207
R71 A.n10 A.n6 5.4492
R72 A.n21 A 4.51815
R73 A.n25 A.n24 3.77267
R74 A.n29 A.n28 3.77267
R75 A.n9 A 3.51423
R76 A.n8 A.n7 2.09615
R77 A.n13 A.n12 2.09615
R78 A.n20 A 1.50638
R79 A.n38 A.n1 1.25789
R80 A A.n2 0.502461
R81 A A.n42 0.502461
R82 A.n23 A.n22 0.41963
R83 VGND.n4 VGND.t0 245.494
R84 VGND.n15 VGND.t7 240.127
R85 VGND.n6 VGND.n5 200.127
R86 VGND.n9 VGND.n8 200.127
R87 VGND.n13 VGND.n2 200.127
R88 VGND.n5 VGND.t6 40.0005
R89 VGND.n5 VGND.t3 40.0005
R90 VGND.n8 VGND.t5 40.0005
R91 VGND.n8 VGND.t2 40.0005
R92 VGND.n2 VGND.t4 40.0005
R93 VGND.n2 VGND.t1 40.0005
R94 VGND.n9 VGND.n7 27.4829
R95 VGND.n13 VGND.n1 22.9652
R96 VGND.n14 VGND.n13 21.4593
R97 VGND.n15 VGND.n14 18.4476
R98 VGND.n9 VGND.n1 16.9417
R99 VGND.n7 VGND.n6 12.424
R100 VGND.n7 VGND.n3 9.3005
R101 VGND.n10 VGND.n9 9.3005
R102 VGND.n11 VGND.n1 9.3005
R103 VGND.n13 VGND.n12 9.3005
R104 VGND.n14 VGND.n0 9.3005
R105 VGND.n16 VGND.n15 7.26269
R106 VGND.n6 VGND.n4 6.80308
R107 VGND.n4 VGND.n3 0.797793
R108 VGND VGND.n16 0.231207
R109 VGND.n16 VGND.n0 0.15127
R110 VGND.n10 VGND.n3 0.120292
R111 VGND.n11 VGND.n10 0.120292
R112 VGND.n12 VGND.n11 0.120292
R113 VGND.n12 VGND.n0 0.120292
R114 Y.n9 Y.n8 317.498
R115 Y.n11 Y.n10 313.452
R116 Y.n19 Y.n18 313.452
R117 Y.n15 Y.n14 313.026
R118 Y.n13 Y.n12 312.618
R119 Y.n17 Y.n16 312.226
R120 Y.n1 Y.n0 207.569
R121 Y.n3 Y.n2 207.569
R122 Y.n5 Y.n4 207.569
R123 Y.n7 Y.n6 207.569
R124 Y.n9 Y.n7 172.8
R125 Y.n20 Y.n1 65.1299
R126 Y.n3 Y.n1 50.4476
R127 Y.n5 Y.n3 50.4476
R128 Y.n7 Y.n5 50.4476
R129 Y.n11 Y.n9 45.177
R130 Y.n13 Y.n11 45.177
R131 Y.n17 Y.n15 44.8005
R132 Y.n19 Y.n17 44.424
R133 Y.n15 Y.n13 44.0476
R134 Y.n0 Y.t6 40.0005
R135 Y.n0 Y.t12 40.0005
R136 Y.n2 Y.t9 40.0005
R137 Y.n2 Y.t11 40.0005
R138 Y.n4 Y.t8 40.0005
R139 Y.n4 Y.t10 40.0005
R140 Y.n6 Y.t7 40.0005
R141 Y.n6 Y.t13 40.0005
R142 Y.n8 Y.t17 26.5955
R143 Y.n8 Y.t0 26.5955
R144 Y.n10 Y.t16 26.5955
R145 Y.n10 Y.t14 26.5955
R146 Y.n12 Y.t19 26.5955
R147 Y.n12 Y.t18 26.5955
R148 Y.n14 Y.t2 26.5955
R149 Y.n14 Y.t1 26.5955
R150 Y.n16 Y.t4 26.5955
R151 Y.n16 Y.t3 26.5955
R152 Y.n18 Y.t5 26.5955
R153 Y.n18 Y.t15 26.5955
R154 Y Y.n19 17.1648
R155 Y.n20 Y 15.4079
R156 Y Y.n20 0.711611
R157 VNB VNB.t7 3602.59
R158 VNB.t6 VNB.t0 1224.6
R159 VNB.t3 VNB.t6 1224.6
R160 VNB.t5 VNB.t3 1224.6
R161 VNB.t2 VNB.t5 1224.6
R162 VNB.t4 VNB.t2 1224.6
R163 VNB.t1 VNB.t4 1224.6
R164 VNB.t7 VNB.t1 1224.6
R165 VPWR.n9 VPWR.t5 349.815
R166 VPWR.n25 VPWR.t0 343.651
R167 VPWR.n17 VPWR.n6 318.558
R168 VPWR.n11 VPWR.n10 318.038
R169 VPWR.n8 VPWR.n7 317.538
R170 VPWR.n23 VPWR.n2 317.058
R171 VPWR.n4 VPWR.n3 317.058
R172 VPWR.n16 VPWR.n15 34.6358
R173 VPWR.n18 VPWR.n4 34.2593
R174 VPWR.n12 VPWR.n11 32.7534
R175 VPWR.n23 VPWR.n22 28.2358
R176 VPWR.n2 VPWR.t9 27.5805
R177 VPWR.n2 VPWR.t6 26.5955
R178 VPWR.n3 VPWR.t10 26.5955
R179 VPWR.n3 VPWR.t8 26.5955
R180 VPWR.n6 VPWR.t1 26.5955
R181 VPWR.n6 VPWR.t11 26.5955
R182 VPWR.n7 VPWR.t3 26.5955
R183 VPWR.n7 VPWR.t2 26.5955
R184 VPWR.n10 VPWR.t7 26.5955
R185 VPWR.n10 VPWR.t4 26.5955
R186 VPWR.n25 VPWR.n24 22.2123
R187 VPWR.n24 VPWR.n23 21.4593
R188 VPWR.n22 VPWR.n4 15.4358
R189 VPWR.n12 VPWR.n8 12.0476
R190 VPWR.n18 VPWR.n17 10.1652
R191 VPWR.n13 VPWR.n12 9.3005
R192 VPWR.n15 VPWR.n14 9.3005
R193 VPWR.n16 VPWR.n5 9.3005
R194 VPWR.n19 VPWR.n18 9.3005
R195 VPWR.n20 VPWR.n4 9.3005
R196 VPWR.n22 VPWR.n21 9.3005
R197 VPWR.n23 VPWR.n1 9.3005
R198 VPWR.n24 VPWR.n0 9.3005
R199 VPWR.n26 VPWR.n25 9.3005
R200 VPWR.n11 VPWR.n9 6.31727
R201 VPWR.n17 VPWR.n16 6.02403
R202 VPWR.n15 VPWR.n8 3.38874
R203 VPWR.n13 VPWR.n9 0.58942
R204 VPWR.n14 VPWR.n13 0.120292
R205 VPWR.n14 VPWR.n5 0.120292
R206 VPWR.n19 VPWR.n5 0.120292
R207 VPWR.n20 VPWR.n19 0.120292
R208 VPWR.n21 VPWR.n20 0.120292
R209 VPWR.n21 VPWR.n1 0.120292
R210 VPWR.n1 VPWR.n0 0.120292
R211 VPWR.n26 VPWR.n0 0.120292
R212 VPWR VPWR.n26 0.0213333
R213 VPB.t9 VPB.t6 251.559
R214 VPB.t7 VPB.t5 248.599
R215 VPB.t4 VPB.t7 248.599
R216 VPB.t3 VPB.t4 248.599
R217 VPB.t2 VPB.t3 248.599
R218 VPB.t1 VPB.t2 248.599
R219 VPB.t11 VPB.t1 248.599
R220 VPB.t10 VPB.t11 248.599
R221 VPB.t8 VPB.t10 248.599
R222 VPB.t6 VPB.t8 248.599
R223 VPB.t0 VPB.t9 248.599
R224 VPB VPB.t0 189.409
C0 Y VGND 0.565628f
C1 VPB A 0.371833f
C2 VPB VPWR 0.137275f
C3 A VPWR 0.257137f
C4 VPB Y 0.028677f
C5 A Y 1.25589f
C6 VPB VGND 0.01291f
C7 VPWR Y 1.08033f
C8 A VGND 0.177761f
C9 VPWR VGND 0.123922f
C10 VGND VNB 0.715601f
C11 Y VNB 0.143222f
C12 VPWR VNB 0.598359f
C13 A VNB 1.15234f
C14 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfbbn_2 VGND VPWR VPB VNB Q Q_N RESET_B SET_B D CLK_N
X0 a_790_47.t0 SET_B.t0 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X1 a_790_47.t2 a_944_21.t2 a_650_21.t0 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2 Q_N.t1 a_1431_21.t4 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X3 a_894_329.t1 a_476_47.t4 a_650_21.t2 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.09 as=0.147 ps=1.23 w=0.84 l=0.15
X4 a_476_47.t2 a_27_47.t2 a_381_47.t1 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND.t10 a_650_21.t4 a_584_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.06705 ps=0.75 w=0.42 l=0.15
X6 VPWR.t3 a_2236_47.t2 Q.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t2 a_650_21.t5 a_560_413.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X8 a_1547_47.t0 a_944_21.t3 a_1431_21.t0 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.83 as=0.0864 ps=0.91 w=0.64 l=0.15
X9 VPWR.t13 CLK_N.t0 a_27_47.t0 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 Q.t0 a_2236_47.t3 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X11 a_381_47.t2 D.t0 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_476_47.t0 a_193_47.t2 a_381_47.t0 VNB.t0 sky130_fd_pr__special_nfet_01v8 ad=0.0702 pd=0.75 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_584_47.t0 a_27_47.t3 a_476_47.t3 VNB.t18 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0702 ps=0.75 w=0.36 l=0.15
X14 VPWR.t0 a_944_21.t4 a_894_329.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2331 pd=1.395 as=0.105 ps=1.09 w=0.84 l=0.15
X15 a_1162_47.t1 a_650_21.t6 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 VGND.t7 a_1431_21.t5 Q_N.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Q.t3 a_2236_47.t4 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X18 VGND.t4 a_1431_21.t6 a_2236_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X19 a_193_47.t1 a_27_47.t4 VGND.t12 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR.t12 RESET_B.t0 a_944_21.t0 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.176 ps=1.83 w=0.64 l=0.15
X21 Q_N.t2 a_1431_21.t7 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X22 VPWR.t9 a_1431_21.t8 a_1343_413# VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X23 VPWR.t1 a_944_21.t5 a_1665_329.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X24 VGND.t9 a_1431_21.t9 a_1366_47.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X25 VGND.t1 a_2236_47.t5 Q.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_1431_21.t3 SET_B.t1 VPWR.t11 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X27 VPWR.t7 a_1431_21.t10 Q_N.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1366_47.t1 a_193_47.t3 a_1257_47# VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X29 a_1665_329.t1 a_1257_47# a_1431_21.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.12285 ps=1.17 w=0.84 l=0.15
X30 a_193_47.t0 a_27_47.t5 VPWR.t14 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X31 a_1257_47# a_27_47.t6 a_1162_47.t0 VNB.t20 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X32 a_650_21.t3 a_476_47.t5 a_790_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X33 a_381_47.t3 D.t1 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X34 a_1431_21.t1 a_1257_47# a_1547_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.1199 ps=1.08 w=0.64 l=0.15
X35 a_650_21.t1 SET_B.t2 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X36 VPWR.t6 a_1431_21.t11 a_2236_47.t0 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X37 VGND.t8 RESET_B.t1 a_944_21.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1113 ps=1.37 w=0.42 l=0.15
X38 a_560_413.t0 a_193_47.t4 a_476_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 VGND.t11 CLK_N.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 SET_B.n0 SET_B.t2 389.618
R1 SET_B.n2 SET_B.t1 387.207
R2 SET_B.n3 SET_B.n2 178.222
R3 SET_B.n3 SET_B.n0 157.042
R4 SET_B.n0 SET_B.t0 143.898
R5 SET_B.n2 SET_B.n1 142.994
R6 SET_B SET_B.n3 5.0092
R7 SET_B.n3 SET_B 3.29747
R8 VGND.n36 VGND.t6 280.51
R9 VGND.n29 VGND.t9 244.153
R10 VGND.n52 VGND.t2 237.877
R11 VGND.n4 VGND.n3 205.707
R12 VGND.n15 VGND.n14 201.488
R13 VGND.n55 VGND.n54 199.739
R14 VGND.n13 VGND.t1 159.758
R15 VGND.n12 VGND.t7 150.457
R16 VGND.n22 VGND.n21 110.672
R17 VGND.n3 VGND.t10 75.7148
R18 VGND.n21 VGND.t8 57.8264
R19 VGND.n14 VGND.t4 54.2862
R20 VGND.n3 VGND.t5 38.5719
R21 VGND.n54 VGND.t12 38.5719
R22 VGND.n54 VGND.t11 38.5719
R23 VGND.n23 VGND.n10 34.6358
R24 VGND.n27 VGND.n10 34.6358
R25 VGND.n28 VGND.n27 34.6358
R26 VGND.n30 VGND.n28 34.6358
R27 VGND.n34 VGND.n8 34.6358
R28 VGND.n35 VGND.n34 34.6358
R29 VGND.n37 VGND.n35 34.6358
R30 VGND.n41 VGND.n6 34.6358
R31 VGND.n42 VGND.n41 34.6358
R32 VGND.n43 VGND.n42 34.6358
R33 VGND.n47 VGND.n46 34.6358
R34 VGND.n48 VGND.n47 34.6358
R35 VGND.n48 VGND.n1 34.6358
R36 VGND.n16 VGND.n15 28.6123
R37 VGND.n16 VGND.n12 27.1064
R38 VGND.n14 VGND.t0 25.9346
R39 VGND.n20 VGND.n12 24.8476
R40 VGND.n21 VGND.t3 24.7418
R41 VGND.n23 VGND.n22 23.3417
R42 VGND.n55 VGND.n53 22.9652
R43 VGND.n53 VGND.n52 22.2123
R44 VGND.n52 VGND.n1 21.4593
R45 VGND.n22 VGND.n20 21.0829
R46 VGND.n43 VGND.n4 18.4476
R47 VGND.n46 VGND.n4 16.1887
R48 VGND.n29 VGND.n8 10.9181
R49 VGND.n53 VGND.n0 9.3005
R50 VGND.n52 VGND.n51 9.3005
R51 VGND.n50 VGND.n1 9.3005
R52 VGND.n49 VGND.n48 9.3005
R53 VGND.n47 VGND.n2 9.3005
R54 VGND.n46 VGND.n45 9.3005
R55 VGND.n44 VGND.n43 9.3005
R56 VGND.n42 VGND.n5 9.3005
R57 VGND.n41 VGND.n40 9.3005
R58 VGND.n39 VGND.n6 9.3005
R59 VGND.n38 VGND.n37 9.3005
R60 VGND.n35 VGND.n7 9.3005
R61 VGND.n34 VGND.n33 9.3005
R62 VGND.n32 VGND.n8 9.3005
R63 VGND.n31 VGND.n30 9.3005
R64 VGND.n28 VGND.n9 9.3005
R65 VGND.n27 VGND.n26 9.3005
R66 VGND.n25 VGND.n10 9.3005
R67 VGND.n24 VGND.n23 9.3005
R68 VGND.n22 VGND.n11 9.3005
R69 VGND.n20 VGND.n19 9.3005
R70 VGND.n18 VGND.n12 9.3005
R71 VGND.n17 VGND.n16 9.3005
R72 VGND.n56 VGND.n55 7.12063
R73 VGND.n15 VGND.n13 6.27324
R74 VGND.n36 VGND.n6 5.27109
R75 VGND.n37 VGND.n36 4.51815
R76 VGND.n30 VGND.n29 4.14168
R77 VGND.n17 VGND.n13 0.689025
R78 VGND.n56 VGND.n0 0.148519
R79 VGND.n18 VGND.n17 0.120292
R80 VGND.n19 VGND.n18 0.120292
R81 VGND.n19 VGND.n11 0.120292
R82 VGND.n24 VGND.n11 0.120292
R83 VGND.n25 VGND.n24 0.120292
R84 VGND.n26 VGND.n25 0.120292
R85 VGND.n26 VGND.n9 0.120292
R86 VGND.n31 VGND.n9 0.120292
R87 VGND.n32 VGND.n31 0.120292
R88 VGND.n33 VGND.n32 0.120292
R89 VGND.n33 VGND.n7 0.120292
R90 VGND.n38 VGND.n7 0.120292
R91 VGND.n39 VGND.n38 0.120292
R92 VGND.n40 VGND.n39 0.120292
R93 VGND.n40 VGND.n5 0.120292
R94 VGND.n44 VGND.n5 0.120292
R95 VGND.n45 VGND.n44 0.120292
R96 VGND.n45 VGND.n2 0.120292
R97 VGND.n49 VGND.n2 0.120292
R98 VGND.n50 VGND.n49 0.120292
R99 VGND.n51 VGND.n50 0.120292
R100 VGND.n51 VGND.n0 0.120292
R101 VGND VGND.n56 0.11354
R102 a_790_47.n0 a_790_47.t2 463.795
R103 a_790_47.t1 a_790_47.n0 49.1523
R104 a_790_47.n0 a_790_47.t0 38.5719
R105 VNB.t12 VNB.t4 2904.85
R106 VNB.t10 VNB.t7 2790.94
R107 VNB.t17 VNB.t11 2733.98
R108 VNB.t16 VNB.t9 2677.02
R109 VNB.t19 VNB.t5 2677.02
R110 VNB.t13 VNB.t8 1566.34
R111 VNB.t20 VNB.t1 1552.1
R112 VNB.t0 VNB.t18 1537.86
R113 VNB.t8 VNB.t14 1423.95
R114 VNB.t11 VNB.t6 1381.23
R115 VNB.t18 VNB.t13 1366.99
R116 VNB.t7 VNB.t2 1352.75
R117 VNB.t1 VNB.t12 1352.75
R118 VNB.t9 VNB.t20 1352.75
R119 VNB.t5 VNB.t0 1352.75
R120 VNB.t2 VNB.t3 1196.12
R121 VNB.t6 VNB.t10 1196.12
R122 VNB.t4 VNB.t17 1196.12
R123 VNB.t14 VNB.t16 1196.12
R124 VNB.t15 VNB.t19 1196.12
R125 VNB VNB.t15 669.256
R126 a_944_21.t0 a_944_21.n3 734.475
R127 a_944_21.n1 a_944_21.t1 287.009
R128 a_944_21.n3 a_944_21.n2 211.846
R129 a_944_21.n0 a_944_21.t3 211.737
R130 a_944_21.n2 a_944_21.t2 210.474
R131 a_944_21.n0 a_944_21.t5 207.404
R132 a_944_21.n2 a_944_21.t4 204.048
R133 a_944_21.n1 a_944_21.n0 152
R134 a_944_21.n3 a_944_21.n1 9.77505
R135 a_650_21.n7 a_650_21.n0 598.178
R136 a_650_21.n8 a_650_21.n7 585
R137 a_650_21.n6 a_650_21.t4 387.961
R138 a_650_21.n3 a_650_21.n2 299.911
R139 a_650_21.n5 a_650_21.n3 215.817
R140 a_650_21.n5 a_650_21.n4 202.456
R141 a_650_21.n7 a_650_21.n6 190.656
R142 a_650_21.n3 a_650_21.t6 167.63
R143 a_650_21.n6 a_650_21.t5 143.746
R144 a_650_21.n1 a_650_21.t1 110.227
R145 a_650_21.n7 a_650_21.n5 81.1737
R146 a_650_21.t2 a_650_21.n0 63.3219
R147 a_650_21.t2 a_650_21.n8 63.3219
R148 a_650_21.n4 a_650_21.t0 25.313
R149 a_650_21.n4 a_650_21.t3 25.313
R150 a_650_21.n1 a_650_21.n0 9.38145
R151 a_650_21.n8 a_650_21.n1 9.38145
R152 a_1431_21.n7 a_1431_21.n6 594.413
R153 a_1431_21.n5 a_1431_21.t9 387.207
R154 a_1431_21.n2 a_1431_21.t4 308.481
R155 a_1431_21.n4 a_1431_21.n2 307.625
R156 a_1431_21.n4 a_1431_21.n3 275.635
R157 a_1431_21.n2 a_1431_21.t7 236.18
R158 a_1431_21.n0 a_1431_21.t11 231.476
R159 a_1431_21.n1 a_1431_21.t10 221.72
R160 a_1431_21.n6 a_1431_21.n5 204.841
R161 a_1431_21.n0 a_1431_21.t6 163.995
R162 a_1431_21.n1 a_1431_21.n0 151.742
R163 a_1431_21.n1 a_1431_21.t5 149.421
R164 a_1431_21.n5 a_1431_21.t8 142.994
R165 a_1431_21.n7 a_1431_21.t3 91.4648
R166 a_1431_21.n2 a_1431_21.n1 85.6894
R167 a_1431_21.t2 a_1431_21.n7 32.8338
R168 a_1431_21.n6 a_1431_21.n4 30.4946
R169 a_1431_21.n3 a_1431_21.t0 25.313
R170 a_1431_21.n3 a_1431_21.t1 25.313
R171 VPWR.n28 VPWR.t1 793.365
R172 VPWR.n21 VPWR.n20 732.75
R173 VPWR.n55 VPWR.t5 667.145
R174 VPWR.n57 VPWR.n1 604.394
R175 VPWR.n49 VPWR.n5 599.485
R176 VPWR.n35 VPWR.n34 585
R177 VPWR.n43 VPWR.t0 353.889
R178 VPWR.n15 VPWR.n14 315.236
R179 VPWR.n19 VPWR.t7 262.498
R180 VPWR.n16 VPWR.t3 255.554
R181 VPWR.n34 VPWR.t11 91.4648
R182 VPWR.n34 VPWR.t9 91.4648
R183 VPWR.n5 VPWR.t10 91.4648
R184 VPWR.n5 VPWR.t2 86.7743
R185 VPWR.n20 VPWR.t12 63.1021
R186 VPWR.n14 VPWR.t6 58.4849
R187 VPWR.n1 VPWR.t14 41.5552
R188 VPWR.n1 VPWR.t13 41.5552
R189 VPWR.n50 VPWR.n3 34.6358
R190 VPWR.n54 VPWR.n3 34.6358
R191 VPWR.n44 VPWR.n6 34.6358
R192 VPWR.n48 VPWR.n6 34.6358
R193 VPWR.n37 VPWR.n36 34.6358
R194 VPWR.n37 VPWR.n8 34.6358
R195 VPWR.n41 VPWR.n8 34.6358
R196 VPWR.n42 VPWR.n41 34.6358
R197 VPWR.n29 VPWR.n10 34.6358
R198 VPWR.n50 VPWR.n49 32.377
R199 VPWR.n14 VPWR.t4 31.831
R200 VPWR.n18 VPWR.n15 28.6123
R201 VPWR.n33 VPWR.n10 28.1331
R202 VPWR.n20 VPWR.t8 27.7871
R203 VPWR.n19 VPWR.n18 27.1064
R204 VPWR.n22 VPWR.n21 24.9229
R205 VPWR.n22 VPWR.n19 24.8476
R206 VPWR.n57 VPWR.n56 22.9652
R207 VPWR.n56 VPWR.n55 22.2123
R208 VPWR.n55 VPWR.n54 21.4593
R209 VPWR.n36 VPWR.n35 19.2758
R210 VPWR.n29 VPWR.n28 14.7581
R211 VPWR.n26 VPWR.n12 10.706
R212 VPWR.n27 VPWR.n26 10.706
R213 VPWR.n18 VPWR.n17 9.3005
R214 VPWR.n19 VPWR.n13 9.3005
R215 VPWR.n23 VPWR.n22 9.3005
R216 VPWR.n24 VPWR.n12 9.3005
R217 VPWR.n26 VPWR.n25 9.3005
R218 VPWR.n27 VPWR.n11 9.3005
R219 VPWR.n30 VPWR.n29 9.3005
R220 VPWR.n31 VPWR.n10 9.3005
R221 VPWR.n33 VPWR.n32 9.3005
R222 VPWR.n36 VPWR.n9 9.3005
R223 VPWR.n38 VPWR.n37 9.3005
R224 VPWR.n39 VPWR.n8 9.3005
R225 VPWR.n41 VPWR.n40 9.3005
R226 VPWR.n42 VPWR.n7 9.3005
R227 VPWR.n45 VPWR.n44 9.3005
R228 VPWR.n46 VPWR.n6 9.3005
R229 VPWR.n48 VPWR.n47 9.3005
R230 VPWR.n49 VPWR.n4 9.3005
R231 VPWR.n51 VPWR.n50 9.3005
R232 VPWR.n52 VPWR.n3 9.3005
R233 VPWR.n54 VPWR.n53 9.3005
R234 VPWR.n55 VPWR.n2 9.3005
R235 VPWR.n56 VPWR.n0 9.3005
R236 VPWR.n49 VPWR.n48 8.28285
R237 VPWR.n58 VPWR.n57 7.12063
R238 VPWR.n16 VPWR.n15 6.27324
R239 VPWR.n43 VPWR.n42 5.27109
R240 VPWR.n44 VPWR.n43 4.51815
R241 VPWR.n28 VPWR.n27 3.49141
R242 VPWR.n35 VPWR.n33 2.09505
R243 VPWR.n17 VPWR.n16 0.689025
R244 VPWR.n21 VPWR.n12 0.349591
R245 VPWR.n58 VPWR.n0 0.148519
R246 VPWR.n17 VPWR.n13 0.120292
R247 VPWR.n23 VPWR.n13 0.120292
R248 VPWR.n24 VPWR.n23 0.120292
R249 VPWR.n25 VPWR.n24 0.120292
R250 VPWR.n25 VPWR.n11 0.120292
R251 VPWR.n30 VPWR.n11 0.120292
R252 VPWR.n31 VPWR.n30 0.120292
R253 VPWR.n32 VPWR.n31 0.120292
R254 VPWR.n32 VPWR.n9 0.120292
R255 VPWR.n38 VPWR.n9 0.120292
R256 VPWR.n39 VPWR.n38 0.120292
R257 VPWR.n40 VPWR.n39 0.120292
R258 VPWR.n40 VPWR.n7 0.120292
R259 VPWR.n45 VPWR.n7 0.120292
R260 VPWR.n46 VPWR.n45 0.120292
R261 VPWR.n47 VPWR.n46 0.120292
R262 VPWR.n47 VPWR.n4 0.120292
R263 VPWR.n51 VPWR.n4 0.120292
R264 VPWR.n52 VPWR.n51 0.120292
R265 VPWR.n53 VPWR.n52 0.120292
R266 VPWR.n53 VPWR.n2 0.120292
R267 VPWR.n2 VPWR.n0 0.120292
R268 VPWR VPWR.n58 0.11354
R269 Q_N Q_N.n0 586.477
R270 Q_N.n3 Q_N.n0 585
R271 Q_N.n2 Q_N.n1 185
R272 Q_N Q_N.n2 80.821
R273 Q_N.n0 Q_N.t0 26.5955
R274 Q_N.n0 Q_N.t1 26.5955
R275 Q_N.n1 Q_N.t3 24.9236
R276 Q_N.n1 Q_N.t2 24.9236
R277 Q_N Q_N.n3 15.262
R278 Q_N.n2 Q_N 6.15435
R279 Q_N.n3 Q_N 1.47742
R280 VPB.t2 VPB.t10 1441.28
R281 VPB.t1 VPB.t14 603.739
R282 VPB.t9 VPB.t8 580.062
R283 VPB.t18 VPB.t7 556.386
R284 VPB.t0 VPB.t3 355.14
R285 VPB.t10 VPB.t13 319.627
R286 VPB.t12 VPB.t15 319.627
R287 VPB.t3 VPB.t12 313.707
R288 VPB.t14 VPB.t11 287.072
R289 VPB.t13 VPB.t6 284.113
R290 VPB.t8 VPB.t5 281.154
R291 VPB.t7 VPB.t17 281.154
R292 VPB.t5 VPB.t4 248.599
R293 VPB.t11 VPB.t9 248.599
R294 VPB.t17 VPB.t0 248.599
R295 VPB.t16 VPB.t18 248.599
R296 VPB.t15 VPB.t2 236.761
R297 VPB.t6 VPB.t1 213.084
R298 VPB VPB.t16 139.097
R299 a_476_47.n3 a_476_47.n2 706.313
R300 a_476_47.n2 a_476_47.n0 287.646
R301 a_476_47.n2 a_476_47.n1 218.335
R302 a_476_47.n1 a_476_47.t5 216.9
R303 a_476_47.n1 a_476_47.t4 210.474
R304 a_476_47.n0 a_476_47.t0 66.6672
R305 a_476_47.n0 a_476_47.t3 63.3338
R306 a_476_47.t1 a_476_47.n3 63.3219
R307 a_476_47.n3 a_476_47.t2 63.3219
R308 a_894_329.t0 a_894_329.t1 58.6315
R309 a_27_47.n2 a_27_47.t2 533.949
R310 a_27_47.t0 a_27_47.n6 420.863
R311 a_27_47.n1 a_27_47.n0 343.399
R312 a_27_47.n1 a_27_47.t6 283.3
R313 a_27_47.n5 a_27_47.t5 263.173
R314 a_27_47.n4 a_27_47.t1 261.099
R315 a_27_47.n5 a_27_47.t4 227.826
R316 a_27_47.n3 a_27_47.n2 164.069
R317 a_27_47.n6 a_27_47.n5 152
R318 a_27_47.n2 a_27_47.t3 141.923
R319 a_27_47.n6 a_27_47.n4 21.4266
R320 a_27_47.n3 a_27_47.n1 12.1819
R321 a_27_47.n4 a_27_47.n3 11.2438
R322 a_381_47.n1 a_381_47.n0 957.008
R323 a_381_47.t1 a_381_47.n1 89.1195
R324 a_381_47.n0 a_381_47.t0 63.3338
R325 a_381_47.n1 a_381_47.t2 63.3219
R326 a_381_47.n0 a_381_47.t3 29.7268
R327 a_584_47.t1 a_584_47.t0 93.5174
R328 a_2236_47.t0 a_2236_47.n2 390.522
R329 a_2236_47.n2 a_2236_47.t1 247.917
R330 a_2236_47.n0 a_2236_47.t2 212.081
R331 a_2236_47.n1 a_2236_47.t3 212.081
R332 a_2236_47.n2 a_2236_47.n1 186.331
R333 a_2236_47.n0 a_2236_47.t5 139.78
R334 a_2236_47.n1 a_2236_47.t4 139.78
R335 a_2236_47.n1 a_2236_47.n0 61.346
R336 Q Q.n0 586.948
R337 Q.n3 Q.n0 585
R338 Q.n2 Q.n1 185
R339 Q Q.n2 76.5674
R340 Q.n0 Q.t1 26.5955
R341 Q.n0 Q.t0 26.5955
R342 Q.n1 Q.t2 24.9236
R343 Q.n1 Q.t3 24.9236
R344 Q Q.n3 16.9744
R345 Q.n2 Q 7.51354
R346 Q.n3 Q 1.94833
R347 a_560_413.t0 a_560_413.t1 211.071
R348 a_1547_47.t0 a_1547_47.t1 508.594
R349 CLK_N.n0 CLK_N.t0 269.921
R350 CLK_N.n0 CLK_N.t1 234.573
R351 CLK_N.n1 CLK_N.n0 152
R352 CLK_N CLK_N.n1 7.57233
R353 CLK_N.n1 CLK_N 4.68782
R354 D.n0 D.t0 331.51
R355 D.n0 D.t1 209.403
R356 D.n1 D.n0 152
R357 D.n1 D 8.58587
R358 D D.n1 2.02977
R359 a_193_47.n1 a_193_47.t3 525.917
R360 a_193_47.t0 a_193_47.n4 366.837
R361 a_193_47.n2 a_193_47.t2 313.505
R362 a_193_47.n2 a_193_47.t4 307.325
R363 a_193_47.n4 a_193_47.t1 300.94
R364 a_193_47.n3 a_193_47.n1 171.565
R365 a_193_47.n1 a_193_47.n0 148.35
R366 a_193_47.n4 a_193_47.n3 10.4403
R367 a_193_47.n3 a_193_47.n2 9.3005
R368 a_1162_47.n1 a_1162_47.n0 67.2005
R369 a_1162_47.n0 a_1162_47.t0 66.6672
R370 a_1162_47.n0 a_1162_47.t1 13.144
R371 RESET_B.n0 RESET_B.t1 201.874
R372 RESET_B.n0 RESET_B.t0 172.953
R373 RESET_B RESET_B.n0 154
R374 a_1665_329.t0 a_1665_329.t1 49.2505
R375 a_1366_47.t0 a_1366_47.t1 93.0601
C0 a_1257_47# RESET_B 4.35e-20
C1 VPB SET_B 0.144443f
C2 RESET_B Q 3.82e-20
C3 a_1257_47# Q_N 9.31e-21
C4 VPB VPWR 0.28939f
C5 a_1115_329# VPWR 0.01609f
C6 CLK_N VPWR 0.017469f
C7 VPB VGND 0.019304f
C8 a_1343_413# VPWR 0.003713f
C9 a_1115_329# VGND 3.84e-19
C10 D VPWR 0.015584f
C11 VPB RESET_B 0.048783f
C12 CLK_N VGND 0.017237f
C13 SET_B VPWR 0.025073f
C14 D VGND 0.013747f
C15 VPB Q_N 0.004352f
C16 a_1257_47# VPB 0.056869f
C17 VPB Q 0.005441f
C18 SET_B VGND 0.290777f
C19 a_1257_47# a_1115_329# 0.004123f
C20 SET_B RESET_B 0.00223f
C21 VPWR VGND 0.124886f
C22 a_1257_47# a_1343_413# 0.009757f
C23 VPWR RESET_B 0.010297f
C24 SET_B Q_N 3.28e-19
C25 a_1257_47# SET_B 0.159109f
C26 VPWR Q_N 0.1383f
C27 SET_B Q 8.77e-20
C28 VGND RESET_B 0.029459f
C29 a_1257_47# VPWR 0.118743f
C30 VPB CLK_N 0.069762f
C31 VGND Q_N 0.134896f
C32 VPWR Q 0.17808f
C33 a_1257_47# VGND 0.13186f
C34 VPB D 0.082544f
C35 RESET_B Q_N 0.001683f
C36 VGND Q 0.112501f
C37 Q VNB 0.02603f
C38 Q_N VNB 0.010197f
C39 RESET_B VNB 0.135273f
C40 VGND VNB 1.4314f
C41 VPWR VNB 1.16512f
C42 SET_B VNB 0.261431f
C43 D VNB 0.125582f
C44 CLK_N VNB 0.195657f
C45 VPB VNB 2.55388f
C46 a_1257_47# VNB 0.119109f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfbbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfbbp_1 VGND VPWR VPB VNB Q Q_N SET_B D CLK
X0 a_788_47.t0 a_942_21.t1 a_648_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 VPWR.t2 RESET_B a_942_21.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1539 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 VGND a_1429_21# a_1364_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X3 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_381_47.t0 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_474_413.t3 a_27_47.t2 a_381_47.t3 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X6 VPWR.t9 a_1429_21# a_2136_47.t0 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_1429_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X8 a_582_47.t0 a_193_47.t2 a_474_413.t1 VNB.t4 sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X9 a_648_21.t3 a_474_413.t4 a_788_47.t2 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X10 a_1341_413.t0 a_193_47.t3 a_1255_47.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1160_47.t0 a_648_21.t4 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X12 a_193_47.t1 a_27_47.t3 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1255_47.t1 a_27_47.t4 a_1113_329.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1743 ps=1.41 w=0.42 l=0.15
X14 Q.t0 a_2136_47.t2 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X15 a_648_21.t2 SET_B.t0 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X16 a_788_47.t1 SET_B.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X17 Q_N.t0 a_1429_21# VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1539 ps=1.335 w=1 l=0.15
X18 Q.t1 a_2136_47.t3 VGND.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X19 VPWR.t1 a_942_21.t2 a_892_329.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2247 pd=1.375 as=0.1134 ps=1.11 w=0.84 l=0.15
X20 a_558_413.t0 a_27_47.t5 a_474_413.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND.t7 a_648_21.t5 a_582_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.06705 ps=0.75 w=0.42 l=0.15
X22 a_892_329.t1 a_474_413.t5 a_648_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X23 VGND.t9 a_1429_21# a_2136_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_193_47.t0 a_27_47.t6 VPWR.t6 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_474_413.t0 a_193_47.t4 a_381_47.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X26 a_1364_47# a_27_47.t7 a_1255_47.t2 VNB.t9 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X27 Q_N.t1 a_1429_21# VGND.t8 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X28 a_1545_47# SET_B.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1199 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 VPWR.t7 a_648_21.t6 a_558_413.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X30 a_381_47.t1 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_1113_329.t1 a_648_21.t7 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1743 pd=1.41 as=0.2247 ps=1.375 w=0.84 l=0.15
X32 VGND.t5 CLK.t1 a_27_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_942_21.t0 a_942_21.n4 740.164
R1 a_942_21.n4 a_942_21.n3 211.846
R2 a_942_21.n2 a_942_21.n1 211.737
R3 a_942_21.n3 a_942_21.t1 210.474
R4 a_942_21.n2 a_942_21.n0 207.404
R5 a_942_21.n3 a_942_21.t2 204.048
R6 a_942_21.n4 a_942_21.n2 161.775
R7 a_648_21.n6 a_648_21.n0 598.178
R8 a_648_21.n7 a_648_21.n6 585
R9 a_648_21.n5 a_648_21.t5 387.961
R10 a_648_21.n2 a_648_21.t7 299.911
R11 a_648_21.n4 a_648_21.n2 215.817
R12 a_648_21.n4 a_648_21.n3 202.456
R13 a_648_21.n6 a_648_21.n5 190.656
R14 a_648_21.n2 a_648_21.t4 167.63
R15 a_648_21.n5 a_648_21.t6 143.746
R16 a_648_21.n1 a_648_21.t2 110.227
R17 a_648_21.n6 a_648_21.n4 81.1737
R18 a_648_21.t1 a_648_21.n0 63.3219
R19 a_648_21.t1 a_648_21.n7 63.3219
R20 a_648_21.n3 a_648_21.t0 25.313
R21 a_648_21.n3 a_648_21.t3 25.313
R22 a_648_21.n1 a_648_21.n0 9.38145
R23 a_648_21.n7 a_648_21.n1 9.38145
R24 a_788_47.t0 a_788_47.n0 468.854
R25 a_788_47.n0 a_788_47.t2 49.1523
R26 a_788_47.n0 a_788_47.t1 38.5719
R27 VNB.t3 VNB.t13 6906.15
R28 VNB.t11 VNB.t9 2904.85
R29 VNB.t13 VNB.t14 2677.02
R30 VNB.t1 VNB.t11 2677.02
R31 VNB.t6 VNB.t0 2677.02
R32 VNB.t9 VNB.t3 2577.35
R33 VNB.t10 VNB.t2 1566.34
R34 VNB.t5 VNB.t4 1509.39
R35 VNB.t2 VNB.t12 1423.95
R36 VNB.t4 VNB.t10 1366.99
R37 VNB.t14 VNB.t7 1352.75
R38 VNB.t0 VNB.t5 1352.75
R39 VNB.t12 VNB.t1 1196.12
R40 VNB.t8 VNB.t6 1196.12
R41 VNB VNB.t8 669.256
R42 VPWR.n14 VPWR.n13 732.75
R43 VPWR.n44 VPWR.t0 666.607
R44 VPWR.n46 VPWR.n1 604.394
R45 VPWR.n38 VPWR.n5 599.485
R46 VPWR.n16 VPWR.n15 321.339
R47 VPWR.n32 VPWR.n8 310.502
R48 VPWR.n5 VPWR.t5 91.4648
R49 VPWR.n5 VPWR.t7 86.7743
R50 VPWR.n8 VPWR.t8 86.7743
R51 VPWR.n13 VPWR.t2 63.1021
R52 VPWR.n15 VPWR.t9 58.4849
R53 VPWR.n1 VPWR.t6 41.5552
R54 VPWR.n1 VPWR.t3 41.5552
R55 VPWR.n8 VPWR.t1 38.6969
R56 VPWR.n39 VPWR.n3 34.6358
R57 VPWR.n43 VPWR.n3 34.6358
R58 VPWR.n33 VPWR.n6 34.6358
R59 VPWR.n37 VPWR.n6 34.6358
R60 VPWR.n26 VPWR.n25 34.6358
R61 VPWR.n26 VPWR.n9 34.6358
R62 VPWR.n30 VPWR.n9 34.6358
R63 VPWR.n31 VPWR.n30 34.6358
R64 VPWR.n20 VPWR.n11 34.6358
R65 VPWR.n15 VPWR.t4 31.831
R66 VPWR.n39 VPWR.n38 31.624
R67 VPWR.n24 VPWR.n11 28.6533
R68 VPWR.n13 VPWR.t10 28.0332
R69 VPWR.n46 VPWR.n45 22.9652
R70 VPWR.n45 VPWR.n44 21.4593
R71 VPWR.n44 VPWR.n43 21.4593
R72 VPWR.n25 VPWR.n24 20.8501
R73 VPWR.n20 VPWR.n19 17.7288
R74 VPWR.n19 VPWR.n18 10.706
R75 VPWR.n18 VPWR.n14 10.1241
R76 VPWR.n18 VPWR.n17 9.3005
R77 VPWR.n19 VPWR.n12 9.3005
R78 VPWR.n21 VPWR.n20 9.3005
R79 VPWR.n22 VPWR.n11 9.3005
R80 VPWR.n24 VPWR.n23 9.3005
R81 VPWR.n25 VPWR.n10 9.3005
R82 VPWR.n27 VPWR.n26 9.3005
R83 VPWR.n28 VPWR.n9 9.3005
R84 VPWR.n30 VPWR.n29 9.3005
R85 VPWR.n31 VPWR.n7 9.3005
R86 VPWR.n34 VPWR.n33 9.3005
R87 VPWR.n35 VPWR.n6 9.3005
R88 VPWR.n37 VPWR.n36 9.3005
R89 VPWR.n38 VPWR.n4 9.3005
R90 VPWR.n40 VPWR.n39 9.3005
R91 VPWR.n41 VPWR.n3 9.3005
R92 VPWR.n43 VPWR.n42 9.3005
R93 VPWR.n44 VPWR.n2 9.3005
R94 VPWR.n45 VPWR.n0 9.3005
R95 VPWR.n38 VPWR.n37 9.03579
R96 VPWR.n16 VPWR.n14 7.84364
R97 VPWR.n47 VPWR.n46 7.12063
R98 VPWR.n32 VPWR.n31 6.02403
R99 VPWR.n33 VPWR.n32 3.76521
R100 VPWR.n17 VPWR.n16 0.211436
R101 VPWR.n47 VPWR.n0 0.148519
R102 VPWR.n17 VPWR.n12 0.120292
R103 VPWR.n21 VPWR.n12 0.120292
R104 VPWR.n22 VPWR.n21 0.120292
R105 VPWR.n23 VPWR.n22 0.120292
R106 VPWR.n23 VPWR.n10 0.120292
R107 VPWR.n27 VPWR.n10 0.120292
R108 VPWR.n28 VPWR.n27 0.120292
R109 VPWR.n29 VPWR.n28 0.120292
R110 VPWR.n29 VPWR.n7 0.120292
R111 VPWR.n34 VPWR.n7 0.120292
R112 VPWR.n35 VPWR.n34 0.120292
R113 VPWR.n36 VPWR.n35 0.120292
R114 VPWR.n36 VPWR.n4 0.120292
R115 VPWR.n40 VPWR.n4 0.120292
R116 VPWR.n41 VPWR.n40 0.120292
R117 VPWR.n42 VPWR.n41 0.120292
R118 VPWR.n42 VPWR.n2 0.120292
R119 VPWR.n2 VPWR.n0 0.120292
R120 VPWR VPWR.n47 0.11354
R121 VPB.t6 VPB.t3 1752.02
R122 VPB.t14 VPB.t15 556.386
R123 VPB.t11 VPB.t0 556.386
R124 VPB.t12 VPB.t9 426.168
R125 VPB.t2 VPB.t12 405.452
R126 VPB.t10 VPB.t13 355.14
R127 VPB.t8 VPB.t5 319.627
R128 VPB.t13 VPB.t8 313.707
R129 VPB.t3 VPB.t14 287.072
R130 VPB.t15 VPB.t7 281.154
R131 VPB.t0 VPB.t1 275.235
R132 VPB.t9 VPB.t6 248.599
R133 VPB.t5 VPB.t2 248.599
R134 VPB.t1 VPB.t10 248.599
R135 VPB.t4 VPB.t11 248.599
R136 VPB VPB.t4 139.097
R137 VGND.n27 VGND.t6 280.51
R138 VGND.n20 VGND.t2 241.294
R139 VGND.n43 VGND.t0 237.47
R140 VGND.n13 VGND.t8 225.673
R141 VGND.n12 VGND.n11 207.585
R142 VGND.n4 VGND.n3 205.707
R143 VGND.n46 VGND.n45 199.739
R144 VGND.n3 VGND.t7 75.7148
R145 VGND.n11 VGND.t9 54.2862
R146 VGND.n3 VGND.t1 38.5719
R147 VGND.n45 VGND.t3 38.5719
R148 VGND.n45 VGND.t5 38.5719
R149 VGND.n14 VGND.n10 34.6358
R150 VGND.n18 VGND.n10 34.6358
R151 VGND.n19 VGND.n18 34.6358
R152 VGND.n21 VGND.n19 34.6358
R153 VGND.n25 VGND.n8 34.6358
R154 VGND.n26 VGND.n25 34.6358
R155 VGND.n28 VGND.n26 34.6358
R156 VGND.n32 VGND.n6 34.6358
R157 VGND.n33 VGND.n32 34.6358
R158 VGND.n34 VGND.n33 34.6358
R159 VGND.n38 VGND.n37 34.6358
R160 VGND.n39 VGND.n38 34.6358
R161 VGND.n39 VGND.n1 34.6358
R162 VGND.n11 VGND.t4 25.9346
R163 VGND.n46 VGND.n44 22.9652
R164 VGND.n43 VGND.n1 21.4593
R165 VGND.n44 VGND.n43 21.4593
R166 VGND.n14 VGND.n13 20.3299
R167 VGND.n34 VGND.n4 19.2005
R168 VGND.n37 VGND.n4 15.4358
R169 VGND.n20 VGND.n8 10.1652
R170 VGND.n15 VGND.n14 9.3005
R171 VGND.n16 VGND.n10 9.3005
R172 VGND.n18 VGND.n17 9.3005
R173 VGND.n19 VGND.n9 9.3005
R174 VGND.n22 VGND.n21 9.3005
R175 VGND.n23 VGND.n8 9.3005
R176 VGND.n25 VGND.n24 9.3005
R177 VGND.n26 VGND.n7 9.3005
R178 VGND.n29 VGND.n28 9.3005
R179 VGND.n30 VGND.n6 9.3005
R180 VGND.n32 VGND.n31 9.3005
R181 VGND.n33 VGND.n5 9.3005
R182 VGND.n35 VGND.n34 9.3005
R183 VGND.n37 VGND.n36 9.3005
R184 VGND.n38 VGND.n2 9.3005
R185 VGND.n40 VGND.n39 9.3005
R186 VGND.n41 VGND.n1 9.3005
R187 VGND.n43 VGND.n42 9.3005
R188 VGND.n44 VGND.n0 9.3005
R189 VGND.n47 VGND.n46 7.12063
R190 VGND.n13 VGND.n12 7.10028
R191 VGND.n28 VGND.n27 5.27109
R192 VGND.n21 VGND.n20 4.89462
R193 VGND.n27 VGND.n6 4.51815
R194 VGND.n15 VGND.n12 0.218617
R195 VGND.n47 VGND.n0 0.148519
R196 VGND.n16 VGND.n15 0.120292
R197 VGND.n17 VGND.n16 0.120292
R198 VGND.n17 VGND.n9 0.120292
R199 VGND.n22 VGND.n9 0.120292
R200 VGND.n23 VGND.n22 0.120292
R201 VGND.n24 VGND.n23 0.120292
R202 VGND.n24 VGND.n7 0.120292
R203 VGND.n29 VGND.n7 0.120292
R204 VGND.n30 VGND.n29 0.120292
R205 VGND.n31 VGND.n30 0.120292
R206 VGND.n31 VGND.n5 0.120292
R207 VGND.n35 VGND.n5 0.120292
R208 VGND.n36 VGND.n35 0.120292
R209 VGND.n36 VGND.n2 0.120292
R210 VGND.n40 VGND.n2 0.120292
R211 VGND.n41 VGND.n40 0.120292
R212 VGND.n42 VGND.n41 0.120292
R213 VGND.n42 VGND.n0 0.120292
R214 VGND VGND.n47 0.11354
R215 CLK.n0 CLK.t0 269.921
R216 CLK.n0 CLK.t1 234.573
R217 CLK.n1 CLK.n0 152
R218 CLK CLK.n1 7.57233
R219 CLK.n1 CLK 4.68782
R220 a_27_47.n2 a_27_47.t7 525.917
R221 a_27_47.t0 a_27_47.n5 385.524
R222 a_27_47.n3 a_27_47.t2 314.259
R223 a_27_47.n3 a_27_47.t5 307.325
R224 a_27_47.n1 a_27_47.t1 282.524
R225 a_27_47.n0 a_27_47.t6 263.173
R226 a_27_47.n0 a_27_47.t3 227.826
R227 a_27_47.n4 a_27_47.n2 171.565
R228 a_27_47.n1 a_27_47.n0 152
R229 a_27_47.n2 a_27_47.t4 148.35
R230 a_27_47.n5 a_27_47.n1 35.3396
R231 a_27_47.n5 a_27_47.n4 10.842
R232 a_27_47.n4 a_27_47.n3 9.3005
R233 D.n0 D.t0 331.51
R234 D.n0 D.t1 209.403
R235 D.n1 D.n0 152
R236 D.n1 D 8.58587
R237 D D.n1 2.02977
R238 a_381_47.n1 a_381_47.n0 958.433
R239 a_381_47.n1 a_381_47.t2 84.4291
R240 a_381_47.n0 a_381_47.t3 63.3338
R241 a_381_47.t0 a_381_47.n1 63.3219
R242 a_381_47.n0 a_381_47.t1 29.7268
R243 a_474_413.n3 a_474_413.n2 706.313
R244 a_474_413.n2 a_474_413.n0 287.646
R245 a_474_413.n2 a_474_413.n1 218.335
R246 a_474_413.n1 a_474_413.t4 216.9
R247 a_474_413.n1 a_474_413.t5 210.474
R248 a_474_413.n0 a_474_413.t1 63.3338
R249 a_474_413.n0 a_474_413.t3 63.3338
R250 a_474_413.n3 a_474_413.t2 63.3219
R251 a_474_413.t0 a_474_413.n3 63.3219
R252 a_2136_47.t0 a_2136_47.n1 384.125
R253 a_2136_47.n1 a_2136_47.t1 243.28
R254 a_2136_47.n0 a_2136_47.t2 239.04
R255 a_2136_47.n1 a_2136_47.n0 175.079
R256 a_2136_47.n0 a_2136_47.t3 166.739
R257 SET_B.n0 SET_B.t0 389.618
R258 SET_B.n2 SET_B.n1 387.207
R259 SET_B.n3 SET_B.n2 178.222
R260 SET_B.n3 SET_B.n0 157.042
R261 SET_B.n0 SET_B.t1 143.898
R262 SET_B.n2 SET_B.t2 142.994
R263 SET_B SET_B.n3 5.0092
R264 SET_B.n3 SET_B 3.29747
R265 a_193_47.n2 a_193_47.t4 533.949
R266 a_193_47.t0 a_193_47.n4 424.863
R267 a_193_47.n1 a_193_47.t3 343.399
R268 a_193_47.n1 a_193_47.n0 283.3
R269 a_193_47.n4 a_193_47.t1 242.915
R270 a_193_47.n3 a_193_47.n2 164.069
R271 a_193_47.n2 a_193_47.t2 141.923
R272 a_193_47.n3 a_193_47.n1 12.1819
R273 a_193_47.n4 a_193_47.n3 10.8242
R274 a_582_47.t1 a_582_47.t0 93.5174
R275 a_1255_47.n4 a_1255_47.n3 692.294
R276 a_1255_47.n3 a_1255_47.t2 337.603
R277 a_1255_47.n2 a_1255_47.n0 241.536
R278 a_1255_47.n3 a_1255_47.n2 235.919
R279 a_1255_47.n2 a_1255_47.n1 196.549
R280 a_1255_47.t0 a_1255_47.n4 63.3219
R281 a_1255_47.n4 a_1255_47.t1 63.3219
R282 a_1160_47.n0 a_1160_47.t0 80.344
R283 a_1113_329.t1 a_1113_329.t0 236.869
R284 Q.n1 Q.t0 353.606
R285 Q.n0 Q.t1 209.923
R286 Q Q.n0 66.6967
R287 Q.n1 Q 9.10538
R288 Q Q.n1 7.47898
R289 Q.n0 Q 6.64665
R290 Q_N.n1 Q_N.t0 353.795
R291 Q_N.n0 Q_N.t1 209.923
R292 Q_N Q_N.n0 71.5041
R293 Q_N.n1 Q_N 8.2361
R294 Q_N Q_N.n1 6.90173
R295 Q_N.n0 Q_N 5.61454
R296 a_892_329.t0 a_892_329.t1 63.3219
R297 a_558_413.t0 a_558_413.t1 211.071
C0 a_1429_21# VPB 0.238464f
C1 RESET_B VPB 0.043004f
C2 a_1545_47# a_1364_47# 4.11e-20
C3 VPB Q_N 0.010057f
C4 CLK VGND 0.017237f
C5 D VPWR 0.015381f
C6 SET_B VPWR 0.025232f
C7 D VGND 0.013539f
C8 VPB Q 0.012256f
C9 a_1545_47# VPB 1.97e-19
C10 SET_B VGND 0.290779f
C11 a_1429_21# SET_B 0.140985f
C12 RESET_B SET_B 0.002256f
C13 a_1663_329# VPWR 0.00506f
C14 VPWR VGND 0.0797f
C15 SET_B Q_N 3.6e-19
C16 a_1429_21# VPWR 0.314499f
C17 RESET_B VPWR 0.009365f
C18 VPWR Q_N 0.061564f
C19 SET_B Q 1.21e-19
C20 a_1429_21# a_1663_329# 0.009453f
C21 a_1429_21# VGND 0.080687f
C22 a_1663_329# Q_N 2.02e-20
C23 RESET_B VGND 0.027687f
C24 a_1545_47# SET_B 0.009502f
C25 VGND Q_N 0.086785f
C26 VPWR Q 0.099216f
C27 a_1429_21# RESET_B 0.087267f
C28 a_1429_21# Q_N 0.123549f
C29 VPB CLK 0.069762f
C30 a_1364_47# SET_B 7.87e-19
C31 RESET_B Q_N 0.001792f
C32 a_1545_47# VPWR 2.86e-19
C33 VGND Q 0.064368f
C34 a_1429_21# Q 0.003171f
C35 a_1545_47# VGND 0.148823f
C36 RESET_B Q 6.25e-20
C37 VPB D 0.081987f
C38 a_1429_21# a_1545_47# 0.039699f
C39 RESET_B a_1545_47# 3.78e-20
C40 VPB SET_B 0.144156f
C41 a_1364_47# VGND 0.001916f
C42 a_1429_21# a_1364_47# 4.2e-20
C43 VPB VPWR 0.253857f
C44 CLK VPWR 0.017469f
C45 VPB VGND 0.015287f
C46 Q VNB 0.094496f
C47 Q_N VNB 0.013395f
C48 VGND VNB 1.30599f
C49 VPWR VNB 1.0532f
C50 SET_B VNB 0.262073f
C51 D VNB 0.12546f
C52 CLK VNB 0.195657f
C53 VPB VNB 2.37668f
C54 a_1545_47# VNB 0.008364f
C55 RESET_B VNB 0.126892f
C56 a_1429_21# VNB 0.391416f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_1 VGND VPWR VPB VNB CLK D RESET_B Q Q_N
X0 Q.t0 a_1283_21.t3 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X1 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VPWR.t2 a_1283_21.t4 a_1847_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_1217_47.t1 a_27_47.t2 a_1108_47.t1 VNB.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4 a_1283_21.t1 a_1108_47.t4 a_1462_47.t0 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413.t1 a_27_47.t3 a_543_47.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 a_1108_47.t2 a_193_47.t2 a_761_289.t0 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND.t1 RESET_B.t0 a_805_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR.t5 CLK.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 Q_N.t1 a_1847_47.t2 VGND.t7 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10 a_448_47.t1 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND.t5 a_1283_21.t5 a_1847_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_761_289.t2 a_543_47.t4 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X13 Q.t1 a_1283_21.t6 VGND.t4 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_193_47.t1 a_27_47.t4 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1108_47.t0 a_27_47.t5 a_761_289.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X16 a_1462_47.t1 RESET_B.t1 VGND.t0 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X17 a_543_47.t0 a_27_47.t6 a_448_47.t0 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X18 a_543_47.t3 a_193_47.t3 a_448_47.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X19 a_448_47.t2 D.t1 VGND.t9 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X20 VPWR.t3 a_1283_21.t7 a_1270_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR.t9 a_1108_47.t5 a_1283_21.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1270_413.t1 a_193_47.t4 a_1108_47.t3 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47.t0 a_27_47.t7 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21.t0 RESET_B.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR.t4 a_761_289.t5 a_651_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X26 a_639_47.t1 a_193_47.t5 a_543_47.t2 VNB.t6 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 Q_N.t0 a_1847_47.t3 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X28 VGND.t3 a_1283_21.t8 a_1217_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X29 a_651_413.t2 RESET_B.t3 VPWR.t11 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X30 VGND.t2 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_761_289.t3 a_543_47.t5 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
R0 a_1283_21.n6 a_1283_21.n5 746.659
R1 a_1283_21.n0 a_1283_21.t7 389.183
R2 a_1283_21.n2 a_1283_21.t4 256.988
R3 a_1283_21.n1 a_1283_21.n0 251.167
R4 a_1283_21.n1 a_1283_21.t1 223.571
R5 a_1283_21.n4 a_1283_21.t3 212.081
R6 a_1283_21.n5 a_1283_21.n4 181.942
R7 a_1283_21.n0 a_1283_21.t8 174.891
R8 a_1283_21.n2 a_1283_21.t5 163.803
R9 a_1283_21.n3 a_1283_21.t6 139.78
R10 a_1283_21.n3 a_1283_21.n2 129.264
R11 a_1283_21.n6 a_1283_21.t2 63.3219
R12 a_1283_21.t0 a_1283_21.n6 63.3219
R13 a_1283_21.n5 a_1283_21.n1 24.6993
R14 a_1283_21.n4 a_1283_21.n3 22.6399
R15 VPWR.n26 VPWR.t8 806.511
R16 VPWR.n2 VPWR.t0 667.778
R17 VPWR.n20 VPWR.n9 604.457
R18 VPWR.n42 VPWR.n1 604.394
R19 VPWR.n29 VPWR.n28 601.679
R20 VPWR.n13 VPWR.n10 585
R21 VPWR.n15 VPWR.n14 585
R22 VPWR.n12 VPWR.n11 251.434
R23 VPWR.n14 VPWR.n13 182.929
R24 VPWR.n9 VPWR.t3 119.608
R25 VPWR.n28 VPWR.t4 93.81
R26 VPWR.n13 VPWR.t9 68.0124
R27 VPWR.n28 VPWR.t11 63.3219
R28 VPWR.n9 VPWR.t6 63.3219
R29 VPWR.n11 VPWR.t2 61.9826
R30 VPWR.n1 VPWR.t7 41.5552
R31 VPWR.n1 VPWR.t5 41.5552
R32 VPWR.n41 VPWR.n40 34.6358
R33 VPWR.n34 VPWR.n4 34.6358
R34 VPWR.n35 VPWR.n34 34.6358
R35 VPWR.n36 VPWR.n35 34.6358
R36 VPWR.n30 VPWR.n27 34.6358
R37 VPWR.n21 VPWR.n7 34.6358
R38 VPWR.n25 VPWR.n7 34.6358
R39 VPWR.n36 VPWR.n2 32.377
R40 VPWR.n26 VPWR.n25 32.0005
R41 VPWR.n11 VPWR.t10 30.1738
R42 VPWR.n20 VPWR.n19 30.1181
R43 VPWR.n14 VPWR.t1 29.316
R44 VPWR.n42 VPWR.n41 22.9652
R45 VPWR.n21 VPWR.n20 20.3299
R46 VPWR.n40 VPWR.n2 18.0711
R47 VPWR.n15 VPWR.n12 17.4004
R48 VPWR.n19 VPWR.n10 12.8758
R49 VPWR.n27 VPWR.n26 9.41227
R50 VPWR.n17 VPWR.n16 9.3005
R51 VPWR.n19 VPWR.n18 9.3005
R52 VPWR.n20 VPWR.n8 9.3005
R53 VPWR.n22 VPWR.n21 9.3005
R54 VPWR.n23 VPWR.n7 9.3005
R55 VPWR.n25 VPWR.n24 9.3005
R56 VPWR.n26 VPWR.n6 9.3005
R57 VPWR.n27 VPWR.n5 9.3005
R58 VPWR.n31 VPWR.n30 9.3005
R59 VPWR.n32 VPWR.n4 9.3005
R60 VPWR.n34 VPWR.n33 9.3005
R61 VPWR.n35 VPWR.n3 9.3005
R62 VPWR.n37 VPWR.n36 9.3005
R63 VPWR.n38 VPWR.n2 9.3005
R64 VPWR.n40 VPWR.n39 9.3005
R65 VPWR.n41 VPWR.n0 9.3005
R66 VPWR.n43 VPWR.n42 7.12063
R67 VPWR.n29 VPWR.n4 6.02403
R68 VPWR.n16 VPWR.n15 5.00414
R69 VPWR.n16 VPWR.n10 4.07323
R70 VPWR.n30 VPWR.n29 3.76521
R71 VPWR.n17 VPWR.n12 0.211448
R72 VPWR.n43 VPWR.n0 0.148519
R73 VPWR.n18 VPWR.n17 0.120292
R74 VPWR.n18 VPWR.n8 0.120292
R75 VPWR.n22 VPWR.n8 0.120292
R76 VPWR.n23 VPWR.n22 0.120292
R77 VPWR.n24 VPWR.n23 0.120292
R78 VPWR.n24 VPWR.n6 0.120292
R79 VPWR.n6 VPWR.n5 0.120292
R80 VPWR.n31 VPWR.n5 0.120292
R81 VPWR.n32 VPWR.n31 0.120292
R82 VPWR.n33 VPWR.n32 0.120292
R83 VPWR.n33 VPWR.n3 0.120292
R84 VPWR.n37 VPWR.n3 0.120292
R85 VPWR.n38 VPWR.n37 0.120292
R86 VPWR.n39 VPWR.n38 0.120292
R87 VPWR.n39 VPWR.n0 0.120292
R88 VPWR VPWR.n43 0.114842
R89 Q Q.t0 246.839
R90 Q Q.t1 148.597
R91 VPB.t10 VPB.t0 790.188
R92 VPB.t3 VPB.t2 648.131
R93 VPB.t14 VPB.t11 583.023
R94 VPB.t12 VPB.t3 485.358
R95 VPB.t8 VPB.t4 414.33
R96 VPB.t1 VPB.t6 319.627
R97 VPB.t11 VPB.t9 292.991
R98 VPB.t7 VPB.t8 292.991
R99 VPB.t2 VPB.t13 287.072
R100 VPB.t4 VPB.t14 287.072
R101 VPB.t0 VPB.t7 272.274
R102 VPB.t9 VPB.t15 254.518
R103 VPB.t6 VPB.t12 248.599
R104 VPB.t15 VPB.t1 248.599
R105 VPB.t5 VPB.t10 248.599
R106 VPB VPB.t5 192.369
R107 a_761_289.n3 a_761_289.n2 647.119
R108 a_761_289.n1 a_761_289.t4 350.253
R109 a_761_289.n2 a_761_289.n0 260.339
R110 a_761_289.n2 a_761_289.n1 246.119
R111 a_761_289.n1 a_761_289.t5 189.588
R112 a_761_289.n3 a_761_289.t1 89.1195
R113 a_761_289.n0 a_761_289.t0 63.3338
R114 a_761_289.t3 a_761_289.n3 41.0422
R115 a_761_289.n0 a_761_289.t2 31.9797
R116 a_639_47.t0 a_639_47.t1 198.571
R117 a_805_47.t0 a_805_47.t1 60.0005
R118 VNB.t9 VNB.t15 3631.07
R119 VNB.t2 VNB.t3 2677.02
R120 VNB.t13 VNB.t2 2677.02
R121 VNB.t6 VNB.t5 2363.75
R122 VNB.t1 VNB.t14 2121.68
R123 VNB.t11 VNB.t12 1879.61
R124 VNB.t7 VNB.t8 1552.1
R125 VNB.t12 VNB.t7 1409.71
R126 VNB.t3 VNB.t4 1381.23
R127 VNB.t8 VNB.t1 1366.99
R128 VNB.t10 VNB.t6 1366.99
R129 VNB.t15 VNB.t10 1352.75
R130 VNB.t14 VNB.t13 1295.79
R131 VNB.t0 VNB.t9 1196.12
R132 VNB.t5 VNB.t11 1025.24
R133 VNB VNB.t0 925.567
R134 a_1847_47.t0 a_1847_47.n1 386.31
R135 a_1847_47.n1 a_1847_47.t1 249.956
R136 a_1847_47.n0 a_1847_47.t3 239.04
R137 a_1847_47.n1 a_1847_47.n0 175.661
R138 a_1847_47.n0 a_1847_47.t2 166.739
R139 a_27_47.n1 a_27_47.t3 530.01
R140 a_27_47.t1 a_27_47.n5 421.021
R141 a_27_47.n0 a_27_47.t5 337.142
R142 a_27_47.n3 a_27_47.t0 280.223
R143 a_27_47.n4 a_27_47.t7 263.173
R144 a_27_47.n4 a_27_47.t4 227.826
R145 a_27_47.n0 a_27_47.t2 199.762
R146 a_27_47.n2 a_27_47.n1 170.81
R147 a_27_47.n2 a_27_47.n0 167.321
R148 a_27_47.n5 a_27_47.n4 152
R149 a_27_47.n1 a_27_47.t6 141.923
R150 a_27_47.n3 a_27_47.n2 10.8376
R151 a_27_47.n5 a_27_47.n3 2.50485
R152 a_1108_47.n3 a_1108_47.n2 636.953
R153 a_1108_47.n1 a_1108_47.t4 366.856
R154 a_1108_47.n2 a_1108_47.n0 300.2
R155 a_1108_47.n2 a_1108_47.n1 225.036
R156 a_1108_47.n1 a_1108_47.t5 174.056
R157 a_1108_47.n0 a_1108_47.t2 70.0005
R158 a_1108_47.t0 a_1108_47.n3 68.0124
R159 a_1108_47.n3 a_1108_47.t3 63.3219
R160 a_1108_47.n0 a_1108_47.t1 61.6672
R161 a_1217_47.t0 a_1217_47.t1 94.7268
R162 a_1462_47.t0 a_1462_47.t1 87.1434
R163 a_543_47.n3 a_543_47.n2 674.338
R164 a_543_47.n1 a_543_47.t5 332.58
R165 a_543_47.n2 a_543_47.n0 284.012
R166 a_543_47.n2 a_543_47.n1 253.648
R167 a_543_47.n1 a_543_47.t4 168.701
R168 a_543_47.t1 a_543_47.n3 96.1553
R169 a_543_47.n3 a_543_47.t3 65.6672
R170 a_543_47.n0 a_543_47.t0 65.0005
R171 a_543_47.n0 a_543_47.t2 45.0005
R172 a_651_413.n0 a_651_413.t2 1327.82
R173 a_651_413.n0 a_651_413.t1 194.655
R174 a_651_413.t0 a_651_413.n0 63.3219
R175 a_193_47.t0 a_193_47.n3 370.026
R176 a_193_47.n0 a_193_47.t2 351.356
R177 a_193_47.n1 a_193_47.t5 334.717
R178 a_193_47.n3 a_193_47.t1 325.971
R179 a_193_47.n1 a_193_47.t3 309.935
R180 a_193_47.n0 a_193_47.t4 305.683
R181 a_193_47.n2 a_193_47.n0 16.879
R182 a_193_47.n3 a_193_47.n2 10.8867
R183 a_193_47.n2 a_193_47.n1 9.3005
R184 RESET_B.n1 RESET_B.t3 408.63
R185 RESET_B.n3 RESET_B.t2 347.577
R186 RESET_B.n3 RESET_B.t1 193.337
R187 RESET_B.n2 RESET_B.n1 167.575
R188 RESET_B.n4 RESET_B.n3 152
R189 RESET_B.n1 RESET_B.t0 132.282
R190 RESET_B RESET_B.n0 14.0185
R191 RESET_B.n4 RESET_B.n2 12.1952
R192 RESET_B.n2 RESET_B.n0 9.38606
R193 RESET_B RESET_B.n4 4.67077
R194 RESET_B.n0 RESET_B 4.53383
R195 VGND.n37 VGND.t9 307.536
R196 VGND.n10 VGND.t4 246.817
R197 VGND.n9 VGND.n8 223.569
R198 VGND.n17 VGND.n16 209.254
R199 VGND.n26 VGND.n25 199.739
R200 VGND.n40 VGND.n39 199.739
R201 VGND.n16 VGND.t0 100.001
R202 VGND.n25 VGND.t1 72.8576
R203 VGND.n16 VGND.t3 70.0005
R204 VGND.n25 VGND.t8 60.5809
R205 VGND.n8 VGND.t5 57.1434
R206 VGND.n39 VGND.t6 38.5719
R207 VGND.n39 VGND.t2 38.5719
R208 VGND.n11 VGND.n7 34.6358
R209 VGND.n15 VGND.n7 34.6358
R210 VGND.n19 VGND.n18 34.6358
R211 VGND.n19 VGND.n5 34.6358
R212 VGND.n23 VGND.n5 34.6358
R213 VGND.n24 VGND.n23 34.6358
R214 VGND.n27 VGND.n3 34.6358
R215 VGND.n31 VGND.n3 34.6358
R216 VGND.n32 VGND.n31 34.6358
R217 VGND.n33 VGND.n32 34.6358
R218 VGND.n33 VGND.n1 34.6358
R219 VGND.n38 VGND.n37 29.7417
R220 VGND.n11 VGND.n10 27.8593
R221 VGND.n8 VGND.t7 25.4291
R222 VGND.n40 VGND.n38 22.9652
R223 VGND.n17 VGND.n15 17.6946
R224 VGND.n37 VGND.n1 14.6829
R225 VGND.n10 VGND.n9 14.3133
R226 VGND.n38 VGND.n0 9.3005
R227 VGND.n37 VGND.n36 9.3005
R228 VGND.n35 VGND.n1 9.3005
R229 VGND.n34 VGND.n33 9.3005
R230 VGND.n32 VGND.n2 9.3005
R231 VGND.n31 VGND.n30 9.3005
R232 VGND.n29 VGND.n3 9.3005
R233 VGND.n28 VGND.n27 9.3005
R234 VGND.n12 VGND.n11 9.3005
R235 VGND.n13 VGND.n7 9.3005
R236 VGND.n15 VGND.n14 9.3005
R237 VGND.n18 VGND.n6 9.3005
R238 VGND.n20 VGND.n19 9.3005
R239 VGND.n21 VGND.n5 9.3005
R240 VGND.n23 VGND.n22 9.3005
R241 VGND.n24 VGND.n4 9.3005
R242 VGND.n27 VGND.n26 7.90638
R243 VGND.n41 VGND.n40 7.12063
R244 VGND.n18 VGND.n17 2.63579
R245 VGND.n26 VGND.n24 1.88285
R246 VGND.n12 VGND.n9 0.211448
R247 VGND.n41 VGND.n0 0.148519
R248 VGND.n13 VGND.n12 0.120292
R249 VGND.n14 VGND.n13 0.120292
R250 VGND.n14 VGND.n6 0.120292
R251 VGND.n20 VGND.n6 0.120292
R252 VGND.n21 VGND.n20 0.120292
R253 VGND.n22 VGND.n21 0.120292
R254 VGND.n22 VGND.n4 0.120292
R255 VGND.n28 VGND.n4 0.120292
R256 VGND.n29 VGND.n28 0.120292
R257 VGND.n30 VGND.n29 0.120292
R258 VGND.n30 VGND.n2 0.120292
R259 VGND.n34 VGND.n2 0.120292
R260 VGND.n35 VGND.n34 0.120292
R261 VGND.n36 VGND.n35 0.120292
R262 VGND.n36 VGND.n0 0.120292
R263 VGND VGND.n41 0.114842
R264 CLK.n0 CLK.t0 294.557
R265 CLK.n0 CLK.t1 211.01
R266 CLK.n1 CLK.n0 152
R267 CLK.n1 CLK 10.4234
R268 CLK CLK.n1 2.01193
R269 Q_N Q_N.t0 400.615
R270 Q_N Q_N.t1 237.101
R271 D.n0 D.t1 333.651
R272 D.n0 D.t0 297.233
R273 D D.n0 196.737
R274 a_448_47.n1 a_448_47.n0 926.024
R275 a_448_47.n1 a_448_47.t3 82.0838
R276 a_448_47.n0 a_448_47.t0 63.3338
R277 a_448_47.t1 a_448_47.n1 63.3219
R278 a_448_47.n0 a_448_47.t2 29.7268
R279 a_1270_413.t0 a_1270_413.t1 126.644
C0 VPB RESET_B 0.138482f
C1 CLK RESET_B 1.09e-19
C2 VPB VPWR 0.235545f
C3 CLK VPWR 0.017406f
C4 D RESET_B 4.72e-19
C5 VPB VGND 0.012976f
C6 CLK VGND 0.017208f
C7 D VPWR 0.081188f
C8 VPB Q 0.014966f
C9 VPB Q_N 0.011751f
C10 D VGND 0.051614f
C11 RESET_B VPWR 0.065186f
C12 RESET_B VGND 0.288101f
C13 VPWR VGND 0.081829f
C14 RESET_B Q 0.001485f
C15 VPWR Q 0.080299f
C16 RESET_B Q_N 2.89e-19
C17 VGND Q 0.091669f
C18 VPWR Q_N 0.085203f
C19 VPB CLK 0.069345f
C20 VGND Q_N 0.066103f
C21 VPB D 0.137565f
C22 Q_N VNB 0.087586f
C23 Q VNB 0.010712f
C24 VGND VNB 1.17272f
C25 VPWR VNB 0.959088f
C26 RESET_B VNB 0.260061f
C27 D VNB 0.159894f
C28 CLK VNB 0.195254f
C29 VPB VNB 2.1109f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_2 VGND VPWR VPB VNB CLK D RESET_B Q_N Q
X0 a_805_47.t0 a_761_289.t4 a_639_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47.t0 a_27_47.t2 a_1108_47.t0 VNB.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21.t2 a_1108_47.t4 a_1462_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 Q_N.t1 a_1659_47.t2 VGND.t11 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_651_413.t0 a_27_47.t3 a_543_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 a_1108_47.t3 a_193_47.t2 a_761_289.t3 VNB.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6 VGND.t4 RESET_B.t0 a_805_47.t1 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 VPWR.t8 a_1283_21.t3 Q.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.155 ps=1.31 w=1 l=0.15
X8 VPWR.t5 CLK.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_448_47.t2 D.t0 VPWR.t10 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR.t9 a_1283_21.t4 a_1659_47.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1522 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_761_289.t1 a_543_47.t4 VGND.t3 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 VGND.t9 a_1283_21.t5 a_1659_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_193_47.t1 a_27_47.t4 VGND.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47.t1 a_27_47.t5 a_761_289.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 VPWR.t12 a_1659_47.t3 Q_N.t3 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1462_47.t0 RESET_B.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X17 a_543_47.t1 a_27_47.t6 a_448_47.t0 VNB.t12 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X18 VGND.t10 a_1659_47.t4 Q_N.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_543_47.t3 a_193_47.t3 a_448_47.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X20 a_448_47.t1 D.t1 VGND.t5 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X21 VPWR.t6 a_1283_21.t6 a_1270_413.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 VPWR.t4 a_1108_47.t5 a_1283_21.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_1270_413.t1 a_193_47.t4 a_1108_47.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 a_193_47.t0 a_27_47.t7 VPWR.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1283_21.t0 RESET_B.t2 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X26 Q.t3 a_1283_21.t7 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10025 ps=0.985 w=0.65 l=0.15
X27 VPWR.t3 a_761_289.t5 a_651_413.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 VGND.t6 a_1283_21.t8 Q.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X29 Q_N.t2 a_1659_47.t5 VPWR.t11 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Q.t0 a_1283_21.t9 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1522 ps=1.335 w=1 l=0.15
X31 a_639_47.t0 a_193_47.t5 a_543_47.t2 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X32 VGND.t8 a_1283_21.t10 a_1217_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X33 a_651_413.t1 RESET_B.t3 VPWR.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X34 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_761_289.t2 a_543_47.t5 VPWR.t13 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
R0 a_761_289.n3 a_761_289.n2 647.119
R1 a_761_289.n1 a_761_289.t4 350.253
R2 a_761_289.n2 a_761_289.n0 260.339
R3 a_761_289.n2 a_761_289.n1 246.119
R4 a_761_289.n1 a_761_289.t5 189.588
R5 a_761_289.n3 a_761_289.t0 89.1195
R6 a_761_289.n0 a_761_289.t3 63.3338
R7 a_761_289.t2 a_761_289.n3 41.0422
R8 a_761_289.n0 a_761_289.t1 31.9797
R9 a_639_47.t1 a_639_47.t0 198.571
R10 a_805_47.t0 a_805_47.t1 60.0005
R11 VNB.t11 VNB.t17 3631.07
R12 VNB.t4 VNB.t7 2677.02
R13 VNB.t1 VNB.t5 2363.75
R14 VNB.t6 VNB.t3 2121.68
R15 VNB.t14 VNB.t13 1879.61
R16 VNB.t15 VNB.t10 1552.1
R17 VNB.t13 VNB.t15 1409.71
R18 VNB.t7 VNB.t8 1381.23
R19 VNB.t10 VNB.t6 1366.99
R20 VNB.t12 VNB.t1 1366.99
R21 VNB.t17 VNB.t12 1352.75
R22 VNB.t8 VNB.t9 1310.03
R23 VNB.t3 VNB.t4 1295.79
R24 VNB.t16 VNB.t2 1196.12
R25 VNB.t9 VNB.t16 1196.12
R26 VNB.t0 VNB.t11 1196.12
R27 VNB.t5 VNB.t14 1025.24
R28 VNB VNB.t0 925.567
R29 a_27_47.n1 a_27_47.t3 530.01
R30 a_27_47.t1 a_27_47.n5 421.021
R31 a_27_47.n0 a_27_47.t5 337.142
R32 a_27_47.n3 a_27_47.t0 280.223
R33 a_27_47.n4 a_27_47.t7 263.173
R34 a_27_47.n4 a_27_47.t4 227.826
R35 a_27_47.n0 a_27_47.t2 199.762
R36 a_27_47.n2 a_27_47.n1 170.81
R37 a_27_47.n2 a_27_47.n0 167.321
R38 a_27_47.n5 a_27_47.n4 152
R39 a_27_47.n1 a_27_47.t6 141.923
R40 a_27_47.n3 a_27_47.n2 10.8376
R41 a_27_47.n5 a_27_47.n3 2.50485
R42 a_1108_47.n3 a_1108_47.n2 636.953
R43 a_1108_47.n1 a_1108_47.t4 366.856
R44 a_1108_47.n2 a_1108_47.n0 300.2
R45 a_1108_47.n2 a_1108_47.n1 225.036
R46 a_1108_47.n1 a_1108_47.t5 174.056
R47 a_1108_47.n0 a_1108_47.t3 70.0005
R48 a_1108_47.t1 a_1108_47.n3 68.0124
R49 a_1108_47.n3 a_1108_47.t2 63.3219
R50 a_1108_47.n0 a_1108_47.t0 61.6672
R51 a_1217_47.t1 a_1217_47.t0 94.7268
R52 a_1462_47.t0 a_1462_47.t1 87.1434
R53 a_1283_21.n6 a_1283_21.n5 695.683
R54 a_1283_21.n3 a_1283_21.t6 389.183
R55 a_1283_21.n2 a_1283_21.t4 257.067
R56 a_1283_21.n4 a_1283_21.n3 254.367
R57 a_1283_21.n4 a_1283_21.t2 223.571
R58 a_1283_21.n0 a_1283_21.t3 212.081
R59 a_1283_21.n1 a_1283_21.t9 212.081
R60 a_1283_21.n5 a_1283_21.n2 189.82
R61 a_1283_21.n2 a_1283_21.t5 176.733
R62 a_1283_21.n3 a_1283_21.t10 174.891
R63 a_1283_21.n0 a_1283_21.t8 139.78
R64 a_1283_21.n1 a_1283_21.t7 139.78
R65 a_1283_21.n2 a_1283_21.n1 70.8399
R66 a_1283_21.n1 a_1283_21.n0 67.1884
R67 a_1283_21.n6 a_1283_21.t1 63.3219
R68 a_1283_21.t0 a_1283_21.n6 63.3219
R69 a_1283_21.n5 a_1283_21.n4 55.019
R70 a_1659_47.t0 a_1659_47.n2 385.462
R71 a_1659_47.n2 a_1659_47.t1 331.031
R72 a_1659_47.n2 a_1659_47.n1 263.92
R73 a_1659_47.n1 a_1659_47.t5 212.081
R74 a_1659_47.n0 a_1659_47.t3 212.081
R75 a_1659_47.n1 a_1659_47.t2 139.78
R76 a_1659_47.n0 a_1659_47.t4 139.78
R77 a_1659_47.n1 a_1659_47.n0 61.346
R78 VGND.n44 VGND.t5 307.536
R79 VGND.n12 VGND.n11 221.142
R80 VGND.n24 VGND.n23 209.254
R81 VGND.n16 VGND.n10 205.698
R82 VGND.n33 VGND.n32 199.739
R83 VGND.n47 VGND.n46 199.739
R84 VGND.n13 VGND.t10 167.999
R85 VGND.n23 VGND.t2 100.001
R86 VGND.n32 VGND.t4 72.8576
R87 VGND.n23 VGND.t8 70.0005
R88 VGND.n32 VGND.t3 60.5809
R89 VGND.n10 VGND.t9 57.1434
R90 VGND.n46 VGND.t1 38.5719
R91 VGND.n46 VGND.t0 38.5719
R92 VGND.n18 VGND.n17 34.6358
R93 VGND.n18 VGND.n7 34.6358
R94 VGND.n22 VGND.n7 34.6358
R95 VGND.n26 VGND.n25 34.6358
R96 VGND.n26 VGND.n5 34.6358
R97 VGND.n30 VGND.n5 34.6358
R98 VGND.n31 VGND.n30 34.6358
R99 VGND.n34 VGND.n3 34.6358
R100 VGND.n38 VGND.n3 34.6358
R101 VGND.n39 VGND.n38 34.6358
R102 VGND.n40 VGND.n39 34.6358
R103 VGND.n40 VGND.n1 34.6358
R104 VGND.n16 VGND.n9 33.1299
R105 VGND.n45 VGND.n44 29.7417
R106 VGND.n12 VGND.n9 26.7299
R107 VGND.n10 VGND.t7 25.4291
R108 VGND.n11 VGND.t11 24.9236
R109 VGND.n11 VGND.t6 24.9236
R110 VGND.n47 VGND.n45 22.9652
R111 VGND.n17 VGND.n16 18.4476
R112 VGND.n24 VGND.n22 17.6946
R113 VGND.n13 VGND.n12 14.8998
R114 VGND.n44 VGND.n1 14.6829
R115 VGND.n45 VGND.n0 9.3005
R116 VGND.n44 VGND.n43 9.3005
R117 VGND.n42 VGND.n1 9.3005
R118 VGND.n41 VGND.n40 9.3005
R119 VGND.n39 VGND.n2 9.3005
R120 VGND.n38 VGND.n37 9.3005
R121 VGND.n36 VGND.n3 9.3005
R122 VGND.n35 VGND.n34 9.3005
R123 VGND.n14 VGND.n9 9.3005
R124 VGND.n16 VGND.n15 9.3005
R125 VGND.n17 VGND.n8 9.3005
R126 VGND.n19 VGND.n18 9.3005
R127 VGND.n20 VGND.n7 9.3005
R128 VGND.n22 VGND.n21 9.3005
R129 VGND.n25 VGND.n6 9.3005
R130 VGND.n27 VGND.n26 9.3005
R131 VGND.n28 VGND.n5 9.3005
R132 VGND.n30 VGND.n29 9.3005
R133 VGND.n31 VGND.n4 9.3005
R134 VGND.n34 VGND.n33 7.90638
R135 VGND.n48 VGND.n47 7.12063
R136 VGND.n25 VGND.n24 2.63579
R137 VGND.n33 VGND.n31 1.88285
R138 VGND.n14 VGND.n13 0.756061
R139 VGND.n48 VGND.n0 0.148519
R140 VGND.n15 VGND.n14 0.120292
R141 VGND.n15 VGND.n8 0.120292
R142 VGND.n19 VGND.n8 0.120292
R143 VGND.n20 VGND.n19 0.120292
R144 VGND.n21 VGND.n20 0.120292
R145 VGND.n21 VGND.n6 0.120292
R146 VGND.n27 VGND.n6 0.120292
R147 VGND.n28 VGND.n27 0.120292
R148 VGND.n29 VGND.n28 0.120292
R149 VGND.n29 VGND.n4 0.120292
R150 VGND.n35 VGND.n4 0.120292
R151 VGND.n36 VGND.n35 0.120292
R152 VGND.n37 VGND.n36 0.120292
R153 VGND.n37 VGND.n2 0.120292
R154 VGND.n41 VGND.n2 0.120292
R155 VGND.n42 VGND.n41 0.120292
R156 VGND.n43 VGND.n42 0.120292
R157 VGND.n43 VGND.n0 0.120292
R158 VGND VGND.n48 0.114842
R159 Q_N Q_N.n0 236.111
R160 Q_N Q_N.n1 119.6
R161 Q_N.n0 Q_N.t3 26.5955
R162 Q_N.n0 Q_N.t2 26.5955
R163 Q_N.n1 Q_N.t0 24.9236
R164 Q_N.n1 Q_N.t1 24.9236
R165 a_543_47.n3 a_543_47.n2 674.338
R166 a_543_47.n1 a_543_47.t5 332.58
R167 a_543_47.n2 a_543_47.n0 284.012
R168 a_543_47.n2 a_543_47.n1 253.648
R169 a_543_47.n1 a_543_47.t4 168.701
R170 a_543_47.t0 a_543_47.n3 96.1553
R171 a_543_47.n3 a_543_47.t3 65.6672
R172 a_543_47.n0 a_543_47.t1 65.0005
R173 a_543_47.n0 a_543_47.t2 45.0005
R174 a_651_413.n0 a_651_413.t1 1327.82
R175 a_651_413.t0 a_651_413.n0 194.655
R176 a_651_413.n0 a_651_413.t2 63.3219
R177 VPB.t1 VPB.t14 790.188
R178 VPB.t5 VPB.t17 583.023
R179 VPB.t7 VPB.t12 577.104
R180 VPB.t3 VPB.t6 414.33
R181 VPB.t11 VPB.t0 319.627
R182 VPB.t17 VPB.t2 292.991
R183 VPB.t8 VPB.t3 292.991
R184 VPB.t12 VPB.t10 287.072
R185 VPB.t6 VPB.t5 287.072
R186 VPB.t10 VPB.t13 272.274
R187 VPB.t14 VPB.t8 272.274
R188 VPB.t2 VPB.t4 254.518
R189 VPB.t15 VPB.t16 248.599
R190 VPB.t13 VPB.t15 248.599
R191 VPB.t0 VPB.t7 248.599
R192 VPB.t4 VPB.t11 248.599
R193 VPB.t9 VPB.t1 248.599
R194 VPB VPB.t9 192.369
R195 a_193_47.t0 a_193_47.n3 370.026
R196 a_193_47.n0 a_193_47.t2 351.356
R197 a_193_47.n1 a_193_47.t5 334.717
R198 a_193_47.n3 a_193_47.t1 325.971
R199 a_193_47.n1 a_193_47.t3 309.935
R200 a_193_47.n0 a_193_47.t4 305.683
R201 a_193_47.n2 a_193_47.n0 16.879
R202 a_193_47.n3 a_193_47.n2 10.8867
R203 a_193_47.n2 a_193_47.n1 9.3005
R204 RESET_B.n1 RESET_B.t3 408.63
R205 RESET_B.n3 RESET_B.t2 347.577
R206 RESET_B.n3 RESET_B.t1 193.337
R207 RESET_B.n2 RESET_B.n1 167.575
R208 RESET_B.n4 RESET_B.n3 152
R209 RESET_B.n1 RESET_B.t0 132.282
R210 RESET_B RESET_B.n0 14.0185
R211 RESET_B.n4 RESET_B.n2 12.1952
R212 RESET_B.n2 RESET_B.n0 9.38606
R213 RESET_B RESET_B.n4 4.67077
R214 RESET_B.n0 RESET_B 4.53383
R215 Q Q.n0 605.824
R216 Q Q.n1 201.621
R217 Q.n0 Q.t1 34.4755
R218 Q.n1 Q.t2 32.3082
R219 Q.n0 Q.t0 26.5955
R220 Q.n1 Q.t3 24.9236
R221 VPWR.n30 VPWR.t13 806.511
R222 VPWR.n2 VPWR.t10 667.778
R223 VPWR.n10 VPWR.t4 667.111
R224 VPWR.n24 VPWR.n9 604.457
R225 VPWR.n46 VPWR.n1 604.394
R226 VPWR.n33 VPWR.n32 601.679
R227 VPWR.n18 VPWR.n12 601.188
R228 VPWR.n14 VPWR.n13 599.74
R229 VPWR.n15 VPWR.t12 278.88
R230 VPWR.n9 VPWR.t6 119.608
R231 VPWR.n32 VPWR.t3 93.81
R232 VPWR.n32 VPWR.t0 63.3219
R233 VPWR.n9 VPWR.t1 63.3219
R234 VPWR.n12 VPWR.t9 61.563
R235 VPWR.n1 VPWR.t2 41.5552
R236 VPWR.n1 VPWR.t5 41.5552
R237 VPWR.n45 VPWR.n44 34.6358
R238 VPWR.n38 VPWR.n4 34.6358
R239 VPWR.n39 VPWR.n38 34.6358
R240 VPWR.n40 VPWR.n39 34.6358
R241 VPWR.n34 VPWR.n31 34.6358
R242 VPWR.n25 VPWR.n7 34.6358
R243 VPWR.n29 VPWR.n7 34.6358
R244 VPWR.n19 VPWR.n10 34.2593
R245 VPWR.n40 VPWR.n2 32.377
R246 VPWR.n30 VPWR.n29 32.0005
R247 VPWR.n12 VPWR.t7 31.0125
R248 VPWR.n24 VPWR.n23 30.1181
R249 VPWR.n18 VPWR.n17 27.1064
R250 VPWR.n13 VPWR.t11 26.5955
R251 VPWR.n13 VPWR.t8 26.5955
R252 VPWR.n46 VPWR.n45 22.9652
R253 VPWR.n25 VPWR.n24 20.3299
R254 VPWR.n44 VPWR.n2 18.0711
R255 VPWR.n19 VPWR.n18 16.5652
R256 VPWR.n17 VPWR.n14 14.3064
R257 VPWR.n31 VPWR.n30 9.41227
R258 VPWR.n17 VPWR.n16 9.3005
R259 VPWR.n18 VPWR.n11 9.3005
R260 VPWR.n20 VPWR.n19 9.3005
R261 VPWR.n21 VPWR.n10 9.3005
R262 VPWR.n23 VPWR.n22 9.3005
R263 VPWR.n24 VPWR.n8 9.3005
R264 VPWR.n26 VPWR.n25 9.3005
R265 VPWR.n27 VPWR.n7 9.3005
R266 VPWR.n29 VPWR.n28 9.3005
R267 VPWR.n30 VPWR.n6 9.3005
R268 VPWR.n31 VPWR.n5 9.3005
R269 VPWR.n35 VPWR.n34 9.3005
R270 VPWR.n36 VPWR.n4 9.3005
R271 VPWR.n38 VPWR.n37 9.3005
R272 VPWR.n39 VPWR.n3 9.3005
R273 VPWR.n41 VPWR.n40 9.3005
R274 VPWR.n42 VPWR.n2 9.3005
R275 VPWR.n44 VPWR.n43 9.3005
R276 VPWR.n45 VPWR.n0 9.3005
R277 VPWR.n23 VPWR.n10 9.03579
R278 VPWR.n47 VPWR.n46 7.12063
R279 VPWR.n15 VPWR.n14 6.77321
R280 VPWR.n33 VPWR.n4 6.02403
R281 VPWR.n34 VPWR.n33 3.76521
R282 VPWR.n16 VPWR.n15 0.816842
R283 VPWR.n47 VPWR.n0 0.148519
R284 VPWR.n16 VPWR.n11 0.120292
R285 VPWR.n20 VPWR.n11 0.120292
R286 VPWR.n21 VPWR.n20 0.120292
R287 VPWR.n22 VPWR.n21 0.120292
R288 VPWR.n22 VPWR.n8 0.120292
R289 VPWR.n26 VPWR.n8 0.120292
R290 VPWR.n27 VPWR.n26 0.120292
R291 VPWR.n28 VPWR.n27 0.120292
R292 VPWR.n28 VPWR.n6 0.120292
R293 VPWR.n6 VPWR.n5 0.120292
R294 VPWR.n35 VPWR.n5 0.120292
R295 VPWR.n36 VPWR.n35 0.120292
R296 VPWR.n37 VPWR.n36 0.120292
R297 VPWR.n37 VPWR.n3 0.120292
R298 VPWR.n41 VPWR.n3 0.120292
R299 VPWR.n42 VPWR.n41 0.120292
R300 VPWR.n43 VPWR.n42 0.120292
R301 VPWR.n43 VPWR.n0 0.120292
R302 VPWR VPWR.n47 0.114842
R303 CLK.n0 CLK.t0 294.557
R304 CLK.n0 CLK.t1 211.01
R305 CLK.n1 CLK.n0 152
R306 CLK.n1 CLK 10.4234
R307 CLK CLK.n1 2.01193
R308 D.n0 D.t1 333.651
R309 D.n0 D.t0 297.233
R310 D D.n0 196.737
R311 a_448_47.n1 a_448_47.n0 926.024
R312 a_448_47.n0 a_448_47.t3 82.0838
R313 a_448_47.n1 a_448_47.t0 63.3338
R314 a_448_47.n0 a_448_47.t2 63.3219
R315 a_448_47.n2 a_448_47.t1 26.3935
R316 a_448_47.n3 a_448_47.n2 14.4005
R317 a_448_47.n2 a_448_47.n1 3.33383
R318 a_1270_413.t0 a_1270_413.t1 126.644
C0 Q Q_N 0.0061f
C1 CLK RESET_B 1.09e-19
C2 D RESET_B 4.72e-19
C3 CLK VPWR 0.017406f
C4 CLK VPB 0.069345f
C5 CLK VGND 0.017208f
C6 D VPWR 0.081188f
C7 D VPB 0.137565f
C8 RESET_B VPWR 0.065186f
C9 D VGND 0.051614f
C10 RESET_B VPB 0.138482f
C11 RESET_B VGND 0.28755f
C12 VPWR VPB 0.250676f
C13 RESET_B Q 8.5e-19
C14 VPWR VGND 0.096782f
C15 VGND VPB 0.013806f
C16 RESET_B Q_N 2.83e-19
C17 VPWR Q 0.014118f
C18 Q VPB 0.002023f
C19 VGND Q 0.114874f
C20 VPWR Q_N 0.157089f
C21 Q_N VPB 0.004225f
C22 VGND Q_N 0.142765f
C23 Q_N VNB 0.025191f
C24 Q VNB 0.003804f
C25 VGND VNB 1.24553f
C26 VPWR VNB 1.02447f
C27 RESET_B VNB 0.260034f
C28 D VNB 0.159894f
C29 CLK VNB 0.195254f
C30 VPB VNB 2.19949f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtn_1 VGND VPWR VPB VNB D RESET_B Q CLK_N
X0 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47.t0 a_193_47.t2 a_1108_47.t1 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21.t1 a_1108_47.t4 a_1462_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413.t0 a_193_47.t3 a_543_47.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47.t3 a_27_47.t2 a_761_289.t3 VNB.t3 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND.t0 RESET_B.t0 a_805_47.t1 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q.t1 a_1283_21.t3 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR.t9 CLK_N.t0 a_27_47.t1 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47.t3 D.t0 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289.t0 a_543_47.t4 VGND.t7 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47.t1 a_27_47.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47.t2 a_193_47.t4 a_761_289.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47.t1 RESET_B.t1 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47.t2 a_193_47.t5 a_448_47.t0 VNB.t13 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47.t0 a_27_47.t4 a_448_47.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47.t2 D.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR.t5 a_1283_21.t4 a_1270_413.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR.t0 a_1108_47.t5 a_1283_21.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413.t0 a_27_47.t5 a_1108_47.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47.t0 a_27_47.t6 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21.t2 RESET_B.t2 VPWR.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR.t7 a_761_289.t5 a_651_413.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q.t0 a_1283_21.t5 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47.t1 a_27_47.t7 a_543_47.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND.t5 a_1283_21.t6 a_1217_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413.t1 RESET_B.t3 VPWR.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND.t2 CLK_N.t1 a_27_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289.t1 a_543_47.t5 VPWR.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
R0 a_761_289.n3 a_761_289.n2 647.119
R1 a_761_289.n1 a_761_289.t4 350.253
R2 a_761_289.n2 a_761_289.n0 260.339
R3 a_761_289.n2 a_761_289.n1 246.119
R4 a_761_289.n1 a_761_289.t5 189.588
R5 a_761_289.n3 a_761_289.t2 89.1195
R6 a_761_289.n0 a_761_289.t3 63.3338
R7 a_761_289.t1 a_761_289.n3 41.0422
R8 a_761_289.n0 a_761_289.t0 31.9797
R9 a_639_47.t0 a_639_47.t1 198.571
R10 a_805_47.t0 a_805_47.t1 60.0005
R11 VNB.t4 VNB.t5 3631.07
R12 VNB.t9 VNB.t7 2961.81
R13 VNB.t11 VNB.t10 2363.75
R14 VNB.t8 VNB.t6 2121.68
R15 VNB.t12 VNB.t0 1879.61
R16 VNB.t3 VNB.t1 1552.1
R17 VNB.t0 VNB.t3 1409.71
R18 VNB.t1 VNB.t8 1366.99
R19 VNB.t13 VNB.t11 1366.99
R20 VNB.t5 VNB.t13 1352.75
R21 VNB.t6 VNB.t9 1295.79
R22 VNB.t2 VNB.t4 1196.12
R23 VNB.t10 VNB.t12 1025.24
R24 VNB VNB.t2 925.567
R25 a_193_47.n1 a_193_47.t3 530.01
R26 a_193_47.t0 a_193_47.n3 421.226
R27 a_193_47.n0 a_193_47.t4 337.142
R28 a_193_47.n3 a_193_47.t1 274.772
R29 a_193_47.n0 a_193_47.t2 199.762
R30 a_193_47.n2 a_193_47.n1 170.81
R31 a_193_47.n2 a_193_47.n0 167.321
R32 a_193_47.n1 a_193_47.t5 141.923
R33 a_193_47.n3 a_193_47.n2 10.476
R34 a_1108_47.n3 a_1108_47.n2 636.953
R35 a_1108_47.n1 a_1108_47.t4 366.856
R36 a_1108_47.n2 a_1108_47.n0 300.2
R37 a_1108_47.n2 a_1108_47.n1 225.036
R38 a_1108_47.n1 a_1108_47.t5 174.056
R39 a_1108_47.n0 a_1108_47.t3 70.0005
R40 a_1108_47.n3 a_1108_47.t2 68.0124
R41 a_1108_47.t0 a_1108_47.n3 63.3219
R42 a_1108_47.n0 a_1108_47.t1 61.6672
R43 a_1217_47.t1 a_1217_47.t0 94.7268
R44 a_1462_47.t0 a_1462_47.t1 87.1434
R45 a_1283_21.n4 a_1283_21.n3 807.871
R46 a_1283_21.n1 a_1283_21.t4 389.183
R47 a_1283_21.n2 a_1283_21.n1 251.167
R48 a_1283_21.n0 a_1283_21.t3 239.04
R49 a_1283_21.n2 a_1283_21.t1 223.571
R50 a_1283_21.n1 a_1283_21.t6 174.891
R51 a_1283_21.n0 a_1283_21.t5 166.739
R52 a_1283_21.n3 a_1283_21.n0 164.161
R53 a_1283_21.t0 a_1283_21.n4 63.3219
R54 a_1283_21.n4 a_1283_21.t2 63.3219
R55 a_1283_21.n3 a_1283_21.n2 37.7195
R56 a_543_47.n3 a_543_47.n2 674.338
R57 a_543_47.n1 a_543_47.t5 332.58
R58 a_543_47.n2 a_543_47.n0 284.012
R59 a_543_47.n2 a_543_47.n1 253.648
R60 a_543_47.n1 a_543_47.t4 168.701
R61 a_543_47.n3 a_543_47.t1 96.1553
R62 a_543_47.t0 a_543_47.n3 65.6672
R63 a_543_47.n0 a_543_47.t2 65.0005
R64 a_543_47.n0 a_543_47.t3 45.0005
R65 a_651_413.n0 a_651_413.t1 1327.82
R66 a_651_413.t0 a_651_413.n0 194.655
R67 a_651_413.n0 a_651_413.t2 63.3219
R68 VPB.t2 VPB.t11 790.188
R69 VPB.t3 VPB.t7 636.293
R70 VPB.t8 VPB.t9 583.023
R71 VPB.t5 VPB.t10 414.33
R72 VPB.t6 VPB.t13 319.627
R73 VPB.t9 VPB.t4 292.991
R74 VPB.t0 VPB.t5 292.991
R75 VPB.t10 VPB.t8 287.072
R76 VPB.t11 VPB.t0 272.274
R77 VPB.t4 VPB.t1 254.518
R78 VPB.t13 VPB.t3 248.599
R79 VPB.t1 VPB.t6 248.599
R80 VPB.t12 VPB.t2 248.599
R81 VPB VPB.t12 192.369
R82 a_27_47.t1 a_27_47.n5 385.682
R83 a_27_47.n2 a_27_47.t2 351.356
R84 a_27_47.n3 a_27_47.t7 334.717
R85 a_27_47.n3 a_27_47.t4 309.935
R86 a_27_47.n2 a_27_47.t5 305.683
R87 a_27_47.n1 a_27_47.t0 282.726
R88 a_27_47.n0 a_27_47.t6 263.173
R89 a_27_47.n0 a_27_47.t3 227.826
R90 a_27_47.n1 a_27_47.n0 152
R91 a_27_47.n5 a_27_47.n1 35.3396
R92 a_27_47.n4 a_27_47.n2 16.879
R93 a_27_47.n5 a_27_47.n4 11.2081
R94 a_27_47.n4 a_27_47.n3 9.3005
R95 RESET_B.n1 RESET_B.t3 408.63
R96 RESET_B.n3 RESET_B.t2 347.577
R97 RESET_B.n3 RESET_B.t1 193.337
R98 RESET_B.n2 RESET_B.n1 167.575
R99 RESET_B.n4 RESET_B.n3 152
R100 RESET_B.n1 RESET_B.t0 132.282
R101 RESET_B RESET_B.n0 14.0185
R102 RESET_B.n4 RESET_B.n2 12.1952
R103 RESET_B.n2 RESET_B.n0 9.38606
R104 RESET_B RESET_B.n4 4.67077
R105 RESET_B.n0 RESET_B 4.53383
R106 VGND.n29 VGND.t4 307.536
R107 VGND.n7 VGND.t6 232.974
R108 VGND.n9 VGND.n8 209.254
R109 VGND.n18 VGND.n17 199.739
R110 VGND.n32 VGND.n31 199.739
R111 VGND.n8 VGND.t1 100.001
R112 VGND.n17 VGND.t0 72.8576
R113 VGND.n8 VGND.t5 70.0005
R114 VGND.n17 VGND.t7 60.5809
R115 VGND.n31 VGND.t3 38.5719
R116 VGND.n31 VGND.t2 38.5719
R117 VGND.n11 VGND.n10 34.6358
R118 VGND.n11 VGND.n5 34.6358
R119 VGND.n15 VGND.n5 34.6358
R120 VGND.n16 VGND.n15 34.6358
R121 VGND.n19 VGND.n3 34.6358
R122 VGND.n23 VGND.n3 34.6358
R123 VGND.n24 VGND.n23 34.6358
R124 VGND.n25 VGND.n24 34.6358
R125 VGND.n25 VGND.n1 34.6358
R126 VGND.n30 VGND.n29 29.7417
R127 VGND.n9 VGND.n7 25.2423
R128 VGND.n32 VGND.n30 22.9652
R129 VGND.n29 VGND.n1 14.6829
R130 VGND.n30 VGND.n0 9.3005
R131 VGND.n29 VGND.n28 9.3005
R132 VGND.n27 VGND.n1 9.3005
R133 VGND.n26 VGND.n25 9.3005
R134 VGND.n24 VGND.n2 9.3005
R135 VGND.n23 VGND.n22 9.3005
R136 VGND.n21 VGND.n3 9.3005
R137 VGND.n20 VGND.n19 9.3005
R138 VGND.n10 VGND.n6 9.3005
R139 VGND.n12 VGND.n11 9.3005
R140 VGND.n13 VGND.n5 9.3005
R141 VGND.n15 VGND.n14 9.3005
R142 VGND.n16 VGND.n4 9.3005
R143 VGND.n19 VGND.n18 7.90638
R144 VGND.n33 VGND.n32 7.12063
R145 VGND.n10 VGND.n9 2.63579
R146 VGND.n18 VGND.n16 1.88285
R147 VGND.n7 VGND.n6 0.199654
R148 VGND.n33 VGND.n0 0.148519
R149 VGND.n12 VGND.n6 0.120292
R150 VGND.n13 VGND.n12 0.120292
R151 VGND.n14 VGND.n13 0.120292
R152 VGND.n14 VGND.n4 0.120292
R153 VGND.n20 VGND.n4 0.120292
R154 VGND.n21 VGND.n20 0.120292
R155 VGND.n22 VGND.n21 0.120292
R156 VGND.n22 VGND.n2 0.120292
R157 VGND.n26 VGND.n2 0.120292
R158 VGND.n27 VGND.n26 0.120292
R159 VGND.n28 VGND.n27 0.120292
R160 VGND.n28 VGND.n0 0.120292
R161 VGND VGND.n33 0.114842
R162 VPWR.n20 VPWR.t6 806.511
R163 VPWR.n2 VPWR.t8 667.778
R164 VPWR.n10 VPWR.t0 667.751
R165 VPWR.n14 VPWR.n9 604.457
R166 VPWR.n36 VPWR.n1 604.394
R167 VPWR.n23 VPWR.n22 601.679
R168 VPWR.n11 VPWR.t4 347.94
R169 VPWR.n9 VPWR.t5 119.608
R170 VPWR.n22 VPWR.t7 93.81
R171 VPWR.n22 VPWR.t2 63.3219
R172 VPWR.n9 VPWR.t1 63.3219
R173 VPWR.n1 VPWR.t3 41.5552
R174 VPWR.n1 VPWR.t9 41.5552
R175 VPWR.n35 VPWR.n34 34.6358
R176 VPWR.n28 VPWR.n4 34.6358
R177 VPWR.n29 VPWR.n28 34.6358
R178 VPWR.n30 VPWR.n29 34.6358
R179 VPWR.n24 VPWR.n21 34.6358
R180 VPWR.n15 VPWR.n7 34.6358
R181 VPWR.n19 VPWR.n7 34.6358
R182 VPWR.n30 VPWR.n2 32.377
R183 VPWR.n20 VPWR.n19 32.0005
R184 VPWR.n14 VPWR.n13 30.1181
R185 VPWR.n36 VPWR.n35 22.9652
R186 VPWR.n15 VPWR.n14 20.3299
R187 VPWR.n34 VPWR.n2 18.0711
R188 VPWR.n21 VPWR.n20 9.41227
R189 VPWR.n13 VPWR.n12 9.3005
R190 VPWR.n14 VPWR.n8 9.3005
R191 VPWR.n16 VPWR.n15 9.3005
R192 VPWR.n17 VPWR.n7 9.3005
R193 VPWR.n19 VPWR.n18 9.3005
R194 VPWR.n20 VPWR.n6 9.3005
R195 VPWR.n21 VPWR.n5 9.3005
R196 VPWR.n25 VPWR.n24 9.3005
R197 VPWR.n26 VPWR.n4 9.3005
R198 VPWR.n28 VPWR.n27 9.3005
R199 VPWR.n29 VPWR.n3 9.3005
R200 VPWR.n31 VPWR.n30 9.3005
R201 VPWR.n32 VPWR.n2 9.3005
R202 VPWR.n34 VPWR.n33 9.3005
R203 VPWR.n35 VPWR.n0 9.3005
R204 VPWR.n13 VPWR.n10 9.03579
R205 VPWR.n37 VPWR.n36 7.12063
R206 VPWR.n11 VPWR.n10 6.33361
R207 VPWR.n23 VPWR.n4 6.02403
R208 VPWR.n24 VPWR.n23 3.76521
R209 VPWR.n12 VPWR.n11 1.75271
R210 VPWR.n37 VPWR.n0 0.148519
R211 VPWR.n12 VPWR.n8 0.120292
R212 VPWR.n16 VPWR.n8 0.120292
R213 VPWR.n17 VPWR.n16 0.120292
R214 VPWR.n18 VPWR.n17 0.120292
R215 VPWR.n18 VPWR.n6 0.120292
R216 VPWR.n6 VPWR.n5 0.120292
R217 VPWR.n25 VPWR.n5 0.120292
R218 VPWR.n26 VPWR.n25 0.120292
R219 VPWR.n27 VPWR.n26 0.120292
R220 VPWR.n27 VPWR.n3 0.120292
R221 VPWR.n31 VPWR.n3 0.120292
R222 VPWR.n32 VPWR.n31 0.120292
R223 VPWR.n33 VPWR.n32 0.120292
R224 VPWR.n33 VPWR.n0 0.120292
R225 VPWR VPWR.n37 0.114842
R226 Q.n1 Q.t1 353.543
R227 Q.n0 Q.t0 209.923
R228 Q Q.n0 47.9019
R229 Q.n0 Q 10.2907
R230 Q.n1 Q 9.28219
R231 Q Q.n1 7.62424
R232 CLK_N.n0 CLK_N.t0 294.557
R233 CLK_N.n0 CLK_N.t1 211.01
R234 CLK_N CLK_N.n0 153.871
R235 D.n0 D.t1 333.651
R236 D.n0 D.t0 297.233
R237 D D.n0 196.737
R238 a_448_47.n1 a_448_47.n0 926.024
R239 a_448_47.t1 a_448_47.n1 82.0838
R240 a_448_47.n0 a_448_47.t0 63.3338
R241 a_448_47.n1 a_448_47.t3 63.3219
R242 a_448_47.n0 a_448_47.t2 29.7268
R243 a_1270_413.t0 a_1270_413.t1 126.644
C0 VPB VGND 0.010245f
C1 D RESET_B 4.72e-19
C2 CLK_N VPWR 0.017406f
C3 VPB Q 0.011004f
C4 D VPWR 0.081188f
C5 CLK_N VGND 0.017208f
C6 D VGND 0.051614f
C7 RESET_B VPWR 0.065186f
C8 RESET_B VGND 0.287765f
C9 VPWR VGND 0.051201f
C10 RESET_B Q 9.12e-19
C11 VPWR Q 0.099692f
C12 VGND Q 0.061585f
C13 VPB CLK_N 0.069345f
C14 VPB D 0.137565f
C15 VPB RESET_B 0.138482f
C16 VPB VPWR 0.216382f
C17 CLK_N RESET_B 1.09e-19
C18 Q VNB 0.089869f
C19 VGND VNB 1.02176f
C20 VPWR VNB 0.831431f
C21 RESET_B VNB 0.263863f
C22 D VNB 0.159894f
C23 CLK_N VNB 0.195254f
C24 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_805_47.t1 a_761_289.t4 a_639_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47.t0 a_27_47.t2 a_1108_47.t1 VNB.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21.t2 a_1108_47.t4 a_1462_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413.t0 a_27_47.t3 a_543_47.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47.t2 a_193_47.t2 a_761_289.t0 VNB.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND.t6 RESET_B.t0 a_805_47.t0 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q.t1 a_1283_21.t3 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR.t7 CLK.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47.t3 D.t0 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289.t2 a_543_47.t4 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47.t1 a_27_47.t4 VGND.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47.t0 a_27_47.t5 a_761_289.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47.t1 RESET_B.t1 VGND.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47.t1 a_27_47.t6 a_448_47.t0 VNB.t7 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47.t2 a_193_47.t3 a_448_47.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47.t2 D.t1 VGND.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR.t2 a_1283_21.t4 a_1270_413.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR.t3 a_1108_47.t5 a_1283_21.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413.t1 a_193_47.t4 a_1108_47.t3 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47.t0 a_27_47.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21.t0 RESET_B.t2 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR.t9 a_761_289.t5 a_651_413.t2 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q.t0 a_1283_21.t5 VGND.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47.t0 a_193_47.t5 a_543_47.t3 VNB.t11 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND.t2 a_1283_21.t6 a_1217_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413.t1 RESET_B.t3 VPWR.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND.t4 CLK.t1 a_27_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289.t3 a_543_47.t5 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
R0 a_761_289.n3 a_761_289.n2 647.119
R1 a_761_289.n1 a_761_289.t4 350.253
R2 a_761_289.n2 a_761_289.n0 260.339
R3 a_761_289.n2 a_761_289.n1 246.119
R4 a_761_289.n1 a_761_289.t5 189.588
R5 a_761_289.n3 a_761_289.t1 89.1195
R6 a_761_289.n0 a_761_289.t0 63.3338
R7 a_761_289.t3 a_761_289.n3 41.0422
R8 a_761_289.n0 a_761_289.t2 31.9797
R9 a_639_47.t1 a_639_47.t0 198.571
R10 a_805_47.t0 a_805_47.t1 60.0005
R11 VNB.t6 VNB.t0 3631.07
R12 VNB.t4 VNB.t2 2961.81
R13 VNB.t11 VNB.t13 2363.75
R14 VNB.t3 VNB.t12 2121.68
R15 VNB.t9 VNB.t10 1879.61
R16 VNB.t1 VNB.t5 1552.1
R17 VNB.t10 VNB.t1 1409.71
R18 VNB.t5 VNB.t3 1366.99
R19 VNB.t7 VNB.t11 1366.99
R20 VNB.t0 VNB.t7 1352.75
R21 VNB.t12 VNB.t4 1295.79
R22 VNB.t8 VNB.t6 1196.12
R23 VNB.t13 VNB.t9 1025.24
R24 VNB VNB.t8 925.567
R25 a_27_47.n1 a_27_47.t3 530.01
R26 a_27_47.t1 a_27_47.n5 421.021
R27 a_27_47.n0 a_27_47.t5 337.142
R28 a_27_47.n3 a_27_47.t0 280.223
R29 a_27_47.n4 a_27_47.t7 263.173
R30 a_27_47.n4 a_27_47.t4 227.826
R31 a_27_47.n0 a_27_47.t2 199.762
R32 a_27_47.n2 a_27_47.n1 170.81
R33 a_27_47.n2 a_27_47.n0 167.321
R34 a_27_47.n5 a_27_47.n4 152
R35 a_27_47.n1 a_27_47.t6 141.923
R36 a_27_47.n3 a_27_47.n2 10.8376
R37 a_27_47.n5 a_27_47.n3 2.50485
R38 a_1108_47.n3 a_1108_47.n2 636.953
R39 a_1108_47.n1 a_1108_47.t4 366.856
R40 a_1108_47.n2 a_1108_47.n0 300.2
R41 a_1108_47.n2 a_1108_47.n1 225.036
R42 a_1108_47.n1 a_1108_47.t5 174.056
R43 a_1108_47.n0 a_1108_47.t2 70.0005
R44 a_1108_47.t0 a_1108_47.n3 68.0124
R45 a_1108_47.n3 a_1108_47.t3 63.3219
R46 a_1108_47.n0 a_1108_47.t1 61.6672
R47 a_1217_47.t1 a_1217_47.t0 94.7268
R48 a_1462_47.t0 a_1462_47.t1 87.1434
R49 a_1283_21.n4 a_1283_21.n3 807.871
R50 a_1283_21.n1 a_1283_21.t4 389.183
R51 a_1283_21.n2 a_1283_21.n1 251.167
R52 a_1283_21.n0 a_1283_21.t3 239.04
R53 a_1283_21.n2 a_1283_21.t2 223.571
R54 a_1283_21.n1 a_1283_21.t6 174.891
R55 a_1283_21.n0 a_1283_21.t5 166.739
R56 a_1283_21.n3 a_1283_21.n0 164.161
R57 a_1283_21.n4 a_1283_21.t1 63.3219
R58 a_1283_21.t0 a_1283_21.n4 63.3219
R59 a_1283_21.n3 a_1283_21.n2 37.7195
R60 a_543_47.n3 a_543_47.n2 674.338
R61 a_543_47.n1 a_543_47.t5 332.58
R62 a_543_47.n2 a_543_47.n0 284.012
R63 a_543_47.n2 a_543_47.n1 253.648
R64 a_543_47.n1 a_543_47.t4 168.701
R65 a_543_47.t0 a_543_47.n3 96.1553
R66 a_543_47.n3 a_543_47.t2 65.6672
R67 a_543_47.n0 a_543_47.t1 65.0005
R68 a_543_47.n0 a_543_47.t3 45.0005
R69 a_651_413.n0 a_651_413.t1 1327.82
R70 a_651_413.t0 a_651_413.n0 194.655
R71 a_651_413.n0 a_651_413.t2 63.3219
R72 VPB.t0 VPB.t10 790.188
R73 VPB.t7 VPB.t5 636.293
R74 VPB.t3 VPB.t12 583.023
R75 VPB.t2 VPB.t13 414.33
R76 VPB.t4 VPB.t6 319.627
R77 VPB.t12 VPB.t1 292.991
R78 VPB.t8 VPB.t2 292.991
R79 VPB.t13 VPB.t3 287.072
R80 VPB.t10 VPB.t8 272.274
R81 VPB.t1 VPB.t9 254.518
R82 VPB.t6 VPB.t7 248.599
R83 VPB.t9 VPB.t4 248.599
R84 VPB.t11 VPB.t0 248.599
R85 VPB VPB.t11 192.369
R86 a_193_47.t0 a_193_47.n3 370.026
R87 a_193_47.n0 a_193_47.t2 351.356
R88 a_193_47.n1 a_193_47.t5 334.717
R89 a_193_47.n3 a_193_47.t1 325.971
R90 a_193_47.n1 a_193_47.t3 309.935
R91 a_193_47.n0 a_193_47.t4 305.683
R92 a_193_47.n2 a_193_47.n0 16.879
R93 a_193_47.n3 a_193_47.n2 10.8867
R94 a_193_47.n2 a_193_47.n1 9.3005
R95 RESET_B.n1 RESET_B.t3 408.63
R96 RESET_B.n3 RESET_B.t2 347.577
R97 RESET_B.n3 RESET_B.t1 193.337
R98 RESET_B.n2 RESET_B.n1 167.575
R99 RESET_B.n4 RESET_B.n3 152
R100 RESET_B.n1 RESET_B.t0 132.282
R101 RESET_B RESET_B.n0 14.0185
R102 RESET_B.n4 RESET_B.n2 12.1952
R103 RESET_B.n2 RESET_B.n0 9.38606
R104 RESET_B RESET_B.n4 4.67077
R105 RESET_B.n0 RESET_B 4.53383
R106 VGND.n29 VGND.t1 307.536
R107 VGND.n7 VGND.t3 232.974
R108 VGND.n9 VGND.n8 209.254
R109 VGND.n18 VGND.n17 199.739
R110 VGND.n32 VGND.n31 199.739
R111 VGND.n8 VGND.t5 100.001
R112 VGND.n17 VGND.t6 72.8576
R113 VGND.n8 VGND.t2 70.0005
R114 VGND.n17 VGND.t7 60.5809
R115 VGND.n31 VGND.t0 38.5719
R116 VGND.n31 VGND.t4 38.5719
R117 VGND.n11 VGND.n10 34.6358
R118 VGND.n11 VGND.n5 34.6358
R119 VGND.n15 VGND.n5 34.6358
R120 VGND.n16 VGND.n15 34.6358
R121 VGND.n19 VGND.n3 34.6358
R122 VGND.n23 VGND.n3 34.6358
R123 VGND.n24 VGND.n23 34.6358
R124 VGND.n25 VGND.n24 34.6358
R125 VGND.n25 VGND.n1 34.6358
R126 VGND.n30 VGND.n29 29.7417
R127 VGND.n9 VGND.n7 25.2423
R128 VGND.n32 VGND.n30 22.9652
R129 VGND.n29 VGND.n1 14.6829
R130 VGND.n30 VGND.n0 9.3005
R131 VGND.n29 VGND.n28 9.3005
R132 VGND.n27 VGND.n1 9.3005
R133 VGND.n26 VGND.n25 9.3005
R134 VGND.n24 VGND.n2 9.3005
R135 VGND.n23 VGND.n22 9.3005
R136 VGND.n21 VGND.n3 9.3005
R137 VGND.n20 VGND.n19 9.3005
R138 VGND.n10 VGND.n6 9.3005
R139 VGND.n12 VGND.n11 9.3005
R140 VGND.n13 VGND.n5 9.3005
R141 VGND.n15 VGND.n14 9.3005
R142 VGND.n16 VGND.n4 9.3005
R143 VGND.n19 VGND.n18 7.90638
R144 VGND.n33 VGND.n32 7.12063
R145 VGND.n10 VGND.n9 2.63579
R146 VGND.n18 VGND.n16 1.88285
R147 VGND.n7 VGND.n6 0.199654
R148 VGND.n33 VGND.n0 0.148519
R149 VGND.n12 VGND.n6 0.120292
R150 VGND.n13 VGND.n12 0.120292
R151 VGND.n14 VGND.n13 0.120292
R152 VGND.n14 VGND.n4 0.120292
R153 VGND.n20 VGND.n4 0.120292
R154 VGND.n21 VGND.n20 0.120292
R155 VGND.n22 VGND.n21 0.120292
R156 VGND.n22 VGND.n2 0.120292
R157 VGND.n26 VGND.n2 0.120292
R158 VGND.n27 VGND.n26 0.120292
R159 VGND.n28 VGND.n27 0.120292
R160 VGND.n28 VGND.n0 0.120292
R161 VGND VGND.n33 0.114842
R162 VPWR.n20 VPWR.t8 806.511
R163 VPWR.n2 VPWR.t6 667.778
R164 VPWR.n10 VPWR.t3 667.751
R165 VPWR.n14 VPWR.n9 604.457
R166 VPWR.n36 VPWR.n1 604.394
R167 VPWR.n23 VPWR.n22 601.679
R168 VPWR.n11 VPWR.t1 347.94
R169 VPWR.n9 VPWR.t2 119.608
R170 VPWR.n22 VPWR.t9 93.81
R171 VPWR.n22 VPWR.t5 63.3219
R172 VPWR.n9 VPWR.t4 63.3219
R173 VPWR.n1 VPWR.t0 41.5552
R174 VPWR.n1 VPWR.t7 41.5552
R175 VPWR.n35 VPWR.n34 34.6358
R176 VPWR.n28 VPWR.n4 34.6358
R177 VPWR.n29 VPWR.n28 34.6358
R178 VPWR.n30 VPWR.n29 34.6358
R179 VPWR.n24 VPWR.n21 34.6358
R180 VPWR.n15 VPWR.n7 34.6358
R181 VPWR.n19 VPWR.n7 34.6358
R182 VPWR.n30 VPWR.n2 32.377
R183 VPWR.n20 VPWR.n19 32.0005
R184 VPWR.n14 VPWR.n13 30.1181
R185 VPWR.n36 VPWR.n35 22.9652
R186 VPWR.n15 VPWR.n14 20.3299
R187 VPWR.n34 VPWR.n2 18.0711
R188 VPWR.n21 VPWR.n20 9.41227
R189 VPWR.n13 VPWR.n12 9.3005
R190 VPWR.n14 VPWR.n8 9.3005
R191 VPWR.n16 VPWR.n15 9.3005
R192 VPWR.n17 VPWR.n7 9.3005
R193 VPWR.n19 VPWR.n18 9.3005
R194 VPWR.n20 VPWR.n6 9.3005
R195 VPWR.n21 VPWR.n5 9.3005
R196 VPWR.n25 VPWR.n24 9.3005
R197 VPWR.n26 VPWR.n4 9.3005
R198 VPWR.n28 VPWR.n27 9.3005
R199 VPWR.n29 VPWR.n3 9.3005
R200 VPWR.n31 VPWR.n30 9.3005
R201 VPWR.n32 VPWR.n2 9.3005
R202 VPWR.n34 VPWR.n33 9.3005
R203 VPWR.n35 VPWR.n0 9.3005
R204 VPWR.n13 VPWR.n10 9.03579
R205 VPWR.n37 VPWR.n36 7.12063
R206 VPWR.n11 VPWR.n10 6.33361
R207 VPWR.n23 VPWR.n4 6.02403
R208 VPWR.n24 VPWR.n23 3.76521
R209 VPWR.n12 VPWR.n11 1.75271
R210 VPWR.n37 VPWR.n0 0.148519
R211 VPWR.n12 VPWR.n8 0.120292
R212 VPWR.n16 VPWR.n8 0.120292
R213 VPWR.n17 VPWR.n16 0.120292
R214 VPWR.n18 VPWR.n17 0.120292
R215 VPWR.n18 VPWR.n6 0.120292
R216 VPWR.n6 VPWR.n5 0.120292
R217 VPWR.n25 VPWR.n5 0.120292
R218 VPWR.n26 VPWR.n25 0.120292
R219 VPWR.n27 VPWR.n26 0.120292
R220 VPWR.n27 VPWR.n3 0.120292
R221 VPWR.n31 VPWR.n3 0.120292
R222 VPWR.n32 VPWR.n31 0.120292
R223 VPWR.n33 VPWR.n32 0.120292
R224 VPWR.n33 VPWR.n0 0.120292
R225 VPWR VPWR.n37 0.114842
R226 Q.n1 Q.t1 353.543
R227 Q.n0 Q.t0 209.923
R228 Q Q.n0 47.9019
R229 Q.n0 Q 10.2907
R230 Q.n1 Q 9.28219
R231 Q Q.n1 7.62424
R232 CLK.n0 CLK.t0 294.557
R233 CLK.n0 CLK.t1 211.01
R234 CLK.n1 CLK.n0 152
R235 CLK.n1 CLK 10.4234
R236 CLK CLK.n1 2.01193
R237 D.n0 D.t1 333.651
R238 D.n0 D.t0 297.233
R239 D D.n0 196.737
R240 a_448_47.n1 a_448_47.n0 926.024
R241 a_448_47.t1 a_448_47.n1 82.0838
R242 a_448_47.n0 a_448_47.t0 63.3338
R243 a_448_47.n1 a_448_47.t3 63.3219
R244 a_448_47.n0 a_448_47.t2 29.7268
R245 a_1270_413.t0 a_1270_413.t1 126.644
C0 VPB CLK 0.069345f
C1 VPB D 0.137565f
C2 VPB RESET_B 0.138482f
C3 CLK RESET_B 1.09e-19
C4 VPB VPWR 0.21644f
C5 CLK VPWR 0.017406f
C6 D RESET_B 4.72e-19
C7 VPB VGND 0.009994f
C8 CLK VGND 0.017208f
C9 D VPWR 0.081188f
C10 VPB Q 0.011004f
C11 RESET_B VPWR 0.065186f
C12 D VGND 0.051614f
C13 RESET_B VGND 0.287765f
C14 RESET_B Q 9.12e-19
C15 VPWR VGND 0.050202f
C16 VPWR Q 0.099692f
C17 VGND Q 0.061585f
C18 Q VNB 0.089869f
C19 VGND VNB 1.02171f
C20 VPWR VNB 0.830843f
C21 RESET_B VNB 0.263863f
C22 D VNB 0.159894f
C23 CLK VNB 0.195254f
C24 VPB VNB 1.84511f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32oi_1 VGND VPWR VPB VNB B2 Y B1 A1 A2 A3
X0 VPWR.t1 A3.t0 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND.t0 A3.t1 a_383_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 a_309_47.t0 A1.t0 Y.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0715 pd=0.87 as=0.15275 ps=1.12 w=0.65 l=0.15
X3 Y.t1 B1.t0 a_109_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.15275 pd=1.12 as=0.07475 ps=0.88 w=0.65 l=0.15
X4 a_27_297.t3 B1.t1 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X5 a_383_47.t1 A2.t0 a_309_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.0715 ps=0.87 w=0.65 l=0.15
X6 a_27_297.t0 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t3 B2.t0 a_27_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR.t2 A1.t1 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X9 a_109_47.t0 B2.t1 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A3.n0 A3.t0 212.154
R1 A3 A3.n0 153.696
R2 A3.n0 A3.t1 150.442
R3 a_27_297.n1 a_27_297.t4 383.798
R4 a_27_297.n2 a_27_297.n1 366.505
R5 a_27_297.n1 a_27_297.n0 287.099
R6 a_27_297.n0 a_27_297.t3 58.1155
R7 a_27_297.n2 a_27_297.t1 28.5655
R8 a_27_297.n0 a_27_297.t2 26.5955
R9 a_27_297.t0 a_27_297.n2 26.5955
R10 VPWR.n1 VPWR.n0 611.934
R11 VPWR.n1 VPWR.t1 248.401
R12 VPWR.n0 VPWR.t0 26.5955
R13 VPWR.n0 VPWR.t2 26.5955
R14 VPWR VPWR.n1 0.772078
R15 VPB.t3 VPB.t2 343.303
R16 VPB.t0 VPB.t1 254.518
R17 VPB.t2 VPB.t0 248.599
R18 VPB.t4 VPB.t3 248.599
R19 VPB VPB.t4 192.369
R20 a_383_47.t0 a_383_47.t1 60.9236
R21 VGND.n0 VGND.t1 289.74
R22 VGND.n0 VGND.t0 155.505
R23 VGND VGND.n0 0.0626155
R24 VNB.t0 VNB.t2 1765.7
R25 VNB.t3 VNB.t1 1366.99
R26 VNB.t4 VNB.t0 1082.2
R27 VNB.t2 VNB.t3 1053.72
R28 VNB VNB.t4 925.567
R29 A1.n0 A1.t1 241.536
R30 A1 A1.n0 193.118
R31 A1.n0 A1.t0 169.237
R32 Y Y.n1 592.864
R33 Y Y.n0 292.235
R34 Y.n0 Y.t0 58.1543
R35 Y.n0 Y.t1 28.6159
R36 Y.n1 Y.t2 26.5955
R37 Y.n1 Y.t3 26.5955
R38 a_309_47.t0 a_309_47.t1 40.6159
R39 B1.n0 B1.t1 236.934
R40 B1 B1.n0 181.048
R41 B1.n0 B1.t0 164.633
R42 a_109_47.t0 a_109_47.t1 42.462
R43 A2.n0 A2.t1 229.397
R44 A2.n0 A2.t0 164.238
R45 A2 A2.n0 155.685
R46 B2.n0 B2.t0 230.155
R47 B2.n0 B2.t1 157.856
R48 B2 B2.n0 155.685
C0 A3 Y 1.48e-19
C1 A2 VPWR 0.020141f
C2 A1 VGND 0.045743f
C3 VPB B2 0.037919f
C4 A2 VGND 0.067977f
C5 A3 VPWR 0.062246f
C6 VPB B1 0.03429f
C7 Y VPWR 0.012009f
C8 A3 VGND 0.054328f
C9 VPB A1 0.027724f
C10 B2 B1 0.059024f
C11 Y VGND 0.067741f
C12 VPB A2 0.026128f
C13 VPWR VGND 0.069526f
C14 VPB A3 0.043195f
C15 B1 A1 0.068965f
C16 B1 A2 0.003228f
C17 VPB Y 0.005864f
C18 B1 A3 6.02e-19
C19 VPB VPWR 0.090295f
C20 A1 A2 0.120956f
C21 B2 Y 0.048092f
C22 B2 VPWR 0.009218f
C23 VPB VGND 0.011889f
C24 A1 A3 2.13e-19
C25 B1 Y 0.100505f
C26 B1 VPWR 0.013386f
C27 A2 A3 0.089769f
C28 B2 VGND 0.032751f
C29 A1 Y 0.043443f
C30 B1 VGND 0.015595f
C31 A1 VPWR 0.018172f
C32 A2 Y 4.37e-19
C33 VGND VNB 0.441169f
C34 VPWR VNB 0.358296f
C35 Y VNB 0.040011f
C36 A3 VNB 0.145342f
C37 A2 VNB 0.097828f
C38 A1 VNB 0.094057f
C39 B1 VNB 0.097928f
C40 B2 VNB 0.14504f
C41 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32oi_2 VNB VPB VGND VPWR B2 B1 Y A1 A2 A3
X0 Y.t7 A1.t0 a_478_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_27_297.t6 A1.t1 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.3775 ps=1.755 w=1 l=0.15
X2 a_27_297.t1 A2.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.305 ps=1.61 w=1 l=0.15
X3 a_27_297.t7 A3.t0 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.335 ps=1.67 w=1 l=0.15
X4 VPWR.t4 A3.t1 a_27_297.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.1375 ps=1.275 w=1 l=0.15
X5 VPWR.t1 A1.t2 a_27_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.3775 pd=1.755 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297.t2 B1.t0 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_478_47.t0 A1.t3 Y.t6 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_478_47.t2 A2.t1 a_730_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t3 A3.t2 a_730_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12025 ps=1.02 w=0.65 l=0.15
X10 Y.t4 B1.t1 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297.t0 B2.t0 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_47.t3 B2.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_47.t1 B1.t2 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y.t1 B1.t3 a_27_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_730_47.t2 A3.t3 VGND.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.20475 ps=1.93 w=0.65 l=0.15
X16 Y.t5 B2.t2 a_27_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VPWR.t5 A2.t2 a_27_297.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND.t1 B2.t3 a_27_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_730_47.t0 A2.t3 a_478_47.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
R0 A1.n2 A1.t2 322.584
R1 A1.n0 A1.t1 221.72
R2 A1.n0 A1.t3 165.488
R3 A1 A1.n0 155.375
R4 A1.n3 A1.n2 152
R5 A1.n1 A1.t0 149.421
R6 A1.n1 A1.n0 58.9116
R7 A1.n3 A1 6.16777
R8 A1 A1.n3 4.53868
R9 A1.n2 A1.n1 1.78569
R10 a_478_47.n0 a_478_47.t1 332.077
R11 a_478_47.n0 a_478_47.t2 331.325
R12 a_478_47.n1 a_478_47.n0 185
R13 a_478_47.t0 a_478_47.n1 26.7697
R14 a_478_47.n1 a_478_47.t3 24.9236
R15 Y.n2 Y.n0 610.225
R16 Y.n2 Y.n1 366.913
R17 Y.n5 Y.n4 241.847
R18 Y.n5 Y.n3 218.506
R19 Y Y.n2 39.1622
R20 Y.n0 Y.t3 26.5955
R21 Y.n0 Y.t4 26.5955
R22 Y.n1 Y.t2 26.5955
R23 Y.n1 Y.t5 26.5955
R24 Y.n4 Y.t6 24.9236
R25 Y.n4 Y.t7 24.9236
R26 Y.n3 Y.t0 24.9236
R27 Y.n3 Y.t1 24.9236
R28 Y Y.n5 1.48887
R29 VNB.t6 VNB.t8 2833.66
R30 VNB.t0 VNB.t4 2833.66
R31 VNB.t8 VNB.t7 1480.91
R32 VNB.t3 VNB.t9 1224.6
R33 VNB.t9 VNB.t6 1196.12
R34 VNB.t4 VNB.t3 1196.12
R35 VNB.t1 VNB.t0 1196.12
R36 VNB.t2 VNB.t1 1196.12
R37 VNB.t5 VNB.t2 1196.12
R38 VNB VNB.t5 911.327
R39 VPWR.n21 VPWR.n20 585
R40 VPWR.n19 VPWR.n0 585
R41 VPWR.n11 VPWR.n2 585
R42 VPWR.n13 VPWR.n12 585
R43 VPWR.n5 VPWR.n4 585
R44 VPWR.n7 VPWR.n6 585
R45 VPWR.n6 VPWR.n5 66.9805
R46 VPWR.n12 VPWR.n11 66.9805
R47 VPWR.n20 VPWR.n19 66.9805
R48 VPWR.n19 VPWR.t1 41.3705
R49 VPWR.n20 VPWR.t2 40.3855
R50 VPWR.n18 VPWR.n17 34.6358
R51 VPWR.n6 VPWR.t3 32.5055
R52 VPWR.n5 VPWR.t4 32.5055
R53 VPWR.n10 VPWR.n9 31.2544
R54 VPWR.n12 VPWR.t0 26.5955
R55 VPWR.n11 VPWR.t5 26.5955
R56 VPWR.n24 VPWR.n0 26.5
R57 VPWR.n13 VPWR.n10 15.1346
R58 VPWR.n17 VPWR.n2 11.3699
R59 VPWR.n9 VPWR.n8 9.3005
R60 VPWR.n10 VPWR.n3 9.3005
R61 VPWR.n15 VPWR.n14 9.3005
R62 VPWR.n17 VPWR.n16 9.3005
R63 VPWR.n18 VPWR.n1 9.3005
R64 VPWR.n23 VPWR.n22 9.3005
R65 VPWR.n8 VPWR.n7 7.99781
R66 VPWR.n7 VPWR.n4 7.91323
R67 VPWR.n21 VPWR.n18 7.60521
R68 VPWR.n22 VPWR.n21 5.70232
R69 VPWR.n14 VPWR.n2 4.53868
R70 VPWR.n14 VPWR.n13 3.37505
R71 VPWR.n9 VPWR.n4 2.32777
R72 VPWR.n22 VPWR.n0 2.21141
R73 VPWR VPWR.n24 0.476158
R74 VPWR.n24 VPWR.n23 0.147154
R75 VPWR.n8 VPWR.n3 0.120292
R76 VPWR.n15 VPWR.n3 0.120292
R77 VPWR.n16 VPWR.n15 0.120292
R78 VPWR.n16 VPWR.n1 0.120292
R79 VPWR.n23 VPWR.n1 0.120292
R80 a_27_297.n1 a_27_297.t7 416.829
R81 a_27_297.n3 a_27_297.t4 388.515
R82 a_27_297.n3 a_27_297.n2 298.673
R83 a_27_297.n1 a_27_297.n0 296.493
R84 a_27_297.n7 a_27_297.n6 296.493
R85 a_27_297.n5 a_27_297.n4 288.601
R86 a_27_297.n6 a_27_297.n5 107.567
R87 a_27_297.n6 a_27_297.n1 91.1064
R88 a_27_297.n5 a_27_297.n3 71.0485
R89 a_27_297.n7 a_27_297.t9 32.5055
R90 a_27_297.n0 a_27_297.t8 27.5805
R91 a_27_297.n2 a_27_297.t3 26.5955
R92 a_27_297.n2 a_27_297.t0 26.5955
R93 a_27_297.n4 a_27_297.t5 26.5955
R94 a_27_297.n4 a_27_297.t2 26.5955
R95 a_27_297.n0 a_27_297.t1 26.5955
R96 a_27_297.t6 a_27_297.n7 26.5955
R97 VPB.t5 VPB.t6 535.67
R98 VPB.t8 VPB.t7 485.358
R99 VPB.t9 VPB.t1 449.844
R100 VPB.t6 VPB.t9 266.356
R101 VPB.t1 VPB.t8 251.559
R102 VPB.t2 VPB.t5 248.599
R103 VPB.t3 VPB.t2 248.599
R104 VPB.t0 VPB.t3 248.599
R105 VPB.t4 VPB.t0 248.599
R106 VPB VPB.t4 189.409
R107 A2.n1 A2.t2 239.742
R108 A2.n4 A2.t0 227.969
R109 A2.n5 A2.n4 152
R110 A2.n2 A2.n0 152
R111 A2.n1 A2.t3 149.421
R112 A2.n3 A2.t1 149.421
R113 A2.n2 A2.n1 56.2338
R114 A2.n4 A2.n3 41.9524
R115 A2.n3 A2.n2 18.7449
R116 A2.n5 A2.n0 7.91323
R117 A2 A2.n5 1.39686
R118 A2.n0 A2 1.39686
R119 A3.n3 A3.t1 275.276
R120 A3.n0 A3.t0 234.952
R121 A3.n0 A3.t2 162.651
R122 A3 A3.n0 152.583
R123 A3.n2 A3.n1 152
R124 A3.n5 A3.n4 152
R125 A3.n3 A3.t3 149.421
R126 A3.n4 A3.n2 60.6968
R127 A3.n2 A3.n0 14.282
R128 A3.n1 A3 7.33141
R129 A3 A3.n5 6.16777
R130 A3.n5 A3 4.53868
R131 A3.n4 A3.n3 4.46346
R132 A3.n1 A3 3.37505
R133 B1.n0 B1.t0 221.72
R134 B1.n1 B1.t1 221.72
R135 B1.n3 B1.n2 152
R136 B1.n0 B1.t2 133.353
R137 B1.n1 B1.t3 133.353
R138 B1.n2 B1.n0 58.7443
R139 B1.n3 B1 14.4213
R140 B1.n4 B1.n3 10.0576
R141 B1.n4 B1 6.5566
R142 B1 B1.n4 6.4005
R143 B1.n2 B1.n1 4.51925
R144 a_730_47.n1 a_730_47.n0 376.865
R145 a_730_47.n0 a_730_47.t3 38.7697
R146 a_730_47.n0 a_730_47.t2 29.539
R147 a_730_47.t1 a_730_47.n1 24.9236
R148 a_730_47.n1 a_730_47.t0 24.9236
R149 VGND.n7 VGND.t2 234.596
R150 VGND.n21 VGND.n1 207.213
R151 VGND.n6 VGND.t3 156.715
R152 VGND.n22 VGND.n21 43.1829
R153 VGND.n9 VGND.n8 34.6358
R154 VGND.n9 VGND.n4 34.6358
R155 VGND.n13 VGND.n4 34.6358
R156 VGND.n14 VGND.n13 34.6358
R157 VGND.n15 VGND.n14 34.6358
R158 VGND.n15 VGND.n2 34.6358
R159 VGND.n19 VGND.n2 34.6358
R160 VGND.n20 VGND.n19 34.6358
R161 VGND.n1 VGND.t0 24.9236
R162 VGND.n1 VGND.t1 24.9236
R163 VGND.n8 VGND.n7 13.9299
R164 VGND.n20 VGND.n0 9.3005
R165 VGND.n19 VGND.n18 9.3005
R166 VGND.n17 VGND.n2 9.3005
R167 VGND.n16 VGND.n15 9.3005
R168 VGND.n14 VGND.n3 9.3005
R169 VGND.n13 VGND.n12 9.3005
R170 VGND.n11 VGND.n4 9.3005
R171 VGND.n10 VGND.n9 9.3005
R172 VGND.n8 VGND.n5 9.3005
R173 VGND.n7 VGND.n6 6.97444
R174 VGND.n21 VGND.n20 0.753441
R175 VGND.n6 VGND.n5 0.592283
R176 VGND.n10 VGND.n5 0.120292
R177 VGND.n11 VGND.n10 0.120292
R178 VGND.n12 VGND.n11 0.120292
R179 VGND.n12 VGND.n3 0.120292
R180 VGND.n16 VGND.n3 0.120292
R181 VGND.n17 VGND.n16 0.120292
R182 VGND.n18 VGND.n17 0.120292
R183 VGND.n18 VGND.n0 0.120292
R184 VGND.n22 VGND.n0 0.120292
R185 VGND VGND.n22 0.0213333
R186 B2.n0 B2.t0 212.081
R187 B2.n2 B2.t2 212.081
R188 B2.n3 B2.n2 173.91
R189 B2.n1 B2 155.048
R190 B2.n0 B2.t1 139.78
R191 B2.n2 B2.t3 139.78
R192 B2.n1 B2.n0 33.5944
R193 B2.n2 B2.n1 27.752
R194 B2.n3 B2 17.6767
R195 B2.n4 B2 11.3783
R196 B2.n4 B2.n3 5.18145
R197 B2 B2.n4 5.18145
R198 a_27_47.t1 a_27_47.n1 340.281
R199 a_27_47.n1 a_27_47.t2 209.018
R200 a_27_47.n1 a_27_47.n0 88.0229
R201 a_27_47.n0 a_27_47.t0 24.9236
R202 a_27_47.n0 a_27_47.t3 24.9236
C0 A1 VPWR 0.043931f
C1 A2 Y 0.001621f
C2 B1 VGND 0.020007f
C3 A2 VPWR 0.041444f
C4 A1 VGND 0.024126f
C5 A3 Y 3.25e-19
C6 VPB B2 0.071827f
C7 A3 VPWR 0.052561f
C8 A2 VGND 0.023678f
C9 VPB B1 0.054491f
C10 A3 VGND 0.079111f
C11 Y VPWR 0.022789f
C12 B2 B1 0.074181f
C13 VPB A1 0.093549f
C14 Y VGND 0.032575f
C15 VPB A2 0.082915f
C16 VPWR VGND 0.120298f
C17 B1 A1 0.040075f
C18 VPB A3 0.103473f
C19 VPB Y 0.008378f
C20 B2 Y 0.061374f
C21 VPB VPWR 0.110151f
C22 A1 A2 0.080213f
C23 B1 Y 0.142741f
C24 VPB VGND 0.007275f
C25 B2 VPWR 0.019567f
C26 B2 VGND 0.031393f
C27 A2 A3 0.085013f
C28 B1 VPWR 0.017326f
C29 A1 Y 0.117312f
C30 VGND VNB 0.702174f
C31 VPWR VNB 0.551414f
C32 Y VNB 0.039152f
C33 A3 VNB 0.292024f
C34 A2 VNB 0.213522f
C35 A1 VNB 0.230324f
C36 B1 VNB 0.181127f
C37 B2 VNB 0.239495f
C38 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32oi_4 VNB VPB VGND VPWR A3 A2 A1 B1 Y B2
X0 a_27_47.t7 B1.t0 Y.t15 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_297.t6 A2.t0 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47.t6 B1.t1 Y.t14 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297.t7 A3.t0 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t11 A1.t0 a_27_297.t19 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.3375 pd=1.675 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1249_47.t7 A3.t1 VGND.t7 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR.t5 A2.t1 a_27_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1249_47.t6 A3.t2 VGND.t6 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t11 B1.t2 a_27_297.t18 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_297.t9 A1.t1 VPWR.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t0 A3.t3 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297.t8 A1.t2 VPWR.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2525 pd=1.505 as=0.3375 ps=1.675 w=1 l=0.15
X12 a_803_47.t7 A2.t2 a_1249_47.t2 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297.t11 B2.t0 Y.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_297.t1 A3.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t10 A1.t3 a_27_297.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X16 a_803_47.t6 A2.t3 a_1249_47.t1 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y.t3 A1.t4 a_803_47.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t5 B2.t1 a_27_297.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR.t2 A3.t5 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 Y.t1 A1.t5 a_803_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_27_297.t13 B2.t2 Y.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1249_47.t3 A2.t4 a_803_47.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13325 ps=1.06 w=0.65 l=0.15
X23 a_27_297.t4 A2.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_47.t0 B2.t3 VGND.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_27_47.t1 B2.t4 VGND.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_1249_47.t0 A2.t6 a_803_47.t4 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR.t3 A2.t7 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2525 ps=1.505 w=1 l=0.15
X28 a_803_47.t1 A1.t6 Y.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_27_297.t17 B1.t3 Y.t10 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X30 a_803_47.t0 A1.t7 Y.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VGND.t2 B2.t5 a_27_47.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 Y.t13 B1.t4 a_27_47.t5 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 Y.t9 B1.t5 a_27_297.t16 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y.t12 B1.t6 a_27_47.t4 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_27_297.t15 B1.t7 Y.t8 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND.t5 A3.t6 a_1249_47.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 Y.t7 B2.t6 a_27_297.t14 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VGND.t4 A3.t7 a_1249_47.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VGND.t3 B2.t7 a_27_47.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n1 B1.t3 212.081
R1 B1.n5 B1.t5 212.081
R2 B1.n7 B1.t7 212.081
R3 B1.n6 B1.t2 212.081
R4 B1 B1.n8 161.31
R5 B1.n3 B1.n2 152
R6 B1.n4 B1.n0 152
R7 B1.n1 B1.t1 139.78
R8 B1.n5 B1.t6 139.78
R9 B1.n7 B1.t0 139.78
R10 B1.n6 B1.t4 139.78
R11 B1.n7 B1.n6 61.346
R12 B1.n4 B1.n3 49.6611
R13 B1.n8 B1.n5 46.7399
R14 B1.n8 B1.n7 14.6066
R15 B1.n2 B1.n0 13.1884
R16 B1.n3 B1.n1 8.76414
R17 B1 B1.n0 3.87929
R18 B1.n5 B1.n4 2.92171
R19 B1.n2 B1 0.776258
R20 Y.n10 Y.n8 334.161
R21 Y.n13 Y.n7 334.161
R22 Y.n10 Y.n9 295.76
R23 Y.n12 Y.n11 293.022
R24 Y.n2 Y.n0 248.248
R25 Y.n2 Y.n1 185
R26 Y.n4 Y.n3 185
R27 Y.n6 Y.n5 185
R28 Y.n4 Y.n2 102.4
R29 Y.n6 Y.n4 63.2476
R30 Y.n8 Y.t6 26.5955
R31 Y.n8 Y.t7 26.5955
R32 Y.n9 Y.t4 26.5955
R33 Y.n9 Y.t5 26.5955
R34 Y.n7 Y.t10 26.5955
R35 Y.n7 Y.t9 26.5955
R36 Y.n11 Y.t8 26.5955
R37 Y.n11 Y.t11 26.5955
R38 Y.n5 Y.t15 24.9236
R39 Y.n5 Y.t13 24.9236
R40 Y.n3 Y.t14 24.9236
R41 Y.n3 Y.t12 24.9236
R42 Y.n1 Y.t0 24.9236
R43 Y.n1 Y.t1 24.9236
R44 Y.n0 Y.t2 24.9236
R45 Y.n0 Y.t3 24.9236
R46 Y Y.n6 23.7278
R47 Y.n13 Y.n10 21.8358
R48 Y.n14 Y 4.26717
R49 Y Y.n14 3.02595
R50 Y.n14 Y.n13 1.97868
R51 Y.n12 Y 1.45813
R52 Y.n13 Y.n12 1.44577
R53 a_27_47.t6 a_27_47.n5 331.325
R54 a_27_47.n1 a_27_47.t3 329.051
R55 a_27_47.n1 a_27_47.n0 201.189
R56 a_27_47.n5 a_27_47.n4 185
R57 a_27_47.n3 a_27_47.n2 185
R58 a_27_47.n3 a_27_47.n1 76.0476
R59 a_27_47.n5 a_27_47.n3 63.2476
R60 a_27_47.n2 a_27_47.t5 24.9236
R61 a_27_47.n2 a_27_47.t1 24.9236
R62 a_27_47.n0 a_27_47.t2 24.9236
R63 a_27_47.n0 a_27_47.t0 24.9236
R64 a_27_47.n4 a_27_47.t4 24.9236
R65 a_27_47.n4 a_27_47.t7 24.9236
R66 VNB.t19 VNB.t0 2677.02
R67 VNB.t17 VNB.t5 2677.02
R68 VNB.t6 VNB.t12 1594.82
R69 VNB.t1 VNB.t3 1196.12
R70 VNB.t2 VNB.t1 1196.12
R71 VNB.t0 VNB.t2 1196.12
R72 VNB.t13 VNB.t19 1196.12
R73 VNB.t14 VNB.t13 1196.12
R74 VNB.t12 VNB.t14 1196.12
R75 VNB.t10 VNB.t6 1196.12
R76 VNB.t4 VNB.t10 1196.12
R77 VNB.t5 VNB.t4 1196.12
R78 VNB.t15 VNB.t17 1196.12
R79 VNB.t18 VNB.t15 1196.12
R80 VNB.t16 VNB.t18 1196.12
R81 VNB.t8 VNB.t16 1196.12
R82 VNB.t9 VNB.t8 1196.12
R83 VNB.t7 VNB.t9 1196.12
R84 VNB.t11 VNB.t7 1196.12
R85 VNB VNB.t11 669.256
R86 A2.n2 A2.t1 205.654
R87 A2.n8 A2.t5 205.654
R88 A2.n9 A2.t7 205.654
R89 A2.n1 A2.t0 205.654
R90 A2.n4 A2.n3 152
R91 A2.n5 A2.n0 152
R92 A2.n7 A2.n6 152
R93 A2.n11 A2.n10 152
R94 A2.n1 A2.t3 144.601
R95 A2.n2 A2.t6 139.78
R96 A2.n8 A2.t2 139.78
R97 A2.n9 A2.t4 139.78
R98 A2.n7 A2.n0 46.8234
R99 A2.n10 A2.n8 45.4462
R100 A2.n3 A2.n2 38.3858
R101 A2.n3 A2.n1 21.5826
R102 A2.n6 A2.n5 19.3427
R103 A2.n11 A2 17.6361
R104 A2 A2.n4 14.2227
R105 A2.n10 A2.n9 12.3948
R106 A2.n4 A2 11.9472
R107 A2.n2 A2.n0 9.6405
R108 A2 A2.n11 8.53383
R109 A2.n5 A2 5.1205
R110 A2.n6 A2 1.70717
R111 A2.n8 A2.n7 1.37764
R112 VPWR.n16 VPWR.n7 599.74
R113 VPWR.n12 VPWR.n9 315.909
R114 VPWR.n18 VPWR.n5 310.502
R115 VPWR.n11 VPWR.n10 310.502
R116 VPWR.n1 VPWR.n0 310.5
R117 VPWR.n25 VPWR.n24 146.25
R118 VPWR.n24 VPWR.t11 66.9805
R119 VPWR.n24 VPWR.t8 65.9955
R120 VPWR.n19 VPWR.n3 34.6358
R121 VPWR.n15 VPWR.n8 34.6358
R122 VPWR.n27 VPWR.n26 30.9811
R123 VPWR.n17 VPWR.n16 28.9887
R124 VPWR.n11 VPWR.n8 27.4829
R125 VPWR.n0 VPWR.t9 26.5955
R126 VPWR.n0 VPWR.t10 26.5955
R127 VPWR.n5 VPWR.t4 26.5955
R128 VPWR.n5 VPWR.t3 26.5955
R129 VPWR.n7 VPWR.t6 26.5955
R130 VPWR.n7 VPWR.t5 26.5955
R131 VPWR.n10 VPWR.t1 26.5955
R132 VPWR.n10 VPWR.t2 26.5955
R133 VPWR.n9 VPWR.t7 26.5955
R134 VPWR.n9 VPWR.t0 26.5955
R135 VPWR.n23 VPWR.n3 25.499
R136 VPWR.n16 VPWR.n15 15.4358
R137 VPWR.n27 VPWR.n1 10.9181
R138 VPWR.n18 VPWR.n17 9.41227
R139 VPWR.n13 VPWR.n8 9.3005
R140 VPWR.n15 VPWR.n14 9.3005
R141 VPWR.n16 VPWR.n6 9.3005
R142 VPWR.n17 VPWR.n4 9.3005
R143 VPWR.n20 VPWR.n19 9.3005
R144 VPWR.n21 VPWR.n3 9.3005
R145 VPWR.n23 VPWR.n22 9.3005
R146 VPWR.n26 VPWR.n2 9.3005
R147 VPWR.n28 VPWR.n27 9.3005
R148 VPWR.n29 VPWR.n1 7.56314
R149 VPWR.n12 VPWR.n11 6.17809
R150 VPWR.n26 VPWR.n25 3.95556
R151 VPWR.n25 VPWR.n23 2.66117
R152 VPWR VPWR.n29 0.936194
R153 VPWR.n13 VPWR.n12 0.653571
R154 VPWR.n19 VPWR.n18 0.376971
R155 VPWR.n29 VPWR.n28 0.147777
R156 VPWR.n14 VPWR.n13 0.120292
R157 VPWR.n14 VPWR.n6 0.120292
R158 VPWR.n6 VPWR.n4 0.120292
R159 VPWR.n20 VPWR.n4 0.120292
R160 VPWR.n21 VPWR.n20 0.120292
R161 VPWR.n22 VPWR.n21 0.120292
R162 VPWR.n22 VPWR.n2 0.120292
R163 VPWR.n28 VPWR.n2 0.120292
R164 a_27_297.n7 a_27_297.t14 917.229
R165 a_27_297.n12 a_27_297.n5 585
R166 a_27_297.n11 a_27_297.n10 585
R167 a_27_297.n9 a_27_297.n8 585
R168 a_27_297.n7 a_27_297.n6 585
R169 a_27_297.n1 a_27_297.t7 404.793
R170 a_27_297.n1 a_27_297.n0 314.952
R171 a_27_297.n15 a_27_297.n2 314.952
R172 a_27_297.n14 a_27_297.n3 314.952
R173 a_27_297.n13 a_27_297.n4 314.952
R174 a_27_297.n17 a_27_297.n16 314.952
R175 a_27_297.n17 a_27_297.t2 129.036
R176 a_27_297.n13 a_27_297.n12 103.153
R177 a_27_297.n16 a_27_297.n1 102.4
R178 a_27_297.n14 a_27_297.n13 93.7417
R179 a_27_297.n15 a_27_297.n14 80.9417
R180 a_27_297.n3 a_27_297.t3 72.8905
R181 a_27_297.n12 a_27_297.n11 63.2476
R182 a_27_297.n11 a_27_297.n9 63.2476
R183 a_27_297.n9 a_27_297.n7 63.2476
R184 a_27_297.n16 a_27_297.n15 63.2476
R185 a_27_297.n5 a_27_297.t10 30.5355
R186 a_27_297.n0 a_27_297.t0 26.5955
R187 a_27_297.n0 a_27_297.t1 26.5955
R188 a_27_297.n2 a_27_297.t5 26.5955
R189 a_27_297.n2 a_27_297.t4 26.5955
R190 a_27_297.n3 a_27_297.t8 26.5955
R191 a_27_297.n4 a_27_297.t19 26.5955
R192 a_27_297.n4 a_27_297.t9 26.5955
R193 a_27_297.n6 a_27_297.t12 26.5955
R194 a_27_297.n6 a_27_297.t13 26.5955
R195 a_27_297.n8 a_27_297.t18 26.5955
R196 a_27_297.n8 a_27_297.t11 26.5955
R197 a_27_297.n10 a_27_297.t16 26.5955
R198 a_27_297.n10 a_27_297.t15 26.5955
R199 a_27_297.n5 a_27_297.t17 26.5955
R200 a_27_297.t6 a_27_297.n17 26.5955
R201 VPB.t6 VPB.t2 556.386
R202 VPB.t19 VPB.t8 488.318
R203 VPB.t8 VPB.t3 387.695
R204 VPB.t17 VPB.t10 260.437
R205 VPB.t0 VPB.t7 248.599
R206 VPB.t1 VPB.t0 248.599
R207 VPB.t2 VPB.t1 248.599
R208 VPB.t5 VPB.t6 248.599
R209 VPB.t4 VPB.t5 248.599
R210 VPB.t3 VPB.t4 248.599
R211 VPB.t9 VPB.t19 248.599
R212 VPB.t10 VPB.t9 248.599
R213 VPB.t16 VPB.t17 248.599
R214 VPB.t15 VPB.t16 248.599
R215 VPB.t18 VPB.t15 248.599
R216 VPB.t11 VPB.t18 248.599
R217 VPB.t12 VPB.t11 248.599
R218 VPB.t13 VPB.t12 248.599
R219 VPB.t14 VPB.t13 248.599
R220 VPB VPB.t14 139.097
R221 A3.n2 A3.t0 212.081
R222 A3.n4 A3.t3 212.081
R223 A3.n5 A3.t4 212.081
R224 A3.n6 A3.t5 212.081
R225 A3.n2 A3.n1 182.069
R226 A3.n3 A3.n0 152
R227 A3.n12 A3.n11 152
R228 A3.n10 A3.n9 152
R229 A3.n8 A3.n7 152
R230 A3.n2 A3.t7 139.78
R231 A3.n4 A3.t2 139.78
R232 A3.n5 A3.t6 139.78
R233 A3.n6 A3.t1 139.78
R234 A3.n11 A3.n10 49.6611
R235 A3.n7 A3.n5 48.2005
R236 A3.n4 A3.n3 39.4369
R237 A3.n1 A3 26.7279
R238 A3.n3 A3.n2 21.9096
R239 A3.n9 A3.n8 21.2298
R240 A3 A3.n0 20.6054
R241 A3.n12 A3 15.6103
R242 A3.n7 A3.n6 13.146
R243 A3 A3.n12 13.1127
R244 A3.n11 A3.n4 10.2247
R245 A3 A3.n0 8.11757
R246 A3.n9 A3 5.62001
R247 A3.n8 A3 1.87367
R248 A3.n10 A3.n5 1.46111
R249 A3.n1 A3 0.62489
R250 A1.n1 A1.t2 230.867
R251 A1.n5 A1.t3 218.048
R252 A1.n11 A1.t0 205.654
R253 A1.n6 A1.t1 205.654
R254 A1.n0 A1.t6 169.867
R255 A1 A1.n0 156.575
R256 A1.n14 A1.n13 152
R257 A1.n10 A1.n9 152
R258 A1.n8 A1.n7 152
R259 A1.n5 A1.n4 152
R260 A1.n3 A1.t5 139.78
R261 A1.n12 A1.t7 139.78
R262 A1.n2 A1.t4 139.78
R263 A1.n6 A1.n5 45.4462
R264 A1.n10 A1.n3 37.1834
R265 A1.n13 A1.n2 31.6748
R266 A1.n13 A1.n12 26.1662
R267 A1.n8 A1.n4 20.7243
R268 A1.n9 A1 18.8957
R269 A1 A1.n14 16.4576
R270 A1.n14 A1 11.5815
R271 A1.n12 A1.n11 11.0176
R272 A1.n2 A1.n1 10.3291
R273 A1.n11 A1.n10 9.6405
R274 A1.n7 A1.n3 9.6405
R275 A1.n9 A1 9.14336
R276 A1.n4 A1 5.48621
R277 A1.n1 A1.n0 1.91614
R278 A1 A1.n8 1.82907
R279 A1.n7 A1.n6 1.37764
R280 VGND.n10 VGND.t4 282.866
R281 VGND.n14 VGND.t7 282.817
R282 VGND.n12 VGND.n11 199.739
R283 VGND.n36 VGND.n2 199.739
R284 VGND.n39 VGND.n38 199.739
R285 VGND.n18 VGND.n8 34.6358
R286 VGND.n19 VGND.n18 34.6358
R287 VGND.n20 VGND.n19 34.6358
R288 VGND.n20 VGND.n6 34.6358
R289 VGND.n24 VGND.n6 34.6358
R290 VGND.n25 VGND.n24 34.6358
R291 VGND.n26 VGND.n25 34.6358
R292 VGND.n26 VGND.n4 34.6358
R293 VGND.n30 VGND.n4 34.6358
R294 VGND.n31 VGND.n30 34.6358
R295 VGND.n32 VGND.n31 34.6358
R296 VGND.n32 VGND.n1 34.6358
R297 VGND.n14 VGND.n8 30.4946
R298 VGND.n36 VGND.n1 28.9887
R299 VGND.n11 VGND.t6 24.9236
R300 VGND.n11 VGND.t5 24.9236
R301 VGND.n2 VGND.t1 24.9236
R302 VGND.n2 VGND.t2 24.9236
R303 VGND.n38 VGND.t0 24.9236
R304 VGND.n38 VGND.t3 24.9236
R305 VGND.n13 VGND.n12 24.4711
R306 VGND.n39 VGND.n37 22.9652
R307 VGND.n37 VGND.n36 15.4358
R308 VGND.n14 VGND.n13 13.9299
R309 VGND.n13 VGND.n9 9.3005
R310 VGND.n15 VGND.n14 9.3005
R311 VGND.n16 VGND.n8 9.3005
R312 VGND.n18 VGND.n17 9.3005
R313 VGND.n19 VGND.n7 9.3005
R314 VGND.n21 VGND.n20 9.3005
R315 VGND.n22 VGND.n6 9.3005
R316 VGND.n24 VGND.n23 9.3005
R317 VGND.n25 VGND.n5 9.3005
R318 VGND.n27 VGND.n26 9.3005
R319 VGND.n28 VGND.n4 9.3005
R320 VGND.n30 VGND.n29 9.3005
R321 VGND.n31 VGND.n3 9.3005
R322 VGND.n33 VGND.n32 9.3005
R323 VGND.n34 VGND.n1 9.3005
R324 VGND.n36 VGND.n35 9.3005
R325 VGND.n37 VGND.n0 9.3005
R326 VGND.n40 VGND.n39 7.12063
R327 VGND.n12 VGND.n10 6.30332
R328 VGND.n10 VGND.n9 0.741903
R329 VGND.n40 VGND.n0 0.148519
R330 VGND.n15 VGND.n9 0.120292
R331 VGND.n16 VGND.n15 0.120292
R332 VGND.n17 VGND.n16 0.120292
R333 VGND.n17 VGND.n7 0.120292
R334 VGND.n21 VGND.n7 0.120292
R335 VGND.n22 VGND.n21 0.120292
R336 VGND.n23 VGND.n22 0.120292
R337 VGND.n23 VGND.n5 0.120292
R338 VGND.n27 VGND.n5 0.120292
R339 VGND.n28 VGND.n27 0.120292
R340 VGND.n29 VGND.n28 0.120292
R341 VGND.n29 VGND.n3 0.120292
R342 VGND.n33 VGND.n3 0.120292
R343 VGND.n34 VGND.n33 0.120292
R344 VGND.n35 VGND.n34 0.120292
R345 VGND.n35 VGND.n0 0.120292
R346 VGND VGND.n40 0.0927068
R347 a_1249_47.n5 a_1249_47.n4 264.435
R348 a_1249_47.n3 a_1249_47.n1 248.248
R349 a_1249_47.n4 a_1249_47.n0 201.189
R350 a_1249_47.n3 a_1249_47.n2 185
R351 a_1249_47.n4 a_1249_47.n3 102.4
R352 a_1249_47.n1 a_1249_47.t2 24.9236
R353 a_1249_47.n1 a_1249_47.t3 24.9236
R354 a_1249_47.n2 a_1249_47.t1 24.9236
R355 a_1249_47.n2 a_1249_47.t0 24.9236
R356 a_1249_47.n0 a_1249_47.t5 24.9236
R357 a_1249_47.n0 a_1249_47.t7 24.9236
R358 a_1249_47.n5 a_1249_47.t4 24.9236
R359 a_1249_47.t6 a_1249_47.n5 24.9236
R360 a_803_47.n4 a_803_47.t2 331.325
R361 a_803_47.n1 a_803_47.t6 331.325
R362 a_803_47.n1 a_803_47.n0 185
R363 a_803_47.n3 a_803_47.n2 185
R364 a_803_47.n5 a_803_47.n4 185
R365 a_803_47.n3 a_803_47.n1 73.7887
R366 a_803_47.n4 a_803_47.n3 63.2476
R367 a_803_47.n2 a_803_47.t5 50.7697
R368 a_803_47.n2 a_803_47.t1 24.9236
R369 a_803_47.n0 a_803_47.t4 24.9236
R370 a_803_47.n0 a_803_47.t7 24.9236
R371 a_803_47.t3 a_803_47.n5 24.9236
R372 a_803_47.n5 a_803_47.t0 24.9236
R373 B2.n0 B2.t0 212.081
R374 B2.n1 B2.t1 212.081
R375 B2.n2 B2.t2 212.081
R376 B2.n5 B2.t6 212.081
R377 B2.n5 B2.n4 182.899
R378 B2.n11 B2.n10 152
R379 B2.n9 B2.n8 152
R380 B2.n7 B2.n6 152
R381 B2.n0 B2.t4 139.78
R382 B2.n1 B2.t5 139.78
R383 B2.n2 B2.t3 139.78
R384 B2.n5 B2.t7 139.78
R385 B2.n1 B2.n0 61.346
R386 B2.n10 B2.n9 49.6611
R387 B2.n6 B2.n2 40.1672
R388 B2.n6 B2.n5 21.1793
R389 B2.n8 B2.n7 18.9222
R390 B2.n4 B2 18.644
R391 B2 B2.n11 13.0788
R392 B2.n11 B2 12.5222
R393 B2.n9 B2.n2 9.49444
R394 B2.n3 B2 8.14595
R395 B2.n8 B2 6.4005
R396 B2.n3 B2 3.89615
R397 B2.n4 B2.n3 3.06137
R398 B2.n10 B2.n1 2.19141
R399 B2.n7 B2 0.278761
C0 B2 B1 0.050963f
C1 VPB A1 0.152006f
C2 Y VGND 0.051987f
C3 VPB A2 0.124033f
C4 VPWR VGND 0.195553f
C5 VPB A3 0.139318f
C6 B1 A1 0.058187f
C7 B1 A2 3.89e-19
C8 VPB Y 0.012377f
C9 B2 Y 0.192765f
C10 B1 A3 4.43e-19
C11 VPB VPWR 0.185164f
C12 A1 A2 0.040203f
C13 B2 VPWR 0.038576f
C14 B1 Y 0.256874f
C15 A1 A3 1.9e-19
C16 VPB VGND 0.014768f
C17 A1 Y 0.138399f
C18 B2 VGND 0.070211f
C19 B1 VPWR 0.02844f
C20 A2 A3 0.025731f
C21 A1 VPWR 0.086596f
C22 A2 Y 8.23e-19
C23 B1 VGND 0.032157f
C24 A3 Y 8.09e-19
C25 A2 VPWR 0.07789f
C26 A1 VGND 0.039157f
C27 VPB B2 0.140779f
C28 A2 VGND 0.037784f
C29 A3 VPWR 0.085763f
C30 VPB B1 0.115432f
C31 A3 VGND 0.095845f
C32 Y VPWR 0.042499f
C33 VGND VNB 1.09159f
C34 VPWR VNB 0.893351f
C35 Y VNB 0.038314f
C36 A3 VNB 0.446533f
C37 A2 VNB 0.373684f
C38 A1 VNB 0.414227f
C39 B1 VNB 0.35759f
C40 B2 VNB 0.441999f
C41 VPB VNB 2.0223f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB
X0 a_465_47.t1 A2.t0 a_381_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t0 A4.t0 a_561_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR.t2 A3.t0 a_297_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297.t3 A2.t1 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297.t1 A4.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR.t4 A1.t0 a_297_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47.t1 A1.t1 a_79_21.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X7 a_297_297.t0 B1.t0 a_79_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR.t0 a_79_21.t3 X.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21.t2 B1.t1 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X10 VGND.t2 a_79_21.t4 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47.t1 A3.t1 a_465_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
R0 A2.n0 A2.t1 241.536
R1 A2.n1 A2.n0 190.109
R2 A2.n0 A2.t0 169.237
R3 A2.n1 A2 14.8762
R4 A2 A2.n1 4.99562
R5 a_381_47.t0 a_381_47.t1 49.8467
R6 a_465_47.t0 a_465_47.t1 60.9236
R7 VNB.t4 VNB.t3 2036.25
R8 VNB.t5 VNB.t4 1836.89
R9 VNB.t0 VNB.t2 1366.99
R10 VNB.t1 VNB.t0 1366.99
R11 VNB.t3 VNB.t1 1196.12
R12 VNB VNB.t5 911.327
R13 A4.n0 A4.t1 230.155
R14 A4.n0 A4.t0 157.856
R15 A4.n1 A4.n0 152
R16 A4.n1 A4 14.3064
R17 A4 A4.n1 2.76128
R18 a_561_47.t0 a_561_47.t1 60.9236
R19 VGND.n1 VGND.n0 209.276
R20 VGND.n1 VGND.t0 156.99
R21 VGND.n0 VGND.t1 51.6928
R22 VGND.n0 VGND.t2 39.6928
R23 VGND VGND.n1 0.157741
R24 A3.n0 A3.t0 241.536
R25 A3.n0 A3.t1 169.237
R26 A3.n1 A3.n0 152
R27 A3 A3.n1 9.6005
R28 A3.n1 A3 1.85313
R29 a_297_297.n1 a_297_297.t1 397.55
R30 a_297_297.n2 a_297_297.n1 361.921
R31 a_297_297.n1 a_297_297.n0 298.673
R32 a_297_297.n0 a_297_297.t2 38.4155
R33 a_297_297.n0 a_297_297.t3 26.5955
R34 a_297_297.n2 a_297_297.t4 26.5955
R35 a_297_297.t0 a_297_297.n2 26.5955
R36 VPWR.n8 VPWR.t0 873.438
R37 VPWR.n4 VPWR.n3 610.235
R38 VPWR.n2 VPWR.n1 604.457
R39 VPWR.n7 VPWR.n6 34.6358
R40 VPWR.n3 VPWR.t1 32.5055
R41 VPWR.n3 VPWR.t2 32.5055
R42 VPWR.n1 VPWR.t3 26.5955
R43 VPWR.n1 VPWR.t4 26.5955
R44 VPWR.n6 VPWR.n2 22.9652
R45 VPWR.n8 VPWR.n7 22.9652
R46 VPWR.n6 VPWR.n5 9.3005
R47 VPWR.n7 VPWR.n0 9.3005
R48 VPWR.n9 VPWR.n8 7.4049
R49 VPWR.n4 VPWR.n2 6.94908
R50 VPWR.n5 VPWR.n4 0.510123
R51 VPWR.n9 VPWR.n0 0.144904
R52 VPWR.n5 VPWR.n0 0.120292
R53 VPWR VPWR.n9 0.117202
R54 VPB.t1 VPB.t0 556.386
R55 VPB.t3 VPB.t2 284.113
R56 VPB.t4 VPB.t3 284.113
R57 VPB.t5 VPB.t4 248.599
R58 VPB.t0 VPB.t5 248.599
R59 VPB VPB.t1 189.409
R60 A1.n0 A1.t0 241.536
R61 A1.n0 A1.t1 169.237
R62 A1 A1.n0 163.417
R63 a_79_21.t0 a_79_21.n2 408.671
R64 a_79_21.n1 a_79_21.t3 235.471
R65 a_79_21.n2 a_79_21.n0 171.476
R66 a_79_21.n1 a_79_21.t4 163.172
R67 a_79_21.n2 a_79_21.n1 152
R68 a_79_21.n0 a_79_21.t1 72.0005
R69 a_79_21.n0 a_79_21.t2 32.3082
R70 B1.n0 B1.t0 229.754
R71 B1.n0 B1.t1 157.453
R72 B1.n1 B1.n0 152
R73 B1.n1 B1 11.055
R74 B1 B1.n1 2.13383
R75 X.n4 X.n3 591.588
R76 X.n4 X.n0 585
R77 X.n5 X.n4 585
R78 X.t1 X 267.276
R79 X.n2 X.t1 261.154
R80 X.n4 X.t0 26.5955
R81 X X.n0 10.5851
R82 X.n5 X 10.5851
R83 X.n2 X.n1 8.12358
R84 X.n1 X 6.64665
R85 X X.n0 6.15435
R86 X X.n5 6.15435
R87 X X.n1 5.08285
R88 X.n3 X 1.96973
R89 X X.n2 1.96973
R90 X.n3 X 1.50638
C0 A3 VPWR 0.024002f
C1 A2 VGND 0.081373f
C2 VPB B1 0.043039f
C3 A3 VGND 0.074439f
C4 A4 VPWR 0.020016f
C5 VPB A1 0.028093f
C6 X VPWR 0.063082f
C7 A4 VGND 0.047952f
C8 B1 A1 0.099069f
C9 VPB A2 0.027392f
C10 X VGND 0.064052f
C11 VPB A3 0.03038f
C12 B1 A2 1.92e-19
C13 VPWR VGND 0.074653f
C14 A1 A2 0.099595f
C15 B1 A3 1.05e-19
C16 VPB A4 0.041818f
C17 B1 A4 6.93e-21
C18 VPB X 0.010526f
C19 A1 A3 0.008128f
C20 VPB VPWR 0.081935f
C21 B1 X 1.21e-19
C22 A2 A3 0.109547f
C23 VPB VGND 0.007308f
C24 B1 VPWR 0.017677f
C25 A3 A4 0.108209f
C26 A1 VPWR 0.019035f
C27 B1 VGND 0.014254f
C28 A1 VGND 0.016977f
C29 A2 VPWR 0.018762f
C30 VGND VNB 0.463871f
C31 VPWR VNB 0.364103f
C32 X VNB 0.092055f
C33 A4 VNB 0.156489f
C34 A3 VNB 0.099237f
C35 A2 VNB 0.096716f
C36 A1 VNB 0.093164f
C37 B1 VNB 0.112609f
C38 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_2 VNB VPB VGND VPWR X A1 A2 A3 A4 B1
X0 a_381_297.t1 A1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR.t3 A2.t0 a_381_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_465_47.t1 A4.t0 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_549_47.t0 A3.t0 a_465_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t5 a_79_21.t3 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t1 a_79_21.t4 X.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47.t1 A2.t1 a_549_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 a_381_297.t0 A3.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t4 A4.t1 a_381_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_381_297.t2 B1.t0 a_79_21.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21.t1 A1.t1 a_665_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t0 B1.t1 a_79_21.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 X.t0 a_79_21.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X.t2 a_79_21.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t0 231.478
R1 A1.n0 A1.t1 159.179
R2 A1.n1 A1.n0 152
R3 A1.n1 A1 16.5823
R4 A1 A1.n1 3.2005
R5 VPWR.n6 VPWR.n3 610.301
R6 VPWR.n5 VPWR.n4 604.457
R7 VPWR.n10 VPWR.t5 342.841
R8 VPWR.n12 VPWR.t0 243.512
R9 VPWR.n9 VPWR.n2 34.6358
R10 VPWR.n4 VPWR.t1 26.5955
R11 VPWR.n4 VPWR.t4 26.5955
R12 VPWR.n3 VPWR.t2 26.5955
R13 VPWR.n3 VPWR.t3 26.5955
R14 VPWR.n10 VPWR.n9 25.977
R15 VPWR.n11 VPWR.n10 24.4711
R16 VPWR.n12 VPWR.n11 19.9534
R17 VPWR.n5 VPWR.n2 19.9534
R18 VPWR.n7 VPWR.n2 9.3005
R19 VPWR.n9 VPWR.n8 9.3005
R20 VPWR.n10 VPWR.n1 9.3005
R21 VPWR.n11 VPWR.n0 9.3005
R22 VPWR.n13 VPWR.n12 9.3005
R23 VPWR.n6 VPWR.n5 7.12603
R24 VPWR.n7 VPWR.n6 0.462921
R25 VPWR.n8 VPWR.n7 0.120292
R26 VPWR.n8 VPWR.n1 0.120292
R27 VPWR.n1 VPWR.n0 0.120292
R28 VPWR.n13 VPWR.n0 0.120292
R29 VPWR VPWR.n13 0.0213333
R30 a_381_297.n1 a_381_297.t1 400.562
R31 a_381_297.n1 a_381_297.n0 361.921
R32 a_381_297.n2 a_381_297.n1 298.673
R33 a_381_297.n2 a_381_297.t3 58.1155
R34 a_381_297.n0 a_381_297.t4 26.5955
R35 a_381_297.n0 a_381_297.t2 26.5955
R36 a_381_297.t0 a_381_297.n2 26.5955
R37 VPB.t6 VPB.t3 556.386
R38 VPB.t1 VPB.t4 343.303
R39 VPB.t4 VPB.t2 248.599
R40 VPB.t5 VPB.t1 248.599
R41 VPB.t3 VPB.t5 248.599
R42 VPB.t0 VPB.t6 248.599
R43 VPB VPB.t0 189.409
R44 A2.n0 A2.t0 241.536
R45 A2.n0 A2.t1 169.237
R46 A2.n1 A2.n0 158.4
R47 A2.n1 A2 16.9679
R48 A2 A2.n1 3.27492
R49 A4.n0 A4.t1 241.536
R50 A4.n0 A4.t0 169.237
R51 A4.n1 A4.n0 152
R52 A4.n1 A4 10.8901
R53 A4 A4.n1 2.10199
R54 VGND.n3 VGND.t1 282.817
R55 VGND.n2 VGND.n1 205.197
R56 VGND.n5 VGND.t2 149.762
R57 VGND.n1 VGND.t3 24.9236
R58 VGND.n1 VGND.t0 24.9236
R59 VGND.n5 VGND.n4 19.9534
R60 VGND.n4 VGND.n3 18.4476
R61 VGND.n6 VGND.n5 9.3005
R62 VGND.n4 VGND.n0 9.3005
R63 VGND.n3 VGND.n2 6.82185
R64 VGND.n2 VGND.n0 0.556872
R65 VGND.n6 VGND.n0 0.120292
R66 VGND VGND.n6 0.0213333
R67 a_465_47.t0 a_465_47.t1 49.8467
R68 VNB.t1 VNB.t0 2677.02
R69 VNB.t3 VNB.t5 1651.78
R70 VNB.t5 VNB.t2 1196.12
R71 VNB.t6 VNB.t3 1196.12
R72 VNB.t0 VNB.t6 1196.12
R73 VNB.t4 VNB.t1 1196.12
R74 VNB VNB.t4 911.327
R75 A3.n0 A3.t1 237.736
R76 A3 A3.n0 181.802
R77 A3.n0 A3.t0 165.435
R78 a_549_47.t0 a_549_47.t1 79.3851
R79 a_79_21.n0 a_79_21.t1 444.642
R80 a_79_21.t2 a_79_21.n3 393.236
R81 a_79_21.n0 a_79_21.t0 267.901
R82 a_79_21.n2 a_79_21.t3 212.081
R83 a_79_21.n1 a_79_21.t5 212.081
R84 a_79_21.n3 a_79_21.n2 177.561
R85 a_79_21.n2 a_79_21.t4 139.78
R86 a_79_21.n1 a_79_21.t6 139.78
R87 a_79_21.n2 a_79_21.n1 61.346
R88 a_79_21.n3 a_79_21.n0 59.1064
R89 X.n0 X 596.789
R90 X.n1 X.n0 585
R91 X X.n2 207.886
R92 X.n0 X.t1 26.5955
R93 X.n0 X.t0 26.5955
R94 X.n2 X.t3 24.9236
R95 X.n2 X.t2 24.9236
R96 X X.n1 11.79
R97 X.n1 X 11.1163
R98 a_665_47.t0 a_665_47.t1 49.8467
R99 B1.n0 B1.t0 228.823
R100 B1.n0 B1.t1 156.524
R101 B1 B1.n0 154.133
C0 VPB VPWR 0.10141f
C1 A4 A2 3.43e-19
C2 B1 VPWR 0.015898f
C3 A3 A2 0.086866f
C4 VPB X 0.004419f
C5 A4 VPWR 0.018796f
C6 VPB VGND 0.008533f
C7 A3 A1 2.59e-20
C8 B1 VGND 0.017962f
C9 A2 A1 0.128076f
C10 A3 VPWR 0.018792f
C11 A2 VPWR 0.021787f
C12 A4 VGND 0.016662f
C13 A3 VGND 0.01123f
C14 A1 VPWR 0.019451f
C15 VPB B1 0.040735f
C16 A2 VGND 0.013186f
C17 VPB A4 0.028835f
C18 A1 VGND 0.013088f
C19 VPWR X 0.158011f
C20 VPB A3 0.032248f
C21 B1 A4 0.07883f
C22 VPWR VGND 0.097843f
C23 VPB A2 0.029744f
C24 X VGND 0.08579f
C25 VPB A1 0.038916f
C26 A4 A3 0.091671f
C27 B1 A2 1.96e-19
C28 VGND VNB 0.50993f
C29 X VNB 0.02808f
C30 VPWR VNB 0.438888f
C31 A1 VNB 0.164498f
C32 A2 VNB 0.097594f
C33 A3 VNB 0.095719f
C34 A4 VNB 0.089541f
C35 B1 VNB 0.112996f
C36 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_4 VNB VPB VGND VPWR A1 A2 A3 A4 X B1
X0 a_639_47.t3 A1.t0 a_79_21.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_639_47.t0 A2.t0 a_889_47.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t3 a_79_21.t6 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR.t11 A3.t0 a_467_297.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.145 ps=1.29 w=1 l=0.15
X4 a_889_47.t2 A2.t1 a_639_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_889_47.t0 A3.t1 a_1079_47.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 X.t2 a_79_21.t7 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t2 B1.t0 a_79_21.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t1 a_79_21.t8 X.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_467_297.t6 A4.t0 VPWR.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t6 a_79_21.t9 X.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t5 a_79_21.t10 X.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_467_297.t2 B1.t1 a_79_21.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X13 a_467_297.t9 A2.t2 VPWR.t10 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t8 A4.t1 a_467_297.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1079_47.t1 A3.t2 a_889_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_79_21.t2 B1.t2 a_467_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_79_21.t0 B1.t3 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X18 a_1079_47.t3 A4.t2 VGND.t7 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR.t9 A2.t3 a_467_297.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 X.t5 a_79_21.t11 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_467_297.t5 A1.t1 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_79_21.t4 A1.t2 a_639_47.t2 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 VPWR.t5 A1.t3 a_467_297.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X24 a_467_297.t0 A3.t3 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X25 VGND.t0 A4.t3 a_1079_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 X.t0 a_79_21.t12 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X.t4 a_79_21.t13 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t1 212.081
R1 A1.n2 A1.t3 212.081
R2 A1 A1.n1 153.745
R3 A1.n4 A1.n3 152
R4 A1.n0 A1.t0 139.78
R5 A1.n2 A1.t2 139.78
R6 A1.n3 A1.n1 49.6611
R7 A1 A1.n4 18.0369
R8 A1.n4 A1 8.72777
R9 A1.n1 A1.n0 7.30353
R10 A1.n3 A1.n2 4.38232
R11 a_79_21.n15 a_79_21.n14 396.277
R12 a_79_21.n2 a_79_21.n1 287.401
R13 a_79_21.n4 a_79_21.t6 212.081
R14 a_79_21.n10 a_79_21.t7 212.081
R15 a_79_21.n5 a_79_21.t8 212.081
R16 a_79_21.n6 a_79_21.t12 212.081
R17 a_79_21.n2 a_79_21.n0 201.941
R18 a_79_21.n8 a_79_21.n7 177.601
R19 a_79_21.n9 a_79_21.n8 152
R20 a_79_21.n11 a_79_21.n3 152
R21 a_79_21.n13 a_79_21.n12 152
R22 a_79_21.n4 a_79_21.t10 139.78
R23 a_79_21.n10 a_79_21.t11 139.78
R24 a_79_21.n5 a_79_21.t9 139.78
R25 a_79_21.n6 a_79_21.t13 139.78
R26 a_79_21.n14 a_79_21.n2 58.7299
R27 a_79_21.n12 a_79_21.n11 49.6611
R28 a_79_21.n10 a_79_21.n9 46.0096
R29 a_79_21.n7 a_79_21.n5 34.3247
R30 a_79_21.n7 a_79_21.n6 27.0217
R31 a_79_21.t1 a_79_21.n15 26.5955
R32 a_79_21.n15 a_79_21.t2 26.5955
R33 a_79_21.n13 a_79_21.n3 25.6005
R34 a_79_21.n8 a_79_21.n3 25.6005
R35 a_79_21.n1 a_79_21.t5 24.9236
R36 a_79_21.n1 a_79_21.t4 24.9236
R37 a_79_21.n0 a_79_21.t3 24.9236
R38 a_79_21.n0 a_79_21.t0 24.9236
R39 a_79_21.n9 a_79_21.n5 15.3369
R40 a_79_21.n14 a_79_21.n13 13.9299
R41 a_79_21.n12 a_79_21.n4 8.03383
R42 a_79_21.n11 a_79_21.n10 3.65202
R43 a_639_47.t2 a_639_47.n1 344.877
R44 a_639_47.n1 a_639_47.t0 326.709
R45 a_639_47.n1 a_639_47.n0 185
R46 a_639_47.n0 a_639_47.t1 24.9236
R47 a_639_47.n0 a_639_47.t3 24.9236
R48 VNB.t1 VNB.t8 2677.02
R49 VNB.t11 VNB.t12 2677.02
R50 VNB.t6 VNB.t3 1253.07
R51 VNB.t0 VNB.t10 1196.12
R52 VNB.t9 VNB.t0 1196.12
R53 VNB.t8 VNB.t9 1196.12
R54 VNB.t2 VNB.t1 1196.12
R55 VNB.t13 VNB.t2 1196.12
R56 VNB.t12 VNB.t13 1196.12
R57 VNB.t3 VNB.t11 1196.12
R58 VNB.t5 VNB.t6 1196.12
R59 VNB.t7 VNB.t5 1196.12
R60 VNB.t4 VNB.t7 1196.12
R61 VNB VNB.t4 911.327
R62 A2.n1 A2.t2 221.72
R63 A2.n2 A2.t3 221.72
R64 A2.n5 A2.n4 152
R65 A2.n3 A2.n0 152
R66 A2.n1 A2.t0 149.421
R67 A2.n2 A2.t1 149.421
R68 A2.n4 A2.n3 60.6968
R69 A2.n5 A2.n0 20.7243
R70 A2.n3 A2.n2 12.4968
R71 A2.n0 A2 6.70526
R72 A2.n4 A2.n1 1.78569
R73 A2 A2.n5 0.610024
R74 a_889_47.n1 a_889_47.n0 472.401
R75 a_889_47.n0 a_889_47.t1 24.9236
R76 a_889_47.n0 a_889_47.t0 24.9236
R77 a_889_47.n1 a_889_47.t3 24.9236
R78 a_889_47.t2 a_889_47.n1 24.9236
R79 X.n5 X.n4 378.199
R80 X.n5 X.n3 314.952
R81 X.n2 X.n1 264.435
R82 X.n2 X.n0 201.189
R83 X.n6 X.n5 33.5064
R84 X.n7 X.n2 33.5064
R85 X.n4 X.t3 26.5955
R86 X.n4 X.t2 26.5955
R87 X.n3 X.t1 26.5955
R88 X.n3 X.t0 26.5955
R89 X.n0 X.t7 24.9236
R90 X.n0 X.t4 24.9236
R91 X.n1 X.t6 24.9236
R92 X.n1 X.t5 24.9236
R93 X.n7 X 22.5887
R94 X X.n6 9.78874
R95 X.n6 X 6.4005
R96 X.n7 X 6.4005
R97 X X.n7 3.01226
R98 VPWR.n31 VPWR.t0 337.096
R99 VPWR.n3 VPWR.t3 336.07
R100 VPWR.n13 VPWR.n10 315.788
R101 VPWR.n29 VPWR.n2 310.502
R102 VPWR.n6 VPWR.n5 310.502
R103 VPWR.n17 VPWR.n8 310.502
R104 VPWR.n12 VPWR.n11 139.048
R105 VPWR.n11 VPWR.t11 72.013
R106 VPWR.n11 VPWR.t4 72.0127
R107 VPWR.n23 VPWR.n22 34.6358
R108 VPWR.n24 VPWR.n23 34.6358
R109 VPWR.n19 VPWR.n18 34.6358
R110 VPWR.n16 VPWR.n9 34.6358
R111 VPWR.n24 VPWR.n3 30.4946
R112 VPWR.n2 VPWR.t2 26.5955
R113 VPWR.n2 VPWR.t1 26.5955
R114 VPWR.n5 VPWR.t6 26.5955
R115 VPWR.n5 VPWR.t5 26.5955
R116 VPWR.n8 VPWR.t10 26.5955
R117 VPWR.n8 VPWR.t9 26.5955
R118 VPWR.n10 VPWR.t7 26.5955
R119 VPWR.n10 VPWR.t8 26.5955
R120 VPWR.n29 VPWR.n28 25.977
R121 VPWR.n31 VPWR.n30 19.9534
R122 VPWR.n30 VPWR.n29 18.4476
R123 VPWR.n28 VPWR.n3 12.424
R124 VPWR.n22 VPWR.n6 9.41227
R125 VPWR.n14 VPWR.n9 9.3005
R126 VPWR.n16 VPWR.n15 9.3005
R127 VPWR.n18 VPWR.n7 9.3005
R128 VPWR.n20 VPWR.n19 9.3005
R129 VPWR.n22 VPWR.n21 9.3005
R130 VPWR.n23 VPWR.n4 9.3005
R131 VPWR.n25 VPWR.n24 9.3005
R132 VPWR.n26 VPWR.n3 9.3005
R133 VPWR.n28 VPWR.n27 9.3005
R134 VPWR.n29 VPWR.n1 9.3005
R135 VPWR.n30 VPWR.n0 9.3005
R136 VPWR.n32 VPWR.n31 9.3005
R137 VPWR.n17 VPWR.n16 6.4005
R138 VPWR.n13 VPWR.n12 5.97266
R139 VPWR.n12 VPWR.n9 4.14168
R140 VPWR.n18 VPWR.n17 3.38874
R141 VPWR.n14 VPWR.n13 0.569425
R142 VPWR.n19 VPWR.n6 0.376971
R143 VPWR.n15 VPWR.n14 0.120292
R144 VPWR.n15 VPWR.n7 0.120292
R145 VPWR.n20 VPWR.n7 0.120292
R146 VPWR.n21 VPWR.n20 0.120292
R147 VPWR.n21 VPWR.n4 0.120292
R148 VPWR.n25 VPWR.n4 0.120292
R149 VPWR.n26 VPWR.n25 0.120292
R150 VPWR.n27 VPWR.n26 0.120292
R151 VPWR.n27 VPWR.n1 0.120292
R152 VPWR.n1 VPWR.n0 0.120292
R153 VPWR.n32 VPWR.n0 0.120292
R154 VPWR VPWR.n32 0.0213333
R155 VPB.t3 VPB.t6 556.386
R156 VPB.t13 VPB.t4 544.548
R157 VPB.t12 VPB.t13 260.437
R158 VPB.t5 VPB.t7 260.437
R159 VPB.t10 VPB.t9 248.599
R160 VPB.t4 VPB.t10 248.599
R161 VPB.t11 VPB.t12 248.599
R162 VPB.t8 VPB.t11 248.599
R163 VPB.t7 VPB.t8 248.599
R164 VPB.t6 VPB.t5 248.599
R165 VPB.t2 VPB.t3 248.599
R166 VPB.t1 VPB.t2 248.599
R167 VPB.t0 VPB.t1 248.599
R168 VPB VPB.t0 189.409
R169 A3.n5 A3.t0 237.787
R170 A3.n1 A3.t3 221.72
R171 A3.n2 A3 168.874
R172 A3.n4 A3.n0 152
R173 A3.n6 A3.n5 152
R174 A3.n1 A3.t2 149.421
R175 A3.n3 A3.t1 149.421
R176 A3.n5 A3.n4 64.2672
R177 A3.n3 A3.n2 51.7709
R178 A3.n2 A3.n1 23.2079
R179 A3.n6 A3.n0 20.946
R180 A3.n4 A3.n3 8.92643
R181 A3 A3.n6 4.07323
R182 A3 A3.n0 2.90959
R183 a_467_297.n1 a_467_297.t6 407.805
R184 a_467_297.n4 a_467_297.t3 402.368
R185 a_467_297.n1 a_467_297.n0 317.964
R186 a_467_297.n5 a_467_297.n2 317.964
R187 a_467_297.n7 a_467_297.n6 317.964
R188 a_467_297.n4 a_467_297.n3 286.329
R189 a_467_297.n6 a_467_297.n1 100.894
R190 a_467_297.n5 a_467_297.n4 94.7937
R191 a_467_297.n6 a_467_297.n5 64.7534
R192 a_467_297.n3 a_467_297.t2 30.5355
R193 a_467_297.n7 a_467_297.t9 30.5355
R194 a_467_297.n0 a_467_297.t7 26.5955
R195 a_467_297.n0 a_467_297.t0 26.5955
R196 a_467_297.n2 a_467_297.t8 26.5955
R197 a_467_297.n2 a_467_297.t5 26.5955
R198 a_467_297.n3 a_467_297.t4 26.5955
R199 a_467_297.t1 a_467_297.n7 26.5955
R200 a_1079_47.n1 a_1079_47.t3 329.805
R201 a_1079_47.t2 a_1079_47.n1 326.709
R202 a_1079_47.n1 a_1079_47.n0 185
R203 a_1079_47.n0 a_1079_47.t0 24.9236
R204 a_1079_47.n0 a_1079_47.t1 24.9236
R205 B1.n0 B1.t1 228.148
R206 B1.n1 B1.t2 212.081
R207 B1.n2 B1 162.615
R208 B1.n2 B1.t3 158.768
R209 B1 B1.n0 155.123
R210 B1.n5 B1.n4 152
R211 B1.n3 B1.t0 139.78
R212 B1.n1 B1.n0 45.2793
R213 B1.n3 B1.n2 42.3581
R214 B1 B1.n5 18.1078
R215 B1.n5 B1 10.6151
R216 B1.n4 B1.n3 7.30353
R217 B1.n4 B1.n1 4.38232
R218 VGND.n6 VGND.t2 282.817
R219 VGND.n15 VGND.t3 282.817
R220 VGND.n5 VGND.n4 206.198
R221 VGND.n13 VGND.n2 199.739
R222 VGND.n9 VGND.n8 198.898
R223 VGND.n9 VGND.n7 30.4946
R224 VGND.n8 VGND.t1 28.6159
R225 VGND.n13 VGND.n1 25.977
R226 VGND.n4 VGND.t7 24.9236
R227 VGND.n4 VGND.t0 24.9236
R228 VGND.n8 VGND.t5 24.9236
R229 VGND.n2 VGND.t4 24.9236
R230 VGND.n2 VGND.t6 24.9236
R231 VGND.n15 VGND.n14 19.9534
R232 VGND.n14 VGND.n13 18.4476
R233 VGND.n9 VGND.n1 12.424
R234 VGND.n6 VGND.n5 9.48347
R235 VGND.n16 VGND.n15 9.3005
R236 VGND.n7 VGND.n3 9.3005
R237 VGND.n10 VGND.n9 9.3005
R238 VGND.n11 VGND.n1 9.3005
R239 VGND.n13 VGND.n12 9.3005
R240 VGND.n14 VGND.n0 9.3005
R241 VGND.n7 VGND.n6 7.90638
R242 VGND.n5 VGND.n3 0.147195
R243 VGND.n10 VGND.n3 0.120292
R244 VGND.n11 VGND.n10 0.120292
R245 VGND.n12 VGND.n11 0.120292
R246 VGND.n12 VGND.n0 0.120292
R247 VGND.n16 VGND.n0 0.120292
R248 VGND VGND.n16 0.0213333
R249 A4.n0 A4.t0 221.72
R250 A4.n1 A4.t1 221.72
R251 A4.n3 A4.n2 152
R252 A4.n0 A4.t2 149.421
R253 A4.n1 A4.t3 149.421
R254 A4.n4 A4.n0 91.1642
R255 A4.n2 A4.n0 58.9116
R256 A4.n4 A4.n3 22.313
R257 A4.n2 A4.n1 16.0672
R258 A4 A4.n4 3.76428
R259 A4.n3 A4 0.582318
C0 A1 VGND 0.018238f
C1 A3 VPWR 0.041449f
C2 A2 VGND 0.01639f
C3 A4 VPWR 0.043098f
C4 VPB B1 0.08154f
C5 A3 VGND 0.021653f
C6 VPB A1 0.056459f
C7 VPWR X 0.321136f
C8 A4 VGND 0.038352f
C9 B1 A1 0.056952f
C10 VPB A2 0.056669f
C11 VPWR VGND 0.159079f
C12 VPB A3 0.086688f
C13 X VGND 0.215542f
C14 A1 A2 0.071049f
C15 VPB A4 0.081231f
C16 A1 A3 2.07e-19
C17 VPB VPWR 0.171447f
C18 VPB X 0.01188f
C19 A2 A3 0.060812f
C20 B1 VPWR 0.021266f
C21 B1 X 9.31e-19
C22 A1 VPWR 0.035154f
C23 VPB VGND 0.017301f
C24 A3 A4 0.063851f
C25 A2 VPWR 0.032986f
C26 B1 VGND 0.033992f
C27 VGND VNB 0.878051f
C28 X VNB 0.070454f
C29 VPWR VNB 0.733692f
C30 A4 VNB 0.250536f
C31 A3 VNB 0.225531f
C32 A2 VNB 0.183848f
C33 A1 VNB 0.183509f
C34 B1 VNB 0.224451f
C35 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_1 VGND VPWR A4 Y B1 A1 A2 A3 VPB VNB
X0 a_236_47.t1 A4.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.163425 ps=1.175 w=0.65 l=0.15
X1 a_428_47.t0 A2.t0 a_336_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_109_297.t1 A1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=2.74 as=0.2125 ps=1.425 w=1 l=0.15
X3 Y.t0 A1.t1 a_428_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.2405 pd=2.04 as=0.138125 ps=1.075 w=0.65 l=0.15
X4 a_336_47.t0 A3.t0 a_236_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5 VPWR.t3 A4.t1 a_109_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.2125 ps=1.425 w=1 l=0.15
X6 a_109_297.t3 B1.t0 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_297.t2 A3.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.205 ps=1.41 w=1 l=0.15
X8 VPWR.t0 A2.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.155 ps=1.31 w=1 l=0.15
X9 VGND.t0 B1.t1 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.163425 pd=1.175 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A4.n0 A4.t1 241.536
R1 A4.n0 A4.t0 169.237
R2 A4.n1 A4.n0 152
R3 A4.n1 A4 12.5798
R4 A4 A4.n1 2.42809
R5 VGND VGND.n0 192.315
R6 VGND.n0 VGND.t1 45.2313
R7 VGND.n0 VGND.t0 44.3082
R8 a_236_47.t0 a_236_47.t1 64.6159
R9 VNB.t1 VNB.t2 1808.41
R10 VNB.t3 VNB.t4 1637.54
R11 VNB.t2 VNB.t0 1423.95
R12 VNB.t0 VNB.t3 1310.03
R13 VNB VNB.t1 911.327
R14 A2.n0 A2.t1 241.536
R15 A2.n0 A2.t0 169.237
R16 A2.n1 A2.n0 152
R17 A2.n1 A2 11.4005
R18 A2 A2.n1 2.2005
R19 a_336_47.t0 a_336_47.t1 57.2313
R20 a_428_47.t0 a_428_47.t1 78.462
R21 A1.n0 A1.t0 230.363
R22 A1.n0 A1.t1 158.064
R23 A1.n1 A1.n0 152
R24 A1.n1 A1 11.9612
R25 A1 A1.n1 2.3087
R26 VPWR.n2 VPWR.n1 607.607
R27 VPWR.n2 VPWR.n0 607.341
R28 VPWR.n0 VPWR.t2 48.2655
R29 VPWR.n1 VPWR.t0 47.2805
R30 VPWR.n1 VPWR.t1 36.4455
R31 VPWR.n0 VPWR.t3 32.5055
R32 VPWR VPWR.n2 0.41385
R33 a_109_297.n1 a_109_297.t1 393.026
R34 a_109_297.n1 a_109_297.n0 372.457
R35 a_109_297.n2 a_109_297.n1 297.769
R36 a_109_297.n0 a_109_297.t3 42.3555
R37 a_109_297.n0 a_109_297.t4 41.3705
R38 a_109_297.n2 a_109_297.t2 32.5055
R39 a_109_297.t0 a_109_297.n2 28.5655
R40 VPB.t0 VPB.t1 340.344
R41 VPB.t3 VPB.t4 340.344
R42 VPB.t4 VPB.t2 331.464
R43 VPB.t2 VPB.t0 272.274
R44 VPB VPB.t3 189.409
R45 Y.n3 Y 593.216
R46 Y.n3 Y.n2 585
R47 Y.n4 Y.n3 585
R48 Y.n1 Y.t0 309.697
R49 Y.n0 Y.t1 209.923
R50 Y.n2 Y.n1 45.5116
R51 Y.n3 Y.t2 26.5955
R52 Y.n1 Y.n0 12.3125
R53 Y.n2 Y 5.92643
R54 Y.n5 Y.n4 5.92289
R55 Y.n4 Y 4.77662
R56 Y.n5 Y 2.84494
R57 Y Y.n5 2.29304
R58 Y.n0 Y 1.2554
R59 A3.n0 A3.t1 241.536
R60 A3.n0 A3.t0 169.237
R61 A3.n1 A3.n0 152
R62 A3.n1 A3 15.2005
R63 A3 A3.n1 2.93383
R64 B1.n0 B1.t0 233.869
R65 B1.n0 B1.t1 161.57
R66 B1 B1.n0 154.934
C0 Y VPWR 0.049972f
C1 A2 A1 0.06459f
C2 Y VPB 0.012692f
C3 Y VGND 0.309318f
C4 VPWR VPB 0.067175f
C5 Y B1 0.111147f
C6 VPWR VGND 0.065018f
C7 VPWR B1 0.016632f
C8 VGND VPB 0.005913f
C9 Y A4 0.035777f
C10 VPB B1 0.037807f
C11 Y A3 0.030276f
C12 VPWR A4 0.018759f
C13 VGND B1 0.01836f
C14 VPB A4 0.031191f
C15 Y A2 0.031025f
C16 VPWR A3 0.014953f
C17 VGND A4 0.012255f
C18 B1 A4 0.101079f
C19 VPB A3 0.029358f
C20 VGND A3 0.010546f
C21 VPWR A2 0.016694f
C22 Y A1 0.037013f
C23 VPB A2 0.030948f
C24 B1 A3 3.7e-19
C25 VGND A2 0.010567f
C26 VPWR A1 0.020081f
C27 VPB A1 0.0449f
C28 A4 A3 0.096005f
C29 VGND A1 0.013547f
C30 A3 A2 0.124345f
C31 VGND VNB 0.389126f
C32 VPWR VNB 0.328737f
C33 Y VNB 0.125749f
C34 A1 VNB 0.160735f
C35 A2 VNB 0.102814f
C36 A3 VNB 0.092102f
C37 A4 VNB 0.092396f
C38 B1 VNB 0.128523f
C39 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_2 VNB VPB VPWR VGND A4 A3 A2 A1 B1 Y
X0 a_149_297.t2 B1.t0 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_757_47.t2 A4.t0 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_757_47.t0 A3.t0 a_567_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t1 A3.t1 a_149_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.145 ps=1.29 w=1 l=0.15
X4 Y.t2 B1.t1 a_149_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 Y.t1 B1.t2 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_567_47.t1 A3.t2 a_757_47.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND.t2 A4.t1 a_757_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t7 A4.t2 a_149_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_149_297.t3 A4.t3 VPWR.t6 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_317_47.t2 A1.t0 Y.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_317_47.t3 A2.t0 a_567_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_149_297.t9 A3.t3 VPWR.t0 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X13 a_149_297.t0 A2.t1 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X14 Y.t4 A1.t1 a_317_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR.t4 A2.t2 a_149_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_567_47.t0 A2.t3 a_317_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_149_297.t8 A1.t2 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND.t0 B1.t3 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR.t3 A1.t3 a_149_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 B1.n0 B1.t0 228.148
R1 B1.n2 B1.t1 212.081
R2 B1 B1.n0 172.293
R3 B1.n3 B1.t2 161.69
R4 B1.n6 B1.n5 152
R5 B1.n3 B1.n1 152
R6 B1.n4 B1.t3 139.78
R7 B1.n2 B1.n0 45.2793
R8 B1.n4 B1.n3 39.4369
R9 B1.n6 B1.n1 21.2298
R10 B1.n5 B1.n4 10.2247
R11 B1.n1 B1 6.5566
R12 B1.n5 B1.n2 4.38232
R13 B1 B1.n6 0.937085
R14 Y.n4 Y.n3 369.356
R15 Y.n2 Y.n1 287.401
R16 Y.n2 Y.n0 201.941
R17 Y.n5 Y.n2 40.6593
R18 Y.n3 Y.t3 26.5955
R19 Y.n3 Y.t2 26.5955
R20 Y.n1 Y.t5 24.9236
R21 Y.n1 Y.t4 24.9236
R22 Y.n0 Y.t0 24.9236
R23 Y.n0 Y.t1 24.9236
R24 Y.n5 Y 21.8358
R25 Y.n4 Y 6.4005
R26 Y.n5 Y 6.4005
R27 Y Y.n5 3.76521
R28 Y Y.n4 0.753441
R29 a_149_297.n3 a_149_297.t3 407.805
R30 a_149_297.n6 a_149_297.t1 400.861
R31 a_149_297.n3 a_149_297.n2 317.964
R32 a_149_297.n4 a_149_297.n1 317.964
R33 a_149_297.n5 a_149_297.n0 317.964
R34 a_149_297.n7 a_149_297.n6 286.329
R35 a_149_297.n4 a_149_297.n3 100.894
R36 a_149_297.n6 a_149_297.n5 94.7937
R37 a_149_297.n5 a_149_297.n4 64.7534
R38 a_149_297.n1 a_149_297.t0 30.5355
R39 a_149_297.n2 a_149_297.t5 26.5955
R40 a_149_297.n2 a_149_297.t9 26.5955
R41 a_149_297.n1 a_149_297.t6 26.5955
R42 a_149_297.n0 a_149_297.t7 26.5955
R43 a_149_297.n0 a_149_297.t8 26.5955
R44 a_149_297.n7 a_149_297.t4 26.5955
R45 a_149_297.t2 a_149_297.n7 26.5955
R46 VPB VPB.t1 553.428
R47 VPB.t6 VPB.t9 544.548
R48 VPB.t0 VPB.t6 260.437
R49 VPB.t5 VPB.t3 248.599
R50 VPB.t9 VPB.t5 248.599
R51 VPB.t7 VPB.t0 248.599
R52 VPB.t8 VPB.t7 248.599
R53 VPB.t4 VPB.t8 248.599
R54 VPB.t2 VPB.t4 248.599
R55 VPB.t1 VPB.t2 248.599
R56 A4.n3 A4.t2 221.72
R57 A4.n1 A4.t3 218.507
R58 A4.n1 A4 209.466
R59 A4.n2 A4.n0 152
R60 A4.n5 A4.n4 152
R61 A4.n3 A4.t1 149.421
R62 A4.n1 A4.t0 146.208
R63 A4.n4 A4.n2 59.8965
R64 A4 A4.n0 17.1641
R65 A4.n5 A4 15.4187
R66 A4.n4 A4.n3 12.4968
R67 A4 A4.n5 10.1823
R68 A4 A4.n0 9.6005
R69 A4.n2 A4.n1 1.66257
R70 VGND.n5 VGND.t1 282.817
R71 VGND.n3 VGND.t0 281.974
R72 VGND.n2 VGND.n1 206.263
R73 VGND.n4 VGND.n3 25.224
R74 VGND.n1 VGND.t3 24.9236
R75 VGND.n1 VGND.t2 24.9236
R76 VGND.n5 VGND.n4 13.177
R77 VGND.n6 VGND.n5 9.3005
R78 VGND.n4 VGND.n0 9.3005
R79 VGND.n3 VGND.n2 6.77219
R80 VGND.n2 VGND.n0 0.160063
R81 VGND.n6 VGND.n0 0.120292
R82 VGND VGND.n6 0.0226354
R83 a_757_47.t2 a_757_47.n1 329.805
R84 a_757_47.n1 a_757_47.t3 326.709
R85 a_757_47.n1 a_757_47.n0 185
R86 a_757_47.n0 a_757_47.t1 24.9236
R87 a_757_47.n0 a_757_47.t0 24.9236
R88 VNB.t4 VNB.t8 2677.02
R89 VNB.t1 VNB.t5 2677.02
R90 VNB.t6 VNB.t7 1196.12
R91 VNB.t3 VNB.t6 1196.12
R92 VNB.t8 VNB.t3 1196.12
R93 VNB.t0 VNB.t4 1196.12
R94 VNB.t9 VNB.t0 1196.12
R95 VNB.t5 VNB.t9 1196.12
R96 VNB.t2 VNB.t1 1196.12
R97 VNB VNB.t2 1181.88
R98 A3.n3 A3.t1 237.787
R99 A3.n0 A3.t3 221.72
R100 A3.n3 A3 159.856
R101 A3 A3.n1 158.109
R102 A3.n5 A3.n4 152
R103 A3.n0 A3.t0 149.421
R104 A3.n2 A3.t2 149.421
R105 A3.n4 A3.n3 64.2672
R106 A3.n2 A3.n1 51.7709
R107 A3.n1 A3.n0 23.2079
R108 A3 A3.n5 13.6732
R109 A3.n5 A3 13.0914
R110 A3.n4 A3.n2 8.92643
R111 a_567_47.n1 a_567_47.n0 472.401
R112 a_567_47.n0 a_567_47.t3 24.9236
R113 a_567_47.n0 a_567_47.t0 24.9236
R114 a_567_47.t2 a_567_47.n1 24.9236
R115 a_567_47.n1 a_567_47.t1 24.9236
R116 VPWR.n8 VPWR.n5 315.728
R117 VPWR.n12 VPWR.n3 310.502
R118 VPWR.n1 VPWR.n0 310.5
R119 VPWR.n7 VPWR.n6 146.25
R120 VPWR.n6 VPWR.t1 77.8155
R121 VPWR.n6 VPWR.t0 73.8755
R122 VPWR.n0 VPWR.t5 26.5955
R123 VPWR.n0 VPWR.t3 26.5955
R124 VPWR.n3 VPWR.t2 26.5955
R125 VPWR.n3 VPWR.t4 26.5955
R126 VPWR.n5 VPWR.t6 26.5955
R127 VPWR.n5 VPWR.t7 26.5955
R128 VPWR.n11 VPWR.n4 25.1944
R129 VPWR.n12 VPWR.n11 23.7181
R130 VPWR.n13 VPWR.n12 20.7064
R131 VPWR.n13 VPWR.n1 17.6946
R132 VPWR.n8 VPWR.n7 11.0018
R133 VPWR.n9 VPWR.n4 9.3005
R134 VPWR.n11 VPWR.n10 9.3005
R135 VPWR.n12 VPWR.n2 9.3005
R136 VPWR.n14 VPWR.n13 9.3005
R137 VPWR.n15 VPWR.n1 7.29417
R138 VPWR.n7 VPWR.n4 2.58926
R139 VPWR.n9 VPWR.n8 0.612196
R140 VPWR VPWR.n15 0.472624
R141 VPWR.n15 VPWR.n14 0.151915
R142 VPWR.n10 VPWR.n9 0.120292
R143 VPWR.n10 VPWR.n2 0.120292
R144 VPWR.n14 VPWR.n2 0.120292
R145 A1.n0 A1.t2 212.081
R146 A1.n1 A1.t3 212.081
R147 A1.n0 A1.t0 139.78
R148 A1.n1 A1.t1 139.78
R149 A1 A1.n2 70.0171
R150 A1.n2 A1.n0 29.8769
R151 A1.n2 A1.n1 24.8667
R152 a_317_47.n0 a_317_47.t1 344.877
R153 a_317_47.n0 a_317_47.t3 326.709
R154 a_317_47.n1 a_317_47.n0 185
R155 a_317_47.n1 a_317_47.t0 24.9236
R156 a_317_47.t2 a_317_47.n1 24.9236
R157 A2.n0 A2.t1 221.72
R158 A2.n1 A2.t2 221.72
R159 A2.n0 A2.t0 149.421
R160 A2.n1 A2.t3 149.421
R161 A2 A2.n2 68.3105
R162 A2.n2 A2.n1 37.1543
R163 A2.n2 A2.n0 28.267
C0 VPB A4 0.082436f
C1 A1 A2 0.071049f
C2 VPB Y 0.027577f
C3 A1 A3 2.07e-19
C4 B1 Y 0.219817f
C5 VPB VPWR 0.12959f
C6 A2 A3 0.060812f
C7 A1 Y 0.04564f
C8 VPB VGND 0.015857f
C9 B1 VPWR 0.019169f
C10 A2 Y 5.21e-19
C11 B1 VGND 0.036803f
C12 A1 VPWR 0.04068f
C13 A3 A4 0.073985f
C14 A1 VGND 0.020431f
C15 A3 Y 2.59e-19
C16 A2 VPWR 0.041001f
C17 A4 Y 1.54e-19
C18 A2 VGND 0.021143f
C19 A3 VPWR 0.047888f
C20 VPB B1 0.084058f
C21 A4 VPWR 0.042665f
C22 A3 VGND 0.025776f
C23 VPB A1 0.056116f
C24 A4 VGND 0.038264f
C25 Y VPWR 0.029531f
C26 VPB A2 0.056669f
C27 B1 A1 0.060918f
C28 Y VGND 0.166597f
C29 VPB A3 0.086688f
C30 VPWR VGND 0.118217f
C31 VGND VNB 0.68764f
C32 VPWR VNB 0.556394f
C33 Y VNB 0.074661f
C34 A4 VNB 0.25588f
C35 A3 VNB 0.22404f
C36 A2 VNB 0.183848f
C37 A1 VNB 0.183054f
C38 B1 VNB 0.25051f
C39 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_4 VNB VPB VGND VPWR A4 A3 A2 A1 Y B1
X0 VPWR.t5 A1.t0 a_27_297# VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.29 ps=1.58 w=1 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.3375 ps=1.675 w=1 l=0.15
X2 Y.t7 A1.t1 a_493_47# VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t6 A1.t2 a_493_47# VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297# A1.t3 VPWR.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR.t6 A2.t0 a_27_297# VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1825 ps=1.365 w=1 l=0.15
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_911_47# A2.t1 a_493_47# VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B1.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.135 ps=1.27 w=1 l=0.15
X14 a_493_47# A1.t4 Y.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_493_47# A1.t5 Y.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_493_47# A2.t2 a_911_47# VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y.t1 B1.t1 a_27_297# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_27_297# B1.t2 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND.t1 B1.t3 Y.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND.t2 B1.t4 Y.t9 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_911_47# A2.t3 a_493_47# VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_27_297# A1.t6 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X27 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X28 Y.t10 B1.t5 VGND.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_27_297# A2.t4 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VPWR.t1 A2.t5 a_27_297# VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.3375 pd=1.675 as=0.135 ps=1.27 w=1 l=0.15
X31 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 Y.t11 B1.t6 a_27_297# VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 VPWR.t2 A1.t7 a_27_297# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 Y.t3 B1.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A1.n11 A1.t0 238.371
R1 A1.n1 A1.t6 212.081
R2 A1.n5 A1.t7 212.081
R3 A1.n0 A1.t3 212.081
R4 A1 A1.n2 159.758
R5 A1.n4 A1.n3 152
R6 A1.n7 A1.n6 152
R7 A1.n9 A1.n8 152
R8 A1.n12 A1.n11 152
R9 A1.n1 A1.t5 139.78
R10 A1.n5 A1.t2 139.78
R11 A1.n0 A1.t4 139.78
R12 A1.n10 A1.t1 139.78
R13 A1.n4 A1.n2 49.6611
R14 A1.n6 A1.n5 46.7399
R15 A1.n9 A1.n0 35.055
R16 A1.n10 A1.n9 26.2914
R17 A1.n11 A1.n10 23.3702
R18 A1.n6 A1.n0 14.6066
R19 A1.n8 A1.n7 13.1884
R20 A1.n3 A1 12.4126
R21 A1.n12 A1 9.30959
R22 A1.n2 A1.n1 8.76414
R23 A1 A1.n12 8.53383
R24 A1.n3 A1 5.4308
R25 A1.n8 A1 3.87929
R26 A1.n5 A1.n4 2.92171
R27 A1.n7 A1 0.776258
R28 VPWR.n13 VPWR.n12 585
R29 VPWR.n15 VPWR.n14 585
R30 VPWR.n3 VPWR.n2 310.502
R31 VPWR.n6 VPWR.n5 310.502
R32 VPWR.n4 VPWR.t1 218.392
R33 VPWR.n14 VPWR.n13 66.9805
R34 VPWR.n7 VPWR.n3 26.7299
R35 VPWR.n13 VPWR.t4 26.5955
R36 VPWR.n14 VPWR.t5 26.5955
R37 VPWR.n2 VPWR.t3 26.5955
R38 VPWR.n2 VPWR.t2 26.5955
R39 VPWR.n5 VPWR.t0 26.5955
R40 VPWR.n5 VPWR.t6 26.5955
R41 VPWR.n12 VPWR.n11 24.5464
R42 VPWR.n7 VPWR.n6 18.824
R43 VPWR.n11 VPWR.n3 17.6946
R44 VPWR.n16 VPWR.n15 10.8154
R45 VPWR.n8 VPWR.n7 9.3005
R46 VPWR.n9 VPWR.n3 9.3005
R47 VPWR.n11 VPWR.n10 9.3005
R48 VPWR.n1 VPWR.n0 9.3005
R49 VPWR.n15 VPWR.n1 7.44777
R50 VPWR.n6 VPWR.n4 6.86272
R51 VPWR VPWR.n16 0.574981
R52 VPWR.n8 VPWR.n4 0.490771
R53 VPWR.n12 VPWR.n1 0.465955
R54 VPWR.n16 VPWR.n0 0.147862
R55 VPWR.n9 VPWR.n8 0.120292
R56 VPWR.n10 VPWR.n9 0.120292
R57 VPWR.n10 VPWR.n0 0.120292
R58 VPB.t8 VPB.t7 449.844
R59 VPB.t0 VPB.t8 432.087
R60 VPB.t6 VPB.t9 304.829
R61 VPB.t3 VPB.t4 248.599
R62 VPB.t9 VPB.t3 248.599
R63 VPB.t5 VPB.t6 248.599
R64 VPB.t7 VPB.t5 248.599
R65 VPB.t1 VPB.t0 248.599
R66 VPB.t2 VPB.t1 248.599
R67 VPB.t10 VPB.t2 248.599
R68 VPB VPB.t10 142.056
R69 A2.n1 A2.n0 218.603
R70 A2.n9 A2.t4 205.654
R71 A2.n6 A2.t0 205.654
R72 A2.n3 A2.t5 203.435
R73 A2 A2.n1 155.048
R74 A2.n6 A2.t1 152.863
R75 A2.n16 A2.n15 152
R76 A2.n13 A2.n12 152
R77 A2.n11 A2.n10 152
R78 A2.n7 A2.n4 152
R79 A2.n14 A2.n2 144.601
R80 A2.n8 A2.t2 139.78
R81 A2.n5 A2.t3 139.78
R82 A2.n15 A2.n1 48.9199
R83 A2.n14 A2.n13 38.8483
R84 A2.n7 A2.n6 29.6091
R85 A2.n10 A2.n5 26.1662
R86 A2.n11 A2.n4 20.7243
R87 A2.n10 A2.n9 18.5919
R88 A2 A2.n16 17.6767
R89 A2.n12 A2 17.6767
R90 A2.n8 A2.n7 15.1491
R91 A2.n9 A2.n8 13.0834
R92 A2.n5 A2.n3 12.2524
R93 A2.n16 A2 10.3624
R94 A2.n12 A2 10.3624
R95 A2.n15 A2.n14 10.0721
R96 A2.n13 A2.n3 7.82251
R97 A2.n4 A2 4.26717
R98 A2 A2.n11 3.04812
R99 Y.n2 Y.n0 333.786
R100 Y.n2 Y.n1 295.712
R101 Y.n5 Y.n4 264.435
R102 Y.n8 Y.n6 248.248
R103 Y.n5 Y.n3 198.177
R104 Y.n8 Y.n7 185
R105 Y.n9 Y.n8 64.377
R106 Y.n9 Y.n5 31.2476
R107 Y Y.n2 27.9536
R108 Y.n0 Y.t2 26.5955
R109 Y.n0 Y.t11 26.5955
R110 Y.n1 Y.t0 26.5955
R111 Y.n1 Y.t1 26.5955
R112 Y.n7 Y.t5 24.9236
R113 Y.n7 Y.t7 24.9236
R114 Y.n6 Y.t4 24.9236
R115 Y.n6 Y.t6 24.9236
R116 Y.n4 Y.t8 24.9236
R117 Y.n4 Y.t3 24.9236
R118 Y.n3 Y.t9 24.9236
R119 Y.n3 Y.t10 24.9236
R120 Y Y.n9 2.61868
R121 VNB.t9 VNB.t4 3047.25
R122 VNB.t6 VNB.t5 1196.12
R123 VNB.t7 VNB.t6 1196.12
R124 VNB.t1 VNB.t7 1196.12
R125 VNB.t3 VNB.t1 1196.12
R126 VNB.t2 VNB.t3 1196.12
R127 VNB.t4 VNB.t2 1196.12
R128 VNB.t10 VNB.t9 1196.12
R129 VNB.t8 VNB.t10 1196.12
R130 VNB.t0 VNB.t8 1196.12
R131 VNB VNB.t0 683.495
R132 A4.n2 A4.n0 212.081
R133 A4.n17 A4.n3 212.081
R134 A4.n8 A4.n6 212.081
R135 A4.n11 A4.n9 212.081
R136 A4 A4.n2 182.694
R137 A4.n19 A4.n18 152
R138 A4.n16 A4.n15 152
R139 A4.n14 A4.n5 152
R140 A4.n13 A4.n12 152
R141 A4.n2 A4.n1 139.78
R142 A4.n17 A4.n4 139.78
R143 A4.n8 A4.n7 139.78
R144 A4.n11 A4.n10 139.78
R145 A4.n16 A4.n5 49.6611
R146 A4.n12 A4.n8 48.2005
R147 A4.n18 A4.n17 39.4369
R148 A4.n18 A4.n2 21.9096
R149 A4.n14 A4.n13 21.2298
R150 A4 A4.n19 20.6054
R151 A4.n15 A4 15.6103
R152 A4.n12 A4.n11 13.146
R153 A4.n15 A4 13.1127
R154 A4.n17 A4.n16 10.2247
R155 A4.n19 A4 8.11757
R156 A4 A4.n14 5.62001
R157 A4.n13 A4 1.87367
R158 A4.n8 A4.n5 1.46111
R159 A3.n7 A3.n5 205.654
R160 A3.n15 A3.n8 205.654
R161 A3.n12 A3.n10 205.654
R162 A3.n2 A3.n0 205.654
R163 A3 A3.n3 168.499
R164 A3.n18 A3.n17 152
R165 A3.n16 A3.n4 152
R166 A3.n14 A3.n13 152
R167 A3.n2 A3.n1 144.601
R168 A3.n7 A3.n6 139.78
R169 A3.n15 A3.n9 139.78
R170 A3.n12 A3.n11 139.78
R171 A3.n17 A3.n16 46.8234
R172 A3.n15 A3.n14 45.4462
R173 A3.n7 A3.n3 38.3858
R174 A3.n3 A3.n2 21.5826
R175 A3.n18 A3.n4 19.3427
R176 A3.n13 A3 15.3605
R177 A3.n14 A3.n12 12.3948
R178 A3.n13 A3 10.8094
R179 A3.n17 A3.n7 9.6405
R180 A3 A3.n4 3.98272
R181 A3 A3.n18 2.84494
R182 A3.n16 A3.n15 1.37764
R183 VGND.n1 VGND.t2 287.877
R184 VGND.n5 VGND.t0 282.596
R185 VGND.n3 VGND.n2 199.739
R186 VGND.n2 VGND.t3 24.9236
R187 VGND.n2 VGND.t1 24.9236
R188 VGND.n5 VGND.n4 19.9534
R189 VGND.n4 VGND.n3 18.4476
R190 VGND VGND.n5 9.3005
R191 VGND.n4 VGND.n0 9.3005
R192 VGND.n3 VGND.n1 6.66294
R193 VGND.n1 VGND.n0 0.687401
R194 VGND VGND.n0 0.120292
R195 B1.n2 B1.t0 212.081
R196 B1.n3 B1.t1 212.081
R197 B1.n8 B1.t2 212.081
R198 B1.n10 B1.t6 212.081
R199 B1.n11 B1.n10 183.731
R200 B1.n5 B1.n4 152
R201 B1.n7 B1.n6 152
R202 B1.n9 B1.n0 152
R203 B1.n2 B1.t4 139.78
R204 B1.n3 B1.t5 139.78
R205 B1.n8 B1.t3 139.78
R206 B1.n10 B1.t7 139.78
R207 B1.n3 B1.n2 61.346
R208 B1.n7 B1.n4 49.6611
R209 B1.n9 B1.n8 40.8975
R210 B1.n10 B1.n9 20.449
R211 B1.n6 B1.n0 18.9222
R212 B1 B1.n11 18.644
R213 B1.n5 B1 13.0788
R214 B1 B1.n5 12.5222
R215 B1.n8 B1.n7 8.76414
R216 B1.n1 B1 8.14595
R217 B1.n6 B1 6.4005
R218 B1.n1 B1 3.89615
R219 B1.n11 B1.n1 3.06137
R220 B1.n4 B1.n3 2.92171
R221 B1 B1.n0 0.278761
C0 a_911_47# A2 0.142014f
C1 a_27_297# A4 0.158745f
C2 a_1269_47# A1 8.47e-20
C3 A2 VGND 0.037703f
C4 A4 Y 9.99e-20
C5 A3 VPWR 0.071877f
C6 VPB B1 0.14505f
C7 a_911_47# A3 0.110107f
C8 a_1269_47# A2 2.35e-19
C9 a_27_297# Y 0.152142f
C10 A4 VPWR 0.084642f
C11 A3 VGND 0.034794f
C12 a_27_297# a_493_47# 0.005466f
C13 a_27_297# VPWR 1.53981f
C14 a_1269_47# A3 0.0336f
C15 a_493_47# Y 0.151685f
C16 VPB A1 0.146413f
C17 A4 VGND 0.069216f
C18 Y VPWR 0.027873f
C19 a_27_297# a_911_47# 0.007284f
C20 a_911_47# Y 0.006967f
C21 B1 A1 0.021277f
C22 a_1269_47# A4 0.154691f
C23 VPB A2 0.150571f
C24 a_493_47# VPWR 0.005481f
C25 a_27_297# VGND 0.028314f
C26 Y VGND 0.251739f
C27 a_27_297# a_1269_47# 0.009832f
C28 a_493_47# a_911_47# 0.150099f
C29 VPB A3 0.115091f
C30 a_911_47# VPWR 0.00522f
C31 a_493_47# VGND 0.3576f
C32 a_1269_47# Y 8.97e-19
C33 VPWR VGND 0.200731f
C34 a_493_47# a_1269_47# 0.013638f
C35 a_1269_47# VPWR 0.006104f
C36 A1 A2 0.066878f
C37 a_911_47# VGND 0.038207f
C38 VPB A4 0.133468f
C39 a_911_47# a_1269_47# 0.165068f
C40 a_27_297# VPB 0.031432f
C41 VPB Y 0.012116f
C42 A1 A3 4.22e-19
C43 a_1269_47# VGND 0.409386f
C44 a_493_47# VPB 1.17e-19
C45 a_27_297# B1 0.062658f
C46 A1 A4 1.24e-19
C47 VPB VPWR 0.184147f
C48 A2 A3 0.05314f
C49 B1 Y 0.317445f
C50 a_911_47# VPB 7.1e-19
C51 a_27_297# A1 0.151459f
C52 A1 Y 0.182736f
C53 VPB VGND 0.014414f
C54 B1 VPWR 0.039633f
C55 a_1269_47# VPB 7.54e-19
C56 a_493_47# A1 0.03619f
C57 a_27_297# A2 0.177699f
C58 A2 Y 0.001388f
C59 A1 VPWR 0.081569f
C60 A3 A4 0.063165f
C61 B1 VGND 0.087659f
C62 a_27_297# A3 0.144626f
C63 a_1269_47# B1 8.46e-21
C64 a_911_47# A1 7.39e-19
C65 a_493_47# A2 0.031821f
C66 A1 VGND 0.04278f
C67 A2 VPWR 0.086738f
C68 A3 Y 2.17e-19
C69 VGND VNB 1.09345f
C70 VPWR VNB 0.889292f
C71 Y VNB 0.057605f
C72 A4 VNB 0.417773f
C73 A3 VNB 0.36098f
C74 A2 VNB 0.409537f
C75 A1 VNB 0.397611f
C76 B1 VNB 0.452916f
C77 VPB VNB 2.0223f
C78 a_1269_47# VNB 0.039686f
C79 a_911_47# VNB 0.015187f
C80 a_493_47# VNB 0.016496f
C81 a_27_297# VNB 0.074581f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221o_4 VNB VPB VPWR VGND A2 X A1 C1 B1 B2
X0 VGND.t6 A2.t0 a_445_47.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t9 B2.t0 a_1053_47.t2 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21.t7 A1.t0 a_445_47.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_445_297# A2.t1 VPWR.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_804_297# C1.t0 a_79_21.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_297# B1.t0 a_804_297# VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t1 a_79_21.t8 X.t7 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1053_47.t1 B2.t1 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_79_21.t3 C1.t1 a_804_297# VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10 a_1053_47.t3 B1.t1 a_79_21.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X.t6 a_79_21.t9 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47.t0 A1.t1 a_79_21.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND.t7 C1.t2 a_79_21.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t3 a_79_21.t10 X.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND.t1 a_79_21.t11 X.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t2 a_79_21.t12 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21.t4 B1.t2 a_1053_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_79_21.t0 C1.t3 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.345 ps=1.69 w=1 l=0.15
X21 X.t1 a_79_21.t13 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_445_47.t1 A2.t2 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_445_297# A1.t2 VPWR.t7 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t4 A2.t3 a_445_297# VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR.t6 A1.t3 a_445_297# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X26 X.t4 a_79_21.t14 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X.t0 a_79_21.t15 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t3 212.081
R1 A2.n1 A2.t1 212.081
R2 A2 A2.n2 153.696
R3 A2.n0 A2.t0 139.78
R4 A2.n1 A2.t2 139.78
R5 A2.n2 A2.n1 40.8975
R6 A2.n2 A2.n0 20.449
R7 a_445_47.n1 a_445_47.n0 323.851
R8 a_445_47.n0 a_445_47.t2 24.9236
R9 a_445_47.n0 a_445_47.t1 24.9236
R10 a_445_47.n1 a_445_47.t3 24.9236
R11 a_445_47.t0 a_445_47.n1 24.9236
R12 VGND.n16 VGND.t6 312.026
R13 VGND.n27 VGND.t4 286.426
R14 VGND.n8 VGND.n7 218.636
R15 VGND.n9 VGND.n6 207.965
R16 VGND.n19 VGND.n18 207.965
R17 VGND.n25 VGND.n1 207.965
R18 VGND.n11 VGND.n10 34.6358
R19 VGND.n11 VGND.n4 34.6358
R20 VGND.n15 VGND.n4 34.6358
R21 VGND.n20 VGND.n17 34.6358
R22 VGND.n24 VGND.n2 34.6358
R23 VGND.n27 VGND.n26 32.377
R24 VGND.n26 VGND.n25 30.8711
R25 VGND.n9 VGND.n8 27.9238
R26 VGND.n7 VGND.t8 24.9236
R27 VGND.n7 VGND.t9 24.9236
R28 VGND.n6 VGND.t0 24.9236
R29 VGND.n6 VGND.t7 24.9236
R30 VGND.n18 VGND.t5 24.9236
R31 VGND.n18 VGND.t2 24.9236
R32 VGND.n1 VGND.t3 24.9236
R33 VGND.n1 VGND.t1 24.9236
R34 VGND.n19 VGND.n2 24.8476
R35 VGND.n17 VGND.n16 18.824
R36 VGND.n16 VGND.n15 15.8123
R37 VGND.n10 VGND.n9 14.3064
R38 VGND.n28 VGND.n27 11.5593
R39 VGND.n20 VGND.n19 9.78874
R40 VGND.n10 VGND.n5 9.3005
R41 VGND.n12 VGND.n11 9.3005
R42 VGND.n13 VGND.n4 9.3005
R43 VGND.n15 VGND.n14 9.3005
R44 VGND.n17 VGND.n3 9.3005
R45 VGND.n21 VGND.n20 9.3005
R46 VGND.n22 VGND.n2 9.3005
R47 VGND.n24 VGND.n23 9.3005
R48 VGND.n26 VGND.n0 9.3005
R49 VGND.n25 VGND.n24 3.76521
R50 VGND.n8 VGND.n5 0.15388
R51 VGND.n12 VGND.n5 0.120292
R52 VGND.n13 VGND.n12 0.120292
R53 VGND.n14 VGND.n13 0.120292
R54 VGND.n14 VGND.n3 0.120292
R55 VGND.n21 VGND.n3 0.120292
R56 VGND.n22 VGND.n21 0.120292
R57 VGND.n23 VGND.n22 0.120292
R58 VGND.n23 VGND.n0 0.120292
R59 VGND.n28 VGND.n0 0.120292
R60 VGND VGND.n28 0.0200312
R61 VNB.t0 VNB.t13 2677.02
R62 VNB.t9 VNB.t6 2677.02
R63 VNB.t13 VNB.t12 1196.12
R64 VNB.t7 VNB.t0 1196.12
R65 VNB.t1 VNB.t7 1196.12
R66 VNB.t10 VNB.t1 1196.12
R67 VNB.t11 VNB.t10 1196.12
R68 VNB.t6 VNB.t11 1196.12
R69 VNB.t8 VNB.t9 1196.12
R70 VNB.t3 VNB.t8 1196.12
R71 VNB.t4 VNB.t3 1196.12
R72 VNB.t2 VNB.t4 1196.12
R73 VNB.t5 VNB.t2 1196.12
R74 VNB VNB.t5 897.087
R75 B2.n5 B2.n4 218.654
R76 B2.n1 B2.n0 212.081
R77 B2 B2.n2 168.153
R78 B2 B2.n5 156.571
R79 B2.n1 B2.t1 152.925
R80 B2.n3 B2.t0 139.78
R81 B2.n3 B2.n2 43.0884
R82 B2.n5 B2.n3 6.57323
R83 B2.n2 B2.n1 5.11262
R84 a_1053_47.t2 a_1053_47.n1 268.077
R85 a_1053_47.n1 a_1053_47.n0 231.278
R86 a_1053_47.n1 a_1053_47.t1 182.636
R87 a_1053_47.n0 a_1053_47.t0 24.9236
R88 a_1053_47.n0 a_1053_47.t3 24.9236
R89 B1.n1 B1.n0 212.081
R90 B1.n3 B1.t0 212.081
R91 B1.n5 B1.n1 209.239
R92 B1.n5 B1.n4 152
R93 B1.n3 B1.t1 141.385
R94 B1.n2 B1.t2 139.78
R95 B1.n4 B1.n3 48.2005
R96 B1 B1.n5 17.3719
R97 B1.n4 B1.n2 11.6853
R98 B1.n2 B1.n1 1.46111
R99 VPB.t5 VPB.t9 559.346
R100 VPB.t1 VPB.t5 251.559
R101 VPB.t4 VPB.t10 248.599
R102 VPB.t9 VPB.t4 248.599
R103 VPB.t2 VPB.t1 248.599
R104 VPB.t3 VPB.t2 248.599
R105 VPB.t6 VPB.t3 248.599
R106 VPB.t7 VPB.t6 248.599
R107 VPB.t8 VPB.t7 248.599
R108 VPB.t0 VPB.t8 248.599
R109 VPB VPB.t0 186.45
R110 A1.n3 A1.t2 216.463
R111 A1.n2 A1.t3 212.081
R112 A1 A1.n0 154.133
R113 A1.n4 A1.n3 152
R114 A1.n0 A1.t0 147.814
R115 A1.n1 A1.t1 139.78
R116 A1.n3 A1.n2 57.6944
R117 A1 A1.n4 55.264
R118 A1.n1 A1.n0 53.3126
R119 A1.n2 A1.n1 13.8763
R120 A1.n4 A1 6.4005
R121 a_79_21.n14 a_79_21.n13 585
R122 a_79_21.n1 a_79_21.t6 328.623
R123 a_79_21.n16 a_79_21.t4 321.599
R124 a_79_21.n14 a_79_21.n12 223.462
R125 a_79_21.n3 a_79_21.t8 212.081
R126 a_79_21.n9 a_79_21.t9 212.081
R127 a_79_21.n4 a_79_21.t10 212.081
R128 a_79_21.n5 a_79_21.t14 212.081
R129 a_79_21.n7 a_79_21.n6 172.725
R130 a_79_21.n8 a_79_21.n7 152
R131 a_79_21.n10 a_79_21.n2 152
R132 a_79_21.n12 a_79_21.n11 152
R133 a_79_21.n3 a_79_21.t12 139.78
R134 a_79_21.n9 a_79_21.t13 139.78
R135 a_79_21.n4 a_79_21.t11 139.78
R136 a_79_21.n5 a_79_21.t15 139.78
R137 a_79_21.n1 a_79_21.n0 88.3446
R138 a_79_21.n17 a_79_21.n16 88.3446
R139 a_79_21.n15 a_79_21.n14 72.9153
R140 a_79_21.n11 a_79_21.n10 49.6611
R141 a_79_21.n15 a_79_21.n1 48.9326
R142 a_79_21.n9 a_79_21.n8 45.2793
R143 a_79_21.n6 a_79_21.n4 33.5944
R144 a_79_21.n6 a_79_21.n5 27.752
R145 a_79_21.n13 a_79_21.t1 26.5955
R146 a_79_21.n13 a_79_21.t3 26.5955
R147 a_79_21.n0 a_79_21.t2 24.9236
R148 a_79_21.n0 a_79_21.t7 24.9236
R149 a_79_21.t5 a_79_21.n17 24.9236
R150 a_79_21.n17 a_79_21.t0 24.9236
R151 a_79_21.n12 a_79_21.n2 20.7243
R152 a_79_21.n7 a_79_21.n2 20.7243
R153 a_79_21.n8 a_79_21.n4 16.0672
R154 a_79_21.n16 a_79_21.n15 12.6659
R155 a_79_21.n11 a_79_21.n3 7.30353
R156 a_79_21.n10 a_79_21.n9 4.38232
R157 VPWR.n7 VPWR.t6 851.475
R158 VPWR.n8 VPWR.n6 606.505
R159 VPWR.n16 VPWR.t2 347.125
R160 VPWR.n14 VPWR.n2 318.293
R161 VPWR.n4 VPWR.n3 318.293
R162 VPWR.n10 VPWR.n9 34.6358
R163 VPWR.n14 VPWR.n13 28.9887
R164 VPWR.n2 VPWR.t0 26.5955
R165 VPWR.n2 VPWR.t3 26.5955
R166 VPWR.n3 VPWR.t5 26.5955
R167 VPWR.n3 VPWR.t1 26.5955
R168 VPWR.n6 VPWR.t7 26.5955
R169 VPWR.n6 VPWR.t4 26.5955
R170 VPWR.n16 VPWR.n15 22.9652
R171 VPWR.n15 VPWR.n14 21.4593
R172 VPWR.n13 VPWR.n4 15.4358
R173 VPWR.n8 VPWR.n7 12.9467
R174 VPWR.n9 VPWR.n8 9.41227
R175 VPWR.n9 VPWR.n5 9.3005
R176 VPWR.n11 VPWR.n10 9.3005
R177 VPWR.n13 VPWR.n12 9.3005
R178 VPWR.n14 VPWR.n1 9.3005
R179 VPWR.n15 VPWR.n0 9.3005
R180 VPWR.n17 VPWR.n16 9.3005
R181 VPWR.n7 VPWR.n5 1.16999
R182 VPWR.n10 VPWR.n4 0.376971
R183 VPWR.n11 VPWR.n5 0.120292
R184 VPWR.n12 VPWR.n11 0.120292
R185 VPWR.n12 VPWR.n1 0.120292
R186 VPWR.n1 VPWR.n0 0.120292
R187 VPWR.n17 VPWR.n0 0.120292
R188 VPWR VPWR.n17 0.0200312
R189 C1.n0 C1.t0 213.738
R190 C1.n1 C1.t1 212.081
R191 C1 C1.n2 164.495
R192 C1.n1 C1.t2 141.375
R193 C1.n0 C1.t3 139.78
R194 C1.n2 C1.n0 35.055
R195 C1.n2 C1.n1 24.8308
R196 X.n5 X.n3 252.931
R197 X.n5 X.n4 208.508
R198 X.n2 X.n0 135.249
R199 X.n2 X.n1 98.982
R200 X X.n5 41.5268
R201 X.n3 X.t7 26.5955
R202 X.n3 X.t6 26.5955
R203 X.n4 X.t5 26.5955
R204 X.n4 X.t4 26.5955
R205 X.n1 X.t3 24.9236
R206 X.n1 X.t0 24.9236
R207 X.n0 X.t2 24.9236
R208 X.n0 X.t1 24.9236
R209 X.n6 X 15.8614
R210 X.n6 X.n2 14.5003
R211 X X.n6 3.06137
C0 a_445_297# VPWR 0.313956f
C1 VPB A2 0.05105f
C2 a_804_297# B2 0.045446f
C3 B1 VGND 0.020198f
C4 a_445_297# a_804_297# 0.341601f
C5 a_804_297# VPWR 0.399874f
C6 a_445_297# X 0.001866f
C7 VPB A1 0.088024f
C8 B2 VGND 0.031133f
C9 VPWR X 0.363863f
C10 a_445_297# VGND 0.006265f
C11 VPB C1 0.056945f
C12 A2 A1 0.064385f
C13 a_804_297# X 2.14e-19
C14 VPWR VGND 0.120854f
C15 a_804_297# VGND 0.008782f
C16 VPB B1 0.073126f
C17 X VGND 0.259694f
C18 VPB B2 0.071336f
C19 A1 C1 0.061904f
C20 a_445_297# VPB 0.016886f
C21 VPB VPWR 0.164277f
C22 a_445_297# A2 0.021453f
C23 a_804_297# VPB 0.0196f
C24 A2 VPWR 0.031225f
C25 C1 B1 0.051191f
C26 VPB X 0.012018f
C27 a_445_297# A1 0.0302f
C28 VPB VGND 0.016447f
C29 A2 X 0.002269f
C30 A1 VPWR 0.029855f
C31 a_804_297# A1 2.37e-19
C32 a_445_297# C1 0.015566f
C33 A2 VGND 0.025311f
C34 C1 VPWR 0.01418f
C35 A1 X 5.46e-19
C36 B1 B2 0.043529f
C37 a_804_297# C1 0.013885f
C38 a_445_297# B1 0.097823f
C39 A1 VGND 0.024175f
C40 C1 X 1.38e-19
C41 B1 VPWR 0.016448f
C42 a_804_297# B1 0.020229f
C43 a_445_297# B2 0.068285f
C44 B1 X 1.48e-20
C45 B2 VPWR 0.019885f
C46 C1 VGND 0.022059f
C47 VGND VNB 0.893778f
C48 X VNB 0.057158f
C49 VPWR VNB 0.733285f
C50 B2 VNB 0.22413f
C51 B1 VNB 0.208694f
C52 C1 VNB 0.168443f
C53 A1 VNB 0.238525f
C54 A2 VNB 0.171429f
C55 VPB VNB 1.57932f
C56 a_804_297# VNB 0.02012f
C57 a_445_297# VNB 0.009773f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221o_2 VPWR VGND VPB VNB C1 B2 B1 A1 A2 X
X0 VPWR.t1 a_27_47.t4 X.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47.t1 A1.t0 a_27_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X.t1 a_27_47.t5 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X3 a_109_297.t0 B1.t0 a_193_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297.t1 B2.t0 a_109_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X.t3 a_27_47.t6 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X6 a_205_47.t0 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR.t3 A2.t0 a_193_297.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297.t3 A1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47.t1 B1.t1 a_205_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X10 VGND.t1 a_27_47.t7 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297.t2 C1.t0 a_27_47.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND.t3 C1.t1 a_27_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND.t4 A2.t1 a_465_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
R0 a_27_47.t3 a_27_47.n4 669.389
R1 a_27_47.n0 a_27_47.t2 326.493
R2 a_27_47.n0 a_27_47.t1 249.615
R3 a_27_47.n1 a_27_47.t0 249.615
R4 a_27_47.n2 a_27_47.t4 212.081
R5 a_27_47.n3 a_27_47.t5 212.081
R6 a_27_47.n4 a_27_47.n3 158.573
R7 a_27_47.n2 a_27_47.t7 139.78
R8 a_27_47.n3 a_27_47.t6 139.78
R9 a_27_47.n4 a_27_47.n1 108.529
R10 a_27_47.n3 a_27_47.n2 61.346
R11 a_27_47.n1 a_27_47.n0 26.6245
R12 X.n0 X 593.784
R13 X.n1 X.n0 585
R14 X X.n2 185.251
R15 X.n3 X.n1 98.9003
R16 X.n0 X.t2 26.5955
R17 X.n0 X.t1 26.5955
R18 X.n2 X.t0 24.9236
R19 X.n2 X.t3 24.9236
R20 X X.n3 11.0708
R21 X.n1 X 8.28285
R22 X.n3 X 8.03187
R23 VPWR.n7 VPWR.t2 838.817
R24 VPWR.n5 VPWR.n3 312.053
R25 VPWR.n4 VPWR.t1 271.707
R26 VPWR.n13 VPWR 37.9123
R27 VPWR.n3 VPWR.t3 35.4605
R28 VPWR.n11 VPWR.n1 34.6358
R29 VPWR.n12 VPWR.n11 34.6358
R30 VPWR.n3 VPWR.t0 26.5955
R31 VPWR.n7 VPWR.n6 22.5887
R32 VPWR.n6 VPWR.n5 21.8358
R33 VPWR.n7 VPWR.n1 19.9534
R34 VPWR.n6 VPWR.n2 9.3005
R35 VPWR.n8 VPWR.n7 9.3005
R36 VPWR.n9 VPWR.n1 9.3005
R37 VPWR.n11 VPWR.n10 9.3005
R38 VPWR.n12 VPWR.n0 9.3005
R39 VPWR.n5 VPWR.n4 6.46279
R40 VPWR VPWR.n12 6.02403
R41 VPWR.n4 VPWR.n2 0.77975
R42 VPWR.n8 VPWR.n2 0.120292
R43 VPWR.n9 VPWR.n8 0.120292
R44 VPWR.n10 VPWR.n9 0.120292
R45 VPWR.n10 VPWR.n0 0.120292
R46 VPWR.n13 VPWR.n0 0.120292
R47 VPWR VPWR.n13 0.0213333
R48 VPB.t4 VPB.t3 556.386
R49 VPB.t3 VPB.t5 284.113
R50 VPB.t5 VPB.t0 275.235
R51 VPB.t0 VPB.t1 248.599
R52 VPB.t2 VPB.t4 248.599
R53 VPB.t6 VPB.t2 248.599
R54 VPB VPB.t6 189.409
R55 A1.n0 A1.t1 236.552
R56 A1.n0 A1.t0 164.251
R57 A1 A1.n0 154.47
R58 a_465_47.t0 a_465_47.t1 60.9236
R59 VNB.t3 VNB.t6 2677.02
R60 VNB.t6 VNB.t5 1366.99
R61 VNB.t4 VNB.t0 1366.99
R62 VNB.t5 VNB.t2 1324.27
R63 VNB.t2 VNB.t1 1196.12
R64 VNB.t0 VNB.t3 1025.24
R65 VNB VNB.t4 911.327
R66 B1.n0 B1.t0 239.505
R67 B1.n0 B1.t1 167.204
R68 B1 B1.n0 157.12
R69 a_193_297.n1 a_193_297.n0 953.038
R70 a_193_297.n0 a_193_297.t2 33.4905
R71 a_193_297.n0 a_193_297.t3 31.5205
R72 a_193_297.t0 a_193_297.n1 26.5955
R73 a_193_297.n1 a_193_297.t1 26.5955
R74 a_109_297.t0 a_109_297.n0 1201.3
R75 a_109_297.n0 a_109_297.t1 26.5955
R76 a_109_297.n0 a_109_297.t2 26.5955
R77 B2.n0 B2.t0 241.536
R78 B2 B2.n0 169.921
R79 B2.n0 B2.t1 169.237
R80 VGND.n12 VGND.n11 202.067
R81 VGND.n4 VGND.n3 200.516
R82 VGND.n2 VGND.t1 159.859
R83 VGND.n11 VGND.t0 36.0005
R84 VGND.n5 VGND.n1 34.6358
R85 VGND.n9 VGND.n1 34.6358
R86 VGND.n10 VGND.n9 34.6358
R87 VGND.n3 VGND.t2 33.2313
R88 VGND.n11 VGND.t3 24.9236
R89 VGND.n3 VGND.t4 24.9236
R90 VGND.n12 VGND.n10 22.9652
R91 VGND.n5 VGND.n4 18.4476
R92 VGND.n6 VGND.n5 9.3005
R93 VGND.n7 VGND.n1 9.3005
R94 VGND.n9 VGND.n8 9.3005
R95 VGND.n10 VGND.n0 9.3005
R96 VGND.n13 VGND.n12 7.12063
R97 VGND.n4 VGND.n2 6.68604
R98 VGND.n12 VGND 3.29747
R99 VGND.n6 VGND.n2 0.727919
R100 VGND.n13 VGND.n0 0.148519
R101 VGND.n7 VGND.n6 0.120292
R102 VGND.n8 VGND.n7 0.120292
R103 VGND.n8 VGND.n0 0.120292
R104 VGND VGND.n13 0.11354
R105 a_205_47.t0 a_205_47.t1 38.7697
R106 A2.n0 A2.t0 241.536
R107 A2.n0 A2.t1 169.237
R108 A2 A2.n0 164.8
R109 C1.n0 C1.t0 231.718
R110 C1 C1.n0 159.619
R111 C1.n0 C1.t1 159.417
C0 B2 B1 0.078429f
C1 VPB A2 0.026961f
C2 C1 A1 1.77e-20
C3 C1 A2 9.03e-21
C4 VPB VPWR 0.094135f
C5 B1 A1 0.060935f
C6 C1 VPWR 0.014042f
C7 VPB X 0.004228f
C8 B2 VPWR 0.00842f
C9 VPB VGND 0.010276f
C10 C1 X 5.03e-20
C11 B2 X 6.77e-20
C12 C1 VGND 0.019751f
C13 B1 VPWR 0.009818f
C14 A1 A2 0.069236f
C15 A1 VPWR 0.01613f
C16 B1 X 9.58e-20
C17 B2 VGND 0.017443f
C18 A1 X 2.77e-19
C19 B1 VGND 0.013269f
C20 A2 VPWR 0.020928f
C21 VPB C1 0.036801f
C22 A2 X 0.001572f
C23 A1 VGND 0.012567f
C24 VPB B2 0.025561f
C25 VPWR X 0.175411f
C26 A2 VGND 0.016752f
C27 VPB B1 0.032075f
C28 C1 B2 0.072571f
C29 VPWR VGND 0.093842f
C30 C1 B1 6.46e-19
C31 VPB A1 0.034297f
C32 X VGND 0.121872f
C33 VGND VNB 0.518524f
C34 X VNB 0.020031f
C35 VPWR VNB 0.443747f
C36 A2 VNB 0.089572f
C37 A1 VNB 0.105908f
C38 B1 VNB 0.108471f
C39 B2 VNB 0.088691f
C40 C1 VNB 0.139355f
C41 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221oi_1 VGND VPWR VPB VNB Y B1 C1 A1 A2 B2
X0 a_465_47.t1 A1.t0 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_109_297.t1 B1.t0 a_193_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297.t2 B2.t0 a_109_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_204_47.t0 B2.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.069875 pd=0.865 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 VGND.t0 A2.t0 a_465_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.099125 ps=0.955 w=0.65 l=0.15
X5 a_193_297.t1 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X6 Y.t0 B1.t1 a_204_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.069875 ps=0.865 w=0.65 l=0.15
X7 VPWR.t0 A2.t1 a_193_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.1525 ps=1.305 w=1 l=0.15
X8 a_109_297.t0 C1.t0 Y.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND.t2 C1.t1 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t1 234.804
R1 A1.n0 A1.t0 162.504
R2 A1 A1.n0 154.762
R3 Y Y.t2 636.313
R4 Y.n0 Y.t1 325.815
R5 Y.n0 Y.t0 249.615
R6 Y.n1 Y.t3 249.615
R7 Y Y.n1 65.0688
R8 Y.n1 Y.n0 26.6245
R9 a_465_47.t0 a_465_47.t1 56.3082
R10 VNB.t0 VNB.t4 2677.02
R11 VNB.t3 VNB.t1 1352.75
R12 VNB.t4 VNB.t2 1295.79
R13 VNB.t1 VNB.t0 1039.48
R14 VNB VNB.t3 925.567
R15 B1.n0 B1.t0 239.04
R16 B1.n0 B1.t1 166.739
R17 B1 B1.n0 156.952
R18 a_193_297.n1 a_193_297.n0 951.119
R19 a_193_297.n0 a_193_297.t3 33.4905
R20 a_193_297.n0 a_193_297.t1 26.5955
R21 a_193_297.t0 a_193_297.n1 26.5955
R22 a_193_297.n1 a_193_297.t2 26.5955
R23 a_109_297.n0 a_109_297.t1 1209.35
R24 a_109_297.n0 a_109_297.t2 26.5955
R25 a_109_297.t0 a_109_297.n0 26.5955
R26 VPB.t1 VPB.t2 556.386
R27 VPB.t2 VPB.t4 269.315
R28 VPB.t3 VPB.t1 248.599
R29 VPB.t0 VPB.t3 248.599
R30 VPB VPB.t0 192.369
R31 B2.n0 B2.t0 241.536
R32 B2.n0 B2.t1 169.237
R33 B2 B2.n0 168.762
R34 VGND.n1 VGND.t0 270.705
R35 VGND.n1 VGND.n0 207.814
R36 VGND.n0 VGND.t1 35.0774
R37 VGND.n0 VGND.t2 24.9236
R38 VGND VGND.n1 0.150974
R39 a_204_47.t0 a_204_47.t1 39.6928
R40 A2.n0 A2.t1 241.536
R41 A2.n0 A2.t0 169.237
R42 A2 A2.n0 159.758
R43 VPWR.n0 VPWR.t1 845.215
R44 VPWR.n0 VPWR.t0 354.211
R45 VPWR VPWR.n0 0.901642
R46 C1.n0 C1.t0 230.155
R47 C1 C1.n0 158.4
R48 C1.n0 C1.t1 157.856
C0 A1 A2 0.077092f
C1 B2 VPWR 0.008783f
C2 B1 Y 0.112632f
C3 C1 VGND 0.019827f
C4 B1 VPWR 0.009821f
C5 B2 VGND 0.017579f
C6 A1 Y 0.094522f
C7 A1 VPWR 0.01682f
C8 B1 VGND 0.013332f
C9 A2 Y 0.103832f
C10 VPB C1 0.038405f
C11 A2 VPWR 0.021049f
C12 A1 VGND 0.013044f
C13 VPB B2 0.025548f
C14 Y VPWR 0.080702f
C15 A2 VGND 0.016f
C16 C1 B2 0.07306f
C17 VPB B1 0.032273f
C18 Y VGND 0.370933f
C19 C1 B1 6.32e-19
C20 VPB A1 0.035145f
C21 VPWR VGND 0.062767f
C22 B2 B1 0.078843f
C23 VPB A2 0.030693f
C24 C1 A2 6.38e-20
C25 VPB Y 0.024108f
C26 C1 Y 0.078818f
C27 B2 A2 6.85e-20
C28 VPB VPWR 0.075926f
C29 B1 A1 0.064319f
C30 B2 Y 0.096707f
C31 VPB VGND 0.007682f
C32 C1 VPWR 0.014165f
C33 B1 A2 1.43e-19
C34 VGND VNB 0.402206f
C35 VPWR VNB 0.346755f
C36 Y VNB 0.146792f
C37 A2 VNB 0.117714f
C38 A1 VNB 0.107316f
C39 B1 VNB 0.108427f
C40 B2 VNB 0.088753f
C41 C1 VNB 0.142368f
C42 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211oi_2 VPWR VGND VPB VNB A2 A1 Y B1 C1
X0 VGND.t4 A2.t0 a_485_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR.t1 A1.t0 a_292_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297.t3 B1.t0 a_292_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y.t5 B1.t1 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47.t2 A2.t1 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297.t5 A2.t2 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND.t0 B1.t2 Y.t4 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR.t2 A2.t3 a_292_297.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47.t1 A1.t1 Y.t7 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND.t2 C1.t0 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y.t0 C1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11 a_37_297.t0 C1.t2 Y.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y.t6 A1.t2 a_485_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13 Y.t2 C1.t3 a_37_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297.t2 A1.t3 VPWR.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297.t0 B1.t3 a_37_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A2.n0 A2.t3 212.081
R1 A2.n1 A2.t2 212.081
R2 A2.n4 A2.n0 182.673
R3 A2.n3 A2.n2 152
R4 A2.n0 A2.t1 139.78
R5 A2.n1 A2.t0 139.78
R6 A2.n2 A2.n1 43.8187
R7 A2.n2 A2.n0 18.9884
R8 A2.n4 A2.n3 12.8005
R9 A2.n4 A2 11.2251
R10 A2.n3 A2 5.1205
R11 A2 A2.n4 2.16665
R12 a_485_47.t0 a_485_47.n1 323.447
R13 a_485_47.n1 a_485_47.t2 273.45
R14 a_485_47.n1 a_485_47.n0 185
R15 a_485_47.n0 a_485_47.t3 25.8467
R16 a_485_47.n0 a_485_47.t1 25.8467
R17 VGND.n4 VGND.t0 281.25
R18 VGND.n10 VGND.t1 241.054
R19 VGND.n5 VGND.n3 205.041
R20 VGND.n8 VGND.n2 199.739
R21 VGND.n3 VGND.t3 25.8467
R22 VGND.n3 VGND.t4 25.8467
R23 VGND.n2 VGND.t5 25.8467
R24 VGND.n2 VGND.t2 25.8467
R25 VGND.n9 VGND.n8 23.7181
R26 VGND.n10 VGND.n9 22.2123
R27 VGND.n8 VGND.n1 20.7064
R28 VGND.n4 VGND.n1 19.2005
R29 VGND.n11 VGND.n10 9.3005
R30 VGND.n6 VGND.n1 9.3005
R31 VGND.n8 VGND.n7 9.3005
R32 VGND.n9 VGND.n0 9.3005
R33 VGND.n5 VGND.n4 7.20769
R34 VGND.n6 VGND.n5 0.167962
R35 VGND.n7 VGND.n6 0.120292
R36 VGND.n7 VGND.n0 0.120292
R37 VGND.n11 VGND.n0 0.120292
R38 VGND VGND.n11 0.0278438
R39 VNB.t0 VNB.t2 2705.5
R40 VNB.t6 VNB.t5 1224.6
R41 VNB.t3 VNB.t6 1224.6
R42 VNB.t2 VNB.t3 1224.6
R43 VNB.t7 VNB.t0 1224.6
R44 VNB.t4 VNB.t7 1224.6
R45 VNB.t1 VNB.t4 1224.6
R46 VNB VNB.t1 1139.16
R47 A1.n1 A1.t0 212.081
R48 A1.n2 A1.t3 212.081
R49 A1.n2 A1.n0 182.673
R50 A1.n4 A1.n3 152
R51 A1.n1 A1.t1 139.78
R52 A1.n2 A1.t2 139.78
R53 A1.n3 A1.n1 43.8187
R54 A1.n3 A1.n2 18.9884
R55 A1.n4 A1.n0 17.4085
R56 A1.n0 A1 5.6325
R57 A1 A1.n4 0.5125
R58 a_292_297.n3 a_292_297.n2 368.567
R59 a_292_297.n2 a_292_297.n0 244.573
R60 a_292_297.n2 a_292_297.n1 206.814
R61 a_292_297.n0 a_292_297.t4 27.5805
R62 a_292_297.n0 a_292_297.t5 27.5805
R63 a_292_297.n1 a_292_297.t3 27.5805
R64 a_292_297.n1 a_292_297.t2 27.5805
R65 a_292_297.n3 a_292_297.t1 27.5805
R66 a_292_297.t0 a_292_297.n3 27.5805
R67 VPWR.n1 VPWR.t2 352.396
R68 VPWR.n5 VPWR.t0 345.884
R69 VPWR.n3 VPWR.n2 318.305
R70 VPWR.n2 VPWR.t3 27.5805
R71 VPWR.n2 VPWR.t1 27.5805
R72 VPWR.n5 VPWR.n4 24.4711
R73 VPWR.n4 VPWR.n3 22.9652
R74 VPWR.n4 VPWR.n0 9.3005
R75 VPWR.n6 VPWR.n5 7.32807
R76 VPWR.n3 VPWR.n1 6.8875
R77 VPWR.n1 VPWR.n0 0.628466
R78 VPWR VPWR.n6 0.59871
R79 VPWR.n6 VPWR.n0 0.15142
R80 VPB.t1 VPB.t4 562.306
R81 VPB.t7 VPB.t6 254.518
R82 VPB.t5 VPB.t7 254.518
R83 VPB.t4 VPB.t5 254.518
R84 VPB.t0 VPB.t1 254.518
R85 VPB.t2 VPB.t0 254.518
R86 VPB.t3 VPB.t2 254.518
R87 VPB VPB.t3 236.761
R88 B1.n0 B1.t0 212.081
R89 B1.n1 B1.t3 212.081
R90 B1 B1.n2 156.864
R91 B1.n0 B1.t2 139.78
R92 B1.n1 B1.t1 139.78
R93 B1.n2 B1.n0 31.4035
R94 B1.n2 B1.n1 31.4035
R95 B1 B1.n3 18.4325
R96 B1.n3 B1 9.30959
R97 B1.n3 B1 5.1205
R98 a_37_297.n0 a_37_297.t1 384.671
R99 a_37_297.n0 a_37_297.t3 373.562
R100 a_37_297.n1 a_37_297.n0 297.55
R101 a_37_297.t2 a_37_297.n1 27.5805
R102 a_37_297.n1 a_37_297.t0 27.5805
R103 Y.n1 Y.n0 292.94
R104 Y.n5 Y.n4 273.32
R105 Y.n7 Y 185.246
R106 Y.n3 Y.n2 185
R107 Y.n8 Y.n7 185
R108 Y.n6 Y.n5 47.6805
R109 Y.n0 Y.t1 27.5805
R110 Y.n0 Y.t2 27.5805
R111 Y.n4 Y.t7 25.8467
R112 Y.n4 Y.t6 25.8467
R113 Y.n2 Y.t4 25.8467
R114 Y.n2 Y.t5 25.8467
R115 Y.n7 Y.t3 25.8467
R116 Y.n7 Y.t0 25.8467
R117 Y Y.n6 15.895
R118 Y Y.n1 12.4213
R119 Y.n3 Y 9.76892
R120 Y.n5 Y.n3 5.72682
R121 Y.n1 Y 3.09135
R122 Y Y.n8 0.229071
R123 Y.n8 Y.n6 0.229071
R124 C1.n0 C1.t2 212.081
R125 C1.n1 C1.t3 212.081
R126 C1.n2 C1.n1 182.673
R127 C1.n0 C1.t0 139.78
R128 C1.n1 C1.t1 139.78
R129 C1.n1 C1.n0 62.8066
R130 C1.n2 C1 11.9612
R131 C1 C1.n2 2.3087
C0 Y VGND 0.27045f
C1 VPB B1 0.062335f
C2 VPWR VGND 0.090196f
C3 C1 B1 0.057966f
C4 VPB A1 0.071138f
C5 VPB A2 0.078568f
C6 B1 A1 0.030811f
C7 VPB Y 0.004207f
C8 B1 A2 0.00174f
C9 VPB VPWR 0.103659f
C10 C1 Y 0.120631f
C11 C1 VPWR 0.020382f
C12 VPB VGND 0.008913f
C13 B1 Y 0.136285f
C14 A1 A2 0.060636f
C15 C1 VGND 0.06149f
C16 B1 VPWR 0.019193f
C17 A1 Y 0.071168f
C18 A2 Y 1.42e-19
C19 B1 VGND 0.034439f
C20 A1 VPWR 0.0448f
C21 A1 VGND 0.022409f
C22 A2 VPWR 0.074628f
C23 Y VPWR 0.012611f
C24 A2 VGND 0.036829f
C25 VPB C1 0.073554f
C26 VGND VNB 0.556493f
C27 VPWR VNB 0.45848f
C28 Y VNB 0.030227f
C29 A2 VNB 0.249907f
C30 A1 VNB 0.207788f
C31 B1 VNB 0.182501f
C32 C1 VNB 0.247888f
C33 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB Y C1 B1 A1 A2
X0 a_56_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR.t1 A2.t0 a_56_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y.t3 C1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47.t1 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297.t0 B1.t0 a_56_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y.t2 C1.t1 a_311_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND.t0 B1.t1 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y.t1 A1.t1 a_139_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 A1.n0 A1.t0 241.536
R1 A1.n0 A1.t1 169.237
R2 A1.n1 A1.n0 152
R3 A1.n2 A1.n1 12.0247
R4 A1.n2 A1 11.7765
R5 A1 A1.n2 4.84898
R6 A1.n1 A1 0.970197
R7 VPWR VPWR.n0 315.284
R8 VPWR.n0 VPWR.t0 27.5805
R9 VPWR.n0 VPWR.t1 27.5805
R10 a_56_297.n0 a_56_297.t2 691.443
R11 a_56_297.n0 a_56_297.t1 27.5805
R12 a_56_297.t0 a_56_297.n0 27.5805
R13 VPB VPB.t2 281.154
R14 VPB.t1 VPB.t3 272.274
R15 VPB.t0 VPB.t1 254.518
R16 VPB.t2 VPB.t0 254.518
R17 A2.n0 A2.t0 228.649
R18 A2.n0 A2.t1 156.35
R19 A2 A2.n0 154.071
R20 C1.n0 C1.t1 231.017
R21 C1.n0 C1.t0 158.716
R22 C1.n1 C1.n0 152
R23 C1.n1 C1 12.1605
R24 C1 C1.n1 2.34717
R25 VGND.n1 VGND.t1 263.68
R26 VGND.n1 VGND.n0 204.78
R27 VGND.n0 VGND.t2 28.6159
R28 VGND.n0 VGND.t0 28.6159
R29 VGND VGND.n1 0.120713
R30 Y.n2 Y.t2 320.08
R31 Y.n1 Y.n0 246.785
R32 Y.n1 Y.t3 210.846
R33 Y.n0 Y.t0 25.8467
R34 Y.n0 Y.t1 25.8467
R35 Y Y.n1 16.7044
R36 Y.n2 Y 5.5408
R37 Y Y.n2 3.24826
R38 VNB VNB.t2 1352.75
R39 VNB.t0 VNB.t3 1310.03
R40 VNB.t1 VNB.t0 1224.6
R41 VNB.t2 VNB.t1 1224.6
R42 a_139_47.t0 a_139_47.t1 51.6928
R43 B1.n0 B1.t0 241.536
R44 B1.n0 B1.t1 169.237
R45 B1.n1 B1.n0 152
R46 B1 B1.n1 13.0788
R47 B1.n1 B1 2.13383
R48 a_311_297.t0 a_311_297.t1 61.0705
C0 VPB A1 0.02657f
C1 Y VGND 0.163399f
C2 VPB B1 0.031109f
C3 A2 A1 0.121006f
C4 A2 B1 4.79e-19
C5 VPB C1 0.041594f
C6 VPB VPWR 0.061754f
C7 A1 B1 0.08485f
C8 A1 C1 3.25e-19
C9 VPB Y 0.02709f
C10 A2 VPWR 0.02132f
C11 VPB VGND 0.007582f
C12 A1 VPWR 0.019745f
C13 B1 C1 0.110271f
C14 A2 VGND 0.049815f
C15 B1 VPWR 0.044975f
C16 A1 Y 0.044115f
C17 C1 VPWR 0.012342f
C18 B1 Y 0.099744f
C19 A1 VGND 0.084314f
C20 B1 VGND 0.017806f
C21 C1 Y 0.131233f
C22 C1 VGND 0.016549f
C23 VPWR Y 0.098999f
C24 VPB A2 0.043825f
C25 VPWR VGND 0.054287f
C26 VGND VNB 0.363898f
C27 Y VNB 0.105029f
C28 VPWR VNB 0.29066f
C29 C1 VNB 0.129395f
C30 B1 VNB 0.092441f
C31 A1 VNB 0.099121f
C32 A2 VNB 0.160478f
C33 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211o_4 VNB VPB VGND VPWR A2 A1 C1 X B1
X0 X.t3 a_79_204.t7 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_473_297# A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X3 X.t7 a_79_204.t8 VGND.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4 VGND.t3 C1.t0 a_79_204.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.104 ps=0.97 w=0.65 l=0.15
X5 a_79_204.t6 B1.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.092625 ps=0.935 w=0.65 l=0.15
X6 VPWR.t5 a_79_204.t9 X.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X7 a_473_297# A2.t0 VPWR.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X8 a_473_297# B1.t1 a_727_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16 ps=1.32 w=1 l=0.15
X9 X.t6 a_79_204.t10 VGND.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VGND.t1 B1.t2 a_79_204.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 a_79_204.t3 C1.t1 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.108875 ps=0.985 w=0.65 l=0.15
X12 VGND.t7 a_79_204.t11 X.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.095875 ps=0.945 w=0.65 l=0.15
X13 a_555_297.t0 B1.t3 a_473_297# VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X14 VPWR.t1 A2.t1 a_473_297# VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X15 VGND.t0 A2.t2 a_1123_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_951_47.t0 A2.t3 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.13975 ps=1.08 w=0.65 l=0.15
X17 VPWR.t4 a_79_204.t12 X.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND.t6 a_79_204.t13 X.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 a_79_204.t0 A1.t1 a_951_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X20 a_79_204.t4 C1.t2 a_555_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 a_727_297.t1 C1.t3 a_79_204.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X22 X.t0 a_79_204.t14 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
R0 a_79_204.n17 a_79_204.n16 693.005
R1 a_79_204.n7 a_79_204.t14 243.483
R2 a_79_204.n14 a_79_204.t11 207.698
R3 a_79_204.n14 a_79_204.t9 204.048
R4 a_79_204.n11 a_79_204.t7 204.048
R5 a_79_204.n5 a_79_204.t12 204.048
R6 a_79_204.n1 a_79_204.t0 203.024
R7 a_79_204.n3 a_79_204.n2 185
R8 a_79_204.n8 a_79_204.n7 167.543
R9 a_79_204.n9 a_79_204.n8 152
R10 a_79_204.n12 a_79_204.n4 152
R11 a_79_204.n15 a_79_204.n14 152
R12 a_79_204.n6 a_79_204.t8 147.814
R13 a_79_204.n10 a_79_204.t13 147.814
R14 a_79_204.n13 a_79_204.t10 147.814
R15 a_79_204.n1 a_79_204.n0 92.5005
R16 a_79_204.n3 a_79_204.n1 53.1664
R17 a_79_204.n16 a_79_204.n3 49.9732
R18 a_79_204.n13 a_79_204.n12 44.549
R19 a_79_204.n0 a_79_204.t3 36.9236
R20 a_79_204.n0 a_79_204.t1 35.0774
R21 a_79_204.n2 a_79_204.t2 33.2313
R22 a_79_204.n10 a_79_204.n9 31.4035
R23 a_79_204.n17 a_79_204.t5 27.5805
R24 a_79_204.t4 a_79_204.n17 27.5805
R25 a_79_204.n9 a_79_204.n5 26.2914
R26 a_79_204.n2 a_79_204.t6 25.8467
R27 a_79_204.n16 a_79_204.n15 23.5434
R28 a_79_204.n7 a_79_204.n6 18.2581
R29 a_79_204.n15 a_79_204.n4 15.5434
R30 a_79_204.n8 a_79_204.n4 15.5434
R31 a_79_204.n12 a_79_204.n11 13.146
R32 a_79_204.n14 a_79_204.n13 5.11262
R33 a_79_204.n11 a_79_204.n10 5.11262
R34 a_79_204.n6 a_79_204.n5 5.11262
R35 VPWR.n7 VPWR.t2 868.366
R36 VPWR.n9 VPWR.n8 598.965
R37 VPWR.n3 VPWR.t5 342.841
R38 VPWR.n23 VPWR.t3 337.2
R39 VPWR.n21 VPWR.n2 310.88
R40 VPWR.n8 VPWR.t0 49.2505
R41 VPWR.n11 VPWR.n10 34.6358
R42 VPWR.n11 VPWR.n5 34.6358
R43 VPWR.n15 VPWR.n5 34.6358
R44 VPWR.n16 VPWR.n15 34.6358
R45 VPWR.n17 VPWR.n16 34.6358
R46 VPWR.n2 VPWR.t6 27.5805
R47 VPWR.n2 VPWR.t4 27.5805
R48 VPWR.n8 VPWR.t1 27.5805
R49 VPWR.n21 VPWR.n20 24.8476
R50 VPWR.n23 VPWR.n22 19.9534
R51 VPWR.n22 VPWR.n21 19.577
R52 VPWR.n10 VPWR.n9 18.824
R53 VPWR.n20 VPWR.n3 15.0593
R54 VPWR.n10 VPWR.n6 9.3005
R55 VPWR.n12 VPWR.n11 9.3005
R56 VPWR.n13 VPWR.n5 9.3005
R57 VPWR.n15 VPWR.n14 9.3005
R58 VPWR.n16 VPWR.n4 9.3005
R59 VPWR.n18 VPWR.n17 9.3005
R60 VPWR.n20 VPWR.n19 9.3005
R61 VPWR.n21 VPWR.n1 9.3005
R62 VPWR.n22 VPWR.n0 9.3005
R63 VPWR.n24 VPWR.n23 9.3005
R64 VPWR.n9 VPWR.n7 6.83865
R65 VPWR.n17 VPWR.n3 0.753441
R66 VPWR.n7 VPWR.n6 0.529382
R67 VPWR.n12 VPWR.n6 0.120292
R68 VPWR.n13 VPWR.n12 0.120292
R69 VPWR.n14 VPWR.n13 0.120292
R70 VPWR.n14 VPWR.n4 0.120292
R71 VPWR.n18 VPWR.n4 0.120292
R72 VPWR.n19 VPWR.n18 0.120292
R73 VPWR.n19 VPWR.n1 0.120292
R74 VPWR.n1 VPWR.n0 0.120292
R75 VPWR.n24 VPWR.n0 0.120292
R76 VPWR VPWR.n24 0.0226354
R77 X.n2 X.n1 362.332
R78 X.n2 X.n0 310.38
R79 X.n5 X.n4 240.959
R80 X.n5 X.n3 198.137
R81 X X.n2 62.9428
R82 X X.n5 39.5794
R83 X.n4 X.t5 28.6159
R84 X.n1 X.t2 27.5805
R85 X.n1 X.t3 27.5805
R86 X.n0 X.t1 27.5805
R87 X.n0 X.t0 27.5805
R88 X.n3 X.t4 25.8467
R89 X.n3 X.t7 25.8467
R90 X.n4 X.t6 25.8467
R91 VPB.t9 VPB.t2 556.386
R92 VPB.t0 VPB.t6 509.034
R93 VPB.t1 VPB.t0 319.627
R94 VPB.t5 VPB.t1 319.627
R95 VPB.t4 VPB.t5 278.193
R96 VPB.t3 VPB.t4 254.518
R97 VPB.t2 VPB.t3 254.518
R98 VPB.t10 VPB.t9 254.518
R99 VPB.t8 VPB.t10 254.518
R100 VPB.t7 VPB.t8 254.518
R101 VPB VPB.t7 192.369
R102 A1.n2 A1.n0 204.048
R103 A1.n3 A1.t0 204.048
R104 A1 A1.n4 154.042
R105 A1.n2 A1.n1 147.814
R106 A1.n3 A1.t1 147.814
R107 A1.n4 A1.n2 49.6611
R108 A1.n4 A1.n3 13.146
R109 VGND.n20 VGND.t9 281.25
R110 VGND.n11 VGND.n5 198.964
R111 VGND.n18 VGND.n2 198.964
R112 VGND.n14 VGND.n13 198.756
R113 VGND.n7 VGND.n6 185
R114 VGND.n8 VGND.t0 157.083
R115 VGND.n6 VGND.t2 46.1543
R116 VGND.n6 VGND.t1 33.2313
R117 VGND.n5 VGND.t4 33.2313
R118 VGND.n11 VGND.n4 33.1299
R119 VGND.n14 VGND.n12 32.7534
R120 VGND.n18 VGND.n1 29.7417
R121 VGND.n5 VGND.t3 28.6159
R122 VGND.n13 VGND.t7 26.7697
R123 VGND.n13 VGND.t5 25.8467
R124 VGND.n2 VGND.t8 25.8467
R125 VGND.n2 VGND.t6 25.8467
R126 VGND.n20 VGND.n19 25.224
R127 VGND.n7 VGND.n4 25.0678
R128 VGND.n19 VGND.n18 14.6829
R129 VGND.n12 VGND.n11 11.2946
R130 VGND.n14 VGND.n1 11.2946
R131 VGND.n19 VGND.n0 9.3005
R132 VGND.n18 VGND.n17 9.3005
R133 VGND.n16 VGND.n1 9.3005
R134 VGND.n15 VGND.n14 9.3005
R135 VGND.n12 VGND.n3 9.3005
R136 VGND.n11 VGND.n10 9.3005
R137 VGND.n9 VGND.n4 9.3005
R138 VGND.n8 VGND.n7 7.55348
R139 VGND.n21 VGND.n20 6.99075
R140 VGND.n9 VGND.n8 0.169562
R141 VGND.n21 VGND.n0 0.150171
R142 VGND.n10 VGND.n9 0.120292
R143 VGND.n10 VGND.n3 0.120292
R144 VGND.n15 VGND.n3 0.120292
R145 VGND.n16 VGND.n15 0.120292
R146 VGND.n17 VGND.n16 0.120292
R147 VGND.n17 VGND.n0 0.120292
R148 VGND VGND.n21 0.113169
R149 VNB.t6 VNB.t0 2449.19
R150 VNB VNB.t10 2050.49
R151 VNB.t1 VNB.t2 1651.78
R152 VNB.t4 VNB.t1 1537.86
R153 VNB.t3 VNB.t4 1381.23
R154 VNB.t5 VNB.t3 1338.51
R155 VNB.t9 VNB.t8 1267.31
R156 VNB.t8 VNB.t5 1238.83
R157 VNB.t2 VNB.t6 1224.6
R158 VNB.t7 VNB.t9 1224.6
R159 VNB.t10 VNB.t7 1224.6
R160 C1.n0 C1.t3 202.44
R161 C1.n1 C1.t2 202.44
R162 C1.n1 C1.t0 145.436
R163 C1.n0 C1.t1 138.173
R164 C1 C1.n2 69.8937
R165 C1.n2 C1.n0 29.9182
R166 C1.n2 C1.n1 21.3278
R167 B1.n1 B1.t1 231.798
R168 B1.n0 B1.t3 231.798
R169 B1 B1.n0 224.472
R170 B1.n0 B1.t0 168.262
R171 B1 B1.n1 163.055
R172 B1.n1 B1.t2 162.127
R173 A2 A2.n0 233.582
R174 A2.n1 A2.t0 231.798
R175 A2.n0 A2.t1 223.036
R176 A2 A2.n1 173.273
R177 A2.n0 A2.t3 168.262
R178 A2.n1 A2.t2 166.51
R179 a_727_297.t0 a_727_297.t1 63.0405
R180 a_555_297.t0 a_555_297.t1 55.1605
R181 a_951_47.t0 a_951_47.t1 51.6928
C0 B1 C1 0.231125f
C1 VPB A2 0.073795f
C2 VPB A1 0.05279f
C3 B1 A2 0.075331f
C4 a_473_297# VPB 0.017146f
C5 B1 A1 1.23e-19
C6 VPB VPWR 0.13389f
C7 a_473_297# B1 0.053189f
C8 VPB X 0.012084f
C9 B1 VPWR 0.02446f
C10 a_473_297# C1 0.017303f
C11 C1 VPWR 0.015804f
C12 B1 X 4.69e-19
C13 VPB VGND 0.009828f
C14 A2 A1 0.203404f
C15 a_473_297# A2 0.182594f
C16 B1 VGND 0.033873f
C17 A2 VPWR 0.046886f
C18 a_473_297# A1 0.027121f
C19 A1 VPWR 0.028419f
C20 C1 VGND 0.030523f
C21 a_473_297# VPWR 0.51593f
C22 A2 VGND 0.069679f
C23 VPWR X 0.349346f
C24 A1 VGND 0.028681f
C25 VPB B1 0.071927f
C26 a_473_297# VGND 0.013604f
C27 VPWR VGND 0.127306f
C28 VPB C1 0.054952f
C29 X VGND 0.243572f
C30 VGND VNB 0.75065f
C31 X VNB 0.0733f
C32 VPWR VNB 0.611806f
C33 A1 VNB 0.169255f
C34 A2 VNB 0.244062f
C35 C1 VNB 0.177791f
C36 B1 VNB 0.198467f
C37 VPB VNB 1.31353f
C38 a_473_297# VNB 0.035689f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211o_2 VNB VPB VGND VPWR X A2 A1 B1 C1
X0 a_79_21.t1 A1.t0 a_348_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.13325 ps=1.06 w=0.65 l=0.15
X1 a_79_21.t0 C1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND.t2 a_79_21.t4 X.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.199875 pd=1.265 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR.t1 a_79_21.t5 X.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21.t2 C1.t1 a_585_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR.t3 A2.t0 a_299_297.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297.t1 A1.t1 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297.t1 B1.t0 a_299_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47.t1 A2.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.199875 ps=1.265 w=0.65 l=0.15
X9 X.t2 a_79_21.t6 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X.t0 a_79_21.t7 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND.t3 B1.t1 a_79_21.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
R0 A1.n0 A1.t1 239.04
R1 A1 A1.n0 168.975
R2 A1.n0 A1.t0 166.739
R3 a_348_47.t0 a_348_47.t1 75.6928
R4 a_79_21.n4 a_79_21.t4 1296.58
R5 a_79_21.t2 a_79_21.n5 492.921
R6 a_79_21.n3 a_79_21.t5 212.081
R7 a_79_21.n2 a_79_21.t6 212.081
R8 a_79_21.n1 a_79_21.t0 182.989
R9 a_79_21.n5 a_79_21.n4 161.641
R10 a_79_21.n2 a_79_21.t7 141.387
R11 a_79_21.n1 a_79_21.n0 98.982
R12 a_79_21.n5 a_79_21.n1 84.1066
R13 a_79_21.n3 a_79_21.n2 62.2897
R14 a_79_21.n0 a_79_21.t3 39.6928
R15 a_79_21.n0 a_79_21.t1 25.8467
R16 a_79_21.n4 a_79_21.n3 19.2805
R17 VNB.t2 VNB.t5 2178.64
R18 VNB.t5 VNB.t3 1594.82
R19 VNB.t3 VNB.t4 1438.19
R20 VNB.t4 VNB.t0 1366.99
R21 VNB.t1 VNB.t2 1224.6
R22 VNB VNB.t1 911.327
R23 C1.n0 C1.t1 230.155
R24 C1.n0 C1.t0 157.856
R25 C1 C1.n0 155.897
R26 VGND.n4 VGND.n2 207.857
R27 VGND.n8 VGND.n7 185
R28 VGND.n6 VGND.n5 185
R29 VGND.n10 VGND.t1 154.322
R30 VGND.n7 VGND.n6 63.6928
R31 VGND.n2 VGND.t0 30.462
R32 VGND.n2 VGND.t3 30.462
R33 VGND.n6 VGND.t4 24.9236
R34 VGND.n7 VGND.t2 24.9236
R35 VGND.n9 VGND.n8 23.1854
R36 VGND.n10 VGND.n9 22.9652
R37 VGND.n5 VGND.n4 10.8893
R38 VGND.n11 VGND.n10 9.3005
R39 VGND.n3 VGND.n1 9.3005
R40 VGND.n9 VGND.n0 9.3005
R41 VGND.n5 VGND.n1 7.36654
R42 VGND.n8 VGND.n1 0.966538
R43 VGND.n4 VGND.n3 0.226386
R44 VGND.n3 VGND.n0 0.120292
R45 VGND.n11 VGND.n0 0.120292
R46 VGND VGND.n11 0.0213333
R47 X.n2 X.n1 286.505
R48 X.n2 X.n0 157.026
R49 X.n1 X.t3 26.5955
R50 X.n1 X.t2 26.5955
R51 X.n0 X.t1 26.2846
R52 X.n0 X.t0 25.4075
R53 X X.n2 15.3326
R54 VPWR.n2 VPWR.n1 607.684
R55 VPWR.n3 VPWR.t1 342.377
R56 VPWR.n5 VPWR.t0 246.309
R57 VPWR.n1 VPWR.t3 39.4005
R58 VPWR.n1 VPWR.t2 37.4305
R59 VPWR.n4 VPWR.n3 23.3417
R60 VPWR.n5 VPWR.n4 22.9652
R61 VPWR.n4 VPWR.n0 9.3005
R62 VPWR.n6 VPWR.n5 9.3005
R63 VPWR.n3 VPWR.n2 6.94396
R64 VPWR.n2 VPWR.n0 0.485703
R65 VPWR.n6 VPWR.n0 0.120292
R66 VPWR VPWR.n6 0.0213333
R67 VPB.t2 VPB.t5 556.386
R68 VPB.t5 VPB.t4 319.627
R69 VPB.t4 VPB.t3 284.113
R70 VPB.t1 VPB.t2 248.599
R71 VPB.t3 VPB.t0 213.084
R72 VPB VPB.t1 189.409
R73 a_585_297.t0 a_585_297.t1 41.3705
R74 A2.n0 A2.t1 929.509
R75 A2.n0 A2.t0 232.214
R76 A2 A2.n0 158.958
R77 a_299_297.n0 a_299_297.t2 671.903
R78 a_299_297.n0 a_299_297.t1 36.4455
R79 a_299_297.t0 a_299_297.n0 28.5655
R80 B1.n0 B1.t0 241.536
R81 B1.n0 B1.t1 169.237
R82 B1 B1.n0 158.123
C0 VPB A1 0.029696f
C1 X VGND 0.107748f
C2 A2 A1 0.064227f
C3 VPB B1 0.025638f
C4 VPB C1 0.036777f
C5 A1 B1 0.069184f
C6 VPB VPWR 0.091679f
C7 VPB X 0.004802f
C8 A2 VPWR 0.015951f
C9 A2 X 9.43e-19
C10 VPB VGND 0.009198f
C11 A1 VPWR 0.015966f
C12 B1 C1 0.079269f
C13 A1 X 3.94e-19
C14 B1 VPWR 0.01195f
C15 A2 VGND 0.015948f
C16 C1 VPWR 0.012939f
C17 A1 VGND 0.014291f
C18 B1 X 9.84e-20
C19 B1 VGND 0.017802f
C20 C1 X 5.87e-20
C21 C1 VGND 0.016465f
C22 VPWR X 0.138423f
C23 VPB A2 0.038628f
C24 VPWR VGND 0.089685f
C25 VGND VNB 0.463866f
C26 X VNB 0.021972f
C27 VPWR VNB 0.397927f
C28 C1 VNB 0.142457f
C29 B1 VNB 0.090574f
C30 A1 VNB 0.094571f
C31 A2 VNB 0.10647f
C32 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR.t2 a_80_21.t4 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21.t1 C1.t0 a_472_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR.t1 A2.t0 a_217_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND.t2 B1.t0 a_80_21.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND.t1 a_80_21.t5 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47.t1 A2.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21.t0 A1.t1 a_300_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297.t0 B1.t1 a_217_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21.t2 C1.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
R0 a_80_21.t1 a_80_21.n3 500.909
R1 a_80_21.n1 a_80_21.t2 270.467
R2 a_80_21.n2 a_80_21.t4 231.017
R3 a_80_21.n1 a_80_21.n0 185
R4 a_80_21.n2 a_80_21.t5 158.716
R5 a_80_21.n3 a_80_21.n2 152
R6 a_80_21.n3 a_80_21.n1 102.07
R7 a_80_21.n0 a_80_21.t3 25.8467
R8 a_80_21.n0 a_80_21.t0 25.8467
R9 X.n1 X.t1 834.038
R10 X X.t1 819.707
R11 X.n0 X.t0 128.258
R12 X.n1 X 7.83334
R13 X X.n0 6.93004
R14 X X.n1 6.168
R15 X.n0 X 5.79322
R16 VPWR.n1 VPWR.n0 604.54
R17 VPWR.n1 VPWR.t2 343.5
R18 VPWR.n0 VPWR.t0 27.5805
R19 VPWR.n0 VPWR.t1 27.5805
R20 VPWR VPWR.n1 0.461646
R21 VPB.t3 VPB.t1 562.306
R22 VPB.t4 VPB.t2 272.274
R23 VPB.t0 VPB.t4 254.518
R24 VPB.t1 VPB.t0 254.518
R25 VPB VPB.t3 201.246
R26 C1.n0 C1.t0 231.017
R27 C1.n0 C1.t1 158.716
R28 C1 C1.n0 154.607
R29 a_472_297.t0 a_472_297.t1 61.0705
R30 A2.n0 A2.t0 231.017
R31 A2.n0 A2.t1 158.716
R32 A2 A2.n0 157.43
R33 a_217_297.n0 a_217_297.t1 658.159
R34 a_217_297.n0 a_217_297.t2 27.5805
R35 a_217_297.t0 a_217_297.n0 27.5805
R36 B1.n0 B1.t1 241.536
R37 B1.n0 B1.t0 169.237
R38 B1 B1.n0 157.042
R39 VGND.n5 VGND.n1 204.948
R40 VGND.n4 VGND.n3 185
R41 VGND.n2 VGND.n0 185
R42 VGND.n3 VGND.n2 66.462
R43 VGND.n3 VGND.t0 40.6159
R44 VGND.n2 VGND.t1 40.6159
R45 VGND.n1 VGND.t3 28.6159
R46 VGND.n1 VGND.t2 28.6159
R47 VGND.n6 VGND.n0 9.40836
R48 VGND.n4 VGND.n0 8.53383
R49 VGND.n5 VGND.n4 7.57682
R50 VGND.n6 VGND.n5 0.250352
R51 VGND VGND.n6 0.122488
R52 VNB.t2 VNB.t1 2705.5
R53 VNB.t3 VNB.t4 1310.03
R54 VNB.t0 VNB.t3 1224.6
R55 VNB.t1 VNB.t0 1224.6
R56 VNB VNB.t2 968.285
R57 a_300_47.t0 a_300_47.t1 51.6928
R58 A1.n0 A1.t0 241.536
R59 A1.n0 A1.t1 169.237
R60 A1 A1.n0 164.024
C0 B1 C1 0.084607f
C1 VPWR VGND 0.066493f
C2 X VPB 0.011762f
C3 X A2 6.82e-19
C4 VPWR VPB 0.075404f
C5 X A1 3.62e-19
C6 VPWR A2 0.016058f
C7 VGND VPB 0.007748f
C8 VGND A2 0.019089f
C9 VPWR A1 0.014884f
C10 X B1 1.18e-19
C11 X C1 7.15e-20
C12 VPWR B1 0.01289f
C13 VGND A1 0.014726f
C14 VPB A2 0.038351f
C15 VPWR C1 0.013731f
C16 VGND B1 0.017479f
C17 VPB A1 0.026604f
C18 VGND C1 0.01758f
C19 VPB B1 0.026706f
C20 A2 A1 0.088064f
C21 VPB C1 0.037912f
C22 A1 B1 0.083391f
C23 X VPWR 0.088406f
C24 X VGND 0.065404f
C25 VGND VNB 0.38475f
C26 VPWR VNB 0.325154f
C27 X VNB 0.08992f
C28 C1 VNB 0.144368f
C29 B1 VNB 0.089926f
C30 A1 VNB 0.090508f
C31 A2 VNB 0.107869f
C32 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47.t0 A1.t0 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X.t1 a_27_47.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297.t2 B1.t0 a_193_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297.t0 B2.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X.t0 a_27_47.t5 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47.t1 B2.t1 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR.t2 A2.t0 a_193_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297.t1 A1.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47.t1 B1.t1 a_205_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297.t1 C1.t0 a_27_47.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND.t1 C1.t1 a_27_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND.t3 A2.t1 a_465_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
R0 A1.n0 A1.t1 236.552
R1 A1.n0 A1.t0 164.251
R2 A1 A1.n0 154.47
R3 a_27_47.t3 a_27_47.n3 669.389
R4 a_27_47.n0 a_27_47.t2 326.493
R5 a_27_47.n0 a_27_47.t1 249.615
R6 a_27_47.n1 a_27_47.t0 249.615
R7 a_27_47.n2 a_27_47.t4 241.536
R8 a_27_47.n2 a_27_47.t5 169.237
R9 a_27_47.n3 a_27_47.n2 152
R10 a_27_47.n3 a_27_47.n1 108.529
R11 a_27_47.n1 a_27_47.n0 26.6245
R12 a_465_47.t0 a_465_47.t1 60.9236
R13 VNB.t2 VNB.t0 2677.02
R14 VNB.t0 VNB.t5 1366.99
R15 VNB.t3 VNB.t4 1366.99
R16 VNB.t5 VNB.t1 1324.27
R17 VNB.t4 VNB.t2 1025.24
R18 VNB VNB.t3 911.327
R19 VPWR.n3 VPWR.t0 838.817
R20 VPWR.n4 VPWR.n2 317.562
R21 VPWR.n9 VPWR 37.9123
R22 VPWR.n2 VPWR.t2 35.4605
R23 VPWR.n7 VPWR.n1 34.6358
R24 VPWR.n8 VPWR.n7 34.6358
R25 VPWR.n2 VPWR.t1 26.5955
R26 VPWR.n3 VPWR.n1 19.9534
R27 VPWR.n5 VPWR.n1 9.3005
R28 VPWR.n7 VPWR.n6 9.3005
R29 VPWR.n8 VPWR.n0 9.3005
R30 VPWR.n4 VPWR.n3 6.63632
R31 VPWR VPWR.n8 6.02403
R32 VPWR.n5 VPWR.n4 0.571201
R33 VPWR.n6 VPWR.n5 0.120292
R34 VPWR.n6 VPWR.n0 0.120292
R35 VPWR.n9 VPWR.n0 0.120292
R36 VPWR VPWR.n9 0.0213333
R37 X.n0 X 593.784
R38 X.n1 X.n0 585
R39 X X.t0 249.867
R40 X.n2 X.n1 98.9003
R41 X.n0 X.t1 26.5955
R42 X X.n2 11.0708
R43 X.n1 X 8.28285
R44 X.n2 X 8.03187
R45 VPB.t3 VPB.t1 556.386
R46 VPB.t1 VPB.t4 284.113
R47 VPB.t4 VPB.t2 275.235
R48 VPB.t0 VPB.t3 248.599
R49 VPB.t5 VPB.t0 248.599
R50 VPB VPB.t5 189.409
R51 B1.n0 B1.t0 239.505
R52 B1.n0 B1.t1 167.204
R53 B1 B1.n0 157.12
R54 a_193_297.n1 a_193_297.n0 953.038
R55 a_193_297.n0 a_193_297.t2 33.4905
R56 a_193_297.n0 a_193_297.t1 31.5205
R57 a_193_297.n1 a_193_297.t3 26.5955
R58 a_193_297.t0 a_193_297.n1 26.5955
R59 a_109_297.n0 a_109_297.t2 1201.3
R60 a_109_297.t0 a_109_297.n0 26.5955
R61 a_109_297.n0 a_109_297.t1 26.5955
R62 B2.n0 B2.t0 241.536
R63 B2 B2.n0 169.921
R64 B2.n0 B2.t1 169.237
R65 VGND.n3 VGND.n0 206.794
R66 VGND.n2 VGND.n1 202.067
R67 VGND.n1 VGND.t2 36.0005
R68 VGND.n0 VGND.t0 33.2313
R69 VGND.n1 VGND.t1 24.9236
R70 VGND.n0 VGND.t3 24.9236
R71 VGND.n3 VGND.n2 5.74703
R72 VGND.n2 VGND 3.29747
R73 VGND VGND.n3 0.148914
R74 a_205_47.t0 a_205_47.t1 38.7697
R75 A2.n0 A2.t0 241.536
R76 A2.n0 A2.t1 169.237
R77 A2 A2.n0 164.8
R78 C1.n0 C1.t0 231.718
R79 C1 C1.n0 159.619
R80 C1.n0 C1.t1 159.417
C0 C1 B2 0.072571f
C1 VPB B1 0.032075f
C2 VPWR VGND 0.072225f
C3 VPB A1 0.034297f
C4 C1 B1 6.46e-19
C5 X VGND 0.061021f
C6 C1 A1 1.77e-20
C7 VPB A2 0.026961f
C8 B2 B1 0.078429f
C9 VPB VPWR 0.079908f
C10 C1 A2 9.03e-21
C11 VPB X 0.011274f
C12 C1 VPWR 0.013943f
C13 B1 A1 0.060935f
C14 B2 VPWR 0.00842f
C15 VPB VGND 0.008441f
C16 C1 X 5.03e-20
C17 B2 X 6.77e-20
C18 C1 VGND 0.019615f
C19 B1 VPWR 0.009818f
C20 A1 A2 0.069236f
C21 B1 X 9.58e-20
C22 A1 VPWR 0.01613f
C23 B2 VGND 0.017443f
C24 A2 VPWR 0.020928f
C25 B1 VGND 0.013269f
C26 A1 X 2.77e-19
C27 VPB C1 0.036702f
C28 A2 X 0.001572f
C29 A1 VGND 0.012567f
C30 VPB B2 0.025561f
C31 A2 VGND 0.016752f
C32 VPWR X 0.089708f
C33 VGND VNB 0.437277f
C34 X VNB 0.091856f
C35 VPWR VNB 0.363959f
C36 A2 VNB 0.089572f
C37 A1 VNB 0.105908f
C38 B1 VNB 0.108471f
C39 B2 VNB 0.088691f
C40 C1 VNB 0.139233f
C41 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211oi_4 VNB VPB B1 VPWR VGND A2 A1 C1 Y
X0 Y.t5 A1.t0 a_109_47.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t9 C1.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t10 A2.t0 a_109_47.t7 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND.t0 B1.t0 Y.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.108875 ps=0.985 w=0.65 l=0.15
X4 VPWR.t3 A1.t1 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297.t2 A1.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t7 A2.t1 a_27_297.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_949_297.t0 B1.t1 a_27_297.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_297.t10 A2.t2 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t1 C1.t1 a_949_297.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X10 a_781_297.t2 C1.t2 Y.t12 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_297.t4 B1.t2 a_781_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND.t3 A2.t3 a_109_47.t4 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y.t4 A1.t3 a_109_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_781_297.t0 B1.t3 a_27_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1301_297.t1 C1.t3 Y.t13 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.15 ps=1.3 w=1 l=0.15
X16 a_27_297.t9 A2.t4 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_109_47.t5 A2.t5 VGND.t4 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_109_47.t1 A1.t4 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y.t9 C1.t4 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VPWR.t1 A1.t5 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_109_47.t0 A1.t6 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t10 C1.t5 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y.t7 B1.t4 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_27_297.t0 A1.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t8 B1.t5 VGND.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X26 VPWR.t4 A2.t6 a_27_297.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 a_27_297.t7 B1.t6 a_1301_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X28 VGND.t6 C1.t6 Y.t11 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X29 a_109_47.t6 A2.t7 VGND.t5 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X30 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.091 ps=0.93 w=0.65 l=0.15
R0 A1.n2 A1.t5 221.72
R1 A1.n1 A1.t7 221.72
R2 A1.n7 A1.t1 221.72
R3 A1.n8 A1.t2 221.72
R4 A1.n4 A1.n3 170.133
R5 A1 A1.n9 161.067
R6 A1.n5 A1.n4 152
R7 A1.n6 A1.n0 152
R8 A1.n2 A1.t6 149.421
R9 A1.n1 A1.t0 149.421
R10 A1.n7 A1.t4 149.421
R11 A1.n8 A1.t3 149.421
R12 A1.n6 A1.n5 60.6968
R13 A1.n9 A1.n7 58.9116
R14 A1.n3 A1.n1 48.2005
R15 A1.n3 A1.n2 26.7783
R16 A1.n4 A1.n0 18.1338
R17 A1.n9 A1.n8 16.0672
R18 A1.n5 A1.n1 12.4968
R19 A1 A1.n0 9.06717
R20 A1.n7 A1.n6 1.78569
R21 a_109_47.n2 a_109_47.n0 248.429
R22 a_109_47.n5 a_109_47.n4 228.008
R23 a_109_47.n4 a_109_47.n3 185
R24 a_109_47.n2 a_109_47.n1 185
R25 a_109_47.n4 a_109_47.n2 43.0085
R26 a_109_47.n1 a_109_47.t2 24.9236
R27 a_109_47.n1 a_109_47.t5 24.9236
R28 a_109_47.n3 a_109_47.t3 24.9236
R29 a_109_47.n3 a_109_47.t1 24.9236
R30 a_109_47.n0 a_109_47.t4 24.9236
R31 a_109_47.n0 a_109_47.t6 24.9236
R32 a_109_47.n5 a_109_47.t7 24.9236
R33 a_109_47.t0 a_109_47.n5 24.9236
R34 Y.n1 Y.n0 636.201
R35 Y.n1 Y.t13 612.581
R36 Y.n11 Y.t10 262.144
R37 Y.n6 Y.n4 241.589
R38 Y.n6 Y.n5 185
R39 Y.n10 Y.n2 96.031
R40 Y.n9 Y.n3 96.031
R41 Y.n8 Y.n7 95.3946
R42 Y Y.n11 94.1213
R43 Y.n8 Y.n6 79.2747
R44 Y Y.n1 48.6498
R45 Y.n11 Y.n10 46.3975
R46 Y.n10 Y.n9 44.4378
R47 Y.n9 Y.n8 39.5815
R48 Y.n7 Y.t6 33.2313
R49 Y.n7 Y.t7 28.6159
R50 Y.n0 Y.t12 27.5805
R51 Y.n0 Y.t1 27.5805
R52 Y.n3 Y.t8 25.8467
R53 Y.n2 Y.t0 24.9236
R54 Y.n2 Y.t9 24.9236
R55 Y.n3 Y.t11 24.9236
R56 Y.n4 Y.t3 24.9236
R57 Y.n4 Y.t4 24.9236
R58 Y.n5 Y.t2 24.9236
R59 Y.n5 Y.t5 24.9236
R60 VNB.t6 VNB.t5 1381.23
R61 VNB.t5 VNB.t7 1224.6
R62 VNB.t7 VNB.t10 1210.36
R63 VNB.t0 VNB.t9 1196.12
R64 VNB.t8 VNB.t0 1196.12
R65 VNB.t10 VNB.t8 1196.12
R66 VNB.t14 VNB.t6 1196.12
R67 VNB.t1 VNB.t14 1196.12
R68 VNB.t4 VNB.t1 1196.12
R69 VNB.t2 VNB.t4 1196.12
R70 VNB.t3 VNB.t2 1196.12
R71 VNB.t12 VNB.t3 1196.12
R72 VNB.t11 VNB.t12 1196.12
R73 VNB.t13 VNB.t11 1196.12
R74 VNB VNB.t13 911.327
R75 C1.n12 C1.t1 218.654
R76 C1.n3 C1.t3 212.081
R77 C1.n2 C1.n1 212.081
R78 C1.n9 C1.t2 212.081
R79 C1.n6 C1.n5 170.133
R80 C1 C1.n12 154.4
R81 C1.n7 C1.n6 152
R82 C1.n10 C1.n0 152
R83 C1.n3 C1.t5 139.78
R84 C1.n11 C1.t6 139.78
R85 C1.n8 C1.t4 139.78
R86 C1.n4 C1.t0 139.78
R87 C1.n11 C1.n10 48.9308
R88 C1.n8 C1.n7 37.246
R89 C1.n5 C1.n3 35.7853
R90 C1.n5 C1.n4 25.5611
R91 C1.n7 C1.n2 19.7187
R92 C1.n6 C1.n0 18.1338
R93 C1 C1.n0 15.7338
R94 C1.n10 C1.n9 6.57323
R95 C1.n9 C1.n8 5.84292
R96 C1.n4 C1.n2 4.38232
R97 C1.n12 C1.n11 0.730803
R98 VGND.n28 VGND.t5 284.291
R99 VGND.n15 VGND.n14 205.707
R100 VGND.n26 VGND.n2 204.609
R101 VGND.n9 VGND.n8 204.302
R102 VGND.n7 VGND.n6 198.964
R103 VGND.n13 VGND.n12 198.964
R104 VGND.n20 VGND.n4 34.6358
R105 VGND.n21 VGND.n20 34.6358
R106 VGND.n22 VGND.n21 34.6358
R107 VGND.n22 VGND.n1 34.6358
R108 VGND.n16 VGND.n13 34.2593
R109 VGND.n26 VGND.n1 32.0005
R110 VGND.n11 VGND.n7 28.9887
R111 VGND.n12 VGND.t2 25.8467
R112 VGND.n12 VGND.t0 25.8467
R113 VGND.n8 VGND.t7 24.9236
R114 VGND.n8 VGND.t9 24.9236
R115 VGND.n6 VGND.t8 24.9236
R116 VGND.n6 VGND.t6 24.9236
R117 VGND.n14 VGND.t1 24.9236
R118 VGND.n14 VGND.t10 24.9236
R119 VGND.n2 VGND.t4 24.9236
R120 VGND.n2 VGND.t3 24.9236
R121 VGND.n28 VGND.n27 22.2123
R122 VGND.n16 VGND.n15 21.8358
R123 VGND.n27 VGND.n26 19.577
R124 VGND.n15 VGND.n4 12.8005
R125 VGND.n13 VGND.n11 10.1652
R126 VGND.n29 VGND.n28 9.3005
R127 VGND.n11 VGND.n10 9.3005
R128 VGND.n13 VGND.n5 9.3005
R129 VGND.n17 VGND.n16 9.3005
R130 VGND.n18 VGND.n4 9.3005
R131 VGND.n20 VGND.n19 9.3005
R132 VGND.n21 VGND.n3 9.3005
R133 VGND.n23 VGND.n22 9.3005
R134 VGND.n24 VGND.n1 9.3005
R135 VGND.n26 VGND.n25 9.3005
R136 VGND.n27 VGND.n0 9.3005
R137 VGND.n9 VGND.n7 6.06983
R138 VGND.n10 VGND.n9 0.645842
R139 VGND.n10 VGND.n5 0.120292
R140 VGND.n17 VGND.n5 0.120292
R141 VGND.n18 VGND.n17 0.120292
R142 VGND.n19 VGND.n18 0.120292
R143 VGND.n19 VGND.n3 0.120292
R144 VGND.n23 VGND.n3 0.120292
R145 VGND.n24 VGND.n23 0.120292
R146 VGND.n25 VGND.n24 0.120292
R147 VGND.n25 VGND.n0 0.120292
R148 VGND.n29 VGND.n0 0.120292
R149 VGND VGND.n29 0.0213333
R150 A2.n1 A2.n0 302.392
R151 A2.n0 A2.t4 241.536
R152 A2.n3 A2.t1 221.72
R153 A2.n5 A2.t2 221.72
R154 A2.n2 A2.t6 221.72
R155 A2.n0 A2.t0 169.237
R156 A2.n4 A2.n1 152
R157 A2.n3 A2.t5 149.421
R158 A2.n5 A2.t3 149.421
R159 A2.n2 A2.t7 149.421
R160 A2 A2.n6 69.2318
R161 A2.n5 A2.n4 58.9116
R162 A2.n6 A2.n2 38.4964
R163 A2.n6 A2.n5 26.582
R164 A2.n4 A2.n3 16.0672
R165 A2 A2.n1 3.25474
R166 B1.n1 B1.t6 241
R167 B1.n6 B1.t2 212.081
R168 B1.n3 B1.t1 212.081
R169 B1.n7 B1.t3 212.081
R170 B1.n10 B1.n1 185.887
R171 B1.n1 B1.n0 168.701
R172 B1.n4 B1.n2 163.569
R173 B1.n9 B1.n8 152.111
R174 B1.n6 B1.n2 152
R175 B1.n3 B1.t5 150.736
R176 B1.n7 B1.t4 139.78
R177 B1.n5 B1.t0 139.78
R178 B1.n8 B1.n6 49.6611
R179 B1.n5 B1.n4 40.1672
R180 B1.n4 B1.n3 11.6853
R181 B1.n8 B1.n7 11.6853
R182 B1.n6 B1.n5 9.49444
R183 B1.n10 B1.n9 9.3005
R184 B1.n9 B1.n2 7.3936
R185 B1 B1.n10 0.0466957
R186 a_27_297.n1 a_27_297.t7 1014.9
R187 a_27_297.n1 a_27_297.n0 585
R188 a_27_297.n6 a_27_297.t8 359.089
R189 a_27_297.n6 a_27_297.n5 296.125
R190 a_27_297.n7 a_27_297.n4 296.125
R191 a_27_297.n9 a_27_297.n8 296.125
R192 a_27_297.n3 a_27_297.n2 289.704
R193 a_27_297.n3 a_27_297.n1 56.7941
R194 a_27_297.n8 a_27_297.n3 40.2779
R195 a_27_297.n8 a_27_297.n7 34.6844
R196 a_27_297.n7 a_27_297.n6 34.6844
R197 a_27_297.n5 a_27_297.t11 26.5955
R198 a_27_297.n5 a_27_297.t10 26.5955
R199 a_27_297.n4 a_27_297.t3 26.5955
R200 a_27_297.n4 a_27_297.t2 26.5955
R201 a_27_297.n2 a_27_297.t5 26.5955
R202 a_27_297.n2 a_27_297.t9 26.5955
R203 a_27_297.n0 a_27_297.t6 26.5955
R204 a_27_297.n0 a_27_297.t4 26.5955
R205 a_27_297.n9 a_27_297.t1 26.5955
R206 a_27_297.t0 a_27_297.n9 26.5955
R207 VPWR.n7 VPWR.n6 604.34
R208 VPWR.n12 VPWR.n1 599.74
R209 VPWR.n10 VPWR.n3 598.965
R210 VPWR.n5 VPWR.n4 598.965
R211 VPWR.n10 VPWR.n9 28.9887
R212 VPWR.n1 VPWR.t6 26.5955
R213 VPWR.n1 VPWR.t4 26.5955
R214 VPWR.n3 VPWR.t2 26.5955
R215 VPWR.n3 VPWR.t7 26.5955
R216 VPWR.n4 VPWR.t0 26.5955
R217 VPWR.n4 VPWR.t3 26.5955
R218 VPWR.n6 VPWR.t5 26.5955
R219 VPWR.n6 VPWR.t1 26.5955
R220 VPWR.n12 VPWR.n11 22.9652
R221 VPWR.n11 VPWR.n10 15.4358
R222 VPWR.n9 VPWR.n5 9.41227
R223 VPWR.n9 VPWR.n8 9.3005
R224 VPWR.n10 VPWR.n2 9.3005
R225 VPWR.n11 VPWR.n0 9.3005
R226 VPWR.n13 VPWR.n12 7.12063
R227 VPWR.n7 VPWR.n5 7.02047
R228 VPWR.n8 VPWR.n7 1.05258
R229 VPWR.n13 VPWR.n0 0.148519
R230 VPWR.n8 VPWR.n2 0.120292
R231 VPWR.n2 VPWR.n0 0.120292
R232 VPWR VPWR.n13 0.11354
R233 VPB.t13 VPB.t12 520.872
R234 VPB.t12 VPB.t4 272.274
R235 VPB.t7 VPB.t14 266.356
R236 VPB.t14 VPB.t13 254.518
R237 VPB.t6 VPB.t7 248.599
R238 VPB.t5 VPB.t6 248.599
R239 VPB.t9 VPB.t5 248.599
R240 VPB.t1 VPB.t9 248.599
R241 VPB.t0 VPB.t1 248.599
R242 VPB.t3 VPB.t0 248.599
R243 VPB.t2 VPB.t3 248.599
R244 VPB.t11 VPB.t2 248.599
R245 VPB.t10 VPB.t11 248.599
R246 VPB.t8 VPB.t10 248.599
R247 VPB VPB.t8 189.409
R248 a_949_297.t0 a_949_297.t1 59.1005
R249 a_781_297.n0 a_781_297.t2 1518.59
R250 a_781_297.t1 a_781_297.n0 26.5955
R251 a_781_297.n0 a_781_297.t0 26.5955
R252 a_1301_297.t0 a_1301_297.t1 61.0705
C0 B1 VPWR 0.144163f
C1 A1 Y 0.127386f
C2 A2 VGND 0.09029f
C3 A1 VGND 0.031603f
C4 C1 VPWR 0.023722f
C5 B1 Y 0.302245f
C6 C1 Y 0.227194f
C7 B1 VGND 0.153083f
C8 C1 VGND 0.062615f
C9 VPWR Y 0.028275f
C10 VPB A2 0.130647f
C11 VPWR VGND 0.084987f
C12 VPB A1 0.115122f
C13 Y VGND 0.468819f
C14 VPB B1 0.127452f
C15 A2 A1 0.286291f
C16 VPB C1 0.123728f
C17 A2 B1 0.112951f
C18 VPB VPWR 0.126377f
C19 A1 B1 3.7e-19
C20 A2 VPWR 0.079684f
C21 VPB Y 0.010302f
C22 VPB VGND 0.007248f
C23 B1 C1 0.228079f
C24 A2 Y 0.045199f
C25 A1 VPWR 0.049361f
C26 VGND VNB 0.826102f
C27 Y VNB 0.090077f
C28 VPWR VNB 0.663483f
C29 C1 VNB 0.356249f
C30 B1 VNB 0.393234f
C31 A1 VNB 0.353022f
C32 A2 VNB 0.409115f
C33 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221oi_2 VNB VPB VGND VPWR A2 A1 B1 B2 Y C1
X0 Y.t4 B1.t0 a_383_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_301_297.t4 B1.t1 a_27_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297.t5 A2.t0 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 B2.t0 a_383_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t2 A1.t0 a_735_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297.t1 B2.t1 a_301_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR.t3 A1.t1 a_301_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t4 A2.t1 a_735_47.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_301_297.t0 A1.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t7 C1.t0 a_27_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND.t5 C1.t1 Y.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y.t0 C1.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1755 ps=1.84 w=0.65 l=0.15
X12 VPWR.t1 A2.t2 a_301_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47.t0 B2.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X14 a_383_47.t1 B1.t2 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_735_47.t0 A2.t3 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X16 a_27_297.t4 C1.t3 Y.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297.t1 B2.t3 a_27_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47.t2 A1.t3 Y.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297.t2 B1.t3 a_301_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 B1.n0 B1.t3 212.081
R1 B1.n1 B1.t1 212.081
R2 B1 B1.n2 153.268
R3 B1.n0 B1.t2 139.78
R4 B1.n1 B1.t0 139.78
R5 B1.n2 B1.n0 30.6732
R6 B1.n2 B1.n1 30.6732
R7 a_383_47.n1 a_383_47.n0 418.873
R8 a_383_47.n0 a_383_47.t3 24.9236
R9 a_383_47.n0 a_383_47.t1 24.9236
R10 a_383_47.n1 a_383_47.t2 24.9236
R11 a_383_47.t0 a_383_47.n1 24.9236
R12 Y Y.n0 323.158
R13 Y.n3 Y.n1 302.935
R14 Y.n3 Y.n2 185
R15 Y.n5 Y.n3 110.797
R16 Y.n5 Y.n4 101.01
R17 Y.n0 Y.t5 26.5955
R18 Y.n0 Y.t7 26.5955
R19 Y.n4 Y.t6 24.9236
R20 Y.n4 Y.t0 24.9236
R21 Y.n2 Y.t3 24.9236
R22 Y.n2 Y.t4 24.9236
R23 Y.n1 Y.t1 24.9236
R24 Y.n1 Y.t2 24.9236
R25 Y Y.n5 14.8485
R26 VNB.t9 VNB.t1 2677.02
R27 VNB.t7 VNB.t6 1423.95
R28 VNB.t2 VNB.t8 1196.12
R29 VNB.t3 VNB.t2 1196.12
R30 VNB.t6 VNB.t3 1196.12
R31 VNB.t4 VNB.t7 1196.12
R32 VNB.t5 VNB.t4 1196.12
R33 VNB.t1 VNB.t5 1196.12
R34 VNB.t0 VNB.t9 1196.12
R35 VNB VNB.t0 939.807
R36 a_27_297.n3 a_27_297.n2 638.836
R37 a_27_297.n2 a_27_297.n1 585
R38 a_27_297.n0 a_27_297.t4 410.938
R39 a_27_297.n0 a_27_297.t5 384.33
R40 a_27_297.n2 a_27_297.n0 64.632
R41 a_27_297.n1 a_27_297.t3 26.5955
R42 a_27_297.n1 a_27_297.t1 26.5955
R43 a_27_297.t0 a_27_297.n3 26.5955
R44 a_27_297.n3 a_27_297.t2 26.5955
R45 a_301_297.n4 a_301_297.t2 877.509
R46 a_301_297.n5 a_301_297.n4 585
R47 a_301_297.n1 a_301_297.n0 301.397
R48 a_301_297.n3 a_301_297.n2 288.089
R49 a_301_297.n1 a_301_297.t5 276.938
R50 a_301_297.n4 a_301_297.n3 65.063
R51 a_301_297.n3 a_301_297.n1 60.3571
R52 a_301_297.n2 a_301_297.t6 34.4755
R53 a_301_297.n2 a_301_297.t1 34.4755
R54 a_301_297.n0 a_301_297.t7 26.5955
R55 a_301_297.n0 a_301_297.t0 26.5955
R56 a_301_297.n5 a_301_297.t3 26.5955
R57 a_301_297.t4 a_301_297.n5 26.5955
R58 VPB.t8 VPB.t2 556.386
R59 VPB.t1 VPB.t6 295.95
R60 VPB.t7 VPB.t5 248.599
R61 VPB.t0 VPB.t7 248.599
R62 VPB.t6 VPB.t0 248.599
R63 VPB.t3 VPB.t1 248.599
R64 VPB.t4 VPB.t3 248.599
R65 VPB.t2 VPB.t4 248.599
R66 VPB.t9 VPB.t8 248.599
R67 VPB VPB.t9 195.327
R68 A2.n2 A2.n0 260.188
R69 A2.n1 A2.t0 241.536
R70 A2.n0 A2.t2 241.536
R71 A2.n1 A2.t1 169.237
R72 A2.n0 A2.t3 169.237
R73 A2.n2 A2.n1 152
R74 A2 A2.n2 23.6805
R75 VPWR.n2 VPWR.n1 613.489
R76 VPWR.n2 VPWR.n0 611.771
R77 VPWR.n0 VPWR.t0 26.5955
R78 VPWR.n0 VPWR.t1 26.5955
R79 VPWR.n1 VPWR.t2 26.5955
R80 VPWR.n1 VPWR.t3 26.5955
R81 VPWR VPWR.n2 1.46107
R82 B2.n1 B2.t1 241.536
R83 B2.n0 B2.t3 241.536
R84 B2.n2 B2.n0 238.481
R85 B2.n1 B2.t2 169.237
R86 B2.n0 B2.t0 169.237
R87 B2.n2 B2.n1 152
R88 B2 B2.n2 6.87457
R89 VGND.n6 VGND.n4 207.965
R90 VGND.n17 VGND.n16 185
R91 VGND.n15 VGND.n14 185
R92 VGND.n5 VGND.t4 174.004
R93 VGND.n19 VGND.t0 154.458
R94 VGND.n16 VGND.n15 96.0005
R95 VGND.n8 VGND.n7 34.6358
R96 VGND.n8 VGND.n2 34.6358
R97 VGND.n4 VGND.t2 33.2313
R98 VGND.n4 VGND.t3 31.3851
R99 VGND.n14 VGND.n2 28.4299
R100 VGND.n7 VGND.n6 27.4829
R101 VGND.n18 VGND.n17 26.924
R102 VGND.n19 VGND.n18 25.224
R103 VGND.n15 VGND.t1 24.9236
R104 VGND.n16 VGND.t5 24.9236
R105 VGND.n6 VGND.n5 14.7279
R106 VGND.n20 VGND.n19 9.3005
R107 VGND.n7 VGND.n3 9.3005
R108 VGND.n9 VGND.n8 9.3005
R109 VGND.n10 VGND.n2 9.3005
R110 VGND.n13 VGND.n12 9.3005
R111 VGND.n11 VGND.n1 9.3005
R112 VGND.n18 VGND.n0 9.3005
R113 VGND.n13 VGND.n1 9.2005
R114 VGND.n17 VGND.n1 0.8005
R115 VGND.n14 VGND.n13 0.4005
R116 VGND.n5 VGND.n3 0.173395
R117 VGND.n9 VGND.n3 0.120292
R118 VGND.n10 VGND.n9 0.120292
R119 VGND.n12 VGND.n10 0.120292
R120 VGND.n12 VGND.n11 0.120292
R121 VGND.n11 VGND.n0 0.120292
R122 VGND.n20 VGND.n0 0.120292
R123 VGND VGND.n20 0.0213333
R124 A1.n0 A1.t1 212.081
R125 A1.n1 A1.t2 212.081
R126 A1 A1.n2 157.12
R127 A1.n0 A1.t3 139.78
R128 A1.n1 A1.t0 139.78
R129 A1.n2 A1.n0 30.6732
R130 A1.n2 A1.n1 30.6732
R131 a_735_47.n1 a_735_47.n0 326.865
R132 a_735_47.n0 a_735_47.t3 24.9236
R133 a_735_47.n0 a_735_47.t0 24.9236
R134 a_735_47.t1 a_735_47.n1 24.9236
R135 a_735_47.n1 a_735_47.t2 24.9236
R136 C1.n0 C1.t3 212.081
R137 C1.n1 C1.t0 212.081
R138 C1.n2 C1.n1 184.864
R139 C1.n0 C1.t1 139.78
R140 C1.n1 C1.t2 139.78
R141 C1.n1 C1.n0 61.346
R142 C1.n2 C1 11.055
R143 C1 C1.n2 2.13383
C0 VPB B2 0.067882f
C1 Y VPWR 0.012872f
C2 A1 VGND 0.017496f
C3 VPB B1 0.050999f
C4 C1 B2 0.0205f
C5 Y VGND 0.258389f
C6 VPB A2 0.070852f
C7 VPWR VGND 0.106412f
C8 VPB A1 0.050973f
C9 B2 B1 0.212706f
C10 B2 A2 0.092645f
C11 VPB Y 0.008117f
C12 C1 Y 0.105935f
C13 VPB VPWR 0.108288f
C14 B2 Y 0.118455f
C15 VPB VGND 0.009915f
C16 C1 VPWR 0.01915f
C17 B1 Y 0.064327f
C18 A2 A1 0.207246f
C19 B2 VPWR 0.022429f
C20 C1 VGND 0.063196f
C21 A2 Y 0.045548f
C22 B1 VPWR 0.015218f
C23 B2 VGND 0.03252f
C24 A1 Y 0.048298f
C25 A2 VPWR 0.045465f
C26 B1 VGND 0.018426f
C27 VPB C1 0.077955f
C28 A2 VGND 0.056836f
C29 A1 VPWR 0.029814f
C30 VGND VNB 0.681558f
C31 VPWR VNB 0.520019f
C32 Y VNB 0.037888f
C33 A1 VNB 0.166288f
C34 A2 VNB 0.230015f
C35 B1 VNB 0.166404f
C36 B2 VNB 0.19461f
C37 C1 VNB 0.254689f
C38 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221oi_4 VNB VPB VPWR VGND C1 Y B2 B1 A2 A1
X0 Y.t12 A1.t0 a_1241_47.t7 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_453_47.t4 B2.t0 VGND.t10 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t6 B1.t0 a_453_47.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X3 Y.t11 A1.t1 a_1241_47.t6 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t7 C1.t0 a_27_297.t11 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_297.t15 A2.t0 VPWR.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X6 Y.t13 B1.t1 a_453_47.t5 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t11 A2.t1 a_1241_47.t3 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t8 C1.t1 VGND.t6 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297.t10 C1.t2 Y.t5 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR.t6 A2.t2 a_471_297.t14 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X11 a_453_47.t6 B1.t2 Y.t14 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_471_297.t7 B2.t1 a_27_297.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND.t9 B2.t2 a_453_47.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_1241_47.t5 A1.t2 Y.t10 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_27_297.t6 B2.t3 a_471_297.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 a_453_47.t7 B1.t3 Y.t15 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_1241_47.t4 A1.t3 Y.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t2 C1.t3 Y.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_1241_47.t2 A2.t3 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y.t1 C1.t4 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 VGND.t4 C1.t5 Y.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR.t5 A2.t4 a_471_297.t13 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_471_297.t5 B2.t4 a_27_297.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X24 a_471_297.t12 A2.t5 VPWR.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_471_297.t3 B1.t4 a_27_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR.t3 A1.t4 a_471_297.t11 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y.t3 C1.t6 a_27_297.t9 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X28 a_27_297.t0 B1.t5 a_471_297.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND.t1 A2.t6 a_1241_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_471_297.t10 A1.t5 VPWR.t2 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_27_297.t3 B1.t6 a_471_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_1241_47.t0 A2.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X33 a_471_297.t0 B1.t7 a_27_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 VPWR.t1 A1.t6 a_471_297.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_27_297.t4 B2.t5 a_471_297.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_471_297.t8 A1.t7 VPWR.t0 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_27_297.t8 C1.t7 Y.t4 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 a_453_47.t2 B2.t6 VGND.t8 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X39 VGND.t7 B2.t7 a_453_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A1.n3 A1.t4 212.081
R1 A1.n5 A1.t5 212.081
R2 A1.n7 A1.t6 212.081
R3 A1.n1 A1.t7 212.081
R4 A1.n4 A1.n0 173.761
R5 A1.n9 A1.n2 173.761
R6 A1.n6 A1.n0 152
R7 A1.n9 A1.n8 152
R8 A1.n3 A1.t3 139.78
R9 A1.n5 A1.t1 139.78
R10 A1.n7 A1.t2 139.78
R11 A1.n1 A1.t0 139.78
R12 A1.n8 A1.n6 49.6611
R13 A1.n7 A1.n2 48.2005
R14 A1.n5 A1.n4 39.4369
R15 A1.n4 A1.n3 21.9096
R16 A1 A1.n0 16.0005
R17 A1.n2 A1.n1 13.146
R18 A1.n6 A1.n5 10.2247
R19 A1 A1.n9 5.7605
R20 A1.n8 A1.n7 1.46111
R21 a_1241_47.n5 a_1241_47.n4 233.874
R22 a_1241_47.n4 a_1241_47.n3 185
R23 a_1241_47.n2 a_1241_47.n0 147.915
R24 a_1241_47.n2 a_1241_47.n1 88.3446
R25 a_1241_47.n4 a_1241_47.n2 53.5212
R26 a_1241_47.n3 a_1241_47.t6 24.9236
R27 a_1241_47.n3 a_1241_47.t5 24.9236
R28 a_1241_47.n1 a_1241_47.t3 24.9236
R29 a_1241_47.n1 a_1241_47.t4 24.9236
R30 a_1241_47.n0 a_1241_47.t1 24.9236
R31 a_1241_47.n0 a_1241_47.t2 24.9236
R32 a_1241_47.n5 a_1241_47.t7 24.9236
R33 a_1241_47.t0 a_1241_47.n5 24.9236
R34 Y.n9 Y.n8 355.233
R35 Y.n9 Y.n7 297.045
R36 Y.n2 Y.n0 246.44
R37 Y.n10 Y.n6 197.315
R38 Y.n2 Y.n1 185
R39 Y.n4 Y.n3 185
R40 Y.n6 Y.n5 185
R41 Y.n13 Y.n11 135.249
R42 Y.n4 Y.n2 121.915
R43 Y.n13 Y.n12 98.982
R44 Y.n6 Y.n4 61.4405
R45 Y.n8 Y.t5 26.5955
R46 Y.n8 Y.t3 26.5955
R47 Y.n7 Y.t4 26.5955
R48 Y.n7 Y.t7 26.5955
R49 Y.n5 Y.t15 24.9236
R50 Y.n5 Y.t6 24.9236
R51 Y.n3 Y.t14 24.9236
R52 Y.n3 Y.t13 24.9236
R53 Y.n1 Y.t10 24.9236
R54 Y.n1 Y.t12 24.9236
R55 Y.n0 Y.t9 24.9236
R56 Y.n0 Y.t11 24.9236
R57 Y.n12 Y.t2 24.9236
R58 Y.n12 Y.t8 24.9236
R59 Y.n11 Y.t0 24.9236
R60 Y.n11 Y.t1 24.9236
R61 Y.n10 Y.n9 21.5346
R62 Y Y.n13 16.2914
R63 Y Y.n10 5.1205
R64 VNB.t10 VNB.t8 2620.06
R65 VNB.t3 VNB.t0 1423.95
R66 VNB.t6 VNB.t2 1253.07
R67 VNB.t7 VNB.t1 1196.12
R68 VNB.t12 VNB.t7 1196.12
R69 VNB.t13 VNB.t12 1196.12
R70 VNB.t15 VNB.t13 1196.12
R71 VNB.t14 VNB.t15 1196.12
R72 VNB.t16 VNB.t14 1196.12
R73 VNB.t0 VNB.t16 1196.12
R74 VNB.t18 VNB.t3 1196.12
R75 VNB.t17 VNB.t18 1196.12
R76 VNB.t19 VNB.t17 1196.12
R77 VNB.t8 VNB.t19 1196.12
R78 VNB.t11 VNB.t10 1196.12
R79 VNB.t2 VNB.t11 1196.12
R80 VNB.t9 VNB.t6 1196.12
R81 VNB.t4 VNB.t9 1196.12
R82 VNB.t5 VNB.t4 1196.12
R83 VNB VNB.t5 968.285
R84 B2 B2.n0 287.952
R85 B2.n0 B2.t4 241.536
R86 B2.n5 B2.t5 216.463
R87 B2.n4 B2.t1 212.081
R88 B2.n2 B2.t3 212.081
R89 B2.n1 B2.t6 201.125
R90 B2 B2.n5 180.817
R91 B2.n0 B2.t7 169.237
R92 B2.n1 B2.t2 139.78
R93 B2.n3 B2.t0 139.78
R94 B2.n5 B2.n4 56.9641
R95 B2.n3 B2.n2 49.6611
R96 B2.n4 B2.n3 11.6853
R97 B2.n2 B2.n1 11.6853
R98 VGND.n36 VGND.n34 243.514
R99 VGND.n13 VGND.n11 207.965
R100 VGND.n21 VGND.n8 207.965
R101 VGND.n43 VGND.n1 207.965
R102 VGND.n36 VGND.n35 185
R103 VGND.n12 VGND.t1 172.655
R104 VGND.n45 VGND.t3 153.107
R105 VGND.n8 VGND.t7 39.6928
R106 VGND.n15 VGND.n14 34.6358
R107 VGND.n15 VGND.n9 34.6358
R108 VGND.n19 VGND.n9 34.6358
R109 VGND.n20 VGND.n19 34.6358
R110 VGND.n22 VGND.n6 34.6358
R111 VGND.n26 VGND.n6 34.6358
R112 VGND.n27 VGND.n26 34.6358
R113 VGND.n28 VGND.n27 34.6358
R114 VGND.n28 VGND.n4 34.6358
R115 VGND.n32 VGND.n4 34.6358
R116 VGND.n33 VGND.n32 34.6358
R117 VGND.n38 VGND.n33 34.6358
R118 VGND.n42 VGND.n2 34.6358
R119 VGND.n44 VGND.n43 32.377
R120 VGND.n14 VGND.n13 29.3652
R121 VGND.n35 VGND.t8 28.6159
R122 VGND.n37 VGND.n2 26.3534
R123 VGND.n11 VGND.t5 24.9236
R124 VGND.n11 VGND.t11 24.9236
R125 VGND.n8 VGND.t0 24.9236
R126 VGND.n35 VGND.t4 24.9236
R127 VGND.n34 VGND.t10 24.9236
R128 VGND.n34 VGND.t9 24.9236
R129 VGND.n1 VGND.t6 24.9236
R130 VGND.n1 VGND.t2 24.9236
R131 VGND.n45 VGND.n44 24.4711
R132 VGND.n37 VGND.n36 22.9652
R133 VGND.n21 VGND.n20 21.8358
R134 VGND.n22 VGND.n21 12.8005
R135 VGND.n13 VGND.n12 12.2291
R136 VGND.n46 VGND.n45 9.3005
R137 VGND.n14 VGND.n10 9.3005
R138 VGND.n16 VGND.n15 9.3005
R139 VGND.n17 VGND.n9 9.3005
R140 VGND.n19 VGND.n18 9.3005
R141 VGND.n20 VGND.n7 9.3005
R142 VGND.n23 VGND.n22 9.3005
R143 VGND.n24 VGND.n6 9.3005
R144 VGND.n26 VGND.n25 9.3005
R145 VGND.n27 VGND.n5 9.3005
R146 VGND.n29 VGND.n28 9.3005
R147 VGND.n30 VGND.n4 9.3005
R148 VGND.n32 VGND.n31 9.3005
R149 VGND.n33 VGND.n3 9.3005
R150 VGND.n39 VGND.n38 9.3005
R151 VGND.n40 VGND.n2 9.3005
R152 VGND.n42 VGND.n41 9.3005
R153 VGND.n44 VGND.n0 9.3005
R154 VGND.n38 VGND.n37 8.28285
R155 VGND.n43 VGND.n42 2.25932
R156 VGND.n12 VGND.n10 0.791449
R157 VGND.n16 VGND.n10 0.120292
R158 VGND.n17 VGND.n16 0.120292
R159 VGND.n18 VGND.n17 0.120292
R160 VGND.n18 VGND.n7 0.120292
R161 VGND.n23 VGND.n7 0.120292
R162 VGND.n24 VGND.n23 0.120292
R163 VGND.n25 VGND.n24 0.120292
R164 VGND.n25 VGND.n5 0.120292
R165 VGND.n29 VGND.n5 0.120292
R166 VGND.n30 VGND.n29 0.120292
R167 VGND.n31 VGND.n30 0.120292
R168 VGND.n31 VGND.n3 0.120292
R169 VGND.n39 VGND.n3 0.120292
R170 VGND.n40 VGND.n39 0.120292
R171 VGND.n41 VGND.n40 0.120292
R172 VGND.n41 VGND.n0 0.120292
R173 VGND.n46 VGND.n0 0.120292
R174 VGND VGND.n46 0.0213333
R175 a_453_47.n6 a_453_47.n5 241.145
R176 a_453_47.n3 a_453_47.n1 233.874
R177 a_453_47.n3 a_453_47.n2 185
R178 a_453_47.n7 a_453_47.n6 185
R179 a_453_47.n4 a_453_47.n0 185
R180 a_453_47.n7 a_453_47.n0 92.3082
R181 a_453_47.n4 a_453_47.n3 48.8732
R182 a_453_47.n6 a_453_47.n4 29.0914
R183 a_453_47.n2 a_453_47.t5 24.9236
R184 a_453_47.n2 a_453_47.t7 24.9236
R185 a_453_47.n1 a_453_47.t1 24.9236
R186 a_453_47.n1 a_453_47.t6 24.9236
R187 a_453_47.n5 a_453_47.t3 24.9236
R188 a_453_47.n5 a_453_47.t2 24.9236
R189 a_453_47.n0 a_453_47.t0 24.9236
R190 a_453_47.t4 a_453_47.n7 24.9236
R191 B1.n2 B1.t5 212.081
R192 B1.n1 B1.t4 212.081
R193 B1.n7 B1.t6 212.081
R194 B1.n8 B1.t7 212.081
R195 B1.n4 B1.n3 167.543
R196 B1 B1.n9 161.601
R197 B1.n5 B1.n4 152
R198 B1.n6 B1.n0 152
R199 B1.n2 B1.t2 139.78
R200 B1.n1 B1.t1 139.78
R201 B1.n7 B1.t3 139.78
R202 B1.n8 B1.t0 139.78
R203 B1.n6 B1.n5 49.6611
R204 B1.n3 B1.n1 48.2005
R205 B1.n9 B1.n7 39.4369
R206 B1.n9 B1.n8 21.9096
R207 B1.n4 B1.n0 15.5434
R208 B1.n3 B1.n2 13.146
R209 B1.n7 B1.n6 10.2247
R210 B1 B1.n0 5.94336
R211 B1.n5 B1.n1 1.46111
R212 C1.n3 C1.t6 212.081
R213 C1.n0 C1.t7 212.081
R214 C1.n1 C1.t0 212.081
R215 C1.n4 C1.t2 212.081
R216 C1 C1.n2 158.4
R217 C1.n3 C1.t4 139.78
R218 C1.n0 C1.t5 139.78
R219 C1.n1 C1.t1 139.78
R220 C1.n4 C1.t3 139.78
R221 C1 C1.n5 85.7128
R222 C1.n1 C1.n0 61.346
R223 C1.n4 C1.n2 37.9763
R224 C1.n5 C1.n4 31.7924
R225 C1.n2 C1.n1 23.3702
R226 C1.n5 C1.n3 22.986
R227 a_27_297.n2 a_27_297.n0 636.201
R228 a_27_297.n2 a_27_297.n1 585
R229 a_27_297.n4 a_27_297.n3 585
R230 a_27_297.n9 a_27_297.n8 300.885
R231 a_27_297.n6 a_27_297.n5 289.288
R232 a_27_297.n8 a_27_297.t9 276.781
R233 a_27_297.n7 a_27_297.t8 214.101
R234 a_27_297.n7 a_27_297.n6 78.7175
R235 a_27_297.n8 a_27_297.n7 67.9256
R236 a_27_297.n4 a_27_297.n2 51.2005
R237 a_27_297.n6 a_27_297.n4 50.1433
R238 a_27_297.n5 a_27_297.t7 26.5955
R239 a_27_297.n5 a_27_297.t6 26.5955
R240 a_27_297.n3 a_27_297.t2 26.5955
R241 a_27_297.n3 a_27_297.t4 26.5955
R242 a_27_297.n1 a_27_297.t1 26.5955
R243 a_27_297.n1 a_27_297.t3 26.5955
R244 a_27_297.n0 a_27_297.t5 26.5955
R245 a_27_297.n0 a_27_297.t0 26.5955
R246 a_27_297.n9 a_27_297.t11 26.5955
R247 a_27_297.t10 a_27_297.n9 26.5955
R248 VPB.t16 VPB.t9 556.386
R249 VPB.t8 VPB.t0 295.95
R250 VPB.t2 VPB.t11 248.599
R251 VPB.t1 VPB.t2 248.599
R252 VPB.t15 VPB.t1 248.599
R253 VPB.t14 VPB.t15 248.599
R254 VPB.t13 VPB.t14 248.599
R255 VPB.t12 VPB.t13 248.599
R256 VPB.t0 VPB.t12 248.599
R257 VPB.t5 VPB.t8 248.599
R258 VPB.t6 VPB.t5 248.599
R259 VPB.t4 VPB.t6 248.599
R260 VPB.t3 VPB.t4 248.599
R261 VPB.t7 VPB.t3 248.599
R262 VPB.t10 VPB.t7 248.599
R263 VPB.t9 VPB.t10 248.599
R264 VPB.t19 VPB.t16 248.599
R265 VPB.t18 VPB.t19 248.599
R266 VPB.t17 VPB.t18 248.599
R267 VPB VPB.t17 201.246
R268 A2.n6 A2.n2 330.041
R269 A2.n2 A2.t2 241.536
R270 A2.n0 A2.t0 212.081
R271 A2.n3 A2.t4 212.081
R272 A2.n4 A2.t5 212.081
R273 A2.n2 A2.t7 169.237
R274 A2.n6 A2.n5 152
R275 A2.n0 A2.t6 139.78
R276 A2.n3 A2.t3 139.78
R277 A2.n4 A2.t1 139.78
R278 A2 A2.n1 83.7928
R279 A2.n5 A2.n3 48.2005
R280 A2.n1 A2.n0 33.2102
R281 A2.n3 A2.n1 21.5682
R282 A2.n5 A2.n4 13.146
R283 A2 A2.n6 8.3205
R284 VPWR.n6 VPWR.n5 585
R285 VPWR.n2 VPWR.n1 585
R286 VPWR.n13 VPWR.n12 585
R287 VPWR.n4 VPWR.n3 334.358
R288 VPWR.n12 VPWR.t0 26.5955
R289 VPWR.n12 VPWR.t6 26.5955
R290 VPWR.n1 VPWR.t2 26.5955
R291 VPWR.n1 VPWR.t1 26.5955
R292 VPWR.n5 VPWR.t4 26.5955
R293 VPWR.n5 VPWR.t3 26.5955
R294 VPWR.n3 VPWR.t7 26.5955
R295 VPWR.n3 VPWR.t5 26.5955
R296 VPWR.n14 VPWR.n13 10.3574
R297 VPWR.n11 VPWR.n10 9.98016
R298 VPWR.n7 VPWR.n6 9.32931
R299 VPWR.n8 VPWR.n7 9.3005
R300 VPWR.n10 VPWR.n9 9.3005
R301 VPWR.n11 VPWR.n0 9.3005
R302 VPWR.n7 VPWR.n2 8.89541
R303 VPWR.n6 VPWR.n4 7.37597
R304 VPWR.n13 VPWR.n11 7.15982
R305 VPWR VPWR.n14 1.55849
R306 VPWR.n10 VPWR.n2 1.08525
R307 VPWR.n8 VPWR.n4 0.750813
R308 VPWR.n14 VPWR.n0 0.148181
R309 VPWR.n9 VPWR.n8 0.120292
R310 VPWR.n9 VPWR.n0 0.120292
R311 a_471_297.n3 a_471_297.n2 585
R312 a_471_297.n5 a_471_297.n4 585
R313 a_471_297.n11 a_471_297.n10 585
R314 a_471_297.n9 a_471_297.n8 585
R315 a_471_297.n13 a_471_297.n12 585
R316 a_471_297.n9 a_471_297.t6 365.832
R317 a_471_297.n1 a_471_297.t15 300.164
R318 a_471_297.n1 a_471_297.n0 297.224
R319 a_471_297.n7 a_471_297.n6 290.341
R320 a_471_297.n12 a_471_297.n7 49.3769
R321 a_471_297.n7 a_471_297.n5 47.6439
R322 a_471_297.n12 a_471_297.n11 43.0085
R323 a_471_297.n11 a_471_297.n9 43.0085
R324 a_471_297.n3 a_471_297.n1 41.3543
R325 a_471_297.n5 a_471_297.n3 41.3543
R326 a_471_297.n6 a_471_297.t14 34.4755
R327 a_471_297.n6 a_471_297.t5 34.4755
R328 a_471_297.n8 a_471_297.t4 26.5955
R329 a_471_297.n8 a_471_297.t7 26.5955
R330 a_471_297.n10 a_471_297.t1 26.5955
R331 a_471_297.n10 a_471_297.t0 26.5955
R332 a_471_297.n4 a_471_297.t9 26.5955
R333 a_471_297.n4 a_471_297.t8 26.5955
R334 a_471_297.n2 a_471_297.t11 26.5955
R335 a_471_297.n2 a_471_297.t10 26.5955
R336 a_471_297.n0 a_471_297.t13 26.5955
R337 a_471_297.n0 a_471_297.t12 26.5955
R338 a_471_297.n13 a_471_297.t2 26.5955
R339 a_471_297.t3 a_471_297.n13 26.5955
C0 VPB C1 0.128784f
C1 A2 VGND 0.08708f
C2 A1 VPWR 0.055217f
C3 VPB B2 0.151139f
C4 Y VPWR 0.025861f
C5 A1 VGND 0.036104f
C6 C1 B2 0.037426f
C7 VPB B1 0.114759f
C8 Y VGND 0.4808f
C9 VPB A2 0.132822f
C10 VPWR VGND 0.185158f
C11 B2 B1 0.294532f
C12 VPB A1 0.114794f
C13 B2 A2 0.092645f
C14 VPB Y 0.012762f
C15 C1 Y 0.289193f
C16 VPB VPWR 0.170347f
C17 B1 A2 5.11e-19
C18 B1 A1 5.76e-19
C19 VPB VGND 0.012903f
C20 C1 VPWR 0.035232f
C21 B2 Y 0.162512f
C22 B2 VPWR 0.03772f
C23 B1 Y 0.139666f
C24 C1 VGND 0.092729f
C25 A2 A1 0.291503f
C26 A2 Y 0.044418f
C27 B2 VGND 0.074372f
C28 B1 VPWR 0.025483f
C29 A1 Y 0.11358f
C30 A2 VPWR 0.082987f
C31 B1 VGND 0.031948f
C32 VGND VNB 1.09533f
C33 VPWR VNB 0.857945f
C34 Y VNB 0.03722f
C35 A1 VNB 0.352953f
C36 A2 VNB 0.404149f
C37 B1 VNB 0.355499f
C38 B2 VNB 0.409277f
C39 C1 VNB 0.400609f
C40 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a222oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a222oi_1 VNB VPB VPWR VGND C2 C1 B1 A2 A1 Y B2
X0 Y.t4 B1.t0 a_393_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1056 pd=0.97 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 VGND.t1 A2.t0 a_561_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1664 pd=1.8 as=0.1056 ps=0.97 w=0.64 l=0.15
X2 VGND.t2 C2.t0 a_109_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.2912 pd=1.55 as=0.0672 ps=0.85 w=0.64 l=0.15
X3 Y.t1 C2.t1 a_109_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t0 A1.t0 a_311_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 a_311_297.t3 A2.t1 VPWR.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X6 a_311_297.t1 B1.t1 a_109_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_297.t3 B2.t0 a_311_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 a_109_297.t0 C1.t0 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_393_47.t1 B2.t1 VGND.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0672 pd=0.85 as=0.2912 ps=1.55 w=0.64 l=0.15
X10 a_109_47.t1 C1.t1 Y.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_561_47.t0 A1.t1 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=0.15
R0 B1.n0 B1.t1 239.929
R1 B1.n0 B1.t0 172.45
R2 B1 B1.n0 155.298
R3 a_393_47.t0 a_393_47.t1 39.3755
R4 Y.n0 Y.t1 827.462
R5 Y.n0 Y.t0 290.8
R6 Y.n2 Y.t2 197.764
R7 Y.n2 Y.n1 158.645
R8 Y Y.n0 44.5244
R9 Y.n1 Y.t3 32.813
R10 Y.n1 Y.t4 29.063
R11 Y Y.n2 20.4805
R12 VNB.t5 VNB.t4 3018.77
R13 VNB.t2 VNB.t0 1366.99
R14 VNB.t3 VNB.t2 1366.99
R15 VNB VNB.t1 1338.51
R16 VNB.t4 VNB.t3 1025.24
R17 VNB.t1 VNB.t5 1025.24
R18 A2.n0 A2.t1 239.929
R19 A2.n0 A2.t0 172.45
R20 A2 A2.n0 155.577
R21 a_561_47.t0 a_561_47.t1 61.8755
R22 VGND.n4 VGND.n3 185
R23 VGND.n2 VGND.n0 185
R24 VGND.n1 VGND.t1 157.065
R25 VGND.n3 VGND.t0 81.563
R26 VGND.n3 VGND.n2 63.7505
R27 VGND.n7 VGND.n0 25.4285
R28 VGND.n2 VGND.t2 25.313
R29 VGND.n4 VGND.n1 13.2007
R30 VGND.n6 VGND.n5 9.3005
R31 VGND.n5 VGND.n4 5.35323
R32 VGND.n5 VGND.n0 2.5605
R33 VGND.n6 VGND.n1 0.160392
R34 VGND VGND.n7 0.159538
R35 VGND.n7 VGND.n6 0.141672
R36 C2.n0 C2.t1 239.929
R37 C2.n0 C2.t0 172.45
R38 C2 C2.n0 154.595
R39 a_109_47.t0 a_109_47.t1 39.3755
R40 a_109_297.n1 a_109_297.n0 989.582
R41 a_109_297.n0 a_109_297.t2 26.5955
R42 a_109_297.n0 a_109_297.t3 26.5955
R43 a_109_297.n1 a_109_297.t1 26.5955
R44 a_109_297.t0 a_109_297.n1 26.5955
R45 VPB.t2 VPB.t4 591.9
R46 VPB.t0 VPB.t5 284.113
R47 VPB VPB.t1 278.193
R48 VPB.t3 VPB.t0 248.599
R49 VPB.t4 VPB.t3 248.599
R50 VPB.t1 VPB.t2 248.599
R51 A1.n0 A1.t0 239.929
R52 A1.n0 A1.t1 172.45
R53 A1 A1.n0 155.298
R54 a_311_297.n0 a_311_297.t2 703.569
R55 a_311_297.n0 a_311_297.t3 288.2
R56 a_311_297.n1 a_311_297.n0 201.549
R57 a_311_297.t0 a_311_297.n1 26.5955
R58 a_311_297.n1 a_311_297.t1 26.5955
R59 VPWR VPWR.n0 329.954
R60 VPWR.n0 VPWR.t1 38.4155
R61 VPWR.n0 VPWR.t0 26.5955
R62 B2.n0 B2.t0 236.129
R63 B2.n0 B2.t1 168.649
R64 B2 B2.n0 155.097
R65 C1.n0 C1.t0 228.548
R66 C1 C1.n0 161.143
R67 C1.n0 C1.t1 161.069
C0 VGND VPB 0.009426f
C1 Y C2 0.109178f
C2 A1 B1 0.081893f
C3 VPWR C1 0.012288f
C4 VPB C1 0.037942f
C5 Y B2 0.067414f
C6 VPWR C2 0.008764f
C7 VGND C1 0.014297f
C8 VPB C2 0.031476f
C9 VPWR B2 0.008595f
C10 VGND C2 0.016538f
C11 Y B1 0.038241f
C12 VPB B2 0.033242f
C13 C1 C2 0.087708f
C14 VPWR B1 0.01154f
C15 VGND B2 0.01589f
C16 VPB B1 0.025462f
C17 VGND B1 0.012999f
C18 A1 A2 0.078822f
C19 C2 B2 0.018479f
C20 A1 Y 0.007758f
C21 A1 VPWR 0.018515f
C22 A2 Y 0.002153f
C23 B2 B1 0.088958f
C24 A1 VPB 0.02637f
C25 A2 VPWR 0.016804f
C26 A1 VGND 0.024359f
C27 A2 VPB 0.030658f
C28 Y VPWR 0.055639f
C29 A2 VGND 0.040274f
C30 Y VPB 0.025848f
C31 Y VGND 0.258587f
C32 VPWR VPB 0.075432f
C33 Y C1 0.106923f
C34 VPWR VGND 0.071744f
C35 VGND VNB 0.463522f
C36 VPWR VNB 0.366504f
C37 Y VNB 0.099097f
C38 A2 VNB 0.131451f
C39 A1 VNB 0.09053f
C40 B1 VNB 0.088501f
C41 B2 VNB 0.101783f
C42 C2 VNB 0.099112f
C43 C1 VNB 0.145879f
C44 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 VNB VPB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_75_199.t1 C1.t0 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X1 a_208_47.t0 A3.t0 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X2 a_315_47.t0 A2.t0 a_208_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 VGND.t0 B1.t0 a_75_199.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_75_199.t3 A1.t0 a_315_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199.t2 C1.t1 a_544_297.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X6 a_544_297.t1 B1.t1 a_201_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X7 VPWR.t3 a_75_199.t4 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297.t0 A3.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X9 VPWR.t1 A2.t1 a_201_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297.t2 A1.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND.t1 a_75_199.t5 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C1.n0 C1.t1 230.363
R1 C1.n0 C1.t0 158.064
R2 C1 C1.n0 154.91
R3 VGND.n2 VGND.n0 206.764
R4 VGND.n2 VGND.n1 205.406
R5 VGND.n0 VGND.t0 38.7697
R6 VGND.n1 VGND.t1 38.7697
R7 VGND.n0 VGND.t2 37.8467
R8 VGND.n1 VGND.t3 24.9236
R9 VGND VGND.n2 0.160517
R10 a_75_199.t2 a_75_199.n3 575.749
R11 a_75_199.n1 a_75_199.t1 360.675
R12 a_75_199.n2 a_75_199.t4 241.536
R13 a_75_199.n1 a_75_199.n0 185
R14 a_75_199.n3 a_75_199.n1 169.448
R15 a_75_199.n2 a_75_199.t5 169.237
R16 a_75_199.n3 a_75_199.n2 152
R17 a_75_199.n0 a_75_199.t3 30.462
R18 a_75_199.n0 a_75_199.t0 29.539
R19 VNB.t2 VNB.t3 1908.09
R20 VNB.t0 VNB.t1 1609.06
R21 VNB.t5 VNB.t2 1523.62
R22 VNB.t4 VNB.t5 1409.71
R23 VNB.t3 VNB.t0 1352.75
R24 VNB VNB.t4 925.567
R25 A3.n0 A3.t1 241.536
R26 A3.n0 A3.t0 169.237
R27 A3 A3.n0 154.91
R28 a_208_47.t0 a_208_47.t1 71.0774
R29 A2.n0 A2.t1 231.017
R30 A2.n0 A2.t0 158.716
R31 A2 A2.n0 155.611
R32 a_315_47.t0 a_315_47.t1 96.0005
R33 B1.n0 B1.t1 241.536
R34 B1.n0 B1.t0 169.237
R35 B1 B1.n0 159.758
R36 A1.n0 A1.t1 241.536
R37 A1.n0 A1.t0 169.237
R38 A1.n1 A1.n0 158.4
R39 A1.n1 A1 15.4952
R40 A1 A1.n1 2.90959
R41 a_544_297.t0 a_544_297.t1 81.7555
R42 VPB.t1 VPB.t2 449.844
R43 VPB.t5 VPB.t3 334.425
R44 VPB.t0 VPB.t1 284.113
R45 VPB.t2 VPB.t5 281.154
R46 VPB.t4 VPB.t0 257.478
R47 VPB VPB.t4 207.166
R48 a_201_297.n1 a_201_297.n0 674.383
R49 a_201_297.t0 a_201_297.n1 34.4755
R50 a_201_297.n0 a_201_297.t2 32.5055
R51 a_201_297.n0 a_201_297.t3 31.5205
R52 a_201_297.n1 a_201_297.t1 30.5355
R53 X.n0 X 593.095
R54 X.n1 X.n0 585
R55 X X.t0 343.892
R56 X.n0 X.t1 31.5205
R57 X X.n1 8.09462
R58 X.n1 X 4.70638
R59 VPWR.n9 VPWR.n1 604.854
R60 VPWR.n3 VPWR.n2 585
R61 VPWR.n5 VPWR.n4 585
R62 VPWR.n4 VPWR.n3 66.9805
R63 VPWR.n1 VPWR.t0 29.5505
R64 VPWR.n4 VPWR.t2 26.5955
R65 VPWR.n3 VPWR.t1 26.5955
R66 VPWR.n1 VPWR.t3 26.5955
R67 VPWR.n8 VPWR.n7 26.5725
R68 VPWR.n9 VPWR.n8 23.3417
R69 VPWR.n6 VPWR.n5 10.2088
R70 VPWR.n7 VPWR.n6 9.3005
R71 VPWR.n8 VPWR.n0 9.3005
R72 VPWR.n5 VPWR.n2 7.91323
R73 VPWR.n10 VPWR.n9 7.4049
R74 VPWR.n7 VPWR.n2 0.233227
R75 VPWR.n10 VPWR.n0 0.144904
R76 VPWR.n6 VPWR.n0 0.120292
R77 VPWR VPWR.n10 0.118504
C0 VPWR B1 0.012527f
C1 VGND A1 0.011328f
C2 X VGND 0.060935f
C3 VGND B1 0.017055f
C4 VPWR VGND 0.07349f
C5 VPB A3 0.026815f
C6 VPB A2 0.037631f
C7 C1 VPB 0.039357f
C8 VPB A1 0.030611f
C9 A3 A2 0.074726f
C10 X VPB 0.010651f
C11 VPB B1 0.029202f
C12 X A3 0.003171f
C13 VPWR VPB 0.074935f
C14 A2 A1 0.068871f
C15 X A2 3.01e-19
C16 VPWR A3 0.018105f
C17 C1 A1 3.21e-19
C18 VGND VPB 0.00772f
C19 C1 X 5.14e-20
C20 X A1 1.2e-19
C21 C1 B1 0.065975f
C22 VGND A3 0.01613f
C23 VPWR A2 0.017412f
C24 C1 VPWR 0.014612f
C25 A1 B1 0.071566f
C26 X B1 7.79e-20
C27 VPWR A1 0.015144f
C28 VGND A2 0.011854f
C29 C1 VGND 0.018145f
C30 X VPWR 0.067555f
C31 VGND VNB 0.436573f
C32 VPWR VNB 0.365173f
C33 X VNB 0.090646f
C34 C1 VNB 0.14827f
C35 B1 VNB 0.094718f
C36 A1 VNB 0.101248f
C37 A2 VNB 0.110292f
C38 A3 VNB 0.090791f
C39 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_2 VPB VNB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_79_21.t1 C1.t0 a_635_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR.t4 A2.t0 a_319_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND.t4 B1.t0 a_79_21.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X3 a_417_47.t1 A2.t1 a_319_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X4 a_79_21.t3 A1.t0 a_417_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X5 a_319_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR.t1 a_79_21.t4 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297.t2 A1.t1 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND.t3 a_79_21.t5 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_319_297.t0 A3.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21.t0 C1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X11 a_635_297.t1 B1.t1 a_319_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X.t2 a_79_21.t6 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X.t0 a_79_21.t7 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 C1.n0 C1.t0 236.934
R1 C1.n0 C1.t1 164.633
R2 C1 C1.n0 154.272
R3 a_635_297.t0 a_635_297.t1 82.7405
R4 a_79_21.t1 a_79_21.n4 582.112
R5 a_79_21.n1 a_79_21.t0 349.38
R6 a_79_21.n3 a_79_21.t4 212.081
R7 a_79_21.n2 a_79_21.t6 212.081
R8 a_79_21.n4 a_79_21.n1 187.107
R9 a_79_21.n1 a_79_21.n0 185
R10 a_79_21.n4 a_79_21.n3 182.673
R11 a_79_21.n3 a_79_21.t5 139.78
R12 a_79_21.n2 a_79_21.t7 139.78
R13 a_79_21.n3 a_79_21.n2 61.346
R14 a_79_21.n0 a_79_21.t3 49.8467
R15 a_79_21.n0 a_79_21.t2 25.8467
R16 VPB.t3 VPB.t0 372.897
R17 VPB.t4 VPB.t1 337.384
R18 VPB.t5 VPB.t4 337.384
R19 VPB.t6 VPB.t5 307.788
R20 VPB.t0 VPB.t6 290.031
R21 VPB.t2 VPB.t3 248.599
R22 VPB VPB.t2 189.409
R23 A2.n0 A2.t0 241.536
R24 A2.n0 A2.t1 169.237
R25 A2 A2.n0 153.423
R26 a_319_297.n1 a_319_297.n0 659.539
R27 a_319_297.n0 a_319_297.t2 50.2355
R28 a_319_297.n1 a_319_297.t3 35.4605
R29 a_319_297.n0 a_319_297.t1 32.5055
R30 a_319_297.t0 a_319_297.n1 31.5205
R31 VPWR.n4 VPWR.n3 605.235
R32 VPWR.n2 VPWR.n1 319.474
R33 VPWR.n8 VPWR.t2 249.901
R34 VPWR.n1 VPWR.t1 55.1605
R35 VPWR.n3 VPWR.t4 40.3855
R36 VPWR.n1 VPWR.t0 39.4005
R37 VPWR.n7 VPWR.n6 34.6358
R38 VPWR.n3 VPWR.t3 32.5055
R39 VPWR.n8 VPWR.n7 25.977
R40 VPWR.n4 VPWR.n2 24.0101
R41 VPWR.n6 VPWR.n5 9.3005
R42 VPWR.n7 VPWR.n0 9.3005
R43 VPWR.n9 VPWR.n8 9.3005
R44 VPWR.n5 VPWR.n4 1.00418
R45 VPWR.n6 VPWR.n2 0.753441
R46 VPWR.n5 VPWR.n0 0.120292
R47 VPWR.n9 VPWR.n0 0.120292
R48 VPWR VPWR.n9 0.0213333
R49 B1.n0 B1.t1 241.536
R50 B1.n0 B1.t0 169.237
R51 B1 B1.n0 161.31
R52 VGND.n2 VGND.n1 206.731
R53 VGND.n4 VGND.n3 199.739
R54 VGND.n6 VGND.t2 155.046
R55 VGND.n3 VGND.t0 48.9236
R56 VGND.n1 VGND.t4 40.6159
R57 VGND.n3 VGND.t3 39.6928
R58 VGND.n1 VGND.t1 38.7697
R59 VGND.n6 VGND.n5 25.977
R60 VGND.n5 VGND.n4 24.4711
R61 VGND.n7 VGND.n6 9.3005
R62 VGND.n5 VGND.n0 9.3005
R63 VGND.n4 VGND.n2 6.92355
R64 VGND.n2 VGND.n0 0.160683
R65 VGND.n7 VGND.n0 0.120292
R66 VGND VGND.n7 0.0213333
R67 VNB.t3 VNB.t0 1794.17
R68 VNB.t4 VNB.t1 1651.78
R69 VNB.t5 VNB.t4 1594.82
R70 VNB.t6 VNB.t5 1480.91
R71 VNB.t0 VNB.t6 1395.47
R72 VNB.t2 VNB.t3 1196.12
R73 VNB VNB.t2 911.327
R74 a_319_47.t0 a_319_47.t1 62.7697
R75 a_417_47.t0 a_417_47.t1 68.3082
R76 A1.n0 A1.t1 241.536
R77 A1.n0 A1.t0 169.237
R78 A1 A1.n0 154.996
R79 A3.n0 A3.t1 241.536
R80 A3.n0 A3.t0 169.237
R81 A3 A3.n0 155.274
R82 X.n3 X 593.34
R83 X.n3 X.n0 585
R84 X.n4 X.n3 585
R85 X.n1 X 186.745
R86 X.n2 X.n1 185
R87 X.n3 X.t3 26.5955
R88 X.n3 X.t2 26.5955
R89 X.n1 X.t1 24.9236
R90 X.n1 X.t0 24.9236
R91 X.n2 X 11.4429
R92 X X.n0 8.33989
R93 X.n4 X 8.33989
R94 X X.n0 4.84898
R95 X X.n4 4.84898
R96 X X.n2 1.74595
C0 A3 A2 0.07643f
C1 VPB A1 0.028933f
C2 VPWR VGND 0.097894f
C3 VPB B1 0.03006f
C4 X VGND 0.108702f
C5 A2 A1 0.089295f
C6 VPB C1 0.034532f
C7 VPB VPWR 0.092365f
C8 VPB X 0.003939f
C9 A1 B1 0.064825f
C10 A3 VPWR 0.017862f
C11 A1 C1 3.24e-19
C12 A2 VPWR 0.013275f
C13 A3 X 9.94e-19
C14 VPB VGND 0.009218f
C15 A3 VGND 0.012278f
C16 A2 X 2.73e-19
C17 A1 VPWR 0.011134f
C18 B1 C1 0.051956f
C19 B1 VPWR 0.012008f
C20 A2 VGND 0.011633f
C21 A1 X 1.43e-19
C22 A1 VGND 0.010045f
C23 B1 X 8.34e-20
C24 C1 VPWR 0.01427f
C25 VPB A3 0.029144f
C26 B1 VGND 0.015441f
C27 C1 X 5.41e-20
C28 VPB A2 0.02793f
C29 C1 VGND 0.017822f
C30 VPWR X 0.159652f
C31 VGND VNB 0.514582f
C32 X VNB 0.024364f
C33 VPWR VNB 0.446583f
C34 C1 VNB 0.139989f
C35 B1 VNB 0.097043f
C36 A1 VNB 0.099082f
C37 A2 VNB 0.093376f
C38 A3 VNB 0.091528f
C39 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_4 VNB VPB VGND VPWR A1 A2 A3 X B1 C1
X0 VPWR.t4 a_109_47.t8 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297.t2 A1.t0 VPWR.t5 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.325 ps=1.65 w=1 l=0.15
X2 X.t2 a_109_47.t9 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_861_47.t3 A3.t0 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.21125 ps=1.3 w=0.65 l=0.15
X4 a_27_297.t1 B1.t0 a_277_297.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1059_47.t3 A2.t0 a_861_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_1059_47.t1 A1.t1 a_109_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_277_297.t3 B1.t1 a_27_297.t0 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t5 a_109_47.t10 X.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X9 a_27_297.t2 C1.t0 a_109_47.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t4 a_109_47.t11 X.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.21125 pd=1.3 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND.t6 A3.t1 a_861_47.t2 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND.t8 C1.t1 a_109_47.t4 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND.t0 B1.t2 a_109_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR.t2 a_109_47.t12 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_109_47.t3 A1.t2 a_1059_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 X.t0 a_109_47.t13 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 X.t5 a_109_47.t14 VGND.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_109_47.t1 B1.t3 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X.t4 a_109_47.t15 VGND.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VPWR.t8 A3.t2 a_277_297.t6 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR.t6 A2.t1 a_277_297.t4 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.325 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47.t7 C1.t2 a_27_297.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VPWR.t7 A1.t3 a_277_297.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 a_277_297.t7 A3.t3 VPWR.t9 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_277_297.t0 A2.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X26 a_109_47.t6 C1.t3 VGND.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 a_861_47.t0 A2.t3 a_1059_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_109_47.n4 a_109_47.n2 463.873
R1 a_109_47.n15 a_109_47.n14 359.384
R2 a_109_47.n7 a_109_47.t12 221.72
R3 a_109_47.n9 a_109_47.t13 221.72
R4 a_109_47.n3 a_109_47.t8 204.173
R5 a_109_47.n1 a_109_47.t9 191.625
R6 a_109_47.n11 a_109_47.t15 179.339
R7 a_109_47.n5 a_109_47.n4 177.601
R8 a_109_47.n4 a_109_47.n3 152
R9 a_109_47.n6 a_109_47.t11 147.99
R10 a_109_47.n10 a_109_47.t10 139.78
R11 a_109_47.n8 a_109_47.t14 139.78
R12 a_109_47.n12 a_109_47.n11 132.935
R13 a_109_47.n12 a_109_47.n0 97.7187
R14 a_109_47.n14 a_109_47.n13 97.7187
R15 a_109_47.n14 a_109_47.n12 63.2476
R16 a_109_47.n9 a_109_47.n8 54.6272
R17 a_109_47.n7 a_109_47.n6 50.1827
R18 a_109_47.n5 a_109_47.n1 42.1718
R19 a_109_47.n11 a_109_47.n10 36.978
R20 a_109_47.n3 a_109_47.n1 29.9942
R21 a_109_47.t5 a_109_47.n15 26.5955
R22 a_109_47.n15 a_109_47.t7 26.5955
R23 a_109_47.n13 a_109_47.t4 24.9236
R24 a_109_47.n13 a_109_47.t6 24.9236
R25 a_109_47.n0 a_109_47.t0 24.9236
R26 a_109_47.n0 a_109_47.t1 24.9236
R27 a_109_47.n2 a_109_47.t2 24.9236
R28 a_109_47.n2 a_109_47.t3 24.9236
R29 a_109_47.n6 a_109_47.n5 15.3493
R30 a_109_47.n8 a_109_47.n7 12.8538
R31 a_109_47.n10 a_109_47.n9 12.8538
R32 X.n4 X.n3 631.307
R33 X.n4 X.n2 587.26
R34 X.n5 X.n0 137.583
R35 X.n5 X.n1 106.377
R36 X.n5 X 42.339
R37 X.n0 X.t4 28.6159
R38 X.n3 X.t3 26.5955
R39 X.n3 X.t2 26.5955
R40 X.n2 X.t1 26.5955
R41 X.n2 X.t0 26.5955
R42 X.n1 X.t6 24.9236
R43 X.n1 X.t5 24.9236
R44 X.n0 X.t7 24.9236
R45 X X.n4 12.1441
R46 X X.n5 2.29794
R47 VPWR.n19 VPWR.t1 868.721
R48 VPWR.n17 VPWR.n2 599.74
R49 VPWR.n4 VPWR.n3 599.74
R50 VPWR.n8 VPWR.n7 599.74
R51 VPWR.n12 VPWR.n6 598.511
R52 VPWR.n9 VPWR.t7 345.015
R53 VPWR.n7 VPWR.t5 101.456
R54 VPWR.n6 VPWR.t0 38.4155
R55 VPWR.n17 VPWR.n16 33.5064
R56 VPWR.n13 VPWR.n12 33.5064
R57 VPWR.n11 VPWR.n8 32.0005
R58 VPWR.n19 VPWR.n18 27.4829
R59 VPWR.n2 VPWR.t3 26.5955
R60 VPWR.n2 VPWR.t2 26.5955
R61 VPWR.n3 VPWR.t9 26.5955
R62 VPWR.n3 VPWR.t4 26.5955
R63 VPWR.n6 VPWR.t8 26.5955
R64 VPWR.n7 VPWR.t6 26.5955
R65 VPWR.n18 VPWR.n17 10.9181
R66 VPWR.n11 VPWR.n10 9.3005
R67 VPWR.n12 VPWR.n5 9.3005
R68 VPWR.n14 VPWR.n13 9.3005
R69 VPWR.n16 VPWR.n15 9.3005
R70 VPWR.n17 VPWR.n1 9.3005
R71 VPWR.n18 VPWR.n0 9.3005
R72 VPWR.n12 VPWR.n11 8.65932
R73 VPWR.n20 VPWR.n19 6.71619
R74 VPWR.n9 VPWR.n8 6.18937
R75 VPWR.n16 VPWR.n4 4.89462
R76 VPWR.n13 VPWR.n4 4.89462
R77 VPWR VPWR.n20 0.582551
R78 VPWR.n10 VPWR.n9 0.295815
R79 VPWR.n20 VPWR.n0 0.160919
R80 VPWR.n10 VPWR.n5 0.120292
R81 VPWR.n14 VPWR.n5 0.120292
R82 VPWR.n15 VPWR.n14 0.120292
R83 VPWR.n15 VPWR.n1 0.120292
R84 VPWR.n1 VPWR.n0 0.120292
R85 VPB.t8 VPB.t1 556.386
R86 VPB.t7 VPB.t6 473.521
R87 VPB.t11 VPB.t0 284.113
R88 VPB.t6 VPB.t9 248.599
R89 VPB.t0 VPB.t7 248.599
R90 VPB.t12 VPB.t11 248.599
R91 VPB.t4 VPB.t12 248.599
R92 VPB.t3 VPB.t4 248.599
R93 VPB.t2 VPB.t3 248.599
R94 VPB.t1 VPB.t2 248.599
R95 VPB.t5 VPB.t8 248.599
R96 VPB.t10 VPB.t5 248.599
R97 VPB.t13 VPB.t10 248.599
R98 VPB VPB.t13 189.409
R99 A1.n1 A1.t3 212.081
R100 A1.n0 A1.t0 212.081
R101 A1 A1.n1 185.674
R102 A1.n1 A1.t1 139.78
R103 A1.n0 A1.t2 139.78
R104 A1.n1 A1.n0 61.346
R105 a_277_297.n3 a_277_297.n2 855.802
R106 a_277_297.n5 a_277_297.n4 388.351
R107 a_277_297.n3 a_277_297.n1 296.493
R108 a_277_297.n4 a_277_297.n0 296.493
R109 a_277_297.n4 a_277_297.n3 67.7652
R110 a_277_297.n1 a_277_297.t6 26.5955
R111 a_277_297.n1 a_277_297.t7 26.5955
R112 a_277_297.n0 a_277_297.t4 26.5955
R113 a_277_297.n0 a_277_297.t0 26.5955
R114 a_277_297.n2 a_277_297.t5 26.5955
R115 a_277_297.n2 a_277_297.t3 26.5955
R116 a_277_297.n5 a_277_297.t1 26.5955
R117 a_277_297.t2 a_277_297.n5 26.5955
R118 A3.n2 A3.t2 194.407
R119 A3.n0 A3.t3 184.768
R120 A3 A3.n2 157.487
R121 A3.n0 A3.t0 149.519
R122 A3.n1 A3.t1 128.534
R123 A3.n1 A3.n0 32.1338
R124 A3.n2 A3.n1 3.21383
R125 VGND.n6 VGND.t6 297.021
R126 VGND.n27 VGND.t9 279.327
R127 VGND.n16 VGND.n4 207.213
R128 VGND.n19 VGND.n18 207.213
R129 VGND.n25 VGND.n1 207.213
R130 VGND.n10 VGND.n9 185
R131 VGND.n8 VGND.n7 185
R132 VGND.n9 VGND.n8 62.7697
R133 VGND.n15 VGND.n5 34.6358
R134 VGND.n20 VGND.n17 34.6358
R135 VGND.n24 VGND.n2 34.6358
R136 VGND.n8 VGND.t7 32.3082
R137 VGND.n7 VGND.n6 30.9984
R138 VGND.n26 VGND.n25 30.8711
R139 VGND.n27 VGND.n26 25.977
R140 VGND.n9 VGND.t4 24.9236
R141 VGND.n4 VGND.t3 24.9236
R142 VGND.n4 VGND.t5 24.9236
R143 VGND.n18 VGND.t2 24.9236
R144 VGND.n18 VGND.t0 24.9236
R145 VGND.n1 VGND.t1 24.9236
R146 VGND.n1 VGND.t8 24.9236
R147 VGND.n19 VGND.n2 24.8476
R148 VGND.n17 VGND.n16 20.3299
R149 VGND.n16 VGND.n15 14.3064
R150 VGND.n20 VGND.n19 9.78874
R151 VGND.n10 VGND.n5 9.63337
R152 VGND.n28 VGND.n27 9.3005
R153 VGND.n12 VGND.n11 9.3005
R154 VGND.n13 VGND.n5 9.3005
R155 VGND.n15 VGND.n14 9.3005
R156 VGND.n17 VGND.n3 9.3005
R157 VGND.n21 VGND.n20 9.3005
R158 VGND.n22 VGND.n2 9.3005
R159 VGND.n24 VGND.n23 9.3005
R160 VGND.n26 VGND.n0 9.3005
R161 VGND.n11 VGND.n10 5.48621
R162 VGND.n25 VGND.n24 3.76521
R163 VGND.n12 VGND.n6 1.44164
R164 VGND.n11 VGND.n7 1.42272
R165 VGND.n13 VGND.n12 0.120292
R166 VGND.n14 VGND.n13 0.120292
R167 VGND.n14 VGND.n3 0.120292
R168 VGND.n21 VGND.n3 0.120292
R169 VGND.n22 VGND.n21 0.120292
R170 VGND.n23 VGND.n22 0.120292
R171 VGND.n23 VGND.n0 0.120292
R172 VGND.n28 VGND.n0 0.120292
R173 VGND VGND.n28 0.0213333
R174 a_861_47.n1 a_861_47.n0 384.507
R175 a_861_47.n0 a_861_47.t1 24.9236
R176 a_861_47.n0 a_861_47.t0 24.9236
R177 a_861_47.t2 a_861_47.n1 24.9236
R178 a_861_47.n1 a_861_47.t3 24.9236
R179 VNB.t10 VNB.t0 2790.94
R180 VNB.t8 VNB.t11 2278.32
R181 VNB.t6 VNB.t9 1253.07
R182 VNB.t1 VNB.t2 1196.12
R183 VNB.t3 VNB.t1 1196.12
R184 VNB.t0 VNB.t3 1196.12
R185 VNB.t11 VNB.t10 1196.12
R186 VNB.t7 VNB.t8 1196.12
R187 VNB.t9 VNB.t7 1196.12
R188 VNB.t4 VNB.t6 1196.12
R189 VNB.t5 VNB.t4 1196.12
R190 VNB.t12 VNB.t5 1196.12
R191 VNB.t13 VNB.t12 1196.12
R192 VNB VNB.t13 911.327
R193 B1.n0 B1.t0 221.72
R194 B1.n1 B1.t1 221.72
R195 B1 B1.n2 168.458
R196 B1.n0 B1.t2 133.353
R197 B1.n1 B1.t3 133.353
R198 B1.n2 B1.n0 58.7443
R199 B1.n2 B1.n1 4.51925
R200 a_27_297.t1 a_27_297.n1 388.517
R201 a_27_297.n1 a_27_297.t3 388.515
R202 a_27_297.n1 a_27_297.n0 298.673
R203 a_27_297.n0 a_27_297.t0 26.5955
R204 a_27_297.n0 a_27_297.t2 26.5955
R205 A2.n3 A2.t2 252.069
R206 A2.n1 A2.t1 221.72
R207 A2.n0 A2.t0 180.661
R208 A2.n0 A2 159.619
R209 A2.n4 A2.n3 152
R210 A2.n2 A2.t3 149.421
R211 A2.n3 A2.n2 37.4894
R212 A2.n1 A2.n0 36.5968
R213 A2.n4 A2 20.1148
R214 A2 A2.n4 7.92431
R215 A2.n2 A2.n1 7.14124
R216 a_1059_47.n1 a_1059_47.t2 319.277
R217 a_1059_47.t1 a_1059_47.n1 192.446
R218 a_1059_47.n1 a_1059_47.n0 97.0637
R219 a_1059_47.n0 a_1059_47.t0 24.9236
R220 a_1059_47.n0 a_1059_47.t3 24.9236
R221 C1.n0 C1.t0 212.081
R222 C1.n1 C1.t2 212.081
R223 C1 C1.n1 186.245
R224 C1.n0 C1.t1 139.78
R225 C1.n1 C1.t3 139.78
R226 C1.n1 C1.n0 61.346
C0 VPB B1 0.063289f
C1 A1 VGND 0.020288f
C2 VPWR X 0.033277f
C3 C1 B1 0.063227f
C4 VPB A3 0.054997f
C5 VPWR VGND 0.148864f
C6 VPB A2 0.074647f
C7 X VGND 0.196358f
C8 VPB A1 0.076968f
C9 VPB VPWR 0.146584f
C10 VPB X 0.007223f
C11 A3 A2 0.047247f
C12 C1 VPWR 0.020713f
C13 B1 VPWR 0.019354f
C14 VPB VGND 0.010844f
C15 A2 A1 0.040851f
C16 A3 VPWR 0.026203f
C17 C1 VGND 0.057974f
C18 B1 X 0.004012f
C19 A3 X 0.001948f
C20 A2 VPWR 0.028252f
C21 B1 VGND 0.030654f
C22 A1 VPWR 0.070356f
C23 A3 VGND 0.033209f
C24 A2 X 4.03e-19
C25 VPB C1 0.071375f
C26 A2 VGND 0.020288f
C27 A1 X 9.42e-20
C28 VGND VNB 0.824179f
C29 X VNB 0.020587f
C30 VPWR VNB 0.691906f
C31 A1 VNB 0.24464f
C32 A2 VNB 0.212885f
C33 A3 VNB 0.190634f
C34 B1 VNB 0.173939f
C35 C1 VNB 0.25621f
C36 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311oi_1 VPB VNB Y C1 B1 A1 A2 A3 VPWR VGND
X0 Y.t2 A1.t0 a_194_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_194_47.t0 A2.t0 a_109_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2 Y.t0 C1.t0 a_376_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1725 ps=1.345 w=1 l=0.15
X3 VPWR.t0 A2.t1 a_109_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 Y.t1 C1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.112125 ps=0.995 w=0.65 l=0.15
X5 VGND.t2 B1.t0 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.115375 ps=1.005 w=0.65 l=0.15
X6 a_109_297.t1 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7 a_376_297.t1 B1.t1 a_109_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.165 ps=1.33 w=1 l=0.15
X8 a_109_297.t2 A3.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47.t1 A3.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t1 241.536
R1 A1 A1.n0 192.868
R2 A1.n0 A1.t0 169.237
R3 a_194_47.t0 a_194_47.t1 51.6928
R4 Y.n5 Y.n4 585
R5 Y.n4 Y.n0 585
R6 Y.n3 Y.n2 245.613
R7 Y.n1 Y.t1 209.923
R8 Y.n5 Y.n3 75.5456
R9 Y.n2 Y.t2 40.6159
R10 Y.n4 Y.t0 26.5955
R11 Y.n3 Y.n1 25.5928
R12 Y.n2 Y.t3 24.9236
R13 Y Y.n0 15.7338
R14 Y.n1 Y 7.05356
R15 Y.n0 Y 2.4005
R16 Y Y.n5 2.4005
R17 VNB.t2 VNB.t4 1438.19
R18 VNB.t4 VNB.t0 1409.71
R19 VNB.t1 VNB.t2 1224.6
R20 VNB.t3 VNB.t1 1210.36
R21 VNB VNB.t3 897.087
R22 A2.n0 A2.t1 241.536
R23 A2.n0 A2.t0 169.237
R24 A2.n1 A2.n0 159.565
R25 A2 A2.n1 15.0979
R26 A2.n1 A2 3.49141
R27 a_109_47.t0 a_109_47.t1 50.7697
R28 C1.n0 C1.t0 230.155
R29 C1.n0 C1.t1 157.856
R30 C1 C1.n0 154.91
R31 a_376_297.t0 a_376_297.t1 67.9655
R32 VPB.t4 VPB.t0 292.991
R33 VPB.t2 VPB.t4 284.113
R34 VPB.t1 VPB.t2 254.518
R35 VPB.t3 VPB.t1 251.559
R36 VPB VPB.t3 186.45
R37 a_109_297.n1 a_109_297.n0 981.556
R38 a_109_297.n0 a_109_297.t3 38.4155
R39 a_109_297.n1 a_109_297.t2 27.5805
R40 a_109_297.n0 a_109_297.t1 26.5955
R41 a_109_297.t0 a_109_297.n1 26.5955
R42 VPWR.n1 VPWR.n0 621.961
R43 VPWR.n1 VPWR.t2 249.887
R44 VPWR.n0 VPWR.t1 28.5655
R45 VPWR.n0 VPWR.t0 26.5955
R46 VPWR VPWR.n1 0.55971
R47 VGND.n1 VGND.n0 206.63
R48 VGND.n1 VGND.t1 156.673
R49 VGND.n0 VGND.t0 33.2313
R50 VGND.n0 VGND.t2 30.462
R51 VGND VGND.n1 0.0714683
R52 B1.n0 B1.t1 241.536
R53 B1 B1.n0 205.737
R54 B1.n0 B1.t0 169.237
R55 A3.n0 A3.t0 212.154
R56 A3.n0 A3.t1 157.856
R57 A3 A3.n0 155.475
C0 A2 Y 3.82e-20
C1 B1 C1 0.052799f
C2 A1 VPWR 0.018604f
C3 A3 VGND 0.053811f
C4 A2 VGND 0.087884f
C5 A1 Y 0.055826f
C6 B1 VPWR 0.05187f
C7 B1 Y 0.15147f
C8 A1 VGND 0.059871f
C9 C1 VPWR 0.014715f
C10 VPB A3 0.038924f
C11 B1 VGND 0.017702f
C12 C1 Y 0.10989f
C13 VPB A2 0.026048f
C14 C1 VGND 0.01826f
C15 VPWR Y 0.034521f
C16 A3 A2 0.093813f
C17 VPB A1 0.026811f
C18 VPWR VGND 0.070009f
C19 VPB B1 0.032473f
C20 Y VGND 0.147695f
C21 A3 B1 5.21e-19
C22 VPB C1 0.042338f
C23 A2 A1 0.141111f
C24 VPB VPWR 0.084745f
C25 A2 B1 6.97e-19
C26 VPB Y 0.018528f
C27 A1 B1 0.074771f
C28 A3 VPWR 0.060382f
C29 A2 VPWR 0.022119f
C30 VPB VGND 0.012869f
C31 A3 Y 1.52e-20
C32 VGND VNB 0.427884f
C33 Y VNB 0.064284f
C34 VPWR VNB 0.369169f
C35 C1 VNB 0.144508f
C36 B1 VNB 0.094127f
C37 A1 VNB 0.093546f
C38 A2 VNB 0.096704f
C39 A3 VNB 0.147815f
C40 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311oi_2 VNB VPB VGND VPWR C1 Y B1 A1 A2 A3
X0 Y.t4 A1.t0 a_277_47.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_641_297.t2 B1.t0 a_109_297.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t5 A1.t1 a_109_297.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297.t5 B1.t1 a_641_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_109_297.t6 A1.t2 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X5 a_277_47.t2 A1.t3 Y.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297.t3 A2.t0 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t1 A3.t0 a_109_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47.t3 A3.t1 VGND.t4 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47.t1 A2.t1 a_277_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND.t3 C1.t0 Y.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X11 VPWR.t2 A2.t2 a_109_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X12 a_641_297.t3 C1.t1 Y.t2 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_277_47.t0 A2.t3 a_27_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t2 B1.t2 Y.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X15 Y.t0 C1.t2 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_109_297.t0 A3.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y.t1 C1.t3 a_641_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X18 VGND.t5 A3.t3 a_27_47.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 Y.t6 B1.t3 VGND.t1 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 A1.n6 A1.t2 220.845
R1 A1.n0 A1.t1 212.081
R2 A1.n2 A1.t0 164.611
R3 A1.n3 A1.n2 152
R4 A1.n5 A1.n4 152
R5 A1.n7 A1.n6 152
R6 A1.n1 A1.t3 139.78
R7 A1.n6 A1.n5 49.6611
R8 A1.n2 A1.n1 36.5157
R9 A1.n4 A1.n3 13.1884
R10 A1.n1 A1.n0 10.2247
R11 A1.n7 A1 8.92171
R12 A1 A1.n7 8.92171
R13 A1.n4 A1 4.26717
R14 A1.n5 A1.n0 2.92171
R15 A1.n3 A1 0.388379
R16 a_277_47.n1 a_277_47.n0 472.401
R17 a_277_47.n0 a_277_47.t3 24.9236
R18 a_277_47.n0 a_277_47.t2 24.9236
R19 a_277_47.n1 a_277_47.t1 24.9236
R20 a_277_47.t0 a_277_47.n1 24.9236
R21 Y.n0 Y 593.34
R22 Y.n1 Y.n0 585
R23 Y.n4 Y.t3 332.83
R24 Y.n6 Y.t0 326.416
R25 Y.n4 Y.n3 202.695
R26 Y.n5 Y.n2 202.695
R27 Y.n2 Y.t5 71.0774
R28 Y.n5 Y.n4 64.0005
R29 Y.n3 Y.t4 28.6159
R30 Y.n3 Y.t7 26.7697
R31 Y.n0 Y.t2 26.5955
R32 Y.n0 Y.t1 26.5955
R33 Y Y.n1 25.3814
R34 Y.n2 Y.t6 24.9236
R35 Y.n6 Y.n5 6.77697
R36 Y.n1 Y 4.84898
R37 Y Y.n6 1.48887
R38 VNB.t4 VNB.t5 2677.02
R39 VNB.t8 VNB.t7 1908.09
R40 VNB.t6 VNB.t9 1281.55
R41 VNB.t7 VNB.t2 1196.12
R42 VNB.t9 VNB.t8 1196.12
R43 VNB.t5 VNB.t6 1196.12
R44 VNB.t3 VNB.t4 1196.12
R45 VNB.t0 VNB.t3 1196.12
R46 VNB.t1 VNB.t0 1196.12
R47 VNB VNB.t1 911.327
R48 B1.n0 B1.t0 212.081
R49 B1.n2 B1.t1 212.081
R50 B1.n1 B1 152.776
R51 B1.n4 B1.n3 152
R52 B1.n0 B1.t3 139.78
R53 B1.n2 B1.t2 139.78
R54 B1.n3 B1.n1 49.6611
R55 B1.n4 B1 12.4126
R56 B1.n1 B1.n0 10.2247
R57 B1 B1.n4 5.4308
R58 B1.n3 B1.n2 1.46111
R59 a_109_297.n3 a_109_297.n2 385.738
R60 a_109_297.n5 a_109_297.n4 378.2
R61 a_109_297.n3 a_109_297.n1 314.952
R62 a_109_297.n4 a_109_297.n0 314.952
R63 a_109_297.n4 a_109_297.n3 65.5064
R64 a_109_297.n0 a_109_297.t2 28.5655
R65 a_109_297.n2 a_109_297.t4 26.5955
R66 a_109_297.n2 a_109_297.t5 26.5955
R67 a_109_297.n1 a_109_297.t7 26.5955
R68 a_109_297.n1 a_109_297.t6 26.5955
R69 a_109_297.n0 a_109_297.t3 26.5955
R70 a_109_297.n5 a_109_297.t1 26.5955
R71 a_109_297.t0 a_109_297.n5 26.5955
R72 a_641_297.n0 a_641_297.t1 912.711
R73 a_641_297.n0 a_641_297.t3 386.286
R74 a_641_297.n1 a_641_297.n0 295.762
R75 a_641_297.n1 a_641_297.t0 55.1605
R76 a_641_297.t2 a_641_297.n1 47.2805
R77 VPB.t9 VPB.t5 556.386
R78 VPB.t6 VPB.t2 396.574
R79 VPB.t3 VPB.t8 260.437
R80 VPB.t4 VPB.t3 254.518
R81 VPB.t2 VPB.t7 248.599
R82 VPB.t5 VPB.t6 248.599
R83 VPB.t8 VPB.t9 248.599
R84 VPB.t1 VPB.t4 248.599
R85 VPB.t0 VPB.t1 248.599
R86 VPB VPB.t0 189.409
R87 VPWR.n5 VPWR.t5 342.274
R88 VPWR.n8 VPWR.n2 310.502
R89 VPWR.n4 VPWR.n3 309.474
R90 VPWR.n10 VPWR.t0 250.463
R91 VPWR.n3 VPWR.t4 30.5355
R92 VPWR.n2 VPWR.t3 26.5955
R93 VPWR.n2 VPWR.t1 26.5955
R94 VPWR.n3 VPWR.t2 26.5955
R95 VPWR.n10 VPWR.n9 25.977
R96 VPWR.n8 VPWR.n7 25.977
R97 VPWR.n9 VPWR.n8 18.4476
R98 VPWR.n7 VPWR.n4 13.177
R99 VPWR.n7 VPWR.n6 9.3005
R100 VPWR.n8 VPWR.n1 9.3005
R101 VPWR.n9 VPWR.n0 9.3005
R102 VPWR.n11 VPWR.n10 9.3005
R103 VPWR.n5 VPWR.n4 6.73206
R104 VPWR.n6 VPWR.n5 0.777878
R105 VPWR.n6 VPWR.n1 0.120292
R106 VPWR.n1 VPWR.n0 0.120292
R107 VPWR.n11 VPWR.n0 0.120292
R108 VPWR VPWR.n11 0.0213333
R109 A2.n0 A2.t2 213.542
R110 A2.n2 A2.t0 212.081
R111 A2 A2.n1 158.982
R112 A2.n4 A2.n3 152
R113 A2.n2 A2.t3 139.78
R114 A2.n0 A2.t1 139.78
R115 A2.n3 A2.n1 49.6611
R116 A2.n4 A2 11.6369
R117 A2.n3 A2.n2 8.76414
R118 A2 A2.n4 6.20656
R119 A2.n1 A2.n0 2.92171
R120 A3.n1 A3.t0 212.081
R121 A3.n2 A3.t2 212.081
R122 A3.n2 A3.n0 183.404
R123 A3.n4 A3.n3 152
R124 A3.n1 A3.t1 139.78
R125 A3.n2 A3.t3 139.78
R126 A3.n3 A3.n1 43.0884
R127 A3.n3 A3.n2 18.2581
R128 A3.n4 A3.n0 13.1884
R129 A3.n0 A3 4.07323
R130 A3 A3.n4 0.582318
R131 VGND.n6 VGND.n5 205.392
R132 VGND.n4 VGND.n3 199.739
R133 VGND.n17 VGND.n16 199.739
R134 VGND.n9 VGND.n8 34.6358
R135 VGND.n10 VGND.n9 34.6358
R136 VGND.n10 VGND.n1 34.6358
R137 VGND.n14 VGND.n1 34.6358
R138 VGND.n15 VGND.n14 34.6358
R139 VGND.n5 VGND.t0 24.9236
R140 VGND.n5 VGND.t3 24.9236
R141 VGND.n3 VGND.t1 24.9236
R142 VGND.n3 VGND.t2 24.9236
R143 VGND.n16 VGND.t4 24.9236
R144 VGND.n16 VGND.t5 24.9236
R145 VGND.n17 VGND.n15 22.9652
R146 VGND.n8 VGND.n4 10.1652
R147 VGND.n8 VGND.n7 9.3005
R148 VGND.n9 VGND.n2 9.3005
R149 VGND.n11 VGND.n10 9.3005
R150 VGND.n12 VGND.n1 9.3005
R151 VGND.n14 VGND.n13 9.3005
R152 VGND.n15 VGND.n0 9.3005
R153 VGND.n6 VGND.n4 7.26311
R154 VGND.n18 VGND.n17 7.12063
R155 VGND.n7 VGND.n6 0.45585
R156 VGND.n18 VGND.n0 0.148519
R157 VGND.n7 VGND.n2 0.120292
R158 VGND.n11 VGND.n2 0.120292
R159 VGND.n12 VGND.n11 0.120292
R160 VGND.n13 VGND.n12 0.120292
R161 VGND.n13 VGND.n0 0.120292
R162 VGND VGND.n18 0.11354
R163 a_27_47.t1 a_27_47.n1 331.325
R164 a_27_47.n1 a_27_47.t2 330.558
R165 a_27_47.n1 a_27_47.n0 202.695
R166 a_27_47.n0 a_27_47.t0 24.9236
R167 a_27_47.n0 a_27_47.t3 24.9236
R168 C1.n3 C1.t1 212.081
R169 C1.n1 C1.t3 212.081
R170 C1.n4 C1.n3 182.899
R171 C1.n2 C1.n0 152
R172 C1.n3 C1.t2 139.78
R173 C1.n1 C1.t0 139.78
R174 C1.n2 C1.n1 40.1672
R175 C1.n3 C1.n2 21.1793
R176 C1.n5 C1.n0 15.7096
R177 C1 C1.n5 14.1622
R178 C1.n0 C1 9.6005
R179 C1.n4 C1 2.99624
R180 C1.n5 C1.n4 1.3622
C0 VPB B1 0.06279f
C1 Y VGND 0.269518f
C2 VPB C1 0.076966f
C3 A2 A1 0.067933f
C4 VPB VPWR 0.12045f
C5 A1 B1 0.060828f
C6 VPB Y 0.010664f
C7 A3 VPWR 0.067955f
C8 VPB VGND 0.010785f
C9 A3 Y 1.7e-19
C10 A2 VPWR 0.039381f
C11 A3 VGND 0.035471f
C12 B1 C1 0.026565f
C13 A1 VPWR 0.040878f
C14 A2 Y 6.28e-19
C15 A1 Y 0.087629f
C16 A2 VGND 0.022434f
C17 B1 VPWR 0.018892f
C18 B1 Y 0.10862f
C19 A1 VGND 0.024796f
C20 C1 VPWR 0.021191f
C21 VPB A3 0.069696f
C22 C1 Y 0.15678f
C23 B1 VGND 0.028967f
C24 VPB A2 0.05465f
C25 C1 VGND 0.036216f
C26 VPWR Y 0.016217f
C27 A3 A2 0.076912f
C28 VPB A1 0.082171f
C29 VPWR VGND 0.108674f
C30 VGND VNB 0.625352f
C31 Y VNB 0.064962f
C32 VPWR VNB 0.55202f
C33 C1 VNB 0.251162f
C34 B1 VNB 0.18139f
C35 A1 VNB 0.225735f
C36 A2 VNB 0.179119f
C37 A3 VNB 0.237402f
C38 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311oi_4 VNB VPB VPWR VGND C1 A3 A2 A1 B1 Y
X0 a_27_47.t3 A2.t0 a_445_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47.t2 A2.t1 a_445_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t3 C1.t0 Y.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.15925 ps=1.14 w=0.65 l=0.15
X3 a_1139_297.t7 B1.t0 a_109_297.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.49 as=0.135 ps=1.27 w=1 l=0.15
X4 a_109_297.t4 A2.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t0 A3.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_109_297.t8 B1.t1 a_1139_297.t6 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t2 C1.t1 VGND.t2 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t1 C1.t2 VGND.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_1139_297.t5 B1.t2 a_109_297.t7 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_445_47.t4 A1.t0 Y.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297.t11 A3.t1 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR.t5 A1.t1 a_109_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_109_297.t6 A1.t2 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_109_297.t10 B1.t3 a_1139_297.t4 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 a_445_47.t5 A1.t3 Y.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VGND.t8 B1.t4 Y.t12 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t8 A3.t2 a_109_297.t12 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR.t10 A1.t4 a_109_297.t14 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_1139_297.t3 C1.t3 Y.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_27_47.t4 A3.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_27_47.t5 A3.t4 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND.t0 C1.t4 Y.t0 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_109_297.t15 A1.t5 VPWR.t11 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y.t6 C1.t5 a_1139_297.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y.t10 A1.t6 a_445_47.t6 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t3 A2.t3 a_109_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_1139_297.t1 C1.t6 Y.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y.t11 A1.t7 a_445_47.t7 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t13 B1.t5 VGND.t9 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 Y.t14 B1.t6 VGND.t10 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.15925 pd=1.14 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VGND.t6 A3.t5 a_27_47.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_445_47.t1 A2.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 a_109_297.t2 A2.t5 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y.t4 C1.t7 a_1139_297.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.49 w=1 l=0.15
X35 a_445_47.t0 A2.t6 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 VPWR.t1 A2.t7 a_109_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VGND.t11 B1.t7 Y.t15 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 a_109_297.t13 A3.t6 VPWR.t9 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X39 VGND.t7 A3.t7 a_27_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n1 A2.t3 212.081
R1 A2.n9 A2.t5 212.081
R2 A2.n2 A2.t7 212.081
R3 A2.n3 A2.t2 212.081
R4 A2.n11 A2.n10 152
R5 A2.n8 A2.n0 152
R6 A2.n7 A2.n6 152
R7 A2.n5 A2.n4 152
R8 A2.n1 A2.t1 139.78
R9 A2.n9 A2.t6 139.78
R10 A2.n2 A2.t0 139.78
R11 A2.n3 A2.t4 139.78
R12 A2.n8 A2.n7 54.0429
R13 A2.n4 A2.n2 52.5823
R14 A2.n10 A2.n9 48.2005
R15 A2.n11 A2.n0 14.352
R16 A2.n10 A2.n1 13.146
R17 A2.n6 A2 12.8005
R18 A2 A2.n5 9.30959
R19 A2.n4 A2.n3 8.76414
R20 A2.n5 A2 8.53383
R21 A2.n9 A2.n8 5.84292
R22 A2.n6 A2 5.04292
R23 A2 A2.n11 1.93989
R24 A2 A2.n0 1.55202
R25 A2.n7 A2.n2 1.46111
R26 a_445_47.n2 a_445_47.n0 248.248
R27 a_445_47.n4 a_445_47.n3 248.248
R28 a_445_47.n2 a_445_47.n1 185
R29 a_445_47.n5 a_445_47.n4 185
R30 a_445_47.n4 a_445_47.n2 102.4
R31 a_445_47.n3 a_445_47.t3 24.9236
R32 a_445_47.n3 a_445_47.t1 24.9236
R33 a_445_47.n1 a_445_47.t7 24.9236
R34 a_445_47.n1 a_445_47.t5 24.9236
R35 a_445_47.n0 a_445_47.t6 24.9236
R36 a_445_47.n0 a_445_47.t4 24.9236
R37 a_445_47.n5 a_445_47.t2 24.9236
R38 a_445_47.t0 a_445_47.n5 24.9236
R39 a_27_47.n2 a_27_47.t7 329.051
R40 a_27_47.n4 a_27_47.t2 322.094
R41 a_27_47.n2 a_27_47.n1 201.189
R42 a_27_47.n3 a_27_47.n0 201.189
R43 a_27_47.n5 a_27_47.n4 185
R44 a_27_47.n4 a_27_47.n3 63.2476
R45 a_27_47.n3 a_27_47.n2 63.2476
R46 a_27_47.n1 a_27_47.t6 24.9236
R47 a_27_47.n1 a_27_47.t4 24.9236
R48 a_27_47.n0 a_27_47.t1 24.9236
R49 a_27_47.n0 a_27_47.t5 24.9236
R50 a_27_47.n5 a_27_47.t0 24.9236
R51 a_27_47.t3 a_27_47.n5 24.9236
R52 VNB.t2 VNB.t13 2677.02
R53 VNB.t18 VNB.t10 1822.65
R54 VNB.t12 VNB.t11 1196.12
R55 VNB.t9 VNB.t12 1196.12
R56 VNB.t10 VNB.t9 1196.12
R57 VNB.t19 VNB.t18 1196.12
R58 VNB.t17 VNB.t19 1196.12
R59 VNB.t16 VNB.t17 1196.12
R60 VNB.t14 VNB.t16 1196.12
R61 VNB.t8 VNB.t14 1196.12
R62 VNB.t15 VNB.t8 1196.12
R63 VNB.t13 VNB.t15 1196.12
R64 VNB.t0 VNB.t2 1196.12
R65 VNB.t3 VNB.t0 1196.12
R66 VNB.t1 VNB.t3 1196.12
R67 VNB.t5 VNB.t1 1196.12
R68 VNB.t6 VNB.t5 1196.12
R69 VNB.t4 VNB.t6 1196.12
R70 VNB.t7 VNB.t4 1196.12
R71 VNB VNB.t7 911.327
R72 C1.n0 C1.t3 212.081
R73 C1.n7 C1.t5 212.081
R74 C1.n1 C1.t6 212.081
R75 C1.n2 C1.t7 212.081
R76 C1 C1.n0 187.774
R77 C1.n9 C1.n8 152
R78 C1.n6 C1.n5 152
R79 C1.n4 C1.n3 152
R80 C1.n0 C1.t2 139.78
R81 C1.n7 C1.t4 139.78
R82 C1.n1 C1.t1 139.78
R83 C1.n2 C1.t0 139.78
R84 C1.n3 C1.n2 54.7732
R85 C1.n6 C1.n1 47.4702
R86 C1.n8 C1.n7 40.1672
R87 C1.n8 C1.n0 21.1793
R88 C1.n7 C1.n6 13.8763
R89 C1.n4 C1 13.3823
R90 C1 C1.n9 11.4429
R91 C1.n5 C1 9.89141
R92 C1.n5 C1 7.95202
R93 C1.n3 C1.n1 6.57323
R94 C1.n9 C1 6.4005
R95 C1 C1.n4 4.46111
R96 Y.n2 Y.n0 334.445
R97 Y.n11 Y.t1 329.051
R98 Y.n6 Y.t9 322.094
R99 Y.n2 Y.n1 296.046
R100 Y.n13 Y.n12 204.589
R101 Y.n11 Y.n10 201.189
R102 Y.n9 Y.n4 201.189
R103 Y.n8 Y.n7 185
R104 Y.n6 Y.n5 185
R105 Y.n12 Y.t3 65.539
R106 Y.n9 Y.n8 63.2476
R107 Y.n8 Y.n6 63.2476
R108 Y.n13 Y.n11 62.1181
R109 Y.n13 Y.n9 56.8476
R110 Y.n0 Y.t7 26.5955
R111 Y.n0 Y.t6 26.5955
R112 Y.n1 Y.t5 26.5955
R113 Y.n1 Y.t4 26.5955
R114 Y.n10 Y.t0 24.9236
R115 Y.n10 Y.t2 24.9236
R116 Y.n5 Y.t8 24.9236
R117 Y.n5 Y.t11 24.9236
R118 Y.n7 Y.t12 24.9236
R119 Y.n7 Y.t10 24.9236
R120 Y.n4 Y.t15 24.9236
R121 Y.n4 Y.t13 24.9236
R122 Y.n12 Y.t14 24.9236
R123 Y.n3 Y.n2 18.0711
R124 Y Y.n3 7.4005
R125 Y.n3 Y 6.2005
R126 Y Y.n13 1.8005
R127 VGND.n13 VGND.n10 205.155
R128 VGND.n12 VGND.n11 199.739
R129 VGND.n16 VGND.n9 199.739
R130 VGND.n19 VGND.n18 199.739
R131 VGND.n35 VGND.n2 199.739
R132 VGND.n38 VGND.n37 199.739
R133 VGND.n23 VGND.n6 34.6358
R134 VGND.n24 VGND.n23 34.6358
R135 VGND.n25 VGND.n24 34.6358
R136 VGND.n25 VGND.n4 34.6358
R137 VGND.n29 VGND.n4 34.6358
R138 VGND.n30 VGND.n29 34.6358
R139 VGND.n31 VGND.n30 34.6358
R140 VGND.n31 VGND.n1 34.6358
R141 VGND.n12 VGND.n8 28.9887
R142 VGND.n35 VGND.n1 28.9887
R143 VGND.n16 VGND.n8 25.977
R144 VGND.n10 VGND.t1 24.9236
R145 VGND.n10 VGND.t0 24.9236
R146 VGND.n11 VGND.t2 24.9236
R147 VGND.n11 VGND.t3 24.9236
R148 VGND.n9 VGND.t10 24.9236
R149 VGND.n9 VGND.t11 24.9236
R150 VGND.n18 VGND.t9 24.9236
R151 VGND.n18 VGND.t8 24.9236
R152 VGND.n2 VGND.t5 24.9236
R153 VGND.n2 VGND.t6 24.9236
R154 VGND.n37 VGND.t4 24.9236
R155 VGND.n37 VGND.t7 24.9236
R156 VGND.n19 VGND.n6 24.4711
R157 VGND.n38 VGND.n36 22.9652
R158 VGND.n19 VGND.n17 19.9534
R159 VGND.n17 VGND.n16 18.4476
R160 VGND.n36 VGND.n35 15.4358
R161 VGND.n14 VGND.n8 9.3005
R162 VGND.n16 VGND.n15 9.3005
R163 VGND.n17 VGND.n7 9.3005
R164 VGND.n20 VGND.n19 9.3005
R165 VGND.n21 VGND.n6 9.3005
R166 VGND.n23 VGND.n22 9.3005
R167 VGND.n24 VGND.n5 9.3005
R168 VGND.n26 VGND.n25 9.3005
R169 VGND.n27 VGND.n4 9.3005
R170 VGND.n29 VGND.n28 9.3005
R171 VGND.n30 VGND.n3 9.3005
R172 VGND.n32 VGND.n31 9.3005
R173 VGND.n33 VGND.n1 9.3005
R174 VGND.n35 VGND.n34 9.3005
R175 VGND.n36 VGND.n0 9.3005
R176 VGND.n39 VGND.n38 7.12063
R177 VGND.n13 VGND.n12 6.06315
R178 VGND.n14 VGND.n13 0.653139
R179 VGND.n39 VGND.n0 0.148519
R180 VGND.n15 VGND.n14 0.120292
R181 VGND.n15 VGND.n7 0.120292
R182 VGND.n20 VGND.n7 0.120292
R183 VGND.n21 VGND.n20 0.120292
R184 VGND.n22 VGND.n21 0.120292
R185 VGND.n22 VGND.n5 0.120292
R186 VGND.n26 VGND.n5 0.120292
R187 VGND.n27 VGND.n26 0.120292
R188 VGND.n28 VGND.n27 0.120292
R189 VGND.n28 VGND.n3 0.120292
R190 VGND.n32 VGND.n3 0.120292
R191 VGND.n33 VGND.n32 0.120292
R192 VGND.n34 VGND.n33 0.120292
R193 VGND.n34 VGND.n0 0.120292
R194 VGND VGND.n39 0.11354
R195 B1.n6 B1.t3 212.081
R196 B1.n1 B1.t0 212.081
R197 B1.n2 B1.t1 212.081
R198 B1.n0 B1.t2 212.081
R199 B1 B1.n3 155.226
R200 B1.n5 B1.n4 152
R201 B1.n7 B1.n6 152
R202 B1.n6 B1.t4 139.78
R203 B1.n1 B1.t6 139.78
R204 B1.n2 B1.t7 139.78
R205 B1.n0 B1.t5 139.78
R206 B1.n2 B1.n1 61.346
R207 B1.n6 B1.n5 54.0429
R208 B1.n3 B1.n0 46.7399
R209 B1.n3 B1.n2 14.6066
R210 B1.n5 B1.n0 7.30353
R211 B1 B1.n7 6.85404
R212 B1.n4 B1 5.03987
R213 B1.n4 B1 4.23357
R214 B1.n7 B1 2.4194
R215 a_109_297.n5 a_109_297.n3 648.247
R216 a_109_297.n5 a_109_297.n4 585
R217 a_109_297.n12 a_109_297.n11 384.224
R218 a_109_297.n8 a_109_297.n2 320.976
R219 a_109_297.n9 a_109_297.n1 320.976
R220 a_109_297.n10 a_109_297.n0 320.976
R221 a_109_297.n13 a_109_297.n12 320.976
R222 a_109_297.n7 a_109_297.n6 296.493
R223 a_109_297.n7 a_109_297.n5 102.4
R224 a_109_297.n8 a_109_297.n7 82.0711
R225 a_109_297.n9 a_109_297.n8 63.2476
R226 a_109_297.n10 a_109_297.n9 63.2476
R227 a_109_297.n12 a_109_297.n10 63.2476
R228 a_109_297.n6 a_109_297.t5 26.5955
R229 a_109_297.n6 a_109_297.t6 26.5955
R230 a_109_297.n4 a_109_297.t7 26.5955
R231 a_109_297.n4 a_109_297.t10 26.5955
R232 a_109_297.n3 a_109_297.t9 26.5955
R233 a_109_297.n3 a_109_297.t8 26.5955
R234 a_109_297.n2 a_109_297.t14 26.5955
R235 a_109_297.n2 a_109_297.t15 26.5955
R236 a_109_297.n1 a_109_297.t3 26.5955
R237 a_109_297.n1 a_109_297.t2 26.5955
R238 a_109_297.n0 a_109_297.t1 26.5955
R239 a_109_297.n0 a_109_297.t4 26.5955
R240 a_109_297.n11 a_109_297.t12 26.5955
R241 a_109_297.n11 a_109_297.t13 26.5955
R242 a_109_297.t0 a_109_297.n13 26.5955
R243 a_109_297.n13 a_109_297.t11 26.5955
R244 a_1139_297.n1 a_1139_297.t4 917.229
R245 a_1139_297.n5 a_1139_297.n4 585
R246 a_1139_297.n3 a_1139_297.n2 585
R247 a_1139_297.n1 a_1139_297.n0 585
R248 a_1139_297.t3 a_1139_297.n5 380.231
R249 a_1139_297.n5 a_1139_297.n3 79.8123
R250 a_1139_297.n2 a_1139_297.t0 69.9355
R251 a_1139_297.n3 a_1139_297.n1 63.2476
R252 a_1139_297.n0 a_1139_297.t6 26.5955
R253 a_1139_297.n0 a_1139_297.t5 26.5955
R254 a_1139_297.n2 a_1139_297.t7 26.5955
R255 a_1139_297.n4 a_1139_297.t2 26.5955
R256 a_1139_297.n4 a_1139_297.t1 26.5955
R257 VPB.t5 VPB.t11 556.386
R258 VPB.t14 VPB.t7 378.817
R259 VPB.t9 VPB.t10 248.599
R260 VPB.t8 VPB.t9 248.599
R261 VPB.t7 VPB.t8 248.599
R262 VPB.t13 VPB.t14 248.599
R263 VPB.t12 VPB.t13 248.599
R264 VPB.t11 VPB.t12 248.599
R265 VPB.t6 VPB.t5 248.599
R266 VPB.t18 VPB.t6 248.599
R267 VPB.t19 VPB.t18 248.599
R268 VPB.t3 VPB.t19 248.599
R269 VPB.t2 VPB.t3 248.599
R270 VPB.t1 VPB.t2 248.599
R271 VPB.t4 VPB.t1 248.599
R272 VPB.t0 VPB.t4 248.599
R273 VPB.t15 VPB.t0 248.599
R274 VPB.t16 VPB.t15 248.599
R275 VPB.t17 VPB.t16 248.599
R276 VPB VPB.t17 189.409
R277 VPWR.n9 VPWR.t5 874.081
R278 VPWR.n23 VPWR.n2 310.502
R279 VPWR.n4 VPWR.n3 310.502
R280 VPWR.n17 VPWR.n6 310.502
R281 VPWR.n8 VPWR.n7 310.502
R282 VPWR.n11 VPWR.n10 310.502
R283 VPWR.n25 VPWR.t9 243.512
R284 VPWR.n16 VPWR.n15 34.6358
R285 VPWR.n18 VPWR.n4 32.0005
R286 VPWR.n12 VPWR.n11 28.9887
R287 VPWR.n2 VPWR.t7 26.5955
R288 VPWR.n2 VPWR.t8 26.5955
R289 VPWR.n3 VPWR.t4 26.5955
R290 VPWR.n3 VPWR.t0 26.5955
R291 VPWR.n6 VPWR.t2 26.5955
R292 VPWR.n6 VPWR.t1 26.5955
R293 VPWR.n7 VPWR.t11 26.5955
R294 VPWR.n7 VPWR.t3 26.5955
R295 VPWR.n10 VPWR.t6 26.5955
R296 VPWR.n10 VPWR.t10 26.5955
R297 VPWR.n23 VPWR.n22 25.977
R298 VPWR.n25 VPWR.n24 19.9534
R299 VPWR.n24 VPWR.n23 18.4476
R300 VPWR.n22 VPWR.n4 12.424
R301 VPWR.n12 VPWR.n8 9.41227
R302 VPWR.n13 VPWR.n12 9.3005
R303 VPWR.n15 VPWR.n14 9.3005
R304 VPWR.n16 VPWR.n5 9.3005
R305 VPWR.n19 VPWR.n18 9.3005
R306 VPWR.n20 VPWR.n4 9.3005
R307 VPWR.n22 VPWR.n21 9.3005
R308 VPWR.n23 VPWR.n1 9.3005
R309 VPWR.n24 VPWR.n0 9.3005
R310 VPWR.n26 VPWR.n25 9.3005
R311 VPWR.n18 VPWR.n17 6.4005
R312 VPWR.n11 VPWR.n9 6.06787
R313 VPWR.n17 VPWR.n16 3.38874
R314 VPWR.n13 VPWR.n9 0.647986
R315 VPWR.n15 VPWR.n8 0.376971
R316 VPWR.n14 VPWR.n13 0.120292
R317 VPWR.n14 VPWR.n5 0.120292
R318 VPWR.n19 VPWR.n5 0.120292
R319 VPWR.n20 VPWR.n19 0.120292
R320 VPWR.n21 VPWR.n20 0.120292
R321 VPWR.n21 VPWR.n1 0.120292
R322 VPWR.n1 VPWR.n0 0.120292
R323 VPWR.n26 VPWR.n0 0.120292
R324 VPWR VPWR.n26 0.0213333
R325 A3.n1 A3.t0 212.081
R326 A3.n4 A3.t1 212.081
R327 A3.n0 A3.t2 212.081
R328 A3.n9 A3.t6 212.081
R329 A3.n10 A3.n9 179.022
R330 A3.n3 A3.n2 152
R331 A3.n6 A3.n5 152
R332 A3.n8 A3.n7 152
R333 A3.n1 A3.t4 139.78
R334 A3.n4 A3.t5 139.78
R335 A3.n0 A3.t3 139.78
R336 A3.n9 A3.t7 139.78
R337 A3.n3 A3.n1 48.9308
R338 A3.n5 A3.n4 41.6278
R339 A3.n8 A3.n0 34.3247
R340 A3.n9 A3.n8 27.0217
R341 A3.n5 A3.n0 19.7187
R342 A3.n7 A3.n6 14.352
R343 A3.n2 A3 12.6066
R344 A3.n10 A3 12.6066
R345 A3.n4 A3.n3 12.4157
R346 A3.n2 A3 5.23686
R347 A3 A3.n10 5.23686
R348 A3.n6 A3 1.74595
R349 A3.n7 A3 1.74595
R350 A1.n10 A1.t5 213.917
R351 A1.n3 A1.t1 205.654
R352 A1.n7 A1.t2 205.654
R353 A1.n11 A1.t4 205.654
R354 A1.n2 A1.t6 200.631
R355 A1.n5 A1.n4 152
R356 A1.n8 A1.n0 152
R357 A1.n13 A1.n12 152
R358 A1.n10 A1.n1 152
R359 A1.n9 A1.t3 139.78
R360 A1.n6 A1.t7 139.78
R361 A1.n2 A1.t0 137.678
R362 A1.n11 A1.n10 49.5776
R363 A1.n9 A1.n8 38.5605
R364 A1.n6 A1.n5 31.6748
R365 A1.n13 A1.n1 14.352
R366 A1.n7 A1.n6 13.7719
R367 A1.n3 A1.n2 13.1979
R368 A1 A1.n0 13.1884
R369 A1.n5 A1.n3 12.3948
R370 A1.n12 A1.n9 12.3948
R371 A1.n4 A1 9.69747
R372 A1.n4 A1 8.14595
R373 A1.n8 A1.n7 5.50907
R374 A1 A1.n0 4.65505
R375 A1.n1 A1 2.32777
R376 A1.n12 A1.n11 1.37764
R377 A1 A1.n13 1.16414
C0 VPB VGND 0.013665f
C1 A3 Y 5.06e-20
C2 A2 VPWR 0.068836f
C3 A3 VGND 0.070183f
C4 B1 C1 0.028082f
C5 A1 VPWR 0.080349f
C6 A2 Y 1.92e-19
C7 A1 Y 0.146498f
C8 A2 VGND 0.035952f
C9 B1 VPWR 0.042932f
C10 C1 VPWR 0.035581f
C11 B1 Y 0.192881f
C12 A1 VGND 0.042978f
C13 VPB A3 0.133909f
C14 B1 VGND 0.070519f
C15 C1 Y 0.346098f
C16 VPB A2 0.116393f
C17 C1 VGND 0.070169f
C18 VPWR Y 0.031502f
C19 VPB A1 0.145173f
C20 A3 A2 0.078238f
C21 VPWR VGND 0.18801f
C22 VPB B1 0.13488f
C23 Y VGND 0.47696f
C24 A3 B1 8.72e-20
C25 A2 A1 0.064307f
C26 VPB C1 0.136883f
C27 A2 B1 2.23e-19
C28 VPB VPWR 0.183013f
C29 A3 VPWR 0.112944f
C30 VPB Y 0.013729f
C31 A1 B1 0.077079f
C32 VGND VNB 1.0288f
C33 Y VNB 0.07536f
C34 VPWR VNB 0.888288f
C35 C1 VNB 0.426141f
C36 B1 VNB 0.365609f
C37 A1 VNB 0.407971f
C38 A2 VNB 0.359141f
C39 A3 VNB 0.420909f
C40 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111o_1 VPB VGND VPWR VNB B1 X D1 A1 A2 C1
X0 VGND.t2 A2.t0 a_660_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1 VGND.t4 C1.t0 a_85_193.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_414_297.t0 C1.t1 a_334_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND.t1 a_85_193.t5 X.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X4 a_334_297.t1 D1.t0 a_85_193.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297.t2 B1.t0 a_414_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297.t1 A2.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47.t0 A1.t0 a_85_193.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8 a_85_193.t3 D1.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9 VPWR.t0 A1.t1 a_516_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193.t2 B1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR.t1 a_85_193.t6 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
R0 A2.n0 A2.t1 235.471
R1 A2.n0 A2.t0 157.785
R2 A2 A2.n0 157.555
R3 a_660_47.t0 a_660_47.t1 47.0774
R4 VGND.n4 VGND.t2 243.331
R5 VGND.n3 VGND.n2 199.841
R6 VGND.n10 VGND.n9 185
R7 VGND.n8 VGND.n0 185
R8 VGND.n9 VGND.n8 63.6928
R9 VGND.n9 VGND.t3 58.1543
R10 VGND.n7 VGND.n6 34.6358
R11 VGND.n8 VGND.t1 34.1543
R12 VGND.n2 VGND.t0 33.2313
R13 VGND.n2 VGND.t4 33.2313
R14 VGND.n11 VGND.n7 26.2788
R15 VGND.n4 VGND.n3 15.0566
R16 VGND.n13 VGND.n0 10.1026
R17 VGND.n12 VGND.n11 9.3005
R18 VGND.n7 VGND.n1 9.3005
R19 VGND.n6 VGND.n5 9.3005
R20 VGND.n10 VGND.n0 7.95726
R21 VGND.n6 VGND.n3 1.12991
R22 VGND.n5 VGND.n4 0.220568
R23 VGND.n13 VGND.n12 0.14286
R24 VGND VGND.n13 0.120574
R25 VGND.n5 VGND.n1 0.120292
R26 VGND.n12 VGND.n1 0.120292
R27 VGND.n11 VGND.n10 0.115815
R28 VNB.t4 VNB.t2 2833.66
R29 VNB.t1 VNB.t0 2050.49
R30 VNB.t5 VNB.t1 1452.43
R31 VNB VNB.t4 1281.55
R32 VNB.t0 VNB.t3 1153.4
R33 VNB.t2 VNB 1124.92
R34 VNB VNB.t5 28.4795
R35 C1.n0 C1.t1 229.754
R36 C1.n0 C1.t0 166.291
R37 C1.n1 C1.n0 152
R38 C1 C1.n1 11.055
R39 C1.n1 C1 2.13383
R40 a_85_193.n3 a_85_193.t5 1784.9
R41 a_85_193.t4 a_85_193.n4 430.851
R42 a_85_193.n2 a_85_193.n0 251.756
R43 a_85_193.n3 a_85_193.t6 223.477
R44 a_85_193.n4 a_85_193.n3 152
R45 a_85_193.n2 a_85_193.n1 95.8789
R46 a_85_193.n0 a_85_193.t0 79.3851
R47 a_85_193.n4 a_85_193.n2 73.7335
R48 a_85_193.n1 a_85_193.t1 31.3851
R49 a_85_193.n1 a_85_193.t3 25.8467
R50 a_85_193.n0 a_85_193.t2 25.8467
R51 a_334_297.t0 a_334_297.t1 49.2505
R52 a_414_297.t0 a_414_297.t1 70.9205
R53 VPB.t2 VPB.t5 648.131
R54 VPB.t4 VPB.t1 420.25
R55 VPB.t0 VPB.t4 301.87
R56 VPB.t1 VPB.t3 248.599
R57 VPB.t5 VPB.t0 236.761
R58 VPB VPB.t2 210.125
R59 X.n1 X 593.534
R60 X.n1 X.n0 585
R61 X.n2 X.n1 585
R62 X X.n4 185.97
R63 X.n4 X.n3 185
R64 X.n4 X.t0 30.462
R65 X.n1 X.t1 28.5655
R66 X X.n3 12.2187
R67 X.n2 X 8.67073
R68 X.n0 X 8.53383
R69 X.n0 X 8.53383
R70 X X.n2 6.4005
R71 X.n3 X 0.970197
R72 D1.n0 D1.t0 234.804
R73 D1.n0 D1.t1 162.504
R74 D1.n1 D1.n0 152
R75 D1 D1.n1 13.5483
R76 D1.n1 D1 1.63771
R77 B1.n0 B1.t0 235.304
R78 B1.n0 B1.t1 157.745
R79 B1.n1 B1.n0 152
R80 B1.n1 B1 13.0291
R81 B1 B1.n1 2.51479
R82 a_516_297.n0 a_516_297.t1 688.063
R83 a_516_297.n0 a_516_297.t2 83.7255
R84 a_516_297.t0 a_516_297.n0 26.5955
R85 VPWR.n1 VPWR.t1 344.568
R86 VPWR.n1 VPWR.n0 326.531
R87 VPWR.n0 VPWR.t2 26.5955
R88 VPWR.n0 VPWR.t0 26.5955
R89 VPWR VPWR.n1 0.154701
R90 A1.n0 A1.t1 1053.26
R91 A1.n0 A1.t0 157.785
R92 A1.n1 A1.n0 152.388
R93 A1.n1 A1 15.9821
R94 A1 A1.n1 8.92171
C0 B1 VPWR 0.043795f
C1 C1 VGND 0.016422f
C2 A1 VPWR 0.02157f
C3 B1 VGND 0.014558f
C4 VPB D1 0.038109f
C5 A2 VPWR 0.021508f
C6 A1 VGND 0.116703f
C7 VPB C1 0.030173f
C8 A2 VGND 0.046422f
C9 X VPWR 0.094258f
C10 D1 C1 0.169347f
C11 VPB B1 0.036936f
C12 X VGND 0.068497f
C13 D1 B1 3.12e-19
C14 VPB A1 0.033363f
C15 VPWR VGND 0.087252f
C16 VPB A2 0.033731f
C17 D1 A1 1.88e-19
C18 C1 B1 0.164685f
C19 VPB X 0.010929f
C20 C1 A1 3.55e-19
C21 B1 A1 0.068882f
C22 D1 X 2.82e-19
C23 VPB VPWR 0.098773f
C24 VPB VGND 0.0102f
C25 B1 A2 3.76e-19
C26 D1 VPWR 0.036977f
C27 D1 VGND 0.015289f
C28 A1 A2 0.083244f
C29 C1 VPWR 0.04987f
C30 VGND VNB 0.505453f
C31 VPWR VNB 0.405283f
C32 X VNB 0.088362f
C33 A2 VNB 0.136216f
C34 A1 VNB 0.114026f
C35 B1 VNB 0.101766f
C36 C1 VNB 0.09306f
C37 D1 VNB 0.10506f
C38 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111o_2 VNB VPB VGND VPWR A2 A1 B1 C1 X D1
X0 VPWR.t3 a_86_235.t5 X.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND.t3 C1.t0 a_86_235.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X.t0 a_86_235.t6 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 a_86_235.t1 D1.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.290875 ps=1.545 w=0.65 l=0.15
X4 X.t3 a_86_235.t7 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_715_47.t0 A1.t0 a_86_235.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.108875 ps=0.985 w=0.65 l=0.15
X6 VGND.t1 A2.t0 a_715_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_499_297.t1 C1.t1 a_427_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND.t4 a_86_235.t8 X.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.290875 pd=1.545 as=0.091 ps=0.93 w=0.65 l=0.15
X9 a_86_235.t0 B1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.121875 ps=1.025 w=0.65 l=0.15
X10 a_607_297.t2 B1.t1 a_499_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X11 a_427_297.t0 D1.t1 a_86_235.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.41 ps=2.82 w=1 l=0.15
X12 VPWR.t0 A1.t1 a_607_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X13 a_607_297.t0 A2.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
R0 a_86_235.t2 a_86_235.n6 393.995
R1 a_86_235.n2 a_86_235.n0 250.077
R2 a_86_235.n3 a_86_235.t6 227.546
R3 a_86_235.n4 a_86_235.t5 212.081
R4 a_86_235.n6 a_86_235.n5 204.244
R5 a_86_235.n2 a_86_235.n1 199.934
R6 a_86_235.n3 a_86_235.t7 139.78
R7 a_86_235.n5 a_86_235.t8 139.78
R8 a_86_235.n6 a_86_235.n2 58.6224
R9 a_86_235.n4 a_86_235.n3 51.1217
R10 a_86_235.n0 a_86_235.t3 36.0005
R11 a_86_235.n0 a_86_235.t0 25.8467
R12 a_86_235.n1 a_86_235.t4 25.8467
R13 a_86_235.n1 a_86_235.t1 25.8467
R14 a_86_235.n5 a_86_235.n4 11.6853
R15 X.n3 X.n2 585
R16 X.n4 X.n3 585
R17 X.n0 X 185.221
R18 X.n1 X.n0 185
R19 X.n3 X.t1 27.5805
R20 X.n3 X.t0 27.5805
R21 X.n0 X.t2 25.8467
R22 X.n0 X.t3 25.8467
R23 X.n1 X 14.7867
R24 X.n4 X 11.6971
R25 X.n2 X 11.6971
R26 X X.n4 3.31084
R27 X.n2 X 3.31084
R28 X X.n1 0.22119
R29 VPWR.n2 VPWR.n1 605.736
R30 VPWR.n5 VPWR.t2 405.423
R31 VPWR.n3 VPWR.t3 251.448
R32 VPWR.n1 VPWR.t1 41.3705
R33 VPWR.n1 VPWR.t0 35.4605
R34 VPWR.n4 VPWR.n3 28.2358
R35 VPWR.n5 VPWR.n4 19.2005
R36 VPWR.n4 VPWR.n0 9.3005
R37 VPWR.n6 VPWR.n5 9.3005
R38 VPWR.n3 VPWR.n2 7.06253
R39 VPWR.n2 VPWR.n0 0.156205
R40 VPWR.n6 VPWR.n0 0.120292
R41 VPWR VPWR.n6 0.0226354
R42 VPB.t6 VPB.t4 665.889
R43 VPB.t1 VPB.t2 319.627
R44 VPB.t0 VPB.t1 319.627
R45 VPB.t3 VPB.t0 319.627
R46 VPB.t5 VPB.t6 254.518
R47 VPB.t4 VPB.t3 213.084
R48 VPB VPB.t5 213.084
R49 C1.n0 C1.t1 236.18
R50 C1.n0 C1.t0 163.881
R51 C1.n1 C1.n0 152
R52 C1 C1.n1 11.7682
R53 C1.n1 C1 2.27147
R54 VGND.n4 VGND.n3 198.964
R55 VGND.n11 VGND.n10 185
R56 VGND.n5 VGND.t1 156.196
R57 VGND.n17 VGND.t5 138.945
R58 VGND.n10 VGND.n9 113.538
R59 VGND.n9 VGND.n1 95.3258
R60 VGND.n3 VGND.t3 35.0774
R61 VGND.n8 VGND.n7 34.6358
R62 VGND.n3 VGND.t0 34.1543
R63 VGND.n16 VGND.n15 30.2886
R64 VGND.n10 VGND.t2 25.8467
R65 VGND.n9 VGND.t4 25.8467
R66 VGND.n17 VGND.n16 19.2005
R67 VGND.n5 VGND.n4 12.7961
R68 VGND.n12 VGND.n1 9.58623
R69 VGND.n18 VGND.n17 9.3005
R70 VGND.n7 VGND.n6 9.3005
R71 VGND.n8 VGND.n2 9.3005
R72 VGND.n13 VGND.n12 9.3005
R73 VGND.n15 VGND.n14 9.3005
R74 VGND.n16 VGND.n0 9.3005
R75 VGND.n11 VGND.n8 8.50305
R76 VGND.n12 VGND.n11 5.67597
R77 VGND.n7 VGND.n4 4.51815
R78 VGND.n15 VGND.n1 1.52334
R79 VGND.n6 VGND.n5 0.222113
R80 VGND.n6 VGND.n2 0.120292
R81 VGND.n13 VGND.n2 0.120292
R82 VGND.n14 VGND.n13 0.120292
R83 VGND.n14 VGND.n0 0.120292
R84 VGND.n18 VGND.n0 0.120292
R85 VGND VGND.n18 0.0226354
R86 VNB.t5 VNB.t2 2976.05
R87 VNB.t3 VNB.t1 1537.86
R88 VNB.t4 VNB.t0 1495.15
R89 VNB.t0 VNB.t3 1381.23
R90 VNB VNB.t6 1253.07
R91 VNB.t2 VNB.t4 1224.6
R92 VNB.t6 VNB.t5 1224.6
R93 D1.n0 D1.t1 236.18
R94 D1.n0 D1.t0 163.881
R95 D1.n1 D1.n0 152
R96 D1 D1.n1 10.9154
R97 D1.n1 D1 1.9032
R98 A1.n0 A1.t1 236.18
R99 A1.n0 A1.t0 161.251
R100 A1.n1 A1.n0 152
R101 A1 A1.n1 8.89806
R102 A1.n1 A1 1.71757
R103 a_715_47.t0 a_715_47.t1 72.0005
R104 A2.n0 A2.t1 236.18
R105 A2.n0 A2.t0 163.881
R106 A2.n1 A2.n0 152
R107 A2.n1 A2 6.4005
R108 A2 A2.n1 1.23559
R109 a_427_297.t0 a_427_297.t1 41.3705
R110 a_499_297.t0 a_499_297.t1 76.8305
R111 B1.n0 B1.t1 236.18
R112 B1.n0 B1.t0 163.881
R113 B1.n1 B1.n0 152
R114 B1.n1 B1 12.5798
R115 B1 B1.n1 2.42809
R116 a_607_297.t0 a_607_297.n0 670.332
R117 a_607_297.n0 a_607_297.t2 39.4005
R118 a_607_297.n0 a_607_297.t1 37.4305
C0 VPB C1 0.031781f
C1 VPWR X 0.176259f
C2 A2 VGND 0.056011f
C3 VPB B1 0.033235f
C4 D1 C1 0.180832f
C5 VPWR VGND 0.109652f
C6 VPB A1 0.034344f
C7 X VGND 0.147354f
C8 VPB A2 0.041352f
C9 C1 B1 0.115714f
C10 D1 A1 2.42e-19
C11 VPB VPWR 0.111903f
C12 C1 A1 9.75e-19
C13 D1 VPWR 0.0384f
C14 C1 A2 2.32e-19
C15 B1 A1 0.112643f
C16 VPB X 0.006459f
C17 VPB VGND 0.009079f
C18 C1 VPWR 0.04356f
C19 D1 VGND 0.01681f
C20 B1 VPWR 0.01524f
C21 A1 A2 0.121755f
C22 C1 VGND 0.01616f
C23 A1 VPWR 0.022645f
C24 B1 VGND 0.013674f
C25 A2 VPWR 0.019029f
C26 VPB D1 0.03576f
C27 A1 VGND 0.115481f
C28 VGND VNB 0.584407f
C29 X VNB 0.027649f
C30 VPWR VNB 0.476066f
C31 A2 VNB 0.153595f
C32 A1 VNB 0.108314f
C33 B1 VNB 0.095357f
C34 C1 VNB 0.097961f
C35 D1 VNB 0.102285f
C36 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111o_4 VNB VPB VGND VPWR D1 C1 B1 A1 A2 X
X0 a_30_297.t2 C1.t0 a_285_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND.t2 C1.t1 a_44_47.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.091 ps=0.93 w=0.65 l=0.15
X2 a_44_47.t1 B1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.2665 ps=1.47 w=0.65 l=0.15
X3 VGND.t9 a_44_47.t10 X.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR.t7 A1.t0 a_477_297.t5 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2575 ps=1.515 w=1 l=0.15
X5 VPWR.t5 a_44_47.t11 X.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 X.t2 a_44_47.t12 VGND.t8 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND.t11 B1.t1 a_44_47.t9 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.2665 pd=1.47 as=0.108875 ps=0.985 w=0.65 l=0.15
X8 X.t1 a_44_47.t13 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 a_477_297.t4 A1.t1 VPWR.t6 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_297.t2 B1.t2 a_477_297.t2 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND.t3 D1.t0 a_44_47.t5 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X12 a_770_47.t1 A2.t0 VGND.t10 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.182 ps=1.86 w=0.65 l=0.15
X13 X.t6 a_44_47.t14 VPWR.t4 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 a_30_297.t0 D1.t1 a_44_47.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VGND.t4 A2.t1 a_770_47.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_44_47.t6 D1.t2 a_30_297.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X17 a_477_297.t1 B1.t3 a_285_297.t3 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2575 pd=1.515 as=0.14 ps=1.28 w=1 l=0.15
X18 a_770_47.t3 A1.t2 a_44_47.t8 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.092625 ps=0.935 w=0.65 l=0.15
X19 a_477_297.t3 A2.t2 VPWR.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR.t3 a_44_47.t15 X.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 a_285_297.t0 C1.t2 a_30_297.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 a_44_47.t7 D1.t3 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_44_47.t4 A1.t3 a_770_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VGND.t6 a_44_47.t16 X.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X25 VPWR.t0 A2.t3 a_477_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 X.t4 a_44_47.t17 VPWR.t2 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 a_44_47.t2 C1.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.102375 ps=0.965 w=0.65 l=0.15
R0 C1.n0 C1.t2 224.069
R1 C1.n3 C1.t0 213.688
R2 C1.n5 C1.n4 152
R3 C1.n2 C1.n1 152
R4 C1.n4 C1.t3 144.971
R5 C1.n0 C1.t1 139.78
R6 C1.n3 C1.n2 40.0436
R7 C1.n1 C1 18.3747
R8 C1.n5 C1 13.4199
R9 C1.n2 C1.n0 13.3482
R10 C1.n4 C1.n3 10.382
R11 C1 C1.n5 5.57469
R12 C1.n1 C1 0.619855
R13 a_285_297.n1 a_285_297.n0 685.479
R14 a_285_297.n0 a_285_297.t3 27.5805
R15 a_285_297.n0 a_285_297.t2 27.5805
R16 a_285_297.n1 a_285_297.t1 27.5805
R17 a_285_297.t0 a_285_297.n1 27.5805
R18 a_30_297.n1 a_30_297.t3 378.591
R19 a_30_297.t2 a_30_297.n1 377.608
R20 a_30_297.n1 a_30_297.n0 212.668
R21 a_30_297.n0 a_30_297.t1 27.5805
R22 a_30_297.n0 a_30_297.t0 27.5805
R23 VPB.t1 VPB.t7 556.386
R24 VPB.t5 VPB.t12 556.386
R25 VPB.t13 VPB.t0 393.615
R26 VPB.t9 VPB.t10 254.518
R27 VPB.t8 VPB.t9 254.518
R28 VPB.t11 VPB.t8 254.518
R29 VPB.t2 VPB.t11 254.518
R30 VPB.t7 VPB.t2 254.518
R31 VPB.t0 VPB.t1 254.518
R32 VPB.t12 VPB.t13 254.518
R33 VPB.t4 VPB.t5 254.518
R34 VPB.t3 VPB.t4 254.518
R35 VPB.t6 VPB.t3 254.518
R36 VPB VPB.t6 204.207
R37 a_44_47.n1 a_44_47.t4 333.87
R38 a_44_47.n18 a_44_47.n17 332.611
R39 a_44_47.n12 a_44_47.n11 240.071
R40 a_44_47.n17 a_44_47.t5 233.145
R41 a_44_47.n8 a_44_47.t11 212.081
R42 a_44_47.n4 a_44_47.t15 212.081
R43 a_44_47.n3 a_44_47.t14 212.081
R44 a_44_47.n9 a_44_47.t17 212.081
R45 a_44_47.n14 a_44_47.n13 201.499
R46 a_44_47.n16 a_44_47.n15 201.139
R47 a_44_47.n6 a_44_47.n5 177.601
R48 a_44_47.n11 a_44_47.n10 152
R49 a_44_47.n8 a_44_47.n2 152
R50 a_44_47.n7 a_44_47.n6 152
R51 a_44_47.n8 a_44_47.t10 139.78
R52 a_44_47.n4 a_44_47.t16 139.78
R53 a_44_47.n3 a_44_47.t12 139.78
R54 a_44_47.n9 a_44_47.t13 139.78
R55 a_44_47.n1 a_44_47.n0 89.7238
R56 a_44_47.n14 a_44_47.n12 88.9268
R57 a_44_47.n8 a_44_47.n7 49.6611
R58 a_44_47.n10 a_44_47.n8 49.6611
R59 a_44_47.n16 a_44_47.n14 45.4742
R60 a_44_47.n5 a_44_47.n3 36.5157
R61 a_44_47.n13 a_44_47.t9 36.0005
R62 a_44_47.t0 a_44_47.n18 27.5805
R63 a_44_47.n18 a_44_47.t6 27.5805
R64 a_44_47.n0 a_44_47.t1 26.7697
R65 a_44_47.n5 a_44_47.n4 26.2914
R66 a_44_47.n15 a_44_47.t3 25.8467
R67 a_44_47.n15 a_44_47.t7 25.8467
R68 a_44_47.n0 a_44_47.t8 25.8467
R69 a_44_47.n13 a_44_47.t2 25.8467
R70 a_44_47.n6 a_44_47.n2 25.6005
R71 a_44_47.n11 a_44_47.n2 25.6005
R72 a_44_47.n17 a_44_47.n16 18.6276
R73 a_44_47.n7 a_44_47.n3 13.146
R74 a_44_47.n10 a_44_47.n9 13.146
R75 a_44_47.n12 a_44_47.n1 5.55539
R76 VGND.n9 VGND.t6 287.683
R77 VGND.n17 VGND.t10 284.471
R78 VGND.n34 VGND.n33 199.739
R79 VGND.n11 VGND.n10 198.964
R80 VGND.n8 VGND.n7 198.964
R81 VGND.n31 VGND.n2 198.964
R82 VGND.n26 VGND.n25 185
R83 VGND.n24 VGND.n23 185
R84 VGND.n25 VGND.n24 96.0005
R85 VGND.n18 VGND.n5 34.6358
R86 VGND.n22 VGND.n5 34.6358
R87 VGND.n2 VGND.t2 33.2313
R88 VGND.n18 VGND.n17 32.7534
R89 VGND.n24 VGND.t0 29.539
R90 VGND.n27 VGND.n1 29.01
R91 VGND.n16 VGND.n8 28.2358
R92 VGND.n32 VGND.n31 27.1064
R93 VGND.n25 VGND.t11 25.8467
R94 VGND.n10 VGND.t8 25.8467
R95 VGND.n10 VGND.t9 25.8467
R96 VGND.n7 VGND.t7 25.8467
R97 VGND.n7 VGND.t4 25.8467
R98 VGND.n33 VGND.t5 25.8467
R99 VGND.n33 VGND.t3 25.8467
R100 VGND.n2 VGND.t1 24.9236
R101 VGND.n12 VGND.n11 23.7181
R102 VGND.n31 VGND.n1 17.3181
R103 VGND.n23 VGND.n22 16.2598
R104 VGND.n12 VGND.n8 16.1887
R105 VGND.n34 VGND.n32 15.8123
R106 VGND.n17 VGND.n16 11.2946
R107 VGND.n26 VGND.n4 9.78163
R108 VGND.n13 VGND.n12 9.3005
R109 VGND.n14 VGND.n8 9.3005
R110 VGND.n16 VGND.n15 9.3005
R111 VGND.n17 VGND.n6 9.3005
R112 VGND.n19 VGND.n18 9.3005
R113 VGND.n20 VGND.n5 9.3005
R114 VGND.n22 VGND.n21 9.3005
R115 VGND.n4 VGND.n3 9.3005
R116 VGND.n28 VGND.n27 9.3005
R117 VGND.n29 VGND.n1 9.3005
R118 VGND.n31 VGND.n30 9.3005
R119 VGND.n32 VGND.n0 9.3005
R120 VGND.n35 VGND.n34 7.45014
R121 VGND.n11 VGND.n9 6.36409
R122 VGND.n23 VGND.n4 2.77786
R123 VGND.n27 VGND.n26 1.3288
R124 VGND.n13 VGND.n9 0.729313
R125 VGND.n35 VGND.n0 0.144329
R126 VGND.n14 VGND.n13 0.120292
R127 VGND.n15 VGND.n14 0.120292
R128 VGND.n15 VGND.n6 0.120292
R129 VGND.n19 VGND.n6 0.120292
R130 VGND.n20 VGND.n19 0.120292
R131 VGND.n21 VGND.n20 0.120292
R132 VGND.n21 VGND.n3 0.120292
R133 VGND.n28 VGND.n3 0.120292
R134 VGND.n29 VGND.n28 0.120292
R135 VGND.n30 VGND.n29 0.120292
R136 VGND.n30 VGND.n0 0.120292
R137 VGND VGND.n35 0.119086
R138 VNB.t3 VNB.t12 2790.94
R139 VNB.t13 VNB.t0 2762.46
R140 VNB.t1 VNB.t13 1381.23
R141 VNB.t2 VNB.t1 1324.27
R142 VNB.t0 VNB.t7 1238.83
R143 VNB.t10 VNB.t8 1224.6
R144 VNB.t11 VNB.t10 1224.6
R145 VNB.t9 VNB.t11 1224.6
R146 VNB.t5 VNB.t9 1224.6
R147 VNB.t12 VNB.t5 1224.6
R148 VNB.t7 VNB.t3 1224.6
R149 VNB.t6 VNB.t2 1224.6
R150 VNB.t4 VNB.t6 1224.6
R151 VNB VNB.t4 1181.88
R152 B1.n0 B1.t3 213.688
R153 B1.n2 B1.t2 213.688
R154 B1.n3 B1.t1 176.115
R155 B1.n0 B1.t0 167.958
R156 B1.n1 B1 159.226
R157 B1.n4 B1.n3 152
R158 B1.n2 B1.n1 54.8743
R159 B1.n3 B1.n2 15.5728
R160 B1.n4 B1 12.3876
R161 B1.n1 B1.n0 8.89896
R162 B1 B1.n4 6.60695
R163 X.n2 X.n1 352.245
R164 X.n2 X.n0 308.212
R165 X.n5 X.n3 255.659
R166 X.n5 X.n4 205.212
R167 X X.n2 31.0561
R168 X.n0 X.t5 27.5805
R169 X.n0 X.t6 27.5805
R170 X.n1 X.t7 27.5805
R171 X.n1 X.t4 27.5805
R172 X.n3 X.t3 25.8467
R173 X.n3 X.t1 25.8467
R174 X.n4 X.t0 25.8467
R175 X.n4 X.t2 25.8467
R176 X X.n5 23.0574
R177 A1.n0 A1.t1 208.868
R178 A1.n2 A1.t0 208.868
R179 A1.n0 A1 166.291
R180 A1.n4 A1.n3 152
R181 A1.n2 A1.t2 145.452
R182 A1.n1 A1.t3 139.78
R183 A1.n3 A1.n1 30.4799
R184 A1.n3 A1.n2 24.8093
R185 A1.n4 A1 19.5205
R186 A1 A1.n4 9.9205
R187 A1.n1 A1.n0 5.67109
R188 a_477_297.t2 a_477_297.n3 388.07
R189 a_477_297.n1 a_477_297.n0 347.283
R190 a_477_297.n1 a_477_297.t4 323.959
R191 a_477_297.n3 a_477_297.n2 289.24
R192 a_477_297.n3 a_477_297.n1 52.4754
R193 a_477_297.n2 a_477_297.t1 51.2205
R194 a_477_297.n2 a_477_297.t5 50.2355
R195 a_477_297.n0 a_477_297.t0 27.5805
R196 a_477_297.n0 a_477_297.t3 27.5805
R197 VPWR.n13 VPWR.t1 868.5
R198 VPWR.n1 VPWR.n0 603.231
R199 VPWR.n5 VPWR.t3 344.798
R200 VPWR.n4 VPWR.n3 311.587
R201 VPWR.n7 VPWR.n6 310.786
R202 VPWR.n14 VPWR.n13 32.7534
R203 VPWR.n12 VPWR.n4 28.2358
R204 VPWR.n0 VPWR.t6 27.5805
R205 VPWR.n0 VPWR.t7 27.5805
R206 VPWR.n3 VPWR.t2 27.5805
R207 VPWR.n3 VPWR.t0 27.5805
R208 VPWR.n6 VPWR.t4 27.5805
R209 VPWR.n6 VPWR.t5 27.5805
R210 VPWR.n8 VPWR.n7 23.7181
R211 VPWR.n8 VPWR.n4 16.1887
R212 VPWR.n14 VPWR.n1 13.177
R213 VPWR.n13 VPWR.n12 11.2946
R214 VPWR.n9 VPWR.n8 9.3005
R215 VPWR.n10 VPWR.n4 9.3005
R216 VPWR.n12 VPWR.n11 9.3005
R217 VPWR.n13 VPWR.n2 9.3005
R218 VPWR.n15 VPWR.n14 9.3005
R219 VPWR.n16 VPWR.n1 7.48186
R220 VPWR.n7 VPWR.n5 6.36409
R221 VPWR VPWR.n16 0.957047
R222 VPWR.n9 VPWR.n5 0.729313
R223 VPWR.n16 VPWR.n15 0.149039
R224 VPWR.n10 VPWR.n9 0.120292
R225 VPWR.n11 VPWR.n10 0.120292
R226 VPWR.n11 VPWR.n2 0.120292
R227 VPWR.n15 VPWR.n2 0.120292
R228 D1.n0 D1.t1 212.081
R229 D1.n2 D1.t2 212.081
R230 D1.n3 D1.n2 184.133
R231 D1.n0 D1.t3 151.811
R232 D1.n1 D1.t0 139.78
R233 D1.n1 D1.n0 52.5823
R234 D1.n3 D1 12.8005
R235 D1.n2 D1.n1 10.2247
R236 D1 D1.n3 2.47068
R237 A2.n0 A2.t3 212.081
R238 A2.n2 A2.t2 212.081
R239 A2.n1 A2 167.041
R240 A2.n3 A2.n2 161.494
R241 A2.n0 A2.t1 139.78
R242 A2.n2 A2.t0 139.78
R243 A2.n2 A2.n1 40.1672
R244 A2 A2.n3 23.3605
R245 A2.n1 A2.n0 22.6399
R246 A2.n3 A2 6.7205
R247 a_770_47.n1 a_770_47.n0 488.762
R248 a_770_47.n0 a_770_47.t2 25.8467
R249 a_770_47.n0 a_770_47.t3 25.8467
R250 a_770_47.n1 a_770_47.t0 25.8467
R251 a_770_47.t1 a_770_47.n1 25.8467
C0 C1 VPB 0.066906f
C1 A2 VPWR 0.036874f
C2 A1 X 3.88e-19
C3 B1 VGND 0.040136f
C4 B1 VPB 0.086422f
C5 C1 D1 0.057444f
C6 A1 VGND 0.02092f
C7 A2 X 0.002923f
C8 A1 VPB 0.07119f
C9 A2 VGND 0.039099f
C10 VPWR X 0.354689f
C11 A2 VPB 0.065638f
C12 VPWR VGND 0.153237f
C13 VPWR VPB 0.156021f
C14 X VGND 0.230147f
C15 VPWR D1 0.019105f
C16 X VPB 0.012057f
C17 C1 B1 0.066677f
C18 VGND VPB 0.011949f
C19 VGND D1 0.036145f
C20 B1 A1 0.040924f
C21 VPB D1 0.076906f
C22 C1 VPWR 0.018747f
C23 B1 VPWR 0.02028f
C24 A1 A2 0.038686f
C25 B1 X 4.01e-20
C26 A1 VPWR 0.03219f
C27 C1 VGND 0.037081f
C28 VGND VNB 0.855865f
C29 X VNB 0.061397f
C30 VPWR VNB 0.723115f
C31 A2 VNB 0.197804f
C32 A1 VNB 0.200042f
C33 B1 VNB 0.23339f
C34 C1 VNB 0.193028f
C35 D1 VNB 0.259318f
C36 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_0 VNB VPB VPWR VGND D1 C1 A2 A1 B1 Y
X0 Y.t1 B1.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1 VPWR.t1 A1.t0 a_313_369.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1216 pd=1.02 as=0.0896 ps=0.92 w=0.64 l=0.15
X2 a_427_47.t0 A1.t1 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_241_369.t1 C1.t0 a_169_369.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.0672 ps=0.85 w=0.64 l=0.15
X4 VGND.t2 C1.t1 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND.t3 A2.t0 a_427_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_169_369.t1 D1.t0 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1888 ps=1.87 w=0.64 l=0.15
X7 Y.t0 D1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.126 ps=1.44 w=0.42 l=0.15
X8 a_313_369.t1 B1.t1 a_241_369.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0896 pd=0.92 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_369.t0 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1952 pd=1.89 as=0.1216 ps=1.02 w=0.64 l=0.15
R0 B1.n0 B1.t1 271.527
R1 B1.n0 B1.t0 218.737
R2 B1.n1 B1.n0 152
R3 B1.n1 B1 8.22907
R4 B1 B1.n1 4.20621
R5 VGND.n7 VGND.t0 249.739
R6 VGND.n3 VGND.t3 244.573
R7 VGND.n2 VGND.n1 198.964
R8 VGND.n1 VGND.t1 51.4291
R9 VGND.n1 VGND.t2 48.5719
R10 VGND.n6 VGND.n5 34.6358
R11 VGND.n8 VGND.n7 13.4417
R12 VGND.n3 VGND.n2 12.6227
R13 VGND.n5 VGND.n4 9.3005
R14 VGND.n6 VGND.n0 9.3005
R15 VGND.n7 VGND.n6 5.64756
R16 VGND.n5 VGND.n2 4.51815
R17 VGND.n4 VGND.n3 0.389715
R18 VGND.n4 VGND.n0 0.120292
R19 VGND.n8 VGND.n0 0.120292
R20 VGND VGND.n8 0.0226354
R21 Y.n0 Y 591.174
R22 Y.n1 Y.n0 585
R23 Y.n5 Y.n4 234.756
R24 Y.n5 Y.n3 194.788
R25 Y.n0 Y.t2 52.3286
R26 Y.n4 Y.t4 40.0005
R27 Y.n4 Y.t1 40.0005
R28 Y.n3 Y.t3 40.0005
R29 Y.n3 Y.t0 40.0005
R30 Y Y.n5 6.28198
R31 Y.n2 Y.n1 4.96991
R32 Y.n1 Y 4.06638
R33 Y Y.n2 2.84494
R34 Y.n2 Y 1.20521
R35 VNB VNB.t0 1580.58
R36 VNB.t2 VNB.t1 1423.95
R37 VNB.t1 VNB.t3 1224.6
R38 VNB.t0 VNB.t2 1224.6
R39 VNB.t3 VNB.t4 1025.24
R40 A1.n1 A1.t1 208.816
R41 A1.n1 A1.t0 200.219
R42 A1.n2 A1.n1 98.3302
R43 A1.n0 A1 14.4598
R44 A1.n0 A1 1.7199
R45 A1.n2 A1.n0 1.48557
R46 A1 A1.n2 0.260964
R47 a_313_369.t0 a_313_369.n0 694.577
R48 a_313_369.n0 a_313_369.t2 43.0943
R49 a_313_369.n0 a_313_369.t1 43.0943
R50 VPWR VPWR.n0 605.673
R51 VPWR.n0 VPWR.t1 64.6411
R52 VPWR.n0 VPWR.t0 52.3286
R53 VPB VPB.t4 369.938
R54 VPB.t2 VPB.t0 313.707
R55 VPB.t1 VPB.t2 254.518
R56 VPB.t3 VPB.t1 213.084
R57 VPB.t4 VPB.t3 213.084
R58 a_427_47.t0 a_427_47.t1 60.0005
R59 C1.n0 C1.t0 270.358
R60 C1.n0 C1.t1 221.867
R61 C1.n1 C1.n0 152
R62 C1 C1.n1 7.78428
R63 C1.n1 C1 3.97888
R64 a_169_369.t0 a_169_369.t1 64.6411
R65 a_241_369.t0 a_241_369.t1 64.6411
R66 A2.n1 A2.t0 285.183
R67 A2.n0 A2.t1 285.07
R68 A2 A2.n0 153.882
R69 A2.n2 A2.n1 152
R70 A2.n1 A2.n0 58.5291
R71 A2 A2.n2 10.9181
R72 A2.n2 A2 1.88285
R73 D1.n1 D1.t0 286.344
R74 D1.n2 D1.t1 182.982
R75 D1.n3 D1.n2 152
R76 D1.n1 D1.n0 152
R77 D1.n2 D1.n1 68.7301
R78 D1.n0 D1 7.6805
R79 D1.n3 D1 6.4005
R80 D1 D1.n3 6.03479
R81 D1.n0 D1 4.75479
C0 VPB Y 0.018054f
C1 D1 Y 0.132027f
C2 VPB VPWR 0.075435f
C3 A1 A2 0.232507f
C4 C1 Y 0.164419f
C5 VPB VGND 0.010724f
C6 D1 VPWR 0.019822f
C7 D1 VGND 0.038081f
C8 C1 VPWR 0.044458f
C9 B1 Y 0.05037f
C10 A1 Y 0.028177f
C11 B1 VPWR 0.015622f
C12 C1 VGND 0.014397f
C13 VPB D1 0.097349f
C14 B1 VGND 0.0141f
C15 A2 Y 0.00255f
C16 A1 VPWR 0.019833f
C17 VPB C1 0.056631f
C18 A1 VGND 0.041712f
C19 A2 VPWR 0.024783f
C20 D1 C1 0.076113f
C21 VPB B1 0.054808f
C22 A2 VGND 0.039777f
C23 VPB A1 0.081929f
C24 Y VPWR 0.0636f
C25 VPB A2 0.102621f
C26 C1 B1 0.16078f
C27 Y VGND 0.201631f
C28 C1 A1 0.00108f
C29 VPWR VGND 0.061517f
C30 B1 A1 0.134443f
C31 C1 A2 4.38e-19
C32 VGND VNB 0.425772f
C33 VPWR VNB 0.332346f
C34 Y VNB 0.060944f
C35 A2 VNB 0.257876f
C36 A1 VNB 0.136357f
C37 B1 VNB 0.109476f
C38 C1 VNB 0.115065f
C39 D1 VNB 0.236403f
C40 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_1 VNB VPWR VGND VPB D1 C1 B1 A1 Y A2
X0 a_316_297.t1 C1.t0 a_217_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.1725 ps=1.345 w=1 l=0.15
X1 Y.t0 D1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND.t2 C1.t1 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 a_420_297.t2 B1.t0 a_316_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR.t0 A1.t0 a_420_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND.t1 A2.t0 a_568_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y.t3 B1.t1 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.24 as=0.12025 ps=1.02 w=0.65 l=0.15
X7 a_420_297.t1 A2.t1 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.1375 ps=1.275 w=1 l=0.15
X8 a_217_297.t1 D1.t1 Y.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47.t1 A1.t1 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.19175 ps=1.24 w=0.65 l=0.15
R0 C1.n0 C1.t0 228.613
R1 C1.n0 C1.t1 161.29
R2 C1.n1 C1.n0 152
R3 C1.n1 C1 10.8901
R4 C1 C1.n1 2.10199
R5 a_217_297.t0 a_217_297.t1 67.9655
R6 a_316_297.t0 a_316_297.t1 72.8905
R7 VPB VPB.t4 511.995
R8 VPB.t0 VPB.t2 432.087
R9 VPB.t1 VPB.t0 307.788
R10 VPB.t4 VPB.t1 292.991
R11 VPB.t2 VPB.t3 251.559
R12 D1.n0 D1.t1 238.59
R13 D1.n0 D1.t0 166.291
R14 D1.n1 D1.n0 152
R15 D1.n1 D1 8.10717
R16 D1 D1.n1 1.56494
R17 VGND.n7 VGND.t0 276.245
R18 VGND.n3 VGND.t1 244.48
R19 VGND.n2 VGND.n1 199.352
R20 VGND.n1 VGND.t3 43.3851
R21 VGND.n6 VGND.n5 34.6358
R22 VGND.n5 VGND.n2 30.1181
R23 VGND.n1 VGND.t2 24.9236
R24 VGND.n8 VGND.n7 15.7005
R25 VGND.n6 VGND.n0 9.3005
R26 VGND.n5 VGND.n4 9.3005
R27 VGND.n3 VGND.n2 6.47776
R28 VGND.n7 VGND.n6 4.51815
R29 VGND.n4 VGND.n3 0.185416
R30 VGND.n4 VGND.n0 0.120292
R31 VGND.n8 VGND.n0 0.120292
R32 VGND VGND.n8 0.0226354
R33 Y Y.n0 590.653
R34 Y.n6 Y.n0 585
R35 Y.n5 Y.n0 585
R36 Y.n3 Y.n1 153.362
R37 Y.n3 Y.n2 97.7818
R38 Y.n0 Y.t1 96.5305
R39 Y.n1 Y.t4 80.3082
R40 Y.n2 Y.t2 41.0927
R41 Y.n4 Y.n3 36.6227
R42 Y.n2 Y.t0 29.984
R43 Y.n1 Y.t3 28.6159
R44 Y Y.n4 10.4732
R45 Y Y.n5 5.81868
R46 Y Y.n6 5.65245
R47 Y.n6 Y 5.65245
R48 Y.n5 Y 5.48621
R49 Y.n4 Y 0.831669
R50 VNB VNB.t0 2349.51
R51 VNB.t3 VNB.t4 2107.44
R52 VNB.t0 VNB.t2 1523.62
R53 VNB.t2 VNB 1338.51
R54 VNB.t4 VNB.t1 1167.64
R55 VNB VNB.t3 142.395
R56 B1.n0 B1.t0 238.25
R57 B1.n0 B1.t1 161.212
R58 B1.n1 B1.n0 152
R59 B1 B1.n1 11.4041
R60 B1.n1 B1 2.13383
R61 a_420_297.n0 a_420_297.t1 698.797
R62 a_420_297.n0 a_420_297.t2 86.6805
R63 a_420_297.t0 a_420_297.n0 27.5805
R64 A1.n0 A1.t0 327.615
R65 A1 A1.n0 157.531
R66 A1.n0 A1.t1 154.554
R67 VPWR VPWR.n0 316.772
R68 VPWR.n0 VPWR.t1 27.5805
R69 VPWR.n0 VPWR.t0 26.5955
R70 A2.n0 A2.t1 235.471
R71 A2.n0 A2.t0 157.785
R72 A2.n1 A2.n0 152
R73 A2 A2.n1 30.2067
R74 A2.n1 A2 4.97828
R75 a_568_47.t0 a_568_47.t1 48.0005
C0 C1 A2 1.74e-19
C1 VPB VPWR 0.076301f
C2 D1 Y 0.162205f
C3 B1 A1 0.072348f
C4 B1 A2 7.88e-19
C5 C1 Y 0.041564f
C6 D1 VPWR 0.065652f
C7 VPB VGND 0.007886f
C8 B1 Y 0.042331f
C9 C1 VPWR 0.049898f
C10 A1 A2 0.086112f
C11 D1 VGND 0.019147f
C12 B1 VPWR 0.043278f
C13 A1 Y 0.008532f
C14 C1 VGND 0.01826f
C15 A1 VPWR 0.020171f
C16 B1 VGND 0.014694f
C17 A2 Y 0.026631f
C18 VPB D1 0.038973f
C19 A2 VPWR 0.022064f
C20 A1 VGND 0.024596f
C21 VPB C1 0.032498f
C22 A2 VGND 0.099038f
C23 Y VPWR 0.074336f
C24 D1 C1 0.146047f
C25 VPB B1 0.035036f
C26 Y VGND 0.273751f
C27 VPB A1 0.036628f
C28 VPWR VGND 0.073379f
C29 D1 A1 1.14e-19
C30 VPB A2 0.034138f
C31 C1 B1 0.167115f
C32 C1 A1 2.99e-19
C33 VPB Y 0.016067f
C34 D1 A2 7.52e-20
C35 VGND VNB 0.474028f
C36 VPWR VNB 0.370362f
C37 Y VNB 0.093275f
C38 A2 VNB 0.149761f
C39 A1 VNB 0.106396f
C40 B1 VNB 0.09744f
C41 C1 VNB 0.096827f
C42 D1 VNB 0.122118f
C43 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_2 VNB VPB VGND VPWR A1 A2 D1 C1 B1 Y
X0 a_467_297.t3 B1.t0 a_28_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X1 a_287_297.t1 D1.t0 Y.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR.t3 A2.t0 a_467_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X3 a_923_47.t1 A2.t1 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 Y.t2 B1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_28_297.t0 B1.t2 a_467_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND.t4 C1.t0 Y.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X7 a_28_297.t2 C1.t1 a_287_297.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X8 Y.t3 A1.t0 a_923_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND.t3 A2.t2 a_684_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17875 ps=1.2 w=0.65 l=0.15
X10 Y.t6 D1.t1 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND.t0 B1.t3 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.105625 ps=0.975 w=0.65 l=0.15
X12 Y.t8 D1.t2 a_115_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_467_297.t1 A1.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.16 ps=1.32 w=1 l=0.15
X14 VGND.t5 D1.t3 Y.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y.t9 C1.t2 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.12675 ps=1.04 w=0.65 l=0.15
X16 VPWR.t1 A1.t2 a_467_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X17 a_115_297.t0 C1.t3 a_28_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X18 a_467_297.t0 A2.t3 VPWR.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_684_47.t0 A1.t3 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.2 as=0.091 ps=0.93 w=0.65 l=0.15
R0 B1.n2 B1.t0 225.226
R1 B1.n0 B1.t2 212.081
R2 B1.n0 B1.t1 172.644
R3 B1 B1.n0 164.8
R4 B1 B1.n2 156.964
R5 B1.n1 B1.t3 139.78
R6 B1.n1 B1.n0 46.0096
R7 B1.n2 B1.n1 3.65202
R8 a_28_297.t0 a_28_297.n1 889.635
R9 a_28_297.n1 a_28_297.n0 585
R10 a_28_297.n1 a_28_297.t3 427.512
R11 a_28_297.n0 a_28_297.t1 35.4605
R12 a_28_297.n0 a_28_297.t2 27.5805
R13 a_467_297.n3 a_467_297.n2 657.684
R14 a_467_297.n1 a_467_297.t1 373.339
R15 a_467_297.n2 a_467_297.t4 318.594
R16 a_467_297.n1 a_467_297.n0 295.32
R17 a_467_297.n2 a_467_297.n1 45.5073
R18 a_467_297.n0 a_467_297.t5 27.5805
R19 a_467_297.n0 a_467_297.t0 27.5805
R20 a_467_297.n3 a_467_297.t2 27.5805
R21 a_467_297.t3 a_467_297.n3 27.5805
R22 VPB.t2 VPB.t4 562.306
R23 VPB.t9 VPB.t1 278.193
R24 VPB.t6 VPB.t3 278.193
R25 VPB.t0 VPB.t9 254.518
R26 VPB.t4 VPB.t0 254.518
R27 VPB.t3 VPB.t2 254.518
R28 VPB.t8 VPB.t6 254.518
R29 VPB.t5 VPB.t8 254.518
R30 VPB.t7 VPB.t5 254.518
R31 VPB VPB.t7 210.125
R32 D1.n0 D1.t0 212.081
R33 D1.n1 D1.t2 212.081
R34 D1.n0 D1.t3 139.78
R35 D1.n1 D1.t1 139.78
R36 D1 D1.n2 71.3012
R37 D1.n2 D1.n0 35.7245
R38 D1.n2 D1.n1 20.8952
R39 Y Y.n0 708.064
R40 Y.n6 Y.t3 304.639
R41 Y.n7 Y.n6 192.284
R42 Y.n8 Y.n7 185
R43 Y.n2 Y.t4 159.696
R44 Y.n2 Y.n1 96.8044
R45 Y.n4 Y.n3 95.698
R46 Y Y.n8 38.0263
R47 Y.n4 Y.n2 37.2875
R48 Y.n5 Y.n4 37.2875
R49 Y.n3 Y.t1 31.3851
R50 Y.n3 Y.t9 28.6159
R51 Y.n0 Y.t7 27.5805
R52 Y.n0 Y.t8 27.5805
R53 Y.n7 Y.t0 25.8467
R54 Y.n7 Y.t2 25.8467
R55 Y.n1 Y.t5 25.8467
R56 Y.n1 Y.t6 25.8467
R57 Y.n6 Y.n5 8.38671
R58 Y.n8 Y.n5 0.441879
R59 a_287_297.t0 a_287_297.t1 55.1605
R60 A2.n1 A2.t0 212.081
R61 A2.n2 A2.t3 212.081
R62 A2 A2.n0 163.57
R63 A2 A2.n3 157.169
R64 A2.n2 A2.t2 141.77
R65 A2.n0 A2.t1 141.052
R66 A2.n3 A2.n1 46.0423
R67 A2.n3 A2.n2 15.8274
R68 A2.n1 A2.n0 2.87811
R69 VPWR.n2 VPWR.n1 604.384
R70 VPWR.n2 VPWR.n0 604.201
R71 VPWR.n1 VPWR.t0 31.5205
R72 VPWR.n1 VPWR.t3 31.5205
R73 VPWR.n0 VPWR.t2 27.5805
R74 VPWR.n0 VPWR.t1 27.5805
R75 VPWR VPWR.n2 1.35132
R76 VGND.n6 VGND.n3 204.96
R77 VGND.n5 VGND.n4 198.964
R78 VGND.n9 VGND.n2 198.964
R79 VGND.n12 VGND.n11 198.964
R80 VGND.n4 VGND.t1 38.7697
R81 VGND.n2 VGND.t7 36.0005
R82 VGND.n2 VGND.t5 36.0005
R83 VGND.n4 VGND.t0 33.2313
R84 VGND.n3 VGND.t2 32.3082
R85 VGND.n3 VGND.t3 31.3851
R86 VGND.n5 VGND.n1 29.7417
R87 VGND.n11 VGND.t6 25.8467
R88 VGND.n11 VGND.t4 25.8467
R89 VGND.n10 VGND.n9 23.7181
R90 VGND.n9 VGND.n1 20.7064
R91 VGND.n12 VGND.n10 20.3299
R92 VGND.n7 VGND.n1 9.3005
R93 VGND.n9 VGND.n8 9.3005
R94 VGND.n10 VGND.n0 9.3005
R95 VGND.n13 VGND.n12 7.25484
R96 VGND.n6 VGND.n5 6.51182
R97 VGND.n7 VGND.n6 0.184042
R98 VGND.n13 VGND.n0 0.146813
R99 VGND.n8 VGND.n7 0.120292
R100 VGND.n8 VGND.n0 0.120292
R101 VGND VGND.n13 0.116571
R102 a_923_47.t0 a_923_47.t1 51.6928
R103 VNB.t0 VNB.t4 1993.53
R104 VNB.t1 VNB.t2 1537.86
R105 VNB.t7 VNB.t9 1537.86
R106 VNB.t4 VNB.t5 1409.71
R107 VNB.t9 VNB.t1 1352.75
R108 VNB.t5 VNB.t3 1224.6
R109 VNB.t2 VNB.t0 1224.6
R110 VNB.t8 VNB.t7 1224.6
R111 VNB.t6 VNB.t8 1224.6
R112 VNB VNB.t6 1011
R113 C1.n0 C1.t1 236.18
R114 C1.n1 C1.t3 229.754
R115 C1 C1.n1 225.797
R116 C1 C1.n0 177.655
R117 C1.n0 C1.t2 163.881
R118 C1.n1 C1.t0 157.453
R119 A1.n0 A1.t1 236.18
R120 A1.n1 A1.t2 229.952
R121 A1 A1.n0 224.511
R122 A1 A1.n1 178.602
R123 A1.n0 A1.t0 163.881
R124 A1.n1 A1.t3 157.653
R125 a_684_47.t0 a_684_47.t1 101.538
R126 a_115_297.t0 a_115_297.t1 55.1605
C0 A1 Y 0.150106f
C1 D1 VGND 0.03078f
C2 B1 VPWR 0.017619f
C3 A1 VPWR 0.04574f
C4 B1 VGND 0.031268f
C5 A2 Y 0.078325f
C6 VPB C1 0.078994f
C7 A1 VGND 0.028794f
C8 A2 VPWR 0.029225f
C9 VPB D1 0.05566f
C10 A2 VGND 0.032887f
C11 Y VPWR 0.028355f
C12 C1 D1 0.214971f
C13 VPB B1 0.06877f
C14 Y VGND 0.575217f
C15 C1 B1 0.071108f
C16 VPB A1 0.084466f
C17 VPWR VGND 0.105161f
C18 VPB A2 0.059575f
C19 VPB Y 0.01406f
C20 VPB VPWR 0.103728f
C21 B1 A1 0.038758f
C22 C1 Y 0.222208f
C23 C1 VPWR 0.023114f
C24 VPB VGND 0.009072f
C25 D1 Y 0.09005f
C26 A1 A2 0.221142f
C27 B1 Y 0.196168f
C28 D1 VPWR 0.014836f
C29 C1 VGND 0.036267f
C30 VGND VNB 0.621187f
C31 VPWR VNB 0.515941f
C32 Y VNB 0.086979f
C33 A2 VNB 0.187789f
C34 A1 VNB 0.260873f
C35 B1 VNB 0.194681f
C36 D1 VNB 0.177744f
C37 C1 VNB 0.256559f
C38 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_4 VNB VPB VGND VPWR A1 Y D1 C1 A2 B1
X0 Y.t3 D1.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_455_297.t3 B1.t0 a_821_297# VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X2 a_28_297.t3 D1.t1 Y.t4 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_821_297# A2.t0 VPWR.t1 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4 a_28_297.t4 C1.t0 a_455_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_455_297.t5 C1.t1 a_28_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND.t4 D1.t2 Y.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND.t10 B1.t1 Y.t13 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR.t0 A2.t1 a_821_297# VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2 ps=1.4 w=1 l=0.15
X9 Y.t7 D1.t3 a_28_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10 Y.t8 C1.t2 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND.t3 D1.t4 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y.t0 D1.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 a_821_297# B1.t2 a_455_297.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 Y.t14 B1.t3 VGND.t11 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y.t6 D1.t6 a_28_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y.t9 C1.t3 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X17 a_1205_47.t3 A2.t2 VGND.t14 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_28_297.t6 C1.t4 a_455_297.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X19 Y.t15 B1.t4 VGND.t12 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X20 a_1205_47.t2 A2.t3 VGND.t15 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND.t8 C1.t5 Y.t10 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VGND.t9 C1.t6 Y.t11 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VPWR.t2 A1.t0 a_821_297# VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X25 a_1205_47.t4 A1.t1 Y.t12 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X26 a_28_297.t0 D1.t7 Y.t5 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND.t0 A2.t4 a_1205_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_455_297.t1 B1.t5 a_821_297# VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X30 a_1205_47.t5 A1.t2 Y.t17 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X31 VGND.t1 A2.t5 a_1205_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.121875 ps=1.025 w=0.65 l=0.15
X32 VPWR.t3 A1.t3 a_821_297# VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X33 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X35 a_455_297.t7 C1.t7 a_28_297.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 a_821_297# B1.t6 a_455_297.t0 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X37 VGND.t13 B1.t7 Y.t16 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.091 ps=0.93 w=0.65 l=0.15
R0 D1.n6 D1.t3 213.542
R1 D1.n3 D1.t6 212.081
R2 D1.n1 D1.t7 212.081
R3 D1.n5 D1.t1 212.081
R4 D1.n4 D1.n0 152
R5 D1.n8 D1.n7 152
R6 D1.n3 D1.t0 139.78
R7 D1.n1 D1.t2 139.78
R8 D1.n5 D1.t4 139.78
R9 D1.n6 D1.t5 139.78
R10 D1.n2 D1.n0 86.3858
R11 D1.n4 D1.n3 49.6611
R12 D1.n7 D1.n5 36.5157
R13 D1.n2 D1.n1 35.7937
R14 D1.n7 D1.n6 24.8308
R15 D1.n3 D1.n2 20.3621
R16 D1.n8 D1.n0 17.0672
R17 D1.n5 D1.n4 13.146
R18 D1 D1.n8 2.5103
R19 VGND.n44 VGND.t2 284.678
R20 VGND.n23 VGND.t13 284.471
R21 VGND.n13 VGND.n12 203.906
R22 VGND.n15 VGND.n14 198.964
R23 VGND.n27 VGND.n8 198.964
R24 VGND.n30 VGND.n29 198.964
R25 VGND.n34 VGND.n5 198.964
R26 VGND.n42 VGND.n2 198.964
R27 VGND.n37 VGND.n36 185
R28 VGND.n36 VGND.t4 40.6159
R29 VGND.n29 VGND.t8 36.9236
R30 VGND.n29 VGND.t12 35.0774
R31 VGND.n17 VGND.n16 34.6358
R32 VGND.n17 VGND.n10 34.6358
R33 VGND.n21 VGND.n10 34.6358
R34 VGND.n22 VGND.n21 34.6358
R35 VGND.n23 VGND.n22 32.377
R36 VGND.n27 VGND.n7 27.8593
R37 VGND.n30 VGND.n28 27.1064
R38 VGND.n34 VGND.n4 27.1064
R39 VGND.n38 VGND.n35 26.4529
R40 VGND.n36 VGND.t7 25.8467
R41 VGND.n12 VGND.t14 25.8467
R42 VGND.n12 VGND.t0 25.8467
R43 VGND.n14 VGND.t15 25.8467
R44 VGND.n14 VGND.t1 25.8467
R45 VGND.n8 VGND.t11 25.8467
R46 VGND.n8 VGND.t10 25.8467
R47 VGND.n5 VGND.t6 25.8467
R48 VGND.n5 VGND.t9 25.8467
R49 VGND.n2 VGND.t5 25.8467
R50 VGND.n2 VGND.t3 25.8467
R51 VGND.n42 VGND.n1 24.0946
R52 VGND.n37 VGND.n1 21.7292
R53 VGND.n43 VGND.n42 20.3299
R54 VGND.n44 VGND.n43 18.4476
R55 VGND.n30 VGND.n4 17.3181
R56 VGND.n35 VGND.n34 17.3181
R57 VGND.n28 VGND.n27 16.5652
R58 VGND.n16 VGND.n15 14.6829
R59 VGND.n23 VGND.n7 11.6711
R60 VGND.n45 VGND.n44 9.3005
R61 VGND.n16 VGND.n11 9.3005
R62 VGND.n18 VGND.n17 9.3005
R63 VGND.n19 VGND.n10 9.3005
R64 VGND.n21 VGND.n20 9.3005
R65 VGND.n22 VGND.n9 9.3005
R66 VGND.n24 VGND.n23 9.3005
R67 VGND.n25 VGND.n7 9.3005
R68 VGND.n27 VGND.n26 9.3005
R69 VGND.n28 VGND.n6 9.3005
R70 VGND.n31 VGND.n30 9.3005
R71 VGND.n32 VGND.n4 9.3005
R72 VGND.n34 VGND.n33 9.3005
R73 VGND.n35 VGND.n3 9.3005
R74 VGND.n39 VGND.n38 9.3005
R75 VGND.n40 VGND.n1 9.3005
R76 VGND.n42 VGND.n41 9.3005
R77 VGND.n43 VGND.n0 9.3005
R78 VGND.n15 VGND.n13 6.82082
R79 VGND.n13 VGND.n11 0.69121
R80 VGND.n38 VGND.n37 0.121255
R81 VGND.n18 VGND.n11 0.120292
R82 VGND.n19 VGND.n18 0.120292
R83 VGND.n20 VGND.n19 0.120292
R84 VGND.n20 VGND.n9 0.120292
R85 VGND.n24 VGND.n9 0.120292
R86 VGND.n25 VGND.n24 0.120292
R87 VGND.n26 VGND.n25 0.120292
R88 VGND.n26 VGND.n6 0.120292
R89 VGND.n31 VGND.n6 0.120292
R90 VGND.n32 VGND.n31 0.120292
R91 VGND.n33 VGND.n32 0.120292
R92 VGND.n33 VGND.n3 0.120292
R93 VGND.n39 VGND.n3 0.120292
R94 VGND.n40 VGND.n39 0.120292
R95 VGND.n41 VGND.n40 0.120292
R96 VGND.n41 VGND.n0 0.120292
R97 VGND.n45 VGND.n0 0.120292
R98 VGND VGND.n45 0.0213333
R99 Y.n2 Y.n0 331.022
R100 Y.n2 Y.n1 298.089
R101 Y.n3 Y.t12 275.599
R102 Y.n3 Y.t17 210.846
R103 Y.n5 Y.n4 185
R104 Y.n7 Y.n6 185
R105 Y.n9 Y.n8 185
R106 Y.n11 Y.n10 185
R107 Y.n13 Y.n12 185
R108 Y.n15 Y.n14 185
R109 Y.n5 Y.n3 102.879
R110 Y Y.n2 73.8471
R111 Y.n13 Y.n11 63.8408
R112 Y.n9 Y.n7 62.0839
R113 Y.n7 Y.n5 57.8173
R114 Y.n11 Y.n9 57.8173
R115 Y.n15 Y.n13 57.6233
R116 Y Y.n15 30.2635
R117 Y.n1 Y.t4 27.5805
R118 Y.n1 Y.t7 27.5805
R119 Y.n0 Y.t5 27.5805
R120 Y.n0 Y.t6 27.5805
R121 Y.n12 Y.t2 25.8467
R122 Y.n12 Y.t3 25.8467
R123 Y.n10 Y.t11 25.8467
R124 Y.n10 Y.t9 25.8467
R125 Y.n8 Y.t10 25.8467
R126 Y.n8 Y.t8 25.8467
R127 Y.n6 Y.t13 25.8467
R128 Y.n6 Y.t15 25.8467
R129 Y.n4 Y.t16 25.8467
R130 Y.n4 Y.t14 25.8467
R131 Y.n14 Y.t1 24.9236
R132 Y.n14 Y.t0 24.9236
R133 VNB.t14 VNB.t17 4015.53
R134 VNB.t17 VNB.t10 2449.19
R135 VNB.t8 VNB.t13 1537.86
R136 VNB.t10 VNB.t1 1495.15
R137 VNB.t4 VNB.t7 1452.43
R138 VNB.t0 VNB.t15 1224.6
R139 VNB.t16 VNB.t0 1224.6
R140 VNB.t1 VNB.t16 1224.6
R141 VNB.t12 VNB.t14 1224.6
R142 VNB.t11 VNB.t12 1224.6
R143 VNB.t13 VNB.t11 1224.6
R144 VNB.t6 VNB.t8 1224.6
R145 VNB.t9 VNB.t6 1224.6
R146 VNB.t7 VNB.t9 1224.6
R147 VNB.t5 VNB.t4 1224.6
R148 VNB.t3 VNB.t5 1224.6
R149 VNB.t2 VNB.t3 1196.12
R150 VNB VNB.t2 968.285
R151 B1.n2 B1.t6 248.595
R152 B1.n4 B1.t5 212.081
R153 B1.n1 B1.t2 212.081
R154 B1.n12 B1.t0 212.081
R155 B1.n7 B1.n2 169.067
R156 B1 B1.n13 160.534
R157 B1.n7 B1.n6 152
R158 B1.n9 B1.n8 152
R159 B1.n11 B1.n0 152
R160 B1.n13 B1.t4 141.242
R161 B1.n10 B1.t1 139.78
R162 B1.n5 B1.t3 139.78
R163 B1.n3 B1.t7 139.78
R164 B1.n13 B1.n12 46.7399
R165 B1.n10 B1.n9 37.9763
R166 B1.n6 B1.n5 24.8308
R167 B1.n6 B1.n4 23.3702
R168 B1.n8 B1.n7 17.0672
R169 B1.n8 B1.n0 17.0672
R170 B1.n4 B1.n3 14.6066
R171 B1.n5 B1.n1 14.6066
R172 B1.n3 B1.n2 11.6853
R173 B1.n11 B1.n10 11.6853
R174 B1.n9 B1.n1 10.2247
R175 B1 B1.n0 8.53383
R176 B1.n12 B1.n11 2.92171
R177 a_455_297.n3 a_455_297.n1 331.17
R178 a_455_297.n4 a_455_297.n0 331.022
R179 a_455_297.n3 a_455_297.n2 298.717
R180 a_455_297.n5 a_455_297.n4 298.717
R181 a_455_297.n4 a_455_297.n3 75.8308
R182 a_455_297.n2 a_455_297.t6 27.5805
R183 a_455_297.n2 a_455_297.t5 27.5805
R184 a_455_297.n1 a_455_297.t4 27.5805
R185 a_455_297.n1 a_455_297.t7 27.5805
R186 a_455_297.n0 a_455_297.t0 27.5805
R187 a_455_297.n0 a_455_297.t1 27.5805
R188 a_455_297.n5 a_455_297.t2 27.5805
R189 a_455_297.t3 a_455_297.n5 27.5805
R190 VPB.t14 VPB.t13 816.822
R191 VPB.t15 VPB.t14 591.9
R192 VPB.t10 VPB.t7 562.306
R193 VPB.t12 VPB.t15 509.034
R194 VPB.t4 VPB.t12 260.437
R195 VPB.t5 VPB.t4 254.518
R196 VPB.t6 VPB.t5 254.518
R197 VPB.t7 VPB.t6 254.518
R198 VPB.t9 VPB.t10 254.518
R199 VPB.t8 VPB.t9 254.518
R200 VPB.t11 VPB.t8 254.518
R201 VPB.t0 VPB.t11 254.518
R202 VPB.t1 VPB.t0 254.518
R203 VPB.t3 VPB.t1 254.518
R204 VPB.t2 VPB.t3 254.518
R205 VPB VPB.t2 195.327
R206 a_28_297.n4 a_28_297.t2 376.236
R207 a_28_297.n2 a_28_297.t6 375.252
R208 a_28_297.n5 a_28_297.n4 296.406
R209 a_28_297.n3 a_28_297.n0 296.406
R210 a_28_297.n2 a_28_297.n1 296.406
R211 a_28_297.n3 a_28_297.n2 57.9373
R212 a_28_297.n4 a_28_297.n3 57.9373
R213 a_28_297.n0 a_28_297.t7 27.5805
R214 a_28_297.n0 a_28_297.t0 27.5805
R215 a_28_297.n1 a_28_297.t5 27.5805
R216 a_28_297.n1 a_28_297.t4 27.5805
R217 a_28_297.n5 a_28_297.t1 27.5805
R218 a_28_297.t3 a_28_297.n5 27.5805
R219 A2.n9 A2.t1 225.957
R220 A2.n4 A2.t0 212.081
R221 A2.n7 A2.n2 212.081
R222 A2.n11 A2.n8 212.081
R223 A2.n9 A2.n1 169.067
R224 A2.n5 A2.n0 152
R225 A2.n15 A2.n14 152
R226 A2.n12 A2.n1 152
R227 A2.n3 A2.t2 139.78
R228 A2.n10 A2.t5 139.78
R229 A2.n13 A2.t3 139.78
R230 A2.n6 A2.t4 139.78
R231 A2.n3 A2.n0 106.746
R232 A2.n5 A2.n4 38.7066
R233 A2.n11 A2.n10 38.7066
R234 A2.n14 A2.n13 26.2914
R235 A2.n14 A2.n7 25.5611
R236 A2.n13 A2.n12 23.3702
R237 A2.n15 A2.n1 17.0672
R238 A2.n6 A2.n5 13.146
R239 A2 A2.n0 12.2985
R240 A2.n4 A2.n3 10.955
R241 A2.n7 A2.n6 10.955
R242 A2.n10 A2.n9 10.2247
R243 A2 A2.n15 4.76913
R244 A2.n12 A2.n11 0.730803
R245 VPWR.n4 VPWR.t1 343.628
R246 VPWR.n8 VPWR.t3 338.533
R247 VPWR.n10 VPWR.t2 338.531
R248 VPWR.n3 VPWR.t0 338.271
R249 VPWR.n7 VPWR.n2 34.6358
R250 VPWR.n9 VPWR.n8 30.8711
R251 VPWR.n4 VPWR.n3 14.2446
R252 VPWR.n8 VPWR.n7 13.5534
R253 VPWR.n5 VPWR.n2 9.3005
R254 VPWR.n7 VPWR.n6 9.3005
R255 VPWR.n8 VPWR.n1 9.3005
R256 VPWR.n9 VPWR.n0 9.3005
R257 VPWR.n10 VPWR.n9 9.03579
R258 VPWR.n11 VPWR.n10 8.35406
R259 VPWR.n3 VPWR.n2 2.25932
R260 VPWR VPWR.n11 1.5595
R261 VPWR.n5 VPWR.n4 0.981597
R262 VPWR.n11 VPWR.n0 0.147187
R263 VPWR.n6 VPWR.n5 0.120292
R264 VPWR.n6 VPWR.n1 0.120292
R265 VPWR.n1 VPWR.n0 0.120292
R266 C1.n13 C1.t7 215.001
R267 C1.n3 C1.t4 212.081
R268 C1.n1 C1.t1 212.081
R269 C1.n10 C1.t0 212.081
R270 C1.n6 C1.n2 170.528
R271 C1 C1.n13 163.546
R272 C1.n6 C1.n5 152
R273 C1.n8 C1.n7 152
R274 C1.n11 C1.n0 152
R275 C1.n12 C1.t3 139.78
R276 C1.n9 C1.t6 139.78
R277 C1.n4 C1.t2 139.78
R278 C1.n2 C1.t5 139.78
R279 C1.n12 C1.n11 40.8975
R280 C1.n5 C1.n3 36.5157
R281 C1.n9 C1.n8 27.752
R282 C1.n8 C1.n1 23.3702
R283 C1.n7 C1.n6 17.0672
R284 C1.n7 C1.n0 17.0672
R285 C1.n5 C1.n4 14.6066
R286 C1.n3 C1.n2 11.6853
R287 C1.n4 C1.n1 11.6853
R288 C1.n10 C1.n9 11.6853
R289 C1.n11 C1.n10 10.2247
R290 C1.n13 C1.n12 8.76414
R291 C1 C1.n0 5.52207
R292 a_1205_47.n1 a_1205_47.t5 345.574
R293 a_1205_47.t3 a_1205_47.n3 273.154
R294 a_1205_47.n1 a_1205_47.n0 185
R295 a_1205_47.n3 a_1205_47.n2 185
R296 a_1205_47.n3 a_1205_47.n1 65.7548
R297 a_1205_47.n0 a_1205_47.t4 42.462
R298 a_1205_47.n0 a_1205_47.t0 26.7697
R299 a_1205_47.n2 a_1205_47.t1 25.8467
R300 a_1205_47.n2 a_1205_47.t2 25.8467
R301 A1.n14 A1.t0 242.754
R302 A1.n5 A1.n4 212.081
R303 A1.n9 A1.t3 212.081
R304 A1.n12 A1.n1 212.081
R305 A1.n7 A1.n6 169.067
R306 A1.n6 A1.t1 157.308
R307 A1.n8 A1.n7 152
R308 A1.n10 A1.n0 152
R309 A1.n16 A1.n15 152
R310 A1.n14 A1.n13 139.78
R311 A1.n11 A1.t2 139.78
R312 A1.n3 A1.n2 139.78
R313 A1.n5 A1.n3 35.055
R314 A1.n12 A1.n11 30.6732
R315 A1.n9 A1.n8 26.2914
R316 A1.n10 A1.n9 23.3702
R317 A1.n15 A1.n14 21.9096
R318 A1 A1.n16 19.577
R319 A1.n7 A1.n0 17.0672
R320 A1.n16 A1.n0 17.0672
R321 A1.n6 A1.n5 10.2247
R322 A1.n15 A1.n12 10.2247
R323 A1.n11 A1.n10 8.76414
R324 A1.n8 A1.n3 4.38232
C0 a_821_297# C1 3.62e-20
C1 A1 Y 0.131455f
C2 C1 VGND 0.071825f
C3 B1 VPWR 0.03286f
C4 a_821_297# B1 0.056036f
C5 A1 VPWR 0.082572f
C6 A2 Y 2.2e-20
C7 B1 VGND 0.073659f
C8 a_821_297# A1 0.211132f
C9 VPB D1 0.122036f
C10 A1 VGND 0.040704f
C11 A2 VPWR 0.0758f
C12 a_821_297# A2 0.2275f
C13 VPB C1 0.135632f
C14 A2 VGND 0.070085f
C15 Y VPWR 0.029487f
C16 a_821_297# Y 0.011009f
C17 D1 C1 0.07096f
C18 VPB B1 0.143868f
C19 Y VGND 0.524494f
C20 a_821_297# VPWR 0.813452f
C21 VPB A1 0.130489f
C22 VPWR VGND 0.194421f
C23 C1 B1 0.059368f
C24 a_821_297# VGND 0.018397f
C25 VPB A2 0.16048f
C26 VPB Y 0.013112f
C27 VPB VPWR 0.18855f
C28 D1 Y 0.321096f
C29 B1 A1 0.051612f
C30 a_821_297# VPB 0.030819f
C31 C1 Y 0.166328f
C32 VPB VGND 0.016846f
C33 D1 VPWR 0.033781f
C34 a_821_297# D1 1.43e-20
C35 C1 VPWR 0.032397f
C36 B1 Y 0.168342f
C37 D1 VGND 0.06905f
C38 A1 A2 0.065368f
C39 VGND VNB 1.09023f
C40 VPWR VNB 0.909091f
C41 Y VNB 0.086884f
C42 A2 VNB 0.45321f
C43 A1 VNB 0.382402f
C44 B1 VNB 0.402276f
C45 C1 VNB 0.381363f
C46 D1 VNB 0.38265f
C47 VPB VNB 2.0223f
C48 a_821_297# VNB 0.02985f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_0 VNB VPB VPWR VGND X B A
X0 VPWR.t1 B.t0 a_40_47.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X.t0 a_40_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X2 VGND.t0 B.t1 a_123_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X.t1 a_40_47.t4 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X4 a_123_47.t0 A.t0 a_40_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 a_40_47.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
R0 B.n0 B.t1 224.304
R1 B.n0 B.t0 218.249
R2 B B.n0 71.0106
R3 a_40_47.n2 a_40_47.n1 682.193
R4 a_40_47.n0 a_40_47.t3 279.142
R5 a_40_47.n1 a_40_47.t1 250.526
R6 a_40_47.n0 a_40_47.t4 145.958
R7 a_40_47.n1 a_40_47.n0 118.642
R8 a_40_47.t0 a_40_47.n2 70.3576
R9 a_40_47.n2 a_40_47.t2 65.6672
R10 VPWR.n1 VPWR.t0 675.346
R11 VPWR.n1 VPWR.n0 218.893
R12 VPWR.n0 VPWR.t1 74.7554
R13 VPWR.n0 VPWR.t2 28.5349
R14 VPWR VPWR.n1 0.282531
R15 VPB.t1 VPB.t2 455.764
R16 VPB.t0 VPB.t1 260.437
R17 VPB VPB.t0 233.802
R18 X.n0 X.t0 356.337
R19 X.n0 X.t1 311.935
R20 X X.n0 1.89668
R21 a_123_47.t0 a_123_47.t1 60.0005
R22 VGND VGND.n0 191.358
R23 VGND.n0 VGND.t1 72.8576
R24 VGND.n0 VGND.t0 58.5719
R25 VNB.t1 VNB.t2 1737.22
R26 VNB VNB.t0 1124.92
R27 VNB.t0 VNB.t1 1025.24
R28 A.n0 A.t0 281.608
R29 A.n0 A.t1 161.374
R30 A A.n0 73.2226
C0 VPWR X 0.111278f
C1 B VGND 0.019565f
C2 VPWR VGND 0.045704f
C3 X VGND 0.105358f
C4 VPB A 0.093286f
C5 VPB B 0.088046f
C6 A B 0.117044f
C7 VPB VPWR 0.062434f
C8 VPB X 0.022086f
C9 A VPWR 0.047791f
C10 A X 1.67e-19
C11 VPB VGND 0.006814f
C12 B VPWR 0.044651f
C13 B X 0.007578f
C14 A VGND 0.017409f
C15 VGND VNB 0.300193f
C16 X VNB 0.10272f
C17 VPWR VNB 0.262881f
C18 B VNB 0.121465f
C19 A VNB 0.194569f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR.t2 B.t0 a_59_75.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X.t0 a_59_75.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND.t1 B.t1 a_145_75.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X.t1 a_59_75.t4 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75.t1 A.t1 a_59_75.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
R0 B.n0 B.t0 261.887
R1 B B.n0 156.864
R2 B.n0 B.t1 155.847
R3 a_59_75.n2 a_59_75.n1 672.948
R4 a_59_75.n1 a_59_75.t2 314.563
R5 a_59_75.n0 a_59_75.t3 236.18
R6 a_59_75.n0 a_59_75.t4 163.881
R7 a_59_75.n1 a_59_75.n0 152
R8 a_59_75.n2 a_59_75.t1 63.3219
R9 a_59_75.t0 a_59_75.n2 63.3219
R10 VPWR.n1 VPWR.t0 682.442
R11 VPWR.n1 VPWR.n0 331.682
R12 VPWR.n0 VPWR.t2 116.341
R13 VPWR.n0 VPWR.t1 28.4453
R14 VPWR VPWR.n1 0.401673
R15 VPB.t2 VPB.t1 319.627
R16 VPB VPB.t0 298.911
R17 VPB.t0 VPB.t2 248.599
R18 X.n0 X 590.984
R19 X.n1 X.n0 585
R20 X X.t1 269.426
R21 X.n0 X.t0 46.2955
R22 X X.n3 11.2645
R23 X X.n2 6.6565
R24 X.n3 X 6.1445
R25 X.n3 X 4.63498
R26 X.n2 X 3.61789
R27 X.n1 X 3.47876
R28 X.n2 X.n1 2.36572
R29 a_145_75.t0 a_145_75.t1 77.1434
R30 VGND VGND.n0 212.421
R31 VGND.n0 VGND.t1 72.8576
R32 VGND.n0 VGND.t0 22.3257
R33 VNB.t1 VNB.t0 1537.86
R34 VNB VNB.t2 1438.19
R35 VNB.t2 VNB.t1 1196.12
R36 A.n0 A.t0 256.07
R37 A.n1 A.n0 152
R38 A.n0 A.t1 150.03
R39 A A.n1 9.22489
R40 A.n1 A 7.6805
C0 VPB A 0.080573f
C1 VPWR A 0.036234f
C2 VPB B 0.06287f
C3 VPB X 0.012653f
C4 VPWR B 0.011747f
C5 VPB VGND 0.007995f
C6 VPWR X 0.111215f
C7 A B 0.097088f
C8 VPWR VGND 0.046078f
C9 A X 1.68e-19
C10 A VGND 0.014715f
C11 B X 0.002761f
C12 B VGND 0.011461f
C13 X VGND 0.099328f
C14 VPB VPWR 0.072934f
C15 VGND VNB 0.311398f
C16 X VNB 0.100184f
C17 B VNB 0.112872f
C18 A VNB 0.173792f
C19 VPWR VNB 0.273451f
C20 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR.t0 B.t0 a_207_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X.t0 a_207_413.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47.t1 a_27_413.t2 a_207_413.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X.t1 a_207_413.t4 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413.t2 a_27_413.t3 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR.t1 A_N.t0 a_27_413.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND.t0 B.t1 a_297_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413.t0 A_N.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 B.n0 B.t1 293.969
R1 B.n1 B.n0 152
R2 B.n0 B.t0 138.338
R3 B B.n1 14.0392
R4 B.n1 B 4.95534
R5 a_207_413.n2 a_207_413.n1 625.684
R6 a_207_413.n1 a_207_413.t1 262.252
R7 a_207_413.n0 a_207_413.t3 240.484
R8 a_207_413.n1 a_207_413.n0 174.924
R9 a_207_413.n0 a_207_413.t4 166.692
R10 a_207_413.t0 a_207_413.n2 68.0124
R11 a_207_413.n2 a_207_413.t2 68.0124
R12 VPWR.n9 VPWR.n1 602.456
R13 VPWR.n3 VPWR.n2 585
R14 VPWR.n5 VPWR.n4 585
R15 VPWR.n4 VPWR.n3 159.476
R16 VPWR.n1 VPWR.t3 96.1553
R17 VPWR.n3 VPWR.t0 86.7743
R18 VPWR.n4 VPWR.t2 66.8398
R19 VPWR.n1 VPWR.t1 63.3219
R20 VPWR.n8 VPWR.n7 27.724
R21 VPWR.n9 VPWR.n8 22.9652
R22 VPWR.n7 VPWR.n6 9.3005
R23 VPWR.n8 VPWR.n0 9.3005
R24 VPWR.n6 VPWR.n5 9.01185
R25 VPWR.n10 VPWR.n9 7.12063
R26 VPWR.n5 VPWR.n2 6.8005
R27 VPWR.n7 VPWR.n2 1.0005
R28 VPWR.n10 VPWR.n0 0.148519
R29 VPWR.n6 VPWR.n0 0.120292
R30 VPWR VPWR.n10 0.114842
R31 VPB.t0 VPB.t2 526.792
R32 VPB.t1 VPB.t3 290.031
R33 VPB.t3 VPB.t0 260.437
R34 VPB VPB.t1 192.369
R35 X.n1 X.t0 358.94
R36 X.n0 X.t1 209.923
R37 X X.n0 79.4838
R38 X.n1 X 7.91583
R39 X.n0 X 6.66717
R40 X X.n1 6.2537
R41 a_27_413.n1 a_27_413.t1 725.558
R42 a_27_413.n0 a_27_413.t3 381.656
R43 a_27_413.t0 a_27_413.n1 243.694
R44 a_27_413.n0 a_27_413.t2 197.62
R45 a_27_413.n1 a_27_413.n0 164.994
R46 a_297_47.t0 a_297_47.t1 68.5719
R47 VNB.t1 VNB.t2 2677.02
R48 VNB.t0 VNB.t3 1395.47
R49 VNB.t2 VNB.t0 1110.68
R50 VNB VNB.t1 925.567
R51 VGND.n1 VGND.t1 247.484
R52 VGND.n1 VGND.n0 206.194
R53 VGND.n0 VGND.t0 58.5719
R54 VGND.n0 VGND.t2 25.4291
R55 VGND VGND.n1 0.0759566
R56 A_N.n0 A_N.t0 327.99
R57 A_N.n0 A_N.t1 199.457
R58 A_N.n1 A_N.n0 152
R59 A_N.n1 A_N 12.1605
R60 A_N A_N.n1 2.34717
C0 VPB A_N 0.080056f
C1 VPB B 0.111061f
C2 VPB VPWR 0.063352f
C3 VPB X 0.012221f
C4 A_N VPWR 0.018219f
C5 B VPWR 0.086692f
C6 VPB VGND 0.007626f
C7 A_N VGND 0.047311f
C8 B X 0.030307f
C9 VPWR X 0.055194f
C10 B VGND 0.01869f
C11 VPWR VGND 0.056424f
C12 X VGND 0.065151f
C13 VGND VNB 0.368472f
C14 X VNB 0.089221f
C15 VPWR VNB 0.291542f
C16 B VNB 0.132317f
C17 A_N VNB 0.201458f
C18 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_4 VNB VPB VGND VPWR A X B
X0 VPWR.t1 B.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1 a_27_47.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 X.t3 a_27_47.t3 VGND.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3 VPWR.t5 a_27_47.t4 X.t7 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND.t0 B.t1 a_110_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 X.t6 a_27_47.t5 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47.t0 A.t1 a_27_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 VPWR.t3 a_27_47.t6 X.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND.t4 a_27_47.t7 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND.t3 a_27_47.t8 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 X.t4 a_27_47.t9 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X11 X.t0 a_27_47.t10 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 B.n0 B.t0 241.536
R1 B.n0 B.t1 169.237
R2 B B.n0 163.249
R3 a_27_47.n11 a_27_47.n10 365.779
R4 a_27_47.n6 a_27_47.t4 212.081
R5 a_27_47.n2 a_27_47.t6 212.081
R6 a_27_47.n1 a_27_47.t5 212.081
R7 a_27_47.n7 a_27_47.t9 212.081
R8 a_27_47.n10 a_27_47.t2 201.811
R9 a_27_47.n4 a_27_47.n3 164.992
R10 a_27_47.n9 a_27_47.n8 152
R11 a_27_47.n6 a_27_47.n0 152
R12 a_27_47.n5 a_27_47.n4 152
R13 a_27_47.n6 a_27_47.t8 139.78
R14 a_27_47.n2 a_27_47.t7 139.78
R15 a_27_47.n1 a_27_47.t10 139.78
R16 a_27_47.n7 a_27_47.t3 139.78
R17 a_27_47.n6 a_27_47.n5 49.6611
R18 a_27_47.n8 a_27_47.n6 49.6611
R19 a_27_47.n3 a_27_47.n1 36.5157
R20 a_27_47.n11 a_27_47.t1 27.5805
R21 a_27_47.t0 a_27_47.n11 27.5805
R22 a_27_47.n3 a_27_47.n2 26.2914
R23 a_27_47.n5 a_27_47.n1 13.146
R24 a_27_47.n8 a_27_47.n7 13.146
R25 a_27_47.n4 a_27_47.n0 12.9915
R26 a_27_47.n9 a_27_47.n0 12.9915
R27 a_27_47.n10 a_27_47.n9 9.36169
R28 VPWR.n5 VPWR.t3 343.55
R29 VPWR.n10 VPWR.t0 338.08
R30 VPWR.n8 VPWR.n2 309.726
R31 VPWR.n4 VPWR.n3 309.726
R32 VPWR.n2 VPWR.t2 35.4605
R33 VPWR.n2 VPWR.t1 34.4755
R34 VPWR.n3 VPWR.t4 27.5805
R35 VPWR.n3 VPWR.t5 27.5805
R36 VPWR.n9 VPWR.n8 22.5887
R37 VPWR.n8 VPWR.n7 21.8358
R38 VPWR.n7 VPWR.n4 21.0829
R39 VPWR.n10 VPWR.n9 19.9534
R40 VPWR.n7 VPWR.n6 9.3005
R41 VPWR.n8 VPWR.n1 9.3005
R42 VPWR.n9 VPWR.n0 9.3005
R43 VPWR.n11 VPWR.n10 9.3005
R44 VPWR.n5 VPWR.n4 6.50634
R45 VPWR.n6 VPWR.n5 0.731956
R46 VPWR.n6 VPWR.n1 0.120292
R47 VPWR.n1 VPWR.n0 0.120292
R48 VPWR.n11 VPWR.n0 0.120292
R49 VPWR VPWR.n11 0.0226354
R50 VPB.t1 VPB.t2 298.911
R51 VPB.t4 VPB.t3 254.518
R52 VPB.t5 VPB.t4 254.518
R53 VPB.t2 VPB.t5 254.518
R54 VPB.t0 VPB.t1 254.518
R55 VPB VPB.t0 195.327
R56 A.n0 A.t0 235.821
R57 A A.n0 163.768
R58 A.n0 A.t1 163.52
R59 VGND.n1 VGND.t4 289.418
R60 VGND.n3 VGND.n2 198.964
R61 VGND.n6 VGND.n5 198.964
R62 VGND.n5 VGND.t1 39.6928
R63 VGND.n5 VGND.t0 38.7697
R64 VGND.n2 VGND.t2 25.8467
R65 VGND.n2 VGND.t3 25.8467
R66 VGND.n6 VGND.n4 24.4711
R67 VGND.n4 VGND.n3 21.0829
R68 VGND.n4 VGND.n0 9.3005
R69 VGND.n7 VGND.n6 6.93132
R70 VGND.n3 VGND.n1 6.50634
R71 VGND.n1 VGND.n0 0.731956
R72 VGND VGND.n7 0.227479
R73 VGND.n7 VGND.n0 0.156225
R74 X.n2 X.n1 360.399
R75 X.n5 X.n4 232.862
R76 X.n2 X.n0 203.161
R77 X.n5 X.n3 95.6721
R78 X X.n2 61.049
R79 X.n0 X.t5 27.5805
R80 X.n0 X.t6 27.5805
R81 X.n1 X.t7 27.5805
R82 X.n1 X.t4 27.5805
R83 X.n4 X.t1 25.8467
R84 X.n4 X.t3 25.8467
R85 X.n3 X.t2 25.8467
R86 X.n3 X.t0 25.8467
R87 X X.n5 22.1918
R88 VNB.t1 VNB.t5 1637.54
R89 VNB.t2 VNB.t4 1224.6
R90 VNB.t3 VNB.t2 1224.6
R91 VNB.t5 VNB.t3 1224.6
R92 VNB.t0 VNB.t1 1025.24
R93 VNB VNB.t0 939.807
R94 a_110_47.t0 a_110_47.t1 38.7697
C0 VPWR VGND 0.066515f
C1 X VGND 0.189539f
C2 VPB A 0.036952f
C3 VPB B 0.027183f
C4 A B 0.092177f
C5 VPB VPWR 0.0747f
C6 VPB X 0.012188f
C7 A VPWR 0.047696f
C8 B VPWR 0.020623f
C9 VPB VGND 0.005697f
C10 A X 2e-19
C11 B X 0.001139f
C12 A VGND 0.014255f
C13 VPWR X 0.325545f
C14 B VGND 0.015936f
C15 VGND VNB 0.394237f
C16 X VNB 0.067157f
C17 VPWR VNB 0.359845f
C18 B VNB 0.091374f
C19 A VNB 0.145451f
C20 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X.t3 a_61_75.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR.t0 a_61_75.t4 X.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR.t2 B.t0 a_61_75.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND.t2 B.t1 a_147_75.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X.t1 a_61_75.t5 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND.t0 a_61_75.t6 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75.t2 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75.t0 A.t1 a_61_75.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
R0 a_61_75.n4 a_61_75.n0 672.948
R1 a_61_75.t0 a_61_75.n4 314.563
R2 a_61_75.n1 a_61_75.t4 212.081
R3 a_61_75.n2 a_61_75.t3 212.081
R4 a_61_75.n4 a_61_75.n3 152
R5 a_61_75.n1 a_61_75.t6 139.78
R6 a_61_75.n2 a_61_75.t5 139.78
R7 a_61_75.n3 a_61_75.n1 65.7278
R8 a_61_75.n0 a_61_75.t1 63.3219
R9 a_61_75.n0 a_61_75.t2 63.3219
R10 a_61_75.n3 a_61_75.n2 13.146
R11 VPWR.n7 VPWR.t3 675.293
R12 VPWR.n2 VPWR.n1 325.627
R13 VPWR.n3 VPWR.t0 273.173
R14 VPWR.n1 VPWR.t2 116.341
R15 VPWR.n6 VPWR.n5 34.6358
R16 VPWR.n1 VPWR.t1 28.4453
R17 VPWR.n8 VPWR.n7 13.4417
R18 VPWR.n3 VPWR.n2 9.85502
R19 VPWR.n7 VPWR.n6 9.41227
R20 VPWR.n5 VPWR.n4 9.3005
R21 VPWR.n6 VPWR.n0 9.3005
R22 VPWR.n5 VPWR.n2 7.15344
R23 VPWR.n4 VPWR.n3 0.516692
R24 VPWR.n4 VPWR.n0 0.120292
R25 VPWR.n8 VPWR.n0 0.120292
R26 VPWR VPWR.n8 0.0226354
R27 X.n0 X 591.116
R28 X.n1 X.n0 585
R29 X X.n3 191.841
R30 X.n3 X.t0 47.0774
R31 X.n0 X.t3 46.2955
R32 X.n0 X.t2 30.5355
R33 X.n3 X.t1 24.9236
R34 X X.n4 11.2645
R35 X X.n2 6.6565
R36 X.n4 X 6.1445
R37 X.n4 X 4.63498
R38 X.n2 X 3.69828
R39 X.n1 X 3.55606
R40 X.n2 X.n1 2.41828
R41 VPB.t1 VPB.t0 319.627
R42 VPB.t2 VPB.t1 319.627
R43 VPB VPB.t3 304.829
R44 VPB.t3 VPB.t2 248.599
R45 B.n0 B.t0 261.887
R46 B B.n0 157.376
R47 B.n0 B.t1 155.847
R48 a_147_75.t0 a_147_75.t1 77.1434
R49 VGND.n1 VGND.n0 211.972
R50 VGND.n1 VGND.t0 163.5
R51 VGND.n0 VGND.t2 72.8576
R52 VGND.n0 VGND.t1 22.3257
R53 VGND VGND.n1 0.494757
R54 VNB.t2 VNB.t1 1537.86
R55 VNB.t3 VNB.t2 1537.86
R56 VNB VNB.t0 1466.67
R57 VNB.t0 VNB.t3 1196.12
R58 A.n0 A.t0 256.07
R59 A.n1 A.n0 152
R60 A.n0 A.t1 150.03
R61 A A.n1 8.05893
R62 A.n1 A 7.1685
C0 VPB A 0.08239f
C1 VPWR A 0.040281f
C2 VPB B 0.064248f
C3 VPB X 0.005513f
C4 VPWR B 0.012524f
C5 VPWR X 0.194597f
C6 A B 0.096585f
C7 A X 1.84e-19
C8 B X 0.002798f
C9 VGND VPB 0.009503f
C10 VGND VPWR 0.07134f
C11 VGND A 0.015556f
C12 VGND B 0.011526f
C13 VPB VPWR 0.090199f
C14 VGND X 0.153129f
C15 VGND VNB 0.390327f
C16 X VNB 0.027496f
C17 B VNB 0.111386f
C18 A VNB 0.177011f
C19 VPWR VNB 0.349659f
C20 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_4 VNB VPB VGND VPWR X A_N B
X0 X.t7 a_27_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.1365 ps=1.07 w=0.65 l=0.15
X1 VGND.t0 B.t0 a_109_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.0715 ps=0.87 w=0.65 l=0.15
X2 VPWR.t0 B.t1 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_199.t1 A_N.t0 VGND.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.10675 ps=1.005 w=0.42 l=0.15
X4 a_33_199.t0 A_N.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.15575 ps=1.355 w=0.42 l=0.15
X5 VPWR.t6 a_27_47.t4 X.t0 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t3 a_27_47.t5 X.t6 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.091 ps=0.93 w=0.65 l=0.15
X7 X.t3 a_27_47.t6 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND.t2 a_27_47.t7 X.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR.t4 a_27_47.t8 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X10 X.t1 a_27_47.t9 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.185 ps=1.37 w=1 l=0.15
X11 a_27_47.t1 a_33_199.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X.t4 a_27_47.t10 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_109_47.t1 a_33_199.t3 a_27_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.0715 pd=0.87 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_47.n11 a_27_47.n10 623.237
R1 a_27_47.n2 a_27_47.t4 212.081
R2 a_27_47.n3 a_27_47.t6 212.081
R3 a_27_47.n6 a_27_47.t8 212.081
R4 a_27_47.n7 a_27_47.t9 212.081
R5 a_27_47.n10 a_27_47.t2 200.643
R6 a_27_47.n5 a_27_47.n0 164.089
R7 a_27_47.n9 a_27_47.n8 152
R8 a_27_47.n1 a_27_47.n0 152
R9 a_27_47.n2 a_27_47.t5 139.78
R10 a_27_47.n7 a_27_47.t3 139.78
R11 a_27_47.n1 a_27_47.t7 139.78
R12 a_27_47.n4 a_27_47.t10 139.78
R13 a_27_47.n3 a_27_47.n2 61.346
R14 a_27_47.n8 a_27_47.n1 49.6611
R15 a_27_47.n6 a_27_47.n5 46.0096
R16 a_27_47.t0 a_27_47.n11 26.5955
R17 a_27_47.n11 a_27_47.t1 26.5955
R18 a_27_47.n5 a_27_47.n4 13.8763
R19 a_27_47.n8 a_27_47.n7 12.4157
R20 a_27_47.n9 a_27_47.n0 12.0894
R21 a_27_47.n10 a_27_47.n9 8.71161
R22 a_27_47.n1 a_27_47.n6 3.65202
R23 a_27_47.n4 a_27_47.n3 1.46111
R24 VGND.n2 VGND.n1 249.274
R25 VGND.n4 VGND.n3 198.964
R26 VGND.n7 VGND.n6 198.964
R27 VGND.n1 VGND.t5 61.4291
R28 VGND.n6 VGND.t4 39.6928
R29 VGND.n6 VGND.t0 37.8467
R30 VGND.n3 VGND.t1 26.7697
R31 VGND.n3 VGND.t2 24.9236
R32 VGND.n7 VGND.n5 24.4711
R33 VGND.n5 VGND.n4 20.7064
R34 VGND.n1 VGND.t3 20.1775
R35 VGND.n5 VGND.n0 9.3005
R36 VGND.n8 VGND.n7 6.93132
R37 VGND.n4 VGND.n2 6.6033
R38 VGND.n2 VGND.n0 0.646617
R39 VGND VGND.n8 0.227479
R40 VGND.n8 VGND.n0 0.156225
R41 X.n2 X.n0 634.035
R42 X.n2 X.n1 585
R43 X.n5 X.n3 235.864
R44 X.n5 X.n4 185
R45 X X.n2 37.7384
R46 X.n0 X.t1 32.5055
R47 X.n3 X.t5 26.7697
R48 X.n1 X.t0 26.5955
R49 X.n1 X.t3 26.5955
R50 X.n0 X.t2 26.5955
R51 X.n4 X.t6 25.8467
R52 X.n4 X.t4 25.8467
R53 X.n3 X.t7 24.9236
R54 X X.n5 1.10395
R55 VNB.t0 VNB.t4 1623.3
R56 VNB.t3 VNB.t5 1438.19
R57 VNB.t1 VNB.t3 1224.6
R58 VNB.t2 VNB.t1 1224.6
R59 VNB.t4 VNB.t2 1224.6
R60 VNB.t6 VNB.t0 1053.72
R61 VNB VNB.t6 925.567
R62 B.n0 B.t1 241.536
R63 B.n0 B.t0 169.237
R64 B B.n0 162.862
R65 a_109_47.t0 a_109_47.t1 40.6159
R66 VPWR.n10 VPWR.t2 868.5
R67 VPWR.n5 VPWR.t6 868.087
R68 VPWR.n8 VPWR.n2 598.965
R69 VPWR.n4 VPWR.n3 598.965
R70 VPWR.t6 VPWR.t1 131.154
R71 VPWR.n2 VPWR.t0 37.4305
R72 VPWR.n2 VPWR.t3 35.4605
R73 VPWR.n3 VPWR.t5 26.5955
R74 VPWR.n3 VPWR.t4 26.5955
R75 VPWR.n9 VPWR.n8 22.5887
R76 VPWR.n7 VPWR.n4 22.2123
R77 VPWR.n8 VPWR.n7 21.8358
R78 VPWR.n10 VPWR.n9 19.9534
R79 VPWR.n7 VPWR.n6 9.3005
R80 VPWR.n8 VPWR.n1 9.3005
R81 VPWR.n9 VPWR.n0 9.3005
R82 VPWR.n11 VPWR.n10 9.3005
R83 VPWR.n5 VPWR.n4 6.49728
R84 VPWR.n6 VPWR.n5 0.667282
R85 VPWR.n6 VPWR.n1 0.120292
R86 VPWR.n1 VPWR.n0 0.120292
R87 VPWR.n11 VPWR.n0 0.120292
R88 VPWR VPWR.n11 0.0226354
R89 VPB.t0 VPB.t3 307.788
R90 VPB.t6 VPB.t1 298.911
R91 VPB.t3 VPB.t4 266.356
R92 VPB.t5 VPB.t6 248.599
R93 VPB.t4 VPB.t5 248.599
R94 VPB.t2 VPB.t0 248.599
R95 VPB VPB.t2 192.369
R96 A_N A_N.n0 154.309
R97 A_N.n0 A_N.t1 143.484
R98 A_N.n0 A_N.t0 129.786
R99 a_33_199.t0 a_33_199.n1 650.668
R100 a_33_199.n1 a_33_199.n0 459.723
R101 a_33_199.n1 a_33_199.t1 295.029
R102 a_33_199.n0 a_33_199.t2 233.01
R103 a_33_199.n0 a_33_199.t3 160.709
C0 VPB B 0.027197f
C1 VPB VPWR 0.08574f
C2 B VPWR 0.016609f
C3 VPB X 0.004239f
C4 B X 4.22e-19
C5 VPB A_N 0.039929f
C6 VPWR X 0.031345f
C7 VPB VGND 0.008054f
C8 B VGND 0.015666f
C9 VPWR A_N 0.011852f
C10 X A_N 0.092307f
C11 VPWR VGND 0.075024f
C12 X VGND 0.107425f
C13 A_N VGND 0.040299f
C14 VGND VNB 0.445737f
C15 A_N VNB 0.124324f
C16 X VNB 0.007246f
C17 VPWR VNB 0.37796f
C18 B VNB 0.091477f
C19 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_2 VNB VPB VPWR VGND A_N X B
X0 VPWR.t1 a_212_413.t3 X.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47.t1 a_27_413.t2 a_212_413.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X.t2 a_212_413.t4 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X.t1 a_212_413.t5 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413.t1 a_27_413.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR.t4 A_N.t0 a_27_413.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR.t3 B.t0 a_212_413.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND.t2 B.t1 a_297_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND.t0 a_212_413.t6 X.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413.t0 A_N.t1 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_212_413.n3 a_212_413.n2 625.684
R1 a_212_413.t0 a_212_413.n3 263.892
R2 a_212_413.n0 a_212_413.t3 212.081
R3 a_212_413.n1 a_212_413.t4 212.081
R4 a_212_413.n3 a_212_413.n1 185.017
R5 a_212_413.n0 a_212_413.t6 136.567
R6 a_212_413.n1 a_212_413.t5 136.567
R7 a_212_413.n2 a_212_413.t2 68.0124
R8 a_212_413.n2 a_212_413.t1 68.0124
R9 a_212_413.n1 a_212_413.n0 59.5417
R10 X X.n0 588.149
R11 X.n3 X.n0 585
R12 X.n2 X.n1 185
R13 X.n3 X.n2 81.8375
R14 X.n0 X.t3 26.5955
R15 X.n0 X.t2 26.5955
R16 X.n1 X.t0 24.9236
R17 X.n1 X.t1 24.9236
R18 X.n2 X 2.17922
R19 X X.n3 1.46935
R20 VPWR.n10 VPWR.n1 602.456
R21 VPWR.n3 VPWR.n2 585
R22 VPWR.n5 VPWR.n4 585
R23 VPWR.n6 VPWR.t1 354.702
R24 VPWR.n4 VPWR.n3 159.476
R25 VPWR.n1 VPWR.t2 107.882
R26 VPWR.n3 VPWR.t3 86.7743
R27 VPWR.n4 VPWR.t0 69.185
R28 VPWR.n1 VPWR.t4 63.3219
R29 VPWR.n9 VPWR.n8 29.1064
R30 VPWR.n10 VPWR.n9 22.9652
R31 VPWR.n8 VPWR.n7 9.3005
R32 VPWR.n9 VPWR.n0 9.3005
R33 VPWR.n6 VPWR.n5 7.81435
R34 VPWR.n11 VPWR.n10 7.12063
R35 VPWR.n5 VPWR.n2 6.8005
R36 VPWR.n8 VPWR.n2 1.5005
R37 VPWR.n7 VPWR.n6 0.562802
R38 VPWR.n11 VPWR.n0 0.148519
R39 VPWR.n7 VPWR.n0 0.120292
R40 VPWR VPWR.n11 0.11354
R41 VPB.t3 VPB.t0 529.751
R42 VPB.t4 VPB.t2 304.829
R43 VPB.t2 VPB.t3 260.437
R44 VPB.t0 VPB.t1 248.599
R45 VPB VPB.t4 189.409
R46 a_27_413.n1 a_27_413.t1 725.837
R47 a_27_413.n0 a_27_413.t3 381.656
R48 a_27_413.t0 a_27_413.n1 244.09
R49 a_27_413.n0 a_27_413.t2 189.588
R50 a_27_413.n1 a_27_413.n0 165.77
R51 a_297_47.t0 a_297_47.t1 77.1434
R52 VNB.t4 VNB.t3 2677.02
R53 VNB.t2 VNB.t1 1395.47
R54 VNB.t1 VNB.t0 1196.12
R55 VNB.t3 VNB.t2 1196.12
R56 VNB VNB.t4 911.327
R57 VGND.n4 VGND.t0 242.849
R58 VGND.n9 VGND.t3 240.833
R59 VGND.n3 VGND.n2 200.041
R60 VGND.n2 VGND.t2 58.5719
R61 VGND.n7 VGND.n1 34.6358
R62 VGND.n8 VGND.n7 34.6358
R63 VGND.n2 VGND.t1 24.9236
R64 VGND.n3 VGND.n1 19.9534
R65 VGND.n9 VGND.n8 19.9534
R66 VGND.n10 VGND.n9 9.3005
R67 VGND.n8 VGND.n0 9.3005
R68 VGND.n7 VGND.n6 9.3005
R69 VGND.n5 VGND.n1 9.3005
R70 VGND.n4 VGND.n3 6.34853
R71 VGND.n5 VGND.n4 0.667593
R72 VGND.n6 VGND.n5 0.120292
R73 VGND.n6 VGND.n0 0.120292
R74 VGND.n10 VGND.n0 0.120292
R75 VGND VGND.n10 0.0213333
R76 A_N.n0 A_N.t0 328.32
R77 A_N.n0 A_N.t1 199.786
R78 A_N.n1 A_N.n0 152
R79 A_N.n1 A_N 13.2272
R80 A_N A_N.n1 1.2805
R81 B.n0 B.t1 293.654
R82 B.n1 B.n0 152
R83 B.n0 B.t0 138.338
R84 B.n1 B 17.5489
R85 B B.n1 4.95534
C0 VPB X 0.007805f
C1 A_N VPWR 0.018071f
C2 VPB VGND 0.009127f
C3 B VPWR 0.08705f
C4 B X 0.030309f
C5 A_N VGND 0.046884f
C6 B VGND 0.018833f
C7 VPWR X 0.112472f
C8 VPWR VGND 0.077171f
C9 X VGND 0.103266f
C10 VPB A_N 0.080843f
C11 VPB B 0.113326f
C12 VPB VPWR 0.078365f
C13 VGND VNB 0.436984f
C14 X VNB 0.036558f
C15 VPWR VNB 0.357551f
C16 B VNB 0.132642f
C17 A_N VNB 0.201516f
C18 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_4 VNB VPB VGND VPWR X A B C
X0 VPWR.t0 A.t0 a_94_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.395 as=0.305 ps=2.61 w=1 l=0.15
X1 a_294_47.t0 B.t0 a_185_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.128375 ps=1.045 w=0.65 l=0.15
X2 a_185_47.t0 A.t1 a_94_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.045 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VPWR.t4 a_94_47.t4 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND.t4 C.t0 a_294_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_94_47.t2 B.t1 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1975 ps=1.395 w=1 l=0.15
X6 X.t2 a_94_47.t5 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X7 X.t7 a_94_47.t6 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR.t6 C.t1 a_94_47.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X9 X.t6 a_94_47.t7 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X10 VGND.t1 a_94_47.t8 X.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VPWR.t2 a_94_47.t9 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND.t0 a_94_47.t10 X.t4 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X.t0 a_94_47.t11 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A.n0 A.t0 241.536
R1 A.n0 A.t1 169.237
R2 A A.n0 158.864
R3 a_94_47.t0 a_94_47.n12 406.841
R4 a_94_47.n12 a_94_47.n11 319.401
R5 a_94_47.n10 a_94_47.t1 237.012
R6 a_94_47.n6 a_94_47.t9 212.081
R7 a_94_47.n2 a_94_47.t4 212.081
R8 a_94_47.n1 a_94_47.t11 212.081
R9 a_94_47.n7 a_94_47.t5 212.081
R10 a_94_47.n4 a_94_47.n3 164.992
R11 a_94_47.n9 a_94_47.n8 152
R12 a_94_47.n6 a_94_47.n0 152
R13 a_94_47.n5 a_94_47.n4 152
R14 a_94_47.n6 a_94_47.t10 139.78
R15 a_94_47.n2 a_94_47.t8 139.78
R16 a_94_47.n1 a_94_47.t6 139.78
R17 a_94_47.n7 a_94_47.t7 139.78
R18 a_94_47.n6 a_94_47.n5 49.6611
R19 a_94_47.n8 a_94_47.n6 49.6611
R20 a_94_47.n12 a_94_47.n10 46.7546
R21 a_94_47.n3 a_94_47.n1 36.5157
R22 a_94_47.n11 a_94_47.t3 27.5805
R23 a_94_47.n11 a_94_47.t2 27.5805
R24 a_94_47.n3 a_94_47.n2 26.2914
R25 a_94_47.n5 a_94_47.n1 13.146
R26 a_94_47.n8 a_94_47.n7 13.146
R27 a_94_47.n4 a_94_47.n0 12.9915
R28 a_94_47.n9 a_94_47.n0 12.9915
R29 a_94_47.n10 a_94_47.n9 9.36169
R30 VPWR.n6 VPWR.t4 343.55
R31 VPWR.n9 VPWR.n3 309.726
R32 VPWR.n5 VPWR.n4 309.726
R33 VPWR.n1 VPWR.n0 305.139
R34 VPWR.n0 VPWR.t0 40.3855
R35 VPWR.n0 VPWR.t5 37.4305
R36 VPWR.n3 VPWR.t3 35.4605
R37 VPWR.n3 VPWR.t6 34.4755
R38 VPWR.n4 VPWR.t1 27.5805
R39 VPWR.n4 VPWR.t2 27.5805
R40 VPWR.n10 VPWR.n9 22.5887
R41 VPWR.n9 VPWR.n8 21.8358
R42 VPWR.n8 VPWR.n5 21.0829
R43 VPWR.n10 VPWR.n1 19.9534
R44 VPWR.n8 VPWR.n7 9.3005
R45 VPWR.n9 VPWR.n2 9.3005
R46 VPWR.n11 VPWR.n10 9.3005
R47 VPWR.n12 VPWR.n1 6.60228
R48 VPWR.n6 VPWR.n5 6.50634
R49 VPWR.n7 VPWR.n6 0.731956
R50 VPWR VPWR.n12 0.222484
R51 VPWR.n12 VPWR.n11 0.161145
R52 VPWR.n7 VPWR.n2 0.120292
R53 VPWR.n11 VPWR.n2 0.120292
R54 VPB VPB.t0 417.291
R55 VPB.t0 VPB.t5 322.587
R56 VPB.t6 VPB.t3 298.911
R57 VPB.t1 VPB.t4 254.518
R58 VPB.t2 VPB.t1 254.518
R59 VPB.t3 VPB.t2 254.518
R60 VPB.t5 VPB.t6 254.518
R61 B.n0 B.t1 235.821
R62 B.n0 B.t0 163.52
R63 B B.n0 156.411
R64 a_185_47.t0 a_185_47.t1 72.9236
R65 a_294_47.t0 a_294_47.t1 38.7697
R66 VNB VNB.t0 2007.77
R67 VNB.t6 VNB.t3 1637.54
R68 VNB.t0 VNB.t5 1552.1
R69 VNB.t4 VNB.t2 1224.6
R70 VNB.t1 VNB.t4 1224.6
R71 VNB.t3 VNB.t1 1224.6
R72 VNB.t5 VNB.t6 1025.24
R73 X.n2 X.n1 360.399
R74 X.n5 X.n4 232.862
R75 X.n2 X.n0 203.161
R76 X.n5 X.n3 95.6721
R77 X X.n2 61.049
R78 X.n0 X.t3 27.5805
R79 X.n0 X.t0 27.5805
R80 X.n1 X.t1 27.5805
R81 X.n1 X.t2 27.5805
R82 X.n4 X.t4 25.8467
R83 X.n4 X.t6 25.8467
R84 X.n3 X.t5 25.8467
R85 X.n3 X.t7 25.8467
R86 X X.n5 22.1918
R87 C.n0 C.t1 241.536
R88 C.n0 C.t0 169.237
R89 C C.n0 163.249
R90 VGND.n1 VGND.t1 289.418
R91 VGND.n3 VGND.n2 198.964
R92 VGND.n6 VGND.n5 198.964
R93 VGND.n5 VGND.t4 44.3082
R94 VGND.n5 VGND.t2 34.1543
R95 VGND.n2 VGND.t3 25.8467
R96 VGND.n2 VGND.t0 25.8467
R97 VGND.n6 VGND.n4 22.2123
R98 VGND.n4 VGND.n3 21.0829
R99 VGND.n4 VGND.n0 9.3005
R100 VGND.n7 VGND.n6 7.06324
R101 VGND.n3 VGND.n1 6.50634
R102 VGND.n1 VGND.n0 0.731956
R103 VGND VGND.n7 0.468986
R104 VGND.n7 VGND.n0 0.155496
C0 VPB C 0.027183f
C1 A B 0.078035f
C2 VPB VPWR 0.091049f
C3 A C 2.62e-19
C4 B C 0.092051f
C5 VPB X 0.012188f
C6 A VPWR 0.049627f
C7 B VPWR 0.022189f
C8 VPB VGND 0.008064f
C9 A VGND 0.024177f
C10 C VPWR 0.020554f
C11 B VGND 0.014333f
C12 C X 0.001026f
C13 C VGND 0.01501f
C14 VPWR X 0.325545f
C15 VPWR VGND 0.08352f
C16 X VGND 0.189572f
C17 VPB A 0.057814f
C18 VPB B 0.030937f
C19 VGND VNB 0.491132f
C20 X VNB 0.067157f
C21 VPWR VNB 0.415096f
C22 C VNB 0.091374f
C23 B VNB 0.103104f
C24 A VNB 0.175032f
C25 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR.t2 a_29_311.t4 X.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t0 a_29_311.t5 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR.t0 A.t0 a_29_311.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND.t1 a_29_311.t6 X.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53.t1 B.t0 a_112_53.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR.t4 C.t0 a_29_311.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X.t2 a_29_311.t7 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53.t0 A.t1 a_29_311.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311.t2 B.t1 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND.t2 C.t1 a_184_53.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
R0 a_29_311.t0 a_29_311.n4 682.33
R1 a_29_311.n3 a_29_311.n2 585
R2 a_29_311.n4 a_29_311.t1 294.425
R3 a_29_311.n1 a_29_311.t4 214.272
R4 a_29_311.n0 a_29_311.t5 212.081
R5 a_29_311.n3 a_29_311.n0 208.171
R6 a_29_311.n0 a_29_311.t7 139.78
R7 a_29_311.n1 a_29_311.t6 139.78
R8 a_29_311.n2 a_29_311.t2 79.5457
R9 a_29_311.n0 a_29_311.n1 61.346
R10 a_29_311.n2 a_29_311.t3 48.5886
R11 a_29_311.n4 a_29_311.n3 16.2697
R12 X.n0 X 593.145
R13 X.n1 X.n0 585
R14 X.n3 X.n2 185
R15 X X.n1 41.1099
R16 X X.n3 29.0306
R17 X.n0 X.t1 26.5955
R18 X.n0 X.t0 26.5955
R19 X.n2 X.t3 24.9236
R20 X.n2 X.t2 24.9236
R21 X.n1 X 7.6805
R22 X.n3 X 5.3765
R23 VPWR.n8 VPWR.n1 600.862
R24 VPWR.n4 VPWR.t2 350.853
R25 VPWR.n3 VPWR.n2 322.551
R26 VPWR.n2 VPWR.t4 98.5005
R27 VPWR.n1 VPWR.t3 63.3219
R28 VPWR.n1 VPWR.t0 63.3219
R29 VPWR.n7 VPWR.n6 33.2275
R30 VPWR.n6 VPWR.n3 30.4946
R31 VPWR.n2 VPWR.t1 26.5955
R32 VPWR VPWR.n8 16.6961
R33 VPWR.n6 VPWR.n5 9.3005
R34 VPWR.n7 VPWR.n0 9.3005
R35 VPWR.n4 VPWR.n3 6.61302
R36 VPWR.n8 VPWR.n7 1.32791
R37 VPWR.n5 VPWR.n4 0.612146
R38 VPWR.n5 VPWR.n0 0.120292
R39 VPWR VPWR.n0 0.120292
R40 VPB.t4 VPB.t1 292.991
R41 VPB.t3 VPB.t4 281.154
R42 VPB.t1 VPB.t2 248.599
R43 VPB.t0 VPB.t3 248.599
R44 VPB VPB.t0 198.287
R45 A.n0 A.t1 186.03
R46 A A.n0 165.132
R47 A.n0 A.t0 160.322
R48 VGND.n1 VGND.t1 240.847
R49 VGND.n1 VGND.n0 210.72
R50 VGND.n0 VGND.t2 88.5937
R51 VGND.n0 VGND.t0 21.907
R52 VGND VGND.n1 0.778402
R53 VNB.t4 VNB.t1 1722.98
R54 VNB.t1 VNB.t2 1196.12
R55 VNB.t0 VNB.t4 1153.4
R56 VNB.t3 VNB.t0 1025.24
R57 VNB VNB.t3 968.285
R58 B.t1 B.t0 398.281
R59 B B.t1 303.034
R60 a_112_53.t0 a_112_53.t1 60.0005
R61 a_184_53.t0 a_184_53.t1 72.8576
R62 C.n0 C.t1 195
R63 C C.n0 164.333
R64 C.n0 C.t0 146.799
C0 X VGND 0.140172f
C1 VPB B 0.092345f
C2 VPB VPWR 0.092909f
C3 VPB A 0.044263f
C4 B VPWR 0.130127f
C5 VPB C 0.035171f
C6 B A 0.083535f
C7 VPB X 0.00641f
C8 B C 0.064888f
C9 VPWR A 0.015648f
C10 B X 8.26e-19
C11 VPWR C 0.008825f
C12 VPB VGND 0.006612f
C13 VPWR X 0.192602f
C14 B VGND 0.007561f
C15 VPWR VGND 0.059136f
C16 A VGND 0.012714f
C17 C X 0.01584f
C18 C VGND 0.071418f
C19 VGND VNB 0.368566f
C20 X VNB 0.039992f
C21 C VNB 0.116494f
C22 A VNB 0.169936f
C23 VPWR VNB 0.335977f
C24 B VNB 0.103283f
C25 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR.t1 A.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR.t3 C.t0 a_27_47.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47.t1 B.t0 a_109_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND.t0 C.t1 a_181_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47.t0 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X.t1 a_27_47.t4 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6 X.t0 a_27_47.t5 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47.t0 A.t1 a_27_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A.n0 A.t0 183.505
R1 A A.n0 155.84
R2 A.n0 A.t1 114.532
R3 a_27_47.n1 a_27_47.t1 699.323
R4 a_27_47.n3 a_27_47.n2 585
R5 a_27_47.n2 a_27_47.n1 374.396
R6 a_27_47.n1 a_27_47.t2 335.384
R7 a_27_47.n0 a_27_47.t4 241.536
R8 a_27_47.n2 a_27_47.n0 182.721
R9 a_27_47.n0 a_27_47.t5 169.237
R10 a_27_47.t0 a_27_47.n3 84.4291
R11 a_27_47.n3 a_27_47.t3 63.3219
R12 VPWR.n2 VPWR.n0 723.785
R13 VPWR.n2 VPWR.n1 615.173
R14 VPWR.n0 VPWR.t3 93.81
R15 VPWR.n1 VPWR.t0 63.3219
R16 VPWR.n1 VPWR.t1 63.3219
R17 VPWR.n0 VPWR.t2 26.9729
R18 VPWR VPWR.n2 0.253242
R19 VPB.t3 VPB.t2 281.154
R20 VPB.t0 VPB.t3 275.235
R21 VPB.t1 VPB.t0 248.599
R22 VPB VPB.t1 192.369
R23 C.n0 C.t1 173.34
R24 C.n1 C.n0 165.189
R25 C.n0 C.t0 162.81
R26 C.n1 C 2.11184
R27 C C.n1 0.970197
R28 B.t1 B.t0 395.01
R29 B B.t1 320.95
R30 a_109_47.t0 a_109_47.t1 60.0005
R31 a_181_47.t0 a_181_47.t1 60.0005
R32 VNB.t1 VNB.t3 1822.65
R33 VNB.t2 VNB.t1 1025.24
R34 VNB.t0 VNB.t2 1025.24
R35 VNB VNB.t0 925.567
R36 VGND VGND.n0 214.873
R37 VGND.n0 VGND.t0 101.43
R38 VGND.n0 VGND.t1 25.9346
R39 X.n0 X 591.75
R40 X.n1 X.n0 585
R41 X.n2 X.t0 209.923
R42 X.n2 X.n1 96.3104
R43 X.n0 X.t1 26.5955
R44 X.n1 X 9.07686
R45 X X.n2 4.18512
C0 VPWR A 0.018456f
C1 VPB X 0.012079f
C2 B C 0.074622f
C3 VPB VGND 0.006035f
C4 B X 0.001105f
C5 VPWR C 0.004639f
C6 VPWR X 0.076623f
C7 B VGND 0.007138f
C8 VPWR VGND 0.047507f
C9 A VGND 0.015376f
C10 C X 0.01492f
C11 C VGND 0.07031f
C12 X VGND 0.070777f
C13 VPB B 0.083634f
C14 VPB VPWR 0.079461f
C15 VPB A 0.042605f
C16 B VPWR 0.128453f
C17 VPB C 0.034705f
C18 B A 0.086925f
C19 VGND VNB 0.300125f
C20 X VNB 0.092275f
C21 C VNB 0.120257f
C22 A VNB 0.174122f
C23 VPWR VNB 0.274246f
C24 B VNB 0.101788f
C25 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR VNB VPB X C B A_N
X0 a_109_53.t1 A_N.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X.t3 a_215_311.t4 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X2 a_109_53.t0 A_N.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND.t0 C.t0 a_373_53.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X4 VGND.t2 a_215_311.t5 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t0 C.t1 a_215_311.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 VPWR.t4 a_215_311.t6 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t0 a_215_311.t7 VPWR.t5 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X8 a_301_53.t1 a_109_53.t2 a_215_311.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_215_311.t1 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53.t1 B.t1 a_301_53.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR.t3 a_109_53.t3 a_215_311.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 A_N A_N.n0 183.971
R1 A_N.n0 A_N.t1 167.094
R2 A_N.n0 A_N.t0 141.387
R3 VPWR.n13 VPWR.t2 688.144
R4 VPWR.n2 VPWR.n1 600.862
R5 VPWR.n4 VPWR.t4 350.38
R6 VPWR.n6 VPWR.n5 324.25
R7 VPWR.n5 VPWR.t0 96.1553
R8 VPWR.n1 VPWR.t1 63.3219
R9 VPWR.n1 VPWR.t3 63.3219
R10 VPWR.n8 VPWR.n7 32.6642
R11 VPWR.n7 VPWR.n6 29.3652
R12 VPWR.n12 VPWR.n11 27.8761
R13 VPWR.n5 VPWR.t5 25.6105
R14 VPWR.n13 VPWR.n12 21.8358
R15 VPWR.n7 VPWR.n3 9.3005
R16 VPWR.n9 VPWR.n8 9.3005
R17 VPWR.n11 VPWR.n10 9.3005
R18 VPWR.n12 VPWR.n0 9.3005
R19 VPWR.n14 VPWR.n13 9.3005
R20 VPWR.n11 VPWR.n2 7.58569
R21 VPWR.n6 VPWR.n4 6.68308
R22 VPWR.n8 VPWR.n2 1.13828
R23 VPWR.n4 VPWR.n3 0.602464
R24 VPWR.n9 VPWR.n3 0.120292
R25 VPWR.n10 VPWR.n9 0.120292
R26 VPWR.n10 VPWR.n0 0.120292
R27 VPWR.n14 VPWR.n0 0.120292
R28 VPWR VPWR.n14 0.0226354
R29 a_109_53.n1 a_109_53.t1 676.715
R30 a_109_53.t0 a_109_53.n1 260.007
R31 a_109_53.n0 a_109_53.t2 186.03
R32 a_109_53.n1 a_109_53.n0 172.314
R33 a_109_53.n0 a_109_53.t3 160.322
R34 VPB.t2 VPB.t5 556.386
R35 VPB.t0 VPB.t4 287.072
R36 VPB.t1 VPB.t0 281.154
R37 VPB.t4 VPB.t3 248.599
R38 VPB.t5 VPB.t1 248.599
R39 VPB VPB.t2 192.369
R40 a_215_311.n0 a_215_311.t2 684.528
R41 a_215_311.n4 a_215_311.n3 599.485
R42 a_215_311.n0 a_215_311.t3 294.425
R43 a_215_311.n1 a_215_311.t6 212.081
R44 a_215_311.n2 a_215_311.t7 212.081
R45 a_215_311.n3 a_215_311.n2 208.876
R46 a_215_311.n1 a_215_311.t5 139.78
R47 a_215_311.n2 a_215_311.t4 139.78
R48 a_215_311.n4 a_215_311.t1 79.5457
R49 a_215_311.n2 a_215_311.n1 61.346
R50 a_215_311.n5 a_215_311.t0 42.96
R51 a_215_311.n6 a_215_311.n5 27.5805
R52 a_215_311.n3 a_215_311.n0 12.8005
R53 a_215_311.n5 a_215_311.n4 5.62907
R54 VGND.n11 VGND.t1 243.008
R55 VGND.n2 VGND.t2 241.667
R56 VGND.n4 VGND.n3 204.905
R57 VGND.n3 VGND.t0 86.3738
R58 VGND.n5 VGND.n1 34.6358
R59 VGND.n9 VGND.n1 34.6358
R60 VGND.n10 VGND.n9 34.6358
R61 VGND.n5 VGND.n4 25.6005
R62 VGND.n11 VGND.n10 25.224
R63 VGND.n3 VGND.t3 22.1912
R64 VGND.n12 VGND.n11 9.3005
R65 VGND.n10 VGND.n0 9.3005
R66 VGND.n9 VGND.n8 9.3005
R67 VGND.n7 VGND.n1 9.3005
R68 VGND.n6 VGND.n5 9.3005
R69 VGND.n4 VGND.n2 6.32311
R70 VGND.n6 VGND.n2 0.668695
R71 VGND.n7 VGND.n6 0.120292
R72 VGND.n8 VGND.n7 0.120292
R73 VGND.n8 VGND.n0 0.120292
R74 VGND.n12 VGND.n0 0.120292
R75 VGND VGND.n12 0.0226354
R76 X.n0 X 592.861
R77 X.n1 X.n0 585
R78 X.n3 X.n2 185
R79 X X.n1 40.9574
R80 X X.n3 29.2858
R81 X.n0 X.t1 26.5955
R82 X.n0 X.t0 26.5955
R83 X.n2 X.t2 24.9236
R84 X.n2 X.t3 24.9236
R85 X.n1 X 7.41103
R86 X.n3 X 5.48621
R87 VNB.t2 VNB.t5 2733.98
R88 VNB.t0 VNB.t4 1694.5
R89 VNB.t4 VNB.t3 1196.12
R90 VNB.t1 VNB.t0 1153.4
R91 VNB.t5 VNB.t1 1025.24
R92 VNB VNB.t2 925.567
R93 C.n0 C.t0 196.549
R94 C C.n0 164.333
R95 C.n0 C.t1 148.35
R96 a_373_53.t0 a_373_53.t1 72.8576
R97 a_301_53.t0 a_301_53.t1 60.0005
R98 B.t0 B.t1 402.005
R99 B B.t0 304.014
C0 VPB VPWR 0.1443f
C1 VPB A_N 0.053476f
C2 B VPWR 0.131796f
C3 VPB C 0.034649f
C4 VPWR A_N 0.036229f
C5 VPB X 0.006463f
C6 B C 0.068381f
C7 VPB VGND 0.011125f
C8 B X 8.71e-19
C9 VPWR C 0.009326f
C10 VPWR X 0.19334f
C11 B VGND 0.00805f
C12 VPWR VGND 0.080155f
C13 C X 0.016079f
C14 A_N VGND 0.043992f
C15 C VGND 0.070559f
C16 X VGND 0.138545f
C17 VPB B 0.092595f
C18 VGND VNB 0.484979f
C19 X VNB 0.040093f
C20 C VNB 0.113927f
C21 A_N VNB 0.187667f
C22 VPWR VNB 0.427551f
C23 B VNB 0.099764f
C24 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93.t1 A_N.t0 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X.t0 a_209_311.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93.t0 A_N.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53.t1 a_109_93.t2 a_209_311.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR.t4 C.t0 a_209_311.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53.t1 B.t0 a_296_53.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X.t1 a_209_311.t5 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311.t0 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR.t3 a_109_93.t3 a_209_311.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND.t2 C.t1 a_368_53.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
R0 A_N.n1 A_N.t1 204.656
R1 A_N.n3 A_N.n2 152
R2 A_N.n1 A_N.n0 152
R3 A_N.n2 A_N.t0 121.109
R4 A_N.n2 A_N.n1 40.9982
R5 A_N A_N.n3 10.7299
R6 A_N.n0 A_N 9.6005
R7 A_N A_N.n0 3.2005
R8 A_N.n3 A_N 2.07109
R9 VGND.n1 VGND.t1 266.767
R10 VGND.n1 VGND.n0 209.524
R11 VGND.n0 VGND.t2 83.899
R12 VGND.n0 VGND.t0 21.795
R13 VGND VGND.n1 0.0556855
R14 a_109_93.t0 a_109_93.n1 712.356
R15 a_109_93.n1 a_109_93.t1 235.934
R16 a_109_93.n0 a_109_93.t2 186.03
R17 a_109_93.n1 a_109_93.n0 176.321
R18 a_109_93.n0 a_109_93.t3 160.322
R19 VNB.t2 VNB.t3 2662.78
R20 VNB.t4 VNB.t0 1651.78
R21 VNB.t1 VNB.t4 1153.4
R22 VNB.t3 VNB.t1 1025.24
R23 VNB VNB.t2 911.327
R24 a_209_311.n1 a_209_311.t1 669.354
R25 a_209_311.n3 a_209_311.n2 585
R26 a_209_311.n1 a_209_311.t2 302.736
R27 a_209_311.n0 a_209_311.t4 241.536
R28 a_209_311.n2 a_209_311.n0 187.637
R29 a_209_311.n0 a_209_311.t5 169.237
R30 a_209_311.n3 a_209_311.t3 51.4029
R31 a_209_311.n4 a_209_311.t0 42.96
R32 a_209_311.n4 a_209_311.n3 33.7719
R33 a_209_311.n5 a_209_311.n4 27.5805
R34 a_209_311.n2 a_209_311.n1 14.3873
R35 VPWR.n4 VPWR.n3 727.241
R36 VPWR.n8 VPWR.t2 669.491
R37 VPWR.n2 VPWR.n1 603.38
R38 VPWR.n3 VPWR.t4 93.81
R39 VPWR.n1 VPWR.t0 63.3219
R40 VPWR.n1 VPWR.t3 63.3219
R41 VPWR.n3 VPWR.t1 28.5169
R42 VPWR.n7 VPWR.n6 26.4678
R43 VPWR.n8 VPWR.n7 25.977
R44 VPWR.n6 VPWR.n5 9.3005
R45 VPWR.n7 VPWR.n0 9.3005
R46 VPWR.n9 VPWR.n8 9.3005
R47 VPWR.n4 VPWR.n2 8.99725
R48 VPWR.n6 VPWR.n2 7.0168
R49 VPWR.n5 VPWR.n4 0.429926
R50 VPWR.n5 VPWR.n0 0.120292
R51 VPWR.n9 VPWR.n0 0.120292
R52 VPWR VPWR.n9 0.0213333
R53 X.n0 X 591.75
R54 X.n1 X.n0 585
R55 X.n2 X.t1 209.923
R56 X.n2 X.n1 96.3104
R57 X.n0 X.t0 26.5955
R58 X.n1 X 9.07686
R59 X X.n2 4.18512
R60 VPB.t2 VPB.t3 538.63
R61 VPB.t4 VPB.t1 281.154
R62 VPB.t0 VPB.t4 281.154
R63 VPB.t3 VPB.t0 248.599
R64 VPB VPB.t2 189.409
R65 a_296_53.t0 a_296_53.t1 60.0005
R66 C.n0 C.t1 196.549
R67 C C.n0 164.333
R68 C.n0 C.t0 148.35
R69 B.t1 B.t0 403.274
R70 B B.t1 303.514
R71 a_368_53.t0 a_368_53.t1 72.8576
C0 A_N B 2.03e-19
C1 VPB C 0.033862f
C2 VPWR B 0.130941f
C3 VPB X 0.011946f
C4 A_N C 7.6e-19
C5 VPB VGND 0.009087f
C6 VPWR C 0.005002f
C7 A_N X 1.44e-19
C8 B C 0.067126f
C9 VPWR X 0.073204f
C10 A_N VGND 0.045011f
C11 VPWR VGND 0.06573f
C12 B X 0.001187f
C13 C X 0.017607f
C14 B VGND 0.007965f
C15 C VGND 0.067785f
C16 X VGND 0.064694f
C17 VPB A_N 0.111271f
C18 VPB VPWR 0.104099f
C19 A_N VPWR 0.051269f
C20 VPB B 0.091418f
C21 VGND VNB 0.439533f
C22 X VNB 0.092491f
C23 C VNB 0.113921f
C24 B VNB 0.1008f
C25 VPWR VNB 0.341582f
C26 A_N VNB 0.196803f
C27 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_4 VNB VPB VGND VPWR A_N X B C
X0 a_98_199.t0 A_N.t0 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1491 pd=1.55 as=0.108375 ps=1.01 w=0.42 l=0.15
X1 X.t3 a_56_297.t4 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR.t6 a_56_297.t5 X.t7 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.15825 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X3 VGND.t1 a_56_297.t6 X.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.108375 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR.t0 a_98_199.t2 a_56_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1875 pd=1.375 as=0.33 ps=2.66 w=1 l=0.15
X5 VPWR.t5 a_56_297.t7 X.t6 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X6 VGND.t2 a_56_297.t8 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_257_47.t0 B.t0 a_152_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.121875 ps=1.025 w=0.65 l=0.15
X8 X.t0 a_56_297.t9 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X9 X.t5 a_56_297.t10 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.1775 ps=1.355 w=1 l=0.15
X10 a_152_47.t0 a_98_199.t3 a_56_297.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.19825 ps=1.91 w=0.65 l=0.15
X11 VPWR.t1 C.t0 a_56_297.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.15 ps=1.3 w=1 l=0.15
X12 a_98_199.t1 A_N.t1 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.15825 ps=1.36 w=0.42 l=0.15
X13 a_56_297.t3 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1875 ps=1.375 w=1 l=0.15
X14 VGND.t5 C.t1 a_257_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.07475 ps=0.88 w=0.65 l=0.15
X15 X.t4 a_56_297.t11 VPWR.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
R0 A_N.n0 A_N.t1 224.934
R1 A_N A_N.n0 152.881
R2 A_N.n0 A_N.t0 131.748
R3 VGND.n2 VGND.n1 204.469
R4 VGND.n4 VGND.n3 198.964
R5 VGND.n7 VGND.n6 198.964
R6 VGND.n1 VGND.t4 62.8576
R7 VGND.n6 VGND.t5 51.6928
R8 VGND.n7 VGND.n5 31.624
R9 VGND.n6 VGND.t3 26.7697
R10 VGND.n3 VGND.t0 25.8467
R11 VGND.n3 VGND.t2 25.8467
R12 VGND.n1 VGND.t1 25.8467
R13 VGND.n5 VGND.n0 9.3005
R14 VGND.n5 VGND.n4 8.65932
R15 VGND.n4 VGND.n2 7.82046
R16 VGND.n8 VGND.n7 6.35761
R17 VGND.n2 VGND.n0 1.00575
R18 VGND VGND.n8 0.45787
R19 VGND.n8 VGND.n0 0.16644
R20 a_98_199.n1 a_98_199.t1 652.038
R21 a_98_199.n1 a_98_199.n0 389.442
R22 a_98_199.t0 a_98_199.n1 309
R23 a_98_199.n0 a_98_199.t2 241.536
R24 a_98_199.n0 a_98_199.t3 169.237
R25 VNB.t7 VNB.t5 1637.54
R26 VNB VNB.t0 1537.86
R27 VNB.t0 VNB.t1 1495.15
R28 VNB.t3 VNB.t6 1452.43
R29 VNB.t2 VNB.t3 1224.6
R30 VNB.t4 VNB.t2 1224.6
R31 VNB.t5 VNB.t4 1224.6
R32 VNB.t1 VNB.t7 1082.2
R33 a_56_297.n10 a_56_297.n9 638.476
R34 a_56_297.t0 a_56_297.n11 383.639
R35 a_56_297.n1 a_56_297.t5 212.081
R36 a_56_297.n2 a_56_297.t11 212.081
R37 a_56_297.n4 a_56_297.t7 212.081
R38 a_56_297.n6 a_56_297.t10 212.081
R39 a_56_297.n3 a_56_297.n0 164.992
R40 a_56_297.n8 a_56_297.n7 152
R41 a_56_297.n5 a_56_297.n0 152
R42 a_56_297.n5 a_56_297.t8 139.78
R43 a_56_297.n1 a_56_297.t6 139.78
R44 a_56_297.n2 a_56_297.t4 139.78
R45 a_56_297.n6 a_56_297.t9 139.78
R46 a_56_297.n11 a_56_297.t1 124.603
R47 a_56_297.n11 a_56_297.n10 110.022
R48 a_56_297.n2 a_56_297.n1 62.8066
R49 a_56_297.n7 a_56_297.n5 49.6611
R50 a_56_297.n4 a_56_297.n3 48.2005
R51 a_56_297.n9 a_56_297.t3 31.5205
R52 a_56_297.n9 a_56_297.t2 27.5805
R53 a_56_297.n3 a_56_297.n2 13.146
R54 a_56_297.n7 a_56_297.n6 13.146
R55 a_56_297.n8 a_56_297.n0 12.9915
R56 a_56_297.n10 a_56_297.n8 9.74378
R57 a_56_297.n5 a_56_297.n4 1.46111
R58 X.n2 X.n0 649
R59 X.n2 X.n1 585
R60 X.n5 X.n4 232.862
R61 X.n5 X.n3 95.6721
R62 X.n6 X.n2 39.6933
R63 X.n0 X.t5 29.5505
R64 X.n0 X.t6 27.5805
R65 X.n1 X.t7 27.5805
R66 X.n1 X.t4 27.5805
R67 X.n4 X.t1 25.8467
R68 X.n4 X.t0 25.8467
R69 X.n3 X.t2 25.8467
R70 X.n3 X.t3 25.8467
R71 X X.n5 6.95702
R72 X X.n6 3.86465
R73 X.n6 X 1.94833
R74 VPWR.n4 VPWR.n3 753.082
R75 VPWR.n2 VPWR.n1 598.965
R76 VPWR.n6 VPWR.n5 598.755
R77 VPWR.n14 VPWR.n13 585
R78 VPWR.n3 VPWR.t7 103.191
R79 VPWR.n13 VPWR.t0 40.3855
R80 VPWR.n1 VPWR.t4 35.4605
R81 VPWR.n1 VPWR.t1 34.4755
R82 VPWR.n7 VPWR.n2 34.2593
R83 VPWR.n3 VPWR.t6 33.5187
R84 VPWR.n13 VPWR.t2 33.4905
R85 VPWR.n12 VPWR.n11 33.1015
R86 VPWR.n5 VPWR.t3 26.5955
R87 VPWR.n5 VPWR.t5 26.5955
R88 VPWR.n15 VPWR.n14 16.3463
R89 VPWR.n11 VPWR.n2 10.1652
R90 VPWR.n8 VPWR.n7 9.3005
R91 VPWR.n9 VPWR.n2 9.3005
R92 VPWR.n11 VPWR.n10 9.3005
R93 VPWR.n12 VPWR.n0 9.3005
R94 VPWR.n7 VPWR.n6 8.65932
R95 VPWR.n6 VPWR.n4 7.44399
R96 VPWR.n14 VPWR.n12 4.46842
R97 VPWR.n8 VPWR.n4 1.00575
R98 VPWR.n15 VPWR.n0 0.141672
R99 VPWR VPWR.n15 0.121778
R100 VPWR.n9 VPWR.n8 0.120292
R101 VPWR.n10 VPWR.n9 0.120292
R102 VPWR.n10 VPWR.n0 0.120292
R103 VPB VPB.t0 319.627
R104 VPB.t0 VPB.t2 310.748
R105 VPB.t6 VPB.t7 301.87
R106 VPB.t1 VPB.t4 298.911
R107 VPB.t2 VPB.t1 266.356
R108 VPB.t4 VPB.t5 260.437
R109 VPB.t3 VPB.t6 254.518
R110 VPB.t5 VPB.t3 248.599
R111 B.n0 B.t1 237.328
R112 B.n0 B.t0 165.029
R113 B B.n0 155.274
R114 a_152_47.t0 a_152_47.t1 69.2313
R115 a_257_47.t0 a_257_47.t1 42.462
R116 C.n0 C.t0 241.536
R117 C.n0 C.t1 169.237
R118 C C.n0 155.897
C0 C X 2.36e-19
C1 VPB C 0.027085f
C2 VPWR X 0.032231f
C3 B C 0.080355f
C4 VPB VPWR 0.102461f
C5 C VGND 0.010125f
C6 VPWR A_N 0.019661f
C7 VPB X 0.004254f
C8 B VPWR 0.01578f
C9 VPWR VGND 0.093036f
C10 X A_N 0.090123f
C11 VPB A_N 0.094623f
C12 B X 2.01e-20
C13 VPB B 0.029539f
C14 X VGND 0.155136f
C15 VPB VGND 0.010729f
C16 A_N VGND 0.040889f
C17 B VGND 0.011224f
C18 C VPWR 0.013159f
C19 VGND VNB 0.54182f
C20 A_N VNB 0.159163f
C21 X VNB 0.010642f
C22 VPWR VNB 0.454083f
C23 C VNB 0.090749f
C24 B VNB 0.094855f
C25 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VPB VNB
X0 a_27_47.t0 C.t0 VPWR.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47.t0 B.t0 a_109_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X.t1 a_27_47.t5 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47.t1 C.t1 a_197_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47.t1 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR.t4 D.t0 a_27_47.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND.t0 D.t1 a_303_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR.t3 B.t1 a_27_47.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X.t0 a_27_47.t6 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47.t1 A.t1 a_27_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 C.n0 C.t0 334.723
R1 C.n0 C.t1 206.19
R2 C C.n0 154.347
R3 VPWR.n6 VPWR.t2 662.841
R4 VPWR.n4 VPWR.n3 599.74
R5 VPWR.n2 VPWR.n1 316.356
R6 VPWR.n1 VPWR.t4 117.451
R7 VPWR.n3 VPWR.t1 86.7743
R8 VPWR.n3 VPWR.t3 86.7743
R9 VPWR.n1 VPWR.t0 42.3555
R10 VPWR.n5 VPWR.n4 28.2358
R11 VPWR.n6 VPWR.n5 19.9534
R12 VPWR.n5 VPWR.n0 9.3005
R13 VPWR.n7 VPWR.n6 9.3005
R14 VPWR.n4 VPWR.n2 6.55
R15 VPWR.n2 VPWR.n0 0.267172
R16 VPWR.n7 VPWR.n0 0.120292
R17 VPWR VPWR.n7 0.0226354
R18 a_27_47.n4 a_27_47.n3 621.865
R19 a_27_47.n1 a_27_47.n0 617.513
R20 a_27_47.n1 a_27_47.t4 315.043
R21 a_27_47.n2 a_27_47.t5 230.793
R22 a_27_47.n3 a_27_47.n2 209.726
R23 a_27_47.n2 a_27_47.t6 158.494
R24 a_27_47.n0 a_27_47.t2 82.0838
R25 a_27_47.n0 a_27_47.t1 82.0838
R26 a_27_47.n4 a_27_47.t3 65.6672
R27 a_27_47.t0 a_27_47.n4 65.6672
R28 a_27_47.n3 a_27_47.n1 64.7534
R29 VPB.t4 VPB.t1 491.277
R30 VPB.t3 VPB.t0 307.788
R31 VPB.t2 VPB.t3 295.95
R32 VPB.t0 VPB.t4 254.518
R33 VPB VPB.t2 192.369
R34 B.n0 B.t1 334.723
R35 B.n0 B.t0 206.19
R36 B B.n0 166.446
R37 a_109_47.t0 a_109_47.t1 82.8576
R38 a_197_47.t0 a_197_47.t1 108.572
R39 VNB.t0 VNB.t3 2363.75
R40 VNB.t1 VNB.t2 1509.39
R41 VNB.t2 VNB.t0 1366.99
R42 VNB.t4 VNB.t1 1253.07
R43 VNB VNB.t4 925.567
R44 X.n4 X.n3 590.082
R45 X.n4 X.n0 585
R46 X.n5 X.n4 585
R47 X.n1 X.t0 129.381
R48 X.n4 X.t1 26.5955
R49 X X.n2 14.7697
R50 X X.n0 10.5851
R51 X.n5 X 10.5851
R52 X X.n1 7.0214
R53 X X.n0 6.15435
R54 X X.n5 6.15435
R55 X.n1 X 5.55208
R56 X.n3 X 3.93896
R57 X.n3 X 3.01226
R58 X.n2 X 1.96973
R59 X.n2 X 1.50638
R60 a_303_47.t0 a_303_47.t1 94.2862
R61 A.n0 A.t0 323.342
R62 A.n0 A.t1 194.809
R63 A A.n0 152.929
R64 D.n0 D.t0 330.12
R65 D.n0 D.t1 201.587
R66 D D.n0 154.514
R67 VGND VGND.n0 120.865
R68 VGND.n0 VGND.t0 108.505
R69 VGND.n0 VGND.t1 38.7697
C0 D VGND 0.089796f
C1 VPWR X 0.094506f
C2 VPB A 0.090662f
C3 VPWR VGND 0.066176f
C4 VPB B 0.064328f
C5 X VGND 0.09025f
C6 A B 0.083909f
C7 VPB C 0.060876f
C8 VPB D 0.078225f
C9 VPB VPWR 0.076952f
C10 B C 0.160614f
C11 VPB X 0.011072f
C12 A VPWR 0.043995f
C13 C D 0.180159f
C14 B VPWR 0.023081f
C15 VPB VGND 0.008524f
C16 A VGND 0.015122f
C17 C VPWR 0.021032f
C18 B VGND 0.045272f
C19 D VPWR 0.020729f
C20 C VGND 0.040816f
C21 D X 0.007457f
C22 VGND VNB 0.39291f
C23 X VNB 0.093317f
C24 VPWR VNB 0.334542f
C25 D VNB 0.130267f
C26 C VNB 0.109828f
C27 B VNB 0.112123f
C28 A VNB 0.220977f
C29 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_2 VNB VPB VGND VPWR X D C B A
X0 VGND.t2 a_27_47.t5 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND.t0 D.t0 a_304_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X.t3 a_27_47.t6 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47.t0 B.t0 a_109_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47.t1 C.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR.t4 a_27_47.t7 X.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47.t1 C.t1 a_198_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47.t0 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR.t0 D.t1 a_27_47.t4 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X.t0 a_27_47.t8 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR.t3 B.t1 a_27_47.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47.t1 A.t1 a_27_47.t3 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 a_27_47.n3 a_27_47.n2 621.865
R1 a_27_47.n5 a_27_47.n4 617.513
R2 a_27_47.n4 a_27_47.t3 315.236
R3 a_27_47.n3 a_27_47.n1 228.357
R4 a_27_47.n0 a_27_47.t7 212.081
R5 a_27_47.n1 a_27_47.t6 212.081
R6 a_27_47.n0 a_27_47.t5 139.78
R7 a_27_47.n1 a_27_47.t8 139.78
R8 a_27_47.t0 a_27_47.n5 84.4291
R9 a_27_47.n5 a_27_47.t2 82.0838
R10 a_27_47.n1 a_27_47.n0 70.1096
R11 a_27_47.n2 a_27_47.t4 65.6672
R12 a_27_47.n2 a_27_47.t1 65.6672
R13 a_27_47.n4 a_27_47.n3 64.7534
R14 X.n3 X 593.216
R15 X.n3 X.n2 585
R16 X.n4 X.n3 585
R17 X.n0 X 186.72
R18 X.n1 X.n0 185
R19 X.n3 X.t2 38.4155
R20 X.n0 X.t1 36.0005
R21 X.n3 X.t3 26.5955
R22 X.n0 X.t0 24.9236
R23 X.n6 X 21.9434
R24 X.n1 X 11.2721
R25 X.n2 X 8.21543
R26 X.n5 X.n4 6.30498
R27 X.n2 X 4.77662
R28 X.n4 X 4.77662
R29 X X.n5 3.65764
R30 X X.n6 2.92621
R31 X.n5 X 1.91095
R32 X X.n1 1.7199
R33 X.n6 X 1.52886
R34 VGND.n1 VGND.t2 149.72
R35 VGND.n1 VGND.n0 128.864
R36 VGND.n0 VGND.t0 121.353
R37 VGND.n0 VGND.t1 16.1729
R38 VGND VGND.n1 0.948592
R39 VNB.t0 VNB.t3 2178.64
R40 VNB.t2 VNB.t5 1509.39
R41 VNB.t3 VNB.t4 1366.99
R42 VNB.t5 VNB.t0 1366.99
R43 VNB.t1 VNB.t2 1267.31
R44 VNB VNB.t1 911.327
R45 D.n0 D.t1 330.12
R46 D.n0 D.t0 201.587
R47 D D.n0 154.708
R48 a_304_47.t0 a_304_47.t1 94.2862
R49 VPWR.n12 VPWR.t1 663.062
R50 VPWR.n10 VPWR.n2 599.74
R51 VPWR.n6 VPWR.t4 349.618
R52 VPWR.n5 VPWR.n4 310.502
R53 VPWR.n4 VPWR.t0 104.645
R54 VPWR.n2 VPWR.t2 86.7743
R55 VPWR.n2 VPWR.t3 86.7743
R56 VPWR.n4 VPWR.t5 42.3555
R57 VPWR.n9 VPWR.n3 34.6358
R58 VPWR.n11 VPWR.n10 28.6123
R59 VPWR.n12 VPWR.n11 19.9534
R60 VPWR.n10 VPWR.n9 15.8123
R61 VPWR.n5 VPWR.n3 12.424
R62 VPWR.n7 VPWR.n3 9.3005
R63 VPWR.n9 VPWR.n8 9.3005
R64 VPWR.n10 VPWR.n1 9.3005
R65 VPWR.n11 VPWR.n0 9.3005
R66 VPWR.n13 VPWR.n12 9.3005
R67 VPWR.n6 VPWR.n5 7.04885
R68 VPWR.n7 VPWR.n6 0.587432
R69 VPWR.n8 VPWR.n7 0.120292
R70 VPWR.n8 VPWR.n1 0.120292
R71 VPWR.n1 VPWR.n0 0.120292
R72 VPWR.n13 VPWR.n0 0.120292
R73 VPWR VPWR.n13 0.0213333
R74 VPB.t0 VPB.t5 452.805
R75 VPB.t3 VPB.t2 307.788
R76 VPB.t1 VPB.t3 298.911
R77 VPB.t5 VPB.t4 284.113
R78 VPB.t2 VPB.t0 254.518
R79 VPB VPB.t1 189.409
R80 B.n0 B.t1 334.723
R81 B.n0 B.t0 206.19
R82 B B.n0 166.243
R83 a_109_47.t0 a_109_47.t1 84.2862
R84 a_198_47.t0 a_198_47.t1 108.572
R85 C.n0 C.t0 334.723
R86 C.n0 C.t1 206.19
R87 C C.n0 154.347
R88 A.n0 A.t0 323.55
R89 A.n0 A.t1 195.017
R90 A A.n0 152.922
C0 D VGND 0.08079f
C1 VPWR X 0.157615f
C2 VPB A 0.090011f
C3 VPWR VGND 0.086668f
C4 VPB B 0.064559f
C5 X VGND 0.131519f
C6 VPB C 0.060875f
C7 A B 0.082601f
C8 VPB D 0.079232f
C9 B C 0.156914f
C10 VPB VPWR 0.092393f
C11 A VPWR 0.040856f
C12 VPB X 0.007046f
C13 C D 0.174741f
C14 B VPWR 0.023068f
C15 VPB VGND 0.010944f
C16 A VGND 0.013622f
C17 C VPWR 0.020869f
C18 D VPWR 0.021477f
C19 B VGND 0.041669f
C20 D X 0.007896f
C21 C VGND 0.037432f
C22 VGND VNB 0.467438f
C23 X VNB 0.036881f
C24 VPWR VNB 0.397956f
C25 D VNB 0.12821f
C26 C VNB 0.109758f
C27 B VNB 0.112394f
C28 A VNB 0.219485f
C29 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
X0 a_226_47.t0 A2_N.t0 a_226_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413.t0 B1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297.t1 A1_N.t0 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR.t2 B2.t0 a_489_413.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413.t1 a_226_47.t3 a_76_199.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199.t1 a_226_47.t4 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND.t1 B1.t1 a_556_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47.t1 B2.t1 a_76_199.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND.t2 A2_N.t1 a_226_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47.t2 A1_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR.t0 a_76_199.t3 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND.t4 a_76_199.t4 X.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2_N.n0 A2_N.t1 206.19
R1 A2_N A2_N.n0 154.429
R2 A2_N.n0 A2_N.t0 142.344
R3 a_226_297.t0 a_226_297.t1 98.5005
R4 a_226_47.t0 a_226_47.n2 710.439
R5 a_226_47.n1 a_226_47.t3 286.32
R6 a_226_47.n2 a_226_47.n0 272.719
R7 a_226_47.n2 a_226_47.n1 152
R8 a_226_47.n1 a_226_47.t4 131.099
R9 a_226_47.n0 a_226_47.t1 38.5719
R10 a_226_47.n0 a_226_47.t2 38.5719
R11 VPB.t2 VPB.t3 565.265
R12 VPB.t0 VPB.t5 346.262
R13 VPB.t4 VPB.t1 248.599
R14 VPB.t3 VPB.t4 248.599
R15 VPB.t5 VPB.t2 213.084
R16 VPB VPB.t0 189.409
R17 B1.n0 B1.t0 327.057
R18 B1.n0 B1.t1 239.768
R19 B1.n1 B1.n0 152
R20 B1.n1 B1 14.0313
R21 B1 B1.n1 2.70819
R22 VPWR.n2 VPWR.n1 612.725
R23 VPWR.n2 VPWR.n0 606.223
R24 VPWR.n0 VPWR.t3 143.06
R25 VPWR.n1 VPWR.t1 63.3219
R26 VPWR.n1 VPWR.t2 63.3219
R27 VPWR.n0 VPWR.t0 25.6105
R28 VPWR VPWR.n2 11.3621
R29 a_489_413.t0 a_489_413.n0 1331.51
R30 a_489_413.n0 a_489_413.t2 63.3219
R31 a_489_413.n0 a_489_413.t1 63.3219
R32 A1_N.n0 A1_N.t1 206.19
R33 A1_N.n1 A1_N.n0 152
R34 A1_N.n0 A1_N.t0 148.35
R35 A1_N.n1 A1_N 11.055
R36 A1_N A1_N.n1 2.13383
R37 B2.n0 B2.t1 305.803
R38 B2.n0 B2.t0 235.109
R39 B2 B2.n0 158.188
R40 a_76_199.t0 a_76_199.n2 648.322
R41 a_76_199.n2 a_76_199.n1 320.529
R42 a_76_199.n2 a_76_199.n0 318.526
R43 a_76_199.n0 a_76_199.t3 241.536
R44 a_76_199.n0 a_76_199.t4 169.237
R45 a_76_199.n1 a_76_199.t2 38.5719
R46 a_76_199.n1 a_76_199.t1 38.5719
R47 VGND.n5 VGND.t1 243.315
R48 VGND.n1 VGND.n0 198.248
R49 VGND.n9 VGND.n8 185
R50 VGND.n7 VGND.n6 185
R51 VGND.n8 VGND.n7 111.43
R52 VGND.n0 VGND.t0 85.7148
R53 VGND.n7 VGND.t3 38.5719
R54 VGND.n8 VGND.t2 38.5719
R55 VGND.n6 VGND.n5 32.5922
R56 VGND.n11 VGND.n10 29.8804
R57 VGND.n0 VGND.t4 25.9346
R58 VGND.n11 VGND.n1 15.4358
R59 VGND VGND.n13 11.0555
R60 VGND.n4 VGND.n3 9.3005
R61 VGND.n10 VGND.n2 9.3005
R62 VGND.n12 VGND.n11 9.3005
R63 VGND.n9 VGND.n3 8.64611
R64 VGND.n13 VGND.n1 4.968
R65 VGND.n13 VGND.n12 2.30116
R66 VGND.n10 VGND.n9 1.68471
R67 VGND.n5 VGND.n4 0.660127
R68 VGND.n4 VGND.n2 0.120292
R69 VGND.n12 VGND.n2 0.120292
R70 VGND.n6 VGND.n3 0.112781
R71 VNB.t2 VNB.t3 2306.8
R72 VNB.t5 VNB.t0 1666.02
R73 VNB.t4 VNB.t1 1196.12
R74 VNB.t3 VNB.t4 1196.12
R75 VNB.t0 VNB.t2 1196.12
R76 VNB VNB.t5 911.327
R77 a_556_47.t0 a_556_47.t1 77.1434
R78 X.t0 X 755.631
R79 X.n1 X.t0 755.481
R80 X.n0 X.t1 209.923
R81 X.n1 X.n0 76.1746
R82 X.n0 X 6.64665
R83 X X.n1 1.23127
C0 VPWR A1_N 0.006721f
C1 B1 VGND 0.047123f
C2 X A2_N 2.55e-19
C3 X VGND 0.062661f
C4 VPWR A2_N 0.004486f
C5 A1_N A2_N 0.10971f
C6 VPWR VGND 0.074322f
C7 VPB B2 0.064546f
C8 A1_N VGND 0.026061f
C9 VPB B1 0.080343f
C10 A2_N VGND 0.017355f
C11 VPB X 0.011346f
C12 B2 B1 0.181843f
C13 VPB VPWR 0.095098f
C14 B2 VPWR 0.016076f
C15 VPB A1_N 0.033866f
C16 VPB A2_N 0.032736f
C17 B1 VPWR 0.018786f
C18 X VPWR 0.058912f
C19 VPB VGND 0.012835f
C20 B2 VGND 0.033524f
C21 X A1_N 0.002114f
C22 VGND VNB 0.461507f
C23 A2_N VNB 0.103283f
C24 A1_N VNB 0.111357f
C25 VPWR VNB 0.368878f
C26 X VNB 0.097534f
C27 B1 VNB 0.206073f
C28 B2 VNB 0.106213f
C29 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_2 VNB VPB VGND VPWR B1 B2 A2_N A1_N X
X0 VPWR.t3 a_82_21.t3 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.435 as=0.135 ps=1.27 w=1 l=0.15
X1 a_646_47.t0 B2.t0 a_82_21.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_574_369.t1 a_313_47.t3 a_82_21.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_574_369.t2 B1.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 VGND.t2 a_82_21.t4 X.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t1 B2.t1 a_574_369.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X6 X.t2 a_82_21.t5 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 X.t0 a_82_21.t6 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8 a_313_47.t1 A2_N.t0 a_313_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_47.t2 A1_N.t0 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 a_313_297.t0 A1_N.t1 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.186 ps=1.435 w=0.64 l=0.15
X11 VGND.t0 A2_N.t1 a_313_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.14175 pd=1.095 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_82_21.t1 a_313_47.t4 VGND.t5 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.14175 ps=1.095 w=0.42 l=0.15
X13 VGND.t3 B1.t1 a_646_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R0 a_82_21.t0 a_82_21.n3 626.556
R1 a_82_21.n3 a_82_21.n1 326.283
R2 a_82_21.n3 a_82_21.n2 318.5
R3 a_82_21.n1 a_82_21.t3 212.081
R4 a_82_21.n0 a_82_21.t6 212.081
R5 a_82_21.n1 a_82_21.t4 139.78
R6 a_82_21.n0 a_82_21.t5 139.78
R7 a_82_21.n1 a_82_21.n0 61.346
R8 a_82_21.n2 a_82_21.t2 38.5719
R9 a_82_21.n2 a_82_21.t1 38.5719
R10 X.n2 X 589.016
R11 X.n3 X.n2 585
R12 X.n1 X.n0 185
R13 X.n3 X.n1 78.1809
R14 X.n2 X.t1 26.5955
R15 X.n2 X.t0 26.5955
R16 X.n0 X.t3 24.9236
R17 X.n0 X.t2 24.9236
R18 X.n1 X 6.77697
R19 X X.n3 1.2554
R20 VPWR.n4 VPWR.n3 748.265
R21 VPWR.n2 VPWR.n1 610.958
R22 VPWR.n0 VPWR.t2 259.964
R23 VPWR.n3 VPWR.t0 93.8833
R24 VPWR.n1 VPWR.t4 41.5552
R25 VPWR.n1 VPWR.t1 41.5552
R26 VPWR.n5 VPWR.n0 31.624
R27 VPWR.n3 VPWR.t3 29.0556
R28 VPWR.n5 VPWR.n4 19.577
R29 VPWR.n7 VPWR.n6 9.42029
R30 VPWR.n6 VPWR.n5 9.3005
R31 VPWR VPWR.n7 7.90638
R32 VPWR.n4 VPWR.n2 7.20206
R33 VPWR.n7 VPWR.n0 3.01226
R34 VPWR.n6 VPWR.n2 0.155249
R35 VPB.t3 VPB.t0 559.346
R36 VPB.t5 VPB.t1 346.262
R37 VPB.t0 VPB.t2 269.315
R38 VPB.t2 VPB.t6 248.599
R39 VPB.t4 VPB.t5 248.599
R40 VPB.t1 VPB.t3 213.084
R41 VPB VPB.t4 213.084
R42 B2.n0 B2.t0 305.803
R43 B2.n0 B2.t1 199.762
R44 B2 B2.n0 158.188
R45 a_646_47.t0 a_646_47.t1 77.1434
R46 VNB.t2 VNB.t0 2349.51
R47 VNB.t4 VNB.t5 1666.02
R48 VNB.t1 VNB.t6 1196.12
R49 VNB.t0 VNB.t1 1196.12
R50 VNB.t5 VNB.t2 1196.12
R51 VNB.t3 VNB.t4 1196.12
R52 VNB VNB.t3 1025.24
R53 a_313_47.t1 a_313_47.n2 683.403
R54 a_313_47.n2 a_313_47.n0 280.248
R55 a_313_47.n1 a_313_47.t3 257.842
R56 a_313_47.n2 a_313_47.n1 152
R57 a_313_47.n1 a_313_47.t4 138.018
R58 a_313_47.n0 a_313_47.t0 38.5719
R59 a_313_47.n0 a_313_47.t2 38.5719
R60 a_574_369.n0 a_574_369.t2 1311.23
R61 a_574_369.n0 a_574_369.t1 52.3286
R62 a_574_369.t0 a_574_369.n0 41.5552
R63 B1.n0 B1.t0 292.324
R64 B1.n0 B1.t1 241.43
R65 B1.n1 B1.n0 152
R66 B1.n1 B1 14.0313
R67 B1 B1.n1 2.70819
R68 VGND.n7 VGND.t3 243.74
R69 VGND.n12 VGND.n11 198.248
R70 VGND.n4 VGND.n3 185
R71 VGND.n6 VGND.n5 185
R72 VGND.n0 VGND.t1 159.48
R73 VGND.n5 VGND.n4 115.715
R74 VGND.n11 VGND.t4 85.7148
R75 VGND.n5 VGND.t5 38.5719
R76 VGND.n4 VGND.t0 38.5719
R77 VGND.n13 VGND.n0 31.624
R78 VGND.n10 VGND.n2 28.5594
R79 VGND.n11 VGND.t2 25.9346
R80 VGND.n13 VGND.n12 19.577
R81 VGND.n12 VGND.n10 17.3181
R82 VGND.n15 VGND.n14 9.42029
R83 VGND.n8 VGND.n2 9.3005
R84 VGND.n10 VGND.n9 9.3005
R85 VGND.n12 VGND.n1 9.3005
R86 VGND.n14 VGND.n13 9.3005
R87 VGND.n6 VGND.n3 9.09524
R88 VGND VGND.n15 7.90638
R89 VGND.n7 VGND.n6 7.26576
R90 VGND.n15 VGND.n0 3.01226
R91 VGND.n3 VGND.n2 1.12331
R92 VGND.n8 VGND.n7 0.26575
R93 VGND.n9 VGND.n8 0.120292
R94 VGND.n9 VGND.n1 0.120292
R95 VGND.n14 VGND.n1 0.120292
R96 A2_N.n0 A2_N.t1 206.19
R97 A2_N.n0 A2_N.t0 177.69
R98 A2_N A2_N.n0 154.429
R99 a_313_297.t0 a_313_297.t1 64.6411
R100 A1_N.n0 A1_N.t0 206.19
R101 A1_N.n0 A1_N.t1 183.696
R102 A1_N.n1 A1_N.n0 152
R103 A1_N.n1 A1_N 11.055
R104 A1_N A1_N.n1 2.13383
C0 VPWR VGND 0.095406f
C1 X A2_N 2.55e-19
C2 A1_N A2_N 0.10971f
C3 X VGND 0.1187f
C4 VPB B2 0.052064f
C5 A1_N VGND 0.027287f
C6 VPB B1 0.065853f
C7 A2_N VGND 0.01755f
C8 B2 B1 0.167345f
C9 VPB VPWR 0.106038f
C10 B2 VPWR 0.016115f
C11 VPB X 0.003829f
C12 B1 VPWR 0.018728f
C13 VPB A1_N 0.033667f
C14 VPB A2_N 0.033422f
C15 VPB VGND 0.013613f
C16 VPWR X 0.144494f
C17 VPWR A1_N 0.008853f
C18 B2 VGND 0.033524f
C19 VPWR A2_N 0.005343f
C20 X A1_N 0.002342f
C21 B1 VGND 0.046692f
C22 VGND VNB 0.540093f
C23 A2_N VNB 0.1055f
C24 A1_N VNB 0.111597f
C25 X VNB 0.026951f
C26 VPWR VNB 0.448052f
C27 B1 VNB 0.200775f
C28 B2 VNB 0.105342f
C29 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_4 VNB VPB VGND VPWR B1 B2 A1_N X A2_N
X0 VGND.t6 a_415_21.t6 a_193_47.t2 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_415_21.t5 A2_N.t0 a_717_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_717_297.t0 A1_N.t0 VPWR.t3 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND.t2 A2_N.t1 a_415_21.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_193_47.t4 a_415_21.t7 a_27_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297.t4 B1.t0 VPWR.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t7 a_193_47.t6 X.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t3 a_193_47.t7 VGND.t10 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t0 B2.t0 a_27_297.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t6 a_193_47.t8 VPWR.t6 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_415_21.t0 A1_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X11 a_415_21.t3 A2_N.t2 VGND.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X.t2 a_193_47.t9 VGND.t9 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297.t1 B2.t1 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_193_47.t0 B2.t2 a_109_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t11 B1.t1 a_109_47.t3 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND.t8 a_193_47.t10 X.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t1 A1_N.t2 a_415_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t7 a_193_47.t11 X.t0 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_109_47.t0 B2.t3 a_193_47.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_193_47.t1 a_415_21.t8 VGND.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR.t5 a_193_47.t12 X.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_27_297.t2 a_415_21.t9 a_193_47.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 X.t4 a_193_47.t13 VPWR.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR.t2 A1_N.t3 a_717_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR.t9 B1.t2 a_27_297.t5 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_717_297.t2 A2_N.t3 a_415_21.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_109_47.t2 B1.t3 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_415_21.n6 a_415_21.n5 690.644
R1 a_415_21.n1 a_415_21.t9 212.081
R2 a_415_21.n0 a_415_21.t7 212.081
R3 a_415_21.n5 a_415_21.n1 195.85
R4 a_415_21.n1 a_415_21.t6 139.78
R5 a_415_21.n0 a_415_21.t8 139.78
R6 a_415_21.n4 a_415_21.n2 135.249
R7 a_415_21.n4 a_415_21.n3 98.982
R8 a_415_21.n1 a_415_21.n0 61.346
R9 a_415_21.n5 a_415_21.n4 52.3982
R10 a_415_21.t4 a_415_21.n6 26.5955
R11 a_415_21.n6 a_415_21.t5 26.5955
R12 a_415_21.n2 a_415_21.t1 24.9236
R13 a_415_21.n2 a_415_21.t3 24.9236
R14 a_415_21.n3 a_415_21.t2 24.9236
R15 a_415_21.n3 a_415_21.t0 24.9236
R16 a_193_47.n13 a_193_47.n12 298.293
R17 a_193_47.n2 a_193_47.n0 263.017
R18 a_193_47.n4 a_193_47.t6 212.081
R19 a_193_47.n6 a_193_47.t8 212.081
R20 a_193_47.n8 a_193_47.t12 212.081
R21 a_193_47.n9 a_193_47.t13 212.081
R22 a_193_47.n5 a_193_47.n3 177.601
R23 a_193_47.n11 a_193_47.n10 152
R24 a_193_47.n7 a_193_47.n3 152
R25 a_193_47.n4 a_193_47.t11 139.78
R26 a_193_47.n6 a_193_47.t9 139.78
R27 a_193_47.n8 a_193_47.t10 139.78
R28 a_193_47.n9 a_193_47.t7 139.78
R29 a_193_47.n2 a_193_47.n1 99.1759
R30 a_193_47.n10 a_193_47.n9 49.6611
R31 a_193_47.n12 a_193_47.n11 40.8242
R32 a_193_47.n12 a_193_47.n2 38.2066
R33 a_193_47.n8 a_193_47.n7 37.9763
R34 a_193_47.n5 a_193_47.n4 35.055
R35 a_193_47.t3 a_193_47.n13 26.5955
R36 a_193_47.n13 a_193_47.t4 26.5955
R37 a_193_47.n6 a_193_47.n5 26.2914
R38 a_193_47.n11 a_193_47.n3 25.6005
R39 a_193_47.n1 a_193_47.t2 24.9236
R40 a_193_47.n1 a_193_47.t1 24.9236
R41 a_193_47.n0 a_193_47.t5 24.9236
R42 a_193_47.n0 a_193_47.t0 24.9236
R43 a_193_47.n7 a_193_47.n6 23.3702
R44 a_193_47.n10 a_193_47.n8 11.6853
R45 VGND.n10 VGND.t7 292.029
R46 VGND.n9 VGND.n8 207.965
R47 VGND.n17 VGND.n16 207.965
R48 VGND.n30 VGND.n29 207.965
R49 VGND.n27 VGND.n26 185
R50 VGND.n25 VGND.n24 185
R51 VGND.n37 VGND.t4 160.8
R52 VGND.n14 VGND.n6 121.451
R53 VGND.n26 VGND.n25 96.0005
R54 VGND.n10 VGND.n9 35.4566
R55 VGND.n13 VGND.n7 34.6358
R56 VGND.n18 VGND.n15 34.6358
R57 VGND.n23 VGND.n4 34.6358
R58 VGND.n31 VGND.n28 34.6358
R59 VGND.n35 VGND.n1 34.6358
R60 VGND.n36 VGND.n35 34.6358
R61 VGND.n37 VGND.n36 32.377
R62 VGND.n25 VGND.t0 24.9236
R63 VGND.n26 VGND.t6 24.9236
R64 VGND.n8 VGND.t9 24.9236
R65 VGND.n8 VGND.t8 24.9236
R66 VGND.n6 VGND.t10 24.9236
R67 VGND.n6 VGND.t1 24.9236
R68 VGND.n16 VGND.t3 24.9236
R69 VGND.n16 VGND.t2 24.9236
R70 VGND.n29 VGND.t5 24.9236
R71 VGND.n29 VGND.t11 24.9236
R72 VGND.n30 VGND.n1 24.8476
R73 VGND.n14 VGND.n13 23.3417
R74 VGND.n18 VGND.n17 17.3181
R75 VGND.n17 VGND.n4 17.3181
R76 VGND.n28 VGND.n27 14.124
R77 VGND.n38 VGND.n37 11.5593
R78 VGND.n15 VGND.n14 11.2946
R79 VGND.n31 VGND.n30 9.78874
R80 VGND.n36 VGND.n0 9.3005
R81 VGND.n35 VGND.n34 9.3005
R82 VGND.n33 VGND.n1 9.3005
R83 VGND.n32 VGND.n31 9.3005
R84 VGND.n28 VGND.n2 9.3005
R85 VGND.n21 VGND.n3 9.3005
R86 VGND.n11 VGND.n7 9.3005
R87 VGND.n13 VGND.n12 9.3005
R88 VGND.n15 VGND.n5 9.3005
R89 VGND.n19 VGND.n18 9.3005
R90 VGND.n20 VGND.n4 9.3005
R91 VGND.n23 VGND.n22 9.3005
R92 VGND.n24 VGND.n23 6.59462
R93 VGND.n24 VGND.n3 6.2005
R94 VGND.n9 VGND.n7 5.27109
R95 VGND.n27 VGND.n3 4.2005
R96 VGND.n11 VGND.n10 1.65809
R97 VGND.n12 VGND.n11 0.120292
R98 VGND.n12 VGND.n5 0.120292
R99 VGND.n19 VGND.n5 0.120292
R100 VGND.n20 VGND.n19 0.120292
R101 VGND.n22 VGND.n20 0.120292
R102 VGND.n22 VGND.n21 0.120292
R103 VGND.n21 VGND.n2 0.120292
R104 VGND.n32 VGND.n2 0.120292
R105 VGND.n33 VGND.n32 0.120292
R106 VGND.n34 VGND.n33 0.120292
R107 VGND.n34 VGND.n0 0.120292
R108 VGND.n38 VGND.n0 0.120292
R109 VGND VGND.n38 0.0213333
R110 VNB.t7 VNB.t0 2677.02
R111 VNB.t10 VNB.t8 1196.12
R112 VNB.t9 VNB.t10 1196.12
R113 VNB.t11 VNB.t9 1196.12
R114 VNB.t1 VNB.t11 1196.12
R115 VNB.t3 VNB.t1 1196.12
R116 VNB.t2 VNB.t3 1196.12
R117 VNB.t0 VNB.t2 1196.12
R118 VNB.t6 VNB.t7 1196.12
R119 VNB.t13 VNB.t6 1196.12
R120 VNB.t12 VNB.t13 1196.12
R121 VNB.t4 VNB.t12 1196.12
R122 VNB.t5 VNB.t4 1196.12
R123 VNB VNB.t5 911.327
R124 A2_N.n0 A2_N.t3 212.081
R125 A2_N.n1 A2_N.t0 212.081
R126 A2_N A2_N.n2 170.881
R127 A2_N.n0 A2_N.t2 139.78
R128 A2_N.n1 A2_N.t1 139.78
R129 A2_N.n2 A2_N.n1 31.4035
R130 A2_N.n2 A2_N.n0 29.9429
R131 a_717_297.n1 a_717_297.n0 935.158
R132 a_717_297.n0 a_717_297.t3 26.5955
R133 a_717_297.n0 a_717_297.t0 26.5955
R134 a_717_297.n1 a_717_297.t1 26.5955
R135 a_717_297.t2 a_717_297.n1 26.5955
R136 VPB.t6 VPB.t0 556.386
R137 VPB.t10 VPB.t11 248.599
R138 VPB.t9 VPB.t10 248.599
R139 VPB.t8 VPB.t9 248.599
R140 VPB.t1 VPB.t8 248.599
R141 VPB.t4 VPB.t1 248.599
R142 VPB.t5 VPB.t4 248.599
R143 VPB.t0 VPB.t5 248.599
R144 VPB.t7 VPB.t6 248.599
R145 VPB.t12 VPB.t7 248.599
R146 VPB.t2 VPB.t12 248.599
R147 VPB.t3 VPB.t2 248.599
R148 VPB.t13 VPB.t3 248.599
R149 VPB VPB.t13 189.409
R150 A1_N.n2 A1_N.n0 259.274
R151 A1_N.n1 A1_N.t3 241.536
R152 A1_N.n0 A1_N.t0 236.18
R153 A1_N.n1 A1_N.t2 169.237
R154 A1_N.n0 A1_N.t1 163.881
R155 A1_N.n2 A1_N.n1 152
R156 A1_N A1_N.n2 1.95606
R157 VPWR.n20 VPWR.t3 873.438
R158 VPWR.n28 VPWR.n1 606.505
R159 VPWR.n26 VPWR.n3 606.505
R160 VPWR.n11 VPWR.n10 604.968
R161 VPWR.n9 VPWR.t7 349.051
R162 VPWR.n13 VPWR.n8 318.293
R163 VPWR.n21 VPWR.n4 34.6358
R164 VPWR.n25 VPWR.n4 34.6358
R165 VPWR.n14 VPWR.n6 34.6358
R166 VPWR.n18 VPWR.n6 34.6358
R167 VPWR.n19 VPWR.n18 34.6358
R168 VPWR.n26 VPWR.n25 32.0005
R169 VPWR.n12 VPWR.n11 30.4946
R170 VPWR.n1 VPWR.t1 26.5955
R171 VPWR.n1 VPWR.t9 26.5955
R172 VPWR.n3 VPWR.t8 26.5955
R173 VPWR.n3 VPWR.t0 26.5955
R174 VPWR.n8 VPWR.t4 26.5955
R175 VPWR.n8 VPWR.t2 26.5955
R176 VPWR.n10 VPWR.t6 26.5955
R177 VPWR.n10 VPWR.t5 26.5955
R178 VPWR.n28 VPWR.n27 25.977
R179 VPWR.n27 VPWR.n26 18.4476
R180 VPWR.n21 VPWR.n20 13.9299
R181 VPWR.n13 VPWR.n12 13.9299
R182 VPWR.n12 VPWR.n7 9.3005
R183 VPWR.n15 VPWR.n14 9.3005
R184 VPWR.n16 VPWR.n6 9.3005
R185 VPWR.n18 VPWR.n17 9.3005
R186 VPWR.n19 VPWR.n5 9.3005
R187 VPWR.n22 VPWR.n21 9.3005
R188 VPWR.n23 VPWR.n4 9.3005
R189 VPWR.n25 VPWR.n24 9.3005
R190 VPWR.n26 VPWR.n2 9.3005
R191 VPWR.n27 VPWR.n0 9.3005
R192 VPWR.n29 VPWR.n28 7.27268
R193 VPWR.n11 VPWR.n9 6.47684
R194 VPWR.n14 VPWR.n13 1.88285
R195 VPWR.n20 VPWR.n19 1.88285
R196 VPWR.n9 VPWR.n7 0.58037
R197 VPWR.n29 VPWR.n0 0.146586
R198 VPWR.n15 VPWR.n7 0.120292
R199 VPWR.n16 VPWR.n15 0.120292
R200 VPWR.n17 VPWR.n16 0.120292
R201 VPWR.n17 VPWR.n5 0.120292
R202 VPWR.n22 VPWR.n5 0.120292
R203 VPWR.n23 VPWR.n22 0.120292
R204 VPWR.n24 VPWR.n23 0.120292
R205 VPWR.n24 VPWR.n2 0.120292
R206 VPWR.n2 VPWR.n0 0.120292
R207 VPWR VPWR.n29 0.115499
R208 a_27_297.n2 a_27_297.t2 889.837
R209 a_27_297.n1 a_27_297.t5 372.416
R210 a_27_297.n1 a_27_297.n0 301.397
R211 a_27_297.n3 a_27_297.n2 191.781
R212 a_27_297.n2 a_27_297.n1 53.1979
R213 a_27_297.n0 a_27_297.t0 26.5955
R214 a_27_297.n0 a_27_297.t1 26.5955
R215 a_27_297.t3 a_27_297.n3 26.5955
R216 a_27_297.n3 a_27_297.t4 26.5955
R217 B1.n2 B1.n0 257.935
R218 B1.n1 B1.t2 241.536
R219 B1.n0 B1.t0 241.536
R220 B1.n1 B1.t3 169.237
R221 B1.n0 B1.t1 169.237
R222 B1.n2 B1.n1 152
R223 B1 B1.n2 6.16346
R224 X.n2 X.n0 350.113
R225 X.n2 X.n1 196.083
R226 X.n5 X.n3 135.249
R227 X.n5 X.n4 98.982
R228 X X.n5 40.5912
R229 X X.n2 29.4632
R230 X.n1 X.t7 26.5955
R231 X.n1 X.t6 26.5955
R232 X.n0 X.t5 26.5955
R233 X.n0 X.t4 26.5955
R234 X.n3 X.t1 24.9236
R235 X.n3 X.t3 24.9236
R236 X.n4 X.t0 24.9236
R237 X.n4 X.t2 24.9236
R238 B2.n0 B2.t0 212.081
R239 B2.n1 B2.t1 212.081
R240 B2 B2.n2 153.304
R241 B2.n0 B2.t3 139.78
R242 B2.n1 B2.t2 139.78
R243 B2.n2 B2.n0 30.6732
R244 B2.n2 B2.n1 30.6732
R245 a_109_47.n1 a_109_47.n0 326.865
R246 a_109_47.n0 a_109_47.t3 24.9236
R247 a_109_47.n0 a_109_47.t0 24.9236
R248 a_109_47.t1 a_109_47.n1 24.9236
R249 a_109_47.n1 a_109_47.t2 24.9236
C0 VPB B2 0.051071f
C1 X VGND 0.28067f
C2 B1 B2 0.203413f
C3 VPB A1_N 0.066853f
C4 VPB A2_N 0.051106f
C5 VPB VPWR 0.163945f
C6 B1 VPWR 0.045458f
C7 VPB X 0.016767f
C8 B2 VPWR 0.033842f
C9 A1_N A2_N 0.219641f
C10 VPB VGND 0.013619f
C11 A1_N VPWR 0.045557f
C12 B1 VGND 0.055357f
C13 B2 VGND 0.018895f
C14 A2_N VPWR 0.011892f
C15 A1_N X 6.08e-19
C16 A2_N X 4.23e-19
C17 A1_N VGND 0.035722f
C18 VPWR X 0.310508f
C19 A2_N VGND 0.020941f
C20 VPB B1 0.065775f
C21 VPWR VGND 0.093434f
C22 VGND VNB 0.864786f
C23 X VNB 0.058656f
C24 VPWR VNB 0.687653f
C25 A2_N VNB 0.166948f
C26 A1_N VNB 0.193418f
C27 B2 VNB 0.167678f
C28 B1 VNB 0.235333f
C29 VPB VNB 1.49072f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2oi_1 VPB VNB VGND VPWR Y A2_N A1_N B2 B1
X0 a_109_47.t1 A2_N.t0 a_109_297.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 a_397_297.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 B2.t0 a_397_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND.t2 A2_N.t1 a_109_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.28275 pd=1.52 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_397_297.t1 a_109_47.t3 Y.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.34 ps=2.68 w=1 l=0.15
X5 a_481_47.t1 B2.t1 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y.t1 a_109_47.t4 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.28275 ps=1.52 w=0.65 l=0.15
X7 VGND.t0 B1.t1 a_481_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_109_297.t1 A1_N.t0 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47.t0 A1_N.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2_N.n0 A2_N.t0 241.536
R1 A2_N.n0 A2_N.t1 169.237
R2 A2_N A2_N.n0 160.695
R3 a_109_297.t0 a_109_297.t1 41.3705
R4 a_109_47.n2 a_109_47.n0 278.741
R5 a_109_47.t1 a_109_47.n2 276.334
R6 a_109_47.n2 a_109_47.n1 212.615
R7 a_109_47.n1 a_109_47.t3 212.081
R8 a_109_47.n1 a_109_47.t4 139.78
R9 a_109_47.n0 a_109_47.t2 24.9236
R10 a_109_47.n0 a_109_47.t0 24.9236
R11 VPB.t1 VPB.t2 639.253
R12 VPB.t3 VPB.t0 248.599
R13 VPB.t2 VPB.t3 248.599
R14 VPB.t4 VPB.t1 213.084
R15 VPB VPB.t4 192.369
R16 B1.n0 B1.t0 236.552
R17 B1.n0 B1.t1 164.251
R18 B1 B1.n0 154.429
R19 VPWR.n1 VPWR.n0 609.931
R20 VPWR.n1 VPWR.t2 344.406
R21 VPWR.n0 VPWR.t0 26.5955
R22 VPWR.n0 VPWR.t1 26.5955
R23 VPWR VPWR.n1 0.0621501
R24 a_397_297.t0 a_397_297.n0 984.596
R25 a_397_297.n0 a_397_297.t2 26.5955
R26 a_397_297.n0 a_397_297.t1 26.5955
R27 B2.n0 B2.t0 241.536
R28 B2.n0 B2.t1 169.237
R29 B2.n1 B2.n0 152
R30 B2.n1 B2 9.99502
R31 B2 B2.n1 1.92927
R32 VGND.n7 VGND.n6 185
R33 VGND.n5 VGND.n4 185
R34 VGND.n3 VGND.t0 156.911
R35 VGND.n9 VGND.t1 149.762
R36 VGND.n5 VGND.t3 72.9236
R37 VGND.n6 VGND.n5 62.7697
R38 VGND.n6 VGND.t2 24.9236
R39 VGND.n8 VGND.n7 22.1206
R40 VGND.n9 VGND.n8 19.9534
R41 VGND.n4 VGND.n3 11.5767
R42 VGND.n10 VGND.n9 9.3005
R43 VGND.n2 VGND.n1 9.3005
R44 VGND.n8 VGND.n0 9.3005
R45 VGND.n4 VGND.n1 6.45615
R46 VGND.n7 VGND.n1 1.11354
R47 VGND.n3 VGND.n2 0.220568
R48 VGND.n2 VGND.n0 0.120292
R49 VGND.n10 VGND.n0 0.120292
R50 VGND VGND.n10 0.0226354
R51 VNB.t3 VNB.t4 2904.85
R52 VNB.t1 VNB.t0 1196.12
R53 VNB.t4 VNB.t1 1196.12
R54 VNB.t2 VNB.t3 1196.12
R55 VNB VNB.t2 925.567
R56 Y.n0 Y.t2 323.373
R57 Y.n3 Y.n2 185
R58 Y.n3 Y.n1 99.7477
R59 Y.n2 Y.t0 24.9236
R60 Y.n2 Y.t1 24.9236
R61 Y.n1 Y 6.02403
R62 Y Y.n3 4.0191
R63 Y.n1 Y.n0 3.36141
R64 Y.n0 Y 2.58064
R65 a_481_47.t0 a_481_47.t1 49.8467
R66 A1_N.n0 A1_N.t0 241.536
R67 A1_N.n0 A1_N.t1 169.237
R68 A1_N.n1 A1_N.n0 152
R69 A1_N.n1 A1_N 9.85996
R70 A1_N A1_N.n1 1.9032
C0 B2 B1 0.118449f
C1 VPB VGND 0.008333f
C2 A2_N VPWR 0.019168f
C3 A1_N VGND 0.049228f
C4 B2 VPWR 0.018426f
C5 A2_N Y 5.53e-19
C6 B1 VPWR 0.017958f
C7 B2 Y 0.077815f
C8 A2_N VGND 0.018747f
C9 B1 Y 0.001119f
C10 B2 VGND 0.067818f
C11 VPWR Y 0.059486f
C12 B1 VGND 0.047865f
C13 VPB A1_N 0.03306f
C14 VPWR VGND 0.068054f
C15 VPB A2_N 0.03082f
C16 Y VGND 0.097822f
C17 VPB B2 0.027236f
C18 A1_N A2_N 0.084163f
C19 VPB B1 0.035037f
C20 VPB VPWR 0.07777f
C21 A1_N VPWR 0.049814f
C22 VPB Y 0.01055f
C23 VGND VNB 0.437984f
C24 Y VNB 0.010219f
C25 VPWR VNB 0.353892f
C26 B1 VNB 0.144942f
C27 B2 VNB 0.096931f
C28 A2_N VNB 0.096924f
C29 A1_N VNB 0.140732f
C30 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2oi_2 VNB VPB VGND VPWR A1_N Y B2 B1 A2_N
X0 a_54_297.t5 B1.t0 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_442_21.t1 A1_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X2 VPWR.t2 B2.t0 a_54_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_442_21.t5 A2_N.t0 VGND.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t5 B2.t1 a_136_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR.t0 A1_N.t1 a_662_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_54_297.t3 B2.t2 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_136_47.t1 B1.t1 VGND.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VGND.t0 A1_N.t2 a_442_21.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND.t2 A2_N.t1 a_442_21.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_136_47.t2 B2.t3 Y.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y.t1 a_442_21.t6 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t4 B1.t2 a_54_297.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_662_297.t3 A2_N.t2 a_442_21.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t6 B1.t3 a_136_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t3 a_442_21.t7 Y.t0 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_442_21.t4 A2_N.t3 a_662_297.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_662_297.t0 A1_N.t3 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_54_297.t0 a_442_21.t8 Y.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 Y.t2 a_442_21.t9 a_54_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R0 B1.n2 B1.n0 244.804
R1 B1.n1 B1.t2 241.536
R2 B1.n0 B1.t0 241.536
R3 B1.n1 B1.t1 169.237
R4 B1.n0 B1.t3 169.237
R5 B1.n2 B1.n1 152
R6 B1 B1.n2 9.48198
R7 VPWR.n3 VPWR.n2 612.919
R8 VPWR.n7 VPWR.n1 606.505
R9 VPWR.n5 VPWR.n4 606.505
R10 VPWR.n6 VPWR.n5 28.6123
R11 VPWR.n1 VPWR.t3 26.5955
R12 VPWR.n1 VPWR.t4 26.5955
R13 VPWR.n4 VPWR.t5 26.5955
R14 VPWR.n4 VPWR.t2 26.5955
R15 VPWR.n2 VPWR.t1 26.5955
R16 VPWR.n2 VPWR.t0 26.5955
R17 VPWR.n7 VPWR.n6 15.8123
R18 VPWR.n6 VPWR.n0 9.3005
R19 VPWR.n8 VPWR.n7 7.65909
R20 VPWR.n5 VPWR.n3 7.03895
R21 VPWR.n3 VPWR.n0 0.158455
R22 VPWR.n8 VPWR.n0 0.141672
R23 VPWR VPWR.n8 0.121778
R24 a_54_297.n1 a_54_297.t0 384.577
R25 a_54_297.t4 a_54_297.n3 372.416
R26 a_54_297.n3 a_54_297.n2 301.397
R27 a_54_297.n1 a_54_297.n0 288.212
R28 a_54_297.n3 a_54_297.n1 57.6089
R29 a_54_297.n0 a_54_297.t1 26.5955
R30 a_54_297.n0 a_54_297.t5 26.5955
R31 a_54_297.n2 a_54_297.t2 26.5955
R32 a_54_297.n2 a_54_297.t3 26.5955
R33 VPB.t2 VPB.t0 556.386
R34 VPB VPB.t6 272.274
R35 VPB.t9 VPB.t8 248.599
R36 VPB.t1 VPB.t9 248.599
R37 VPB.t0 VPB.t1 248.599
R38 VPB.t3 VPB.t2 248.599
R39 VPB.t7 VPB.t3 248.599
R40 VPB.t4 VPB.t7 248.599
R41 VPB.t5 VPB.t4 248.599
R42 VPB.t6 VPB.t5 248.599
R43 A1_N.n0 A1_N.t3 212.081
R44 A1_N.n1 A1_N.t1 212.081
R45 A1_N A1_N.n2 152.787
R46 A1_N.n0 A1_N.t2 139.78
R47 A1_N.n1 A1_N.t0 139.78
R48 A1_N.n2 A1_N.n0 32.1338
R49 A1_N.n2 A1_N.n1 29.2126
R50 VGND.n7 VGND.n6 207.965
R51 VGND.n18 VGND.n3 207.965
R52 VGND.n16 VGND.n15 185
R53 VGND.n14 VGND.n13 185
R54 VGND.n8 VGND.t2 170.091
R55 VGND.n25 VGND.t5 160.8
R56 VGND.n15 VGND.n14 96.0005
R57 VGND.n19 VGND.n1 34.6358
R58 VGND.n23 VGND.n1 34.6358
R59 VGND.n24 VGND.n23 34.6358
R60 VGND.n18 VGND.n17 34.2593
R61 VGND.n12 VGND.n5 30.7652
R62 VGND.n7 VGND.n5 27.4829
R63 VGND.n14 VGND.t1 24.9236
R64 VGND.n15 VGND.t3 24.9236
R65 VGND.n6 VGND.t7 24.9236
R66 VGND.n6 VGND.t0 24.9236
R67 VGND.n3 VGND.t4 24.9236
R68 VGND.n3 VGND.t6 24.9236
R69 VGND.n17 VGND.n16 24.2887
R70 VGND.n25 VGND.n24 22.2123
R71 VGND.n26 VGND.n25 21.724
R72 VGND.n8 VGND.n7 14.0525
R73 VGND.n24 VGND.n0 9.3005
R74 VGND.n23 VGND.n22 9.3005
R75 VGND.n21 VGND.n1 9.3005
R76 VGND.n20 VGND.n19 9.3005
R77 VGND.n17 VGND.n2 9.3005
R78 VGND.n10 VGND.n4 9.3005
R79 VGND.n9 VGND.n5 9.3005
R80 VGND.n12 VGND.n11 9.3005
R81 VGND.n13 VGND.n4 8.9005
R82 VGND.n16 VGND.n4 1.5005
R83 VGND.n9 VGND.n8 0.850429
R84 VGND.n19 VGND.n18 0.376971
R85 VGND.n13 VGND.n12 0.3005
R86 VGND.n11 VGND.n9 0.120292
R87 VGND.n11 VGND.n10 0.120292
R88 VGND.n10 VGND.n2 0.120292
R89 VGND.n20 VGND.n2 0.120292
R90 VGND.n21 VGND.n20 0.120292
R91 VGND.n22 VGND.n21 0.120292
R92 VGND.n22 VGND.n0 0.120292
R93 VGND.n26 VGND.n0 0.120292
R94 VGND VGND.n26 0.0226354
R95 a_442_21.n3 a_442_21.n0 433.293
R96 a_442_21.n2 a_442_21.t8 212.081
R97 a_442_21.n1 a_442_21.t9 212.081
R98 a_442_21.n3 a_442_21.n2 182.673
R99 a_442_21.n2 a_442_21.t7 139.78
R100 a_442_21.n1 a_442_21.t6 139.78
R101 a_442_21.n5 a_442_21.n4 135.249
R102 a_442_21.n6 a_442_21.n5 98.982
R103 a_442_21.n2 a_442_21.n1 61.346
R104 a_442_21.n5 a_442_21.n3 60.6375
R105 a_442_21.n0 a_442_21.t3 26.5955
R106 a_442_21.n0 a_442_21.t4 26.5955
R107 a_442_21.n4 a_442_21.t2 24.9236
R108 a_442_21.n4 a_442_21.t5 24.9236
R109 a_442_21.n6 a_442_21.t0 24.9236
R110 a_442_21.t1 a_442_21.n6 24.9236
R111 VNB.t5 VNB.t1 2677.02
R112 VNB VNB.t8 1310.03
R113 VNB.t9 VNB.t2 1196.12
R114 VNB.t0 VNB.t9 1196.12
R115 VNB.t1 VNB.t0 1196.12
R116 VNB.t6 VNB.t5 1196.12
R117 VNB.t7 VNB.t6 1196.12
R118 VNB.t4 VNB.t7 1196.12
R119 VNB.t3 VNB.t4 1196.12
R120 VNB.t8 VNB.t3 1196.12
R121 B2.n0 B2.t0 212.081
R122 B2.n1 B2.t2 212.081
R123 B2 B2.n2 162.881
R124 B2.n0 B2.t3 139.78
R125 B2.n1 B2.t1 139.78
R126 B2.n2 B2.n0 30.6732
R127 B2.n2 B2.n1 30.6732
R128 A2_N.n0 A2_N.t2 212.081
R129 A2_N.n1 A2_N.t3 212.081
R130 A2_N A2_N.n2 155.84
R131 A2_N.n0 A2_N.t1 139.78
R132 A2_N.n1 A2_N.t0 139.78
R133 A2_N.n2 A2_N.n1 32.1338
R134 A2_N.n2 A2_N.n0 29.2126
R135 a_136_47.n1 a_136_47.n0 326.865
R136 a_136_47.n0 a_136_47.t0 24.9236
R137 a_136_47.n0 a_136_47.t2 24.9236
R138 a_136_47.n1 a_136_47.t3 24.9236
R139 a_136_47.t1 a_136_47.n1 24.9236
R140 Y Y.n0 304.445
R141 Y.n3 Y.n1 259.257
R142 Y.n3 Y.n2 98.982
R143 Y Y.n3 27.3259
R144 Y.n0 Y.t3 26.5955
R145 Y.n0 Y.t2 26.5955
R146 Y.n2 Y.t0 24.9236
R147 Y.n2 Y.t1 24.9236
R148 Y.n1 Y.t4 24.9236
R149 Y.n1 Y.t5 24.9236
R150 a_662_297.t1 a_662_297.n1 382.622
R151 a_662_297.n1 a_662_297.t3 292.2
R152 a_662_297.n1 a_662_297.n0 288.212
R153 a_662_297.n0 a_662_297.t2 26.5955
R154 a_662_297.n0 a_662_297.t0 26.5955
C0 B1 B2 0.200396f
C1 VPB A1_N 0.057413f
C2 VPB A2_N 0.060649f
C3 VPB VPWR 0.117192f
C4 VPB Y 0.004864f
C5 B1 VPWR 0.048488f
C6 B1 Y 0.077163f
C7 B2 VPWR 0.03265f
C8 VPB VGND 0.011177f
C9 A1_N A2_N 0.064839f
C10 B1 VGND 0.058251f
C11 A1_N VPWR 0.033738f
C12 B2 Y 0.050033f
C13 A1_N Y 8.27e-19
C14 A2_N VPWR 0.021178f
C15 B2 VGND 0.018564f
C16 A1_N VGND 0.030248f
C17 A2_N Y 1.2e-19
C18 VPWR Y 0.011998f
C19 A2_N VGND 0.054931f
C20 VPB B1 0.070943f
C21 VPWR VGND 0.108246f
C22 VPB B2 0.051071f
C23 Y VGND 0.142952f
C24 VGND VNB 0.682533f
C25 Y VNB 0.015285f
C26 VPWR VNB 0.518318f
C27 A2_N VNB 0.210481f
C28 A1_N VNB 0.179878f
C29 B2 VNB 0.167865f
C30 B1 VNB 0.236366f
C31 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2oi_4 VNB VPB VGND VPWR Y B1 A2_N B2 A1_N
X0 Y.t3 B2.t0 a_109_47.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND.t3 B1.t0 a_109_47.t7 VNB.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND.t12 a_751_21.t12 Y.t4 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_751_21.t0 A2_N.t0 a_1139_297.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_1139_297.t5 A1_N.t0 VPWR.t7 VPB.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t11 B2.t1 a_27_297.t11 VPB.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t8 A2_N.t1 a_751_21.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_297.t10 B2.t2 VPWR.t10 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t6 A1_N.t1 a_1139_297.t6 VPB.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y.t5 a_751_21.t13 VGND.t13 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_1139_297.t7 A1_N.t2 VPWR.t5 VPB.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR.t3 B1.t1 a_27_297.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_297.t3 a_751_21.t14 Y.t6 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 Y.t7 a_751_21.t15 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t4 A1_N.t3 a_1139_297.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 a_751_21.t3 A1_N.t4 VGND.t6 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X16 a_27_297.t6 B1.t2 VPWR.t2 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297.t1 a_751_21.t16 Y.t8 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND.t2 B1.t3 a_109_47.t6 VNB.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y.t2 B2.t3 a_109_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y.t9 a_751_21.t17 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_1139_297.t2 A2_N.t2 a_751_21.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X22 a_751_21.t7 A2_N.t3 a_1139_297.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297.t5 B1.t4 VPWR.t1 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND.t7 A1_N.t5 a_751_21.t4 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VGND.t4 A1_N.t6 a_751_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_109_47.t5 B1.t5 VGND.t1 VNB.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VGND.t9 A2_N.t4 a_751_21.t8 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_109_47.t2 B2.t4 Y.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 VPWR.t9 B2.t5 a_27_297.t9 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_109_47.t1 B2.t6 Y.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 Y.t10 a_751_21.t18 VGND.t14 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_27_297.t8 B2.t7 VPWR.t8 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_751_21.t2 A1_N.t7 VGND.t5 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 a_751_21.t9 A2_N.t5 VGND.t10 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 VPWR.t0 B1.t6 a_27_297.t4 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 a_1139_297.t0 A2_N.t6 a_751_21.t10 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_109_47.t0 B1.t7 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 VGND.t15 a_751_21.t19 Y.t11 VNB.t16 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_751_21.t11 A2_N.t7 VGND.t11 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B2.n3 B2.t7 212.081
R1 B2.n1 B2.t5 212.081
R2 B2.n5 B2.t1 212.081
R3 B2.n6 B2.t2 212.081
R4 B2 B2.n7 158.4
R5 B2.n4 B2.n0 152
R6 B2.n3 B2.t0 139.78
R7 B2.n1 B2.t6 139.78
R8 B2.n5 B2.t4 139.78
R9 B2.n6 B2.t3 139.78
R10 B2.n2 B2.n0 92.1128
R11 B2.n4 B2.n3 49.6611
R12 B2.n7 B2.n5 37.9763
R13 B2.n2 B2.n1 34.6708
R14 B2.n7 B2.n6 23.3702
R15 B2.n3 B2.n2 20.1075
R16 B2 B2.n0 15.3605
R17 B2.n5 B2.n4 11.6853
R18 a_109_47.n2 a_109_47.n0 233.874
R19 a_109_47.n2 a_109_47.n1 185
R20 a_109_47.n5 a_109_47.n4 147.913
R21 a_109_47.n4 a_109_47.n3 88.3446
R22 a_109_47.n4 a_109_47.n2 53.5212
R23 a_109_47.n3 a_109_47.t3 24.9236
R24 a_109_47.n3 a_109_47.t5 24.9236
R25 a_109_47.n1 a_109_47.t4 24.9236
R26 a_109_47.n1 a_109_47.t2 24.9236
R27 a_109_47.n0 a_109_47.t7 24.9236
R28 a_109_47.n0 a_109_47.t1 24.9236
R29 a_109_47.n5 a_109_47.t6 24.9236
R30 a_109_47.t0 a_109_47.n5 24.9236
R31 Y.n10 Y.n9 303.473
R32 Y.n8 Y.n7 302.166
R33 Y.n5 Y.n3 226.355
R34 Y.n5 Y.n4 185
R35 Y.n2 Y.n1 135.391
R36 Y.n2 Y.n0 98.8627
R37 Y.n6 Y.n5 69.9629
R38 Y.n8 Y.n6 45.9299
R39 Y.n10 Y.n8 37.1205
R40 Y.n9 Y.t6 26.5955
R41 Y.n9 Y.t7 26.5955
R42 Y.n7 Y.t8 26.5955
R43 Y.n7 Y.t9 26.5955
R44 Y.n3 Y.t1 24.9236
R45 Y.n3 Y.t2 24.9236
R46 Y.n4 Y.t0 24.9236
R47 Y.n4 Y.t3 24.9236
R48 Y.n1 Y.t11 24.9236
R49 Y.n1 Y.t5 24.9236
R50 Y.n0 Y.t4 24.9236
R51 Y.n0 Y.t10 24.9236
R52 Y.n6 Y.n2 5.88122
R53 Y Y.n10 4.07323
R54 VNB.t16 VNB.t7 2677.02
R55 VNB.t12 VNB.t9 1196.12
R56 VNB.t10 VNB.t12 1196.12
R57 VNB.t11 VNB.t10 1196.12
R58 VNB.t1 VNB.t11 1196.12
R59 VNB.t2 VNB.t1 1196.12
R60 VNB.t8 VNB.t2 1196.12
R61 VNB.t7 VNB.t8 1196.12
R62 VNB.t14 VNB.t16 1196.12
R63 VNB.t13 VNB.t14 1196.12
R64 VNB.t15 VNB.t13 1196.12
R65 VNB.t19 VNB.t15 1196.12
R66 VNB.t3 VNB.t19 1196.12
R67 VNB.t6 VNB.t3 1196.12
R68 VNB.t4 VNB.t6 1196.12
R69 VNB.t5 VNB.t4 1196.12
R70 VNB.t17 VNB.t5 1196.12
R71 VNB.t18 VNB.t17 1196.12
R72 VNB.t0 VNB.t18 1196.12
R73 VNB VNB.t0 911.327
R74 B1.n3 B1.n2 326.37
R75 B1.n2 B1.t4 241.536
R76 B1.n1 B1.t1 212.081
R77 B1.n6 B1.t2 212.081
R78 B1.n7 B1.t6 212.081
R79 B1.n2 B1.t0 169.237
R80 B1.n4 B1.n3 152
R81 B1.n5 B1.n0 152
R82 B1.n9 B1.n8 152
R83 B1.n1 B1.t5 139.78
R84 B1.n6 B1.t3 139.78
R85 B1.n7 B1.t7 139.78
R86 B1.n5 B1.n4 49.6611
R87 B1.n8 B1.n6 48.9308
R88 B1 B1.n9 24.6862
R89 B1.n3 B1.n0 20.7243
R90 B1.n9 B1.n0 20.7243
R91 B1.n8 B1.n7 12.4157
R92 B1.n4 B1.n1 10.955
R93 B1.n6 B1.n5 0.730803
R94 VGND.n13 VGND.t8 298.442
R95 VGND.n14 VGND.n12 207.965
R96 VGND.n17 VGND.n16 207.965
R97 VGND.n23 VGND.n9 207.965
R98 VGND.n34 VGND.n6 207.965
R99 VGND.n37 VGND.n36 207.965
R100 VGND.n49 VGND.n1 207.965
R101 VGND.n28 VGND.n27 185
R102 VGND.n26 VGND.n25 185
R103 VGND.n51 VGND.t0 160.8
R104 VGND.n27 VGND.n26 96.0005
R105 VGND.n18 VGND.n15 34.6358
R106 VGND.n22 VGND.n10 34.6358
R107 VGND.n38 VGND.n35 34.6358
R108 VGND.n42 VGND.n4 34.6358
R109 VGND.n43 VGND.n42 34.6358
R110 VGND.n44 VGND.n43 34.6358
R111 VGND.n44 VGND.n2 34.6358
R112 VGND.n48 VGND.n2 34.6358
R113 VGND.n24 VGND.n23 33.8829
R114 VGND.n51 VGND.n50 32.377
R115 VGND.n50 VGND.n49 30.8711
R116 VGND.n33 VGND.n7 30.4887
R117 VGND.n17 VGND.n10 27.8593
R118 VGND.n34 VGND.n33 27.8593
R119 VGND.n26 VGND.t6 24.9236
R120 VGND.n27 VGND.t15 24.9236
R121 VGND.n12 VGND.t11 24.9236
R122 VGND.n12 VGND.t9 24.9236
R123 VGND.n16 VGND.t10 24.9236
R124 VGND.n16 VGND.t4 24.9236
R125 VGND.n9 VGND.t5 24.9236
R126 VGND.n9 VGND.t7 24.9236
R127 VGND.n6 VGND.t13 24.9236
R128 VGND.n6 VGND.t12 24.9236
R129 VGND.n36 VGND.t14 24.9236
R130 VGND.n36 VGND.t3 24.9236
R131 VGND.n1 VGND.t1 24.9236
R132 VGND.n1 VGND.t2 24.9236
R133 VGND.n25 VGND.n24 24.6652
R134 VGND.n15 VGND.n14 21.8358
R135 VGND.n38 VGND.n37 21.8358
R136 VGND.n14 VGND.n13 19.5226
R137 VGND.n37 VGND.n4 12.8005
R138 VGND.n52 VGND.n51 11.5593
R139 VGND.n50 VGND.n0 9.3005
R140 VGND.n48 VGND.n47 9.3005
R141 VGND.n46 VGND.n2 9.3005
R142 VGND.n45 VGND.n44 9.3005
R143 VGND.n43 VGND.n3 9.3005
R144 VGND.n42 VGND.n41 9.3005
R145 VGND.n40 VGND.n4 9.3005
R146 VGND.n39 VGND.n38 9.3005
R147 VGND.n35 VGND.n5 9.3005
R148 VGND.n33 VGND.n32 9.3005
R149 VGND.n31 VGND.n7 9.3005
R150 VGND.n30 VGND.n29 9.3005
R151 VGND.n15 VGND.n11 9.3005
R152 VGND.n19 VGND.n18 9.3005
R153 VGND.n20 VGND.n10 9.3005
R154 VGND.n22 VGND.n21 9.3005
R155 VGND.n24 VGND.n8 9.3005
R156 VGND.n29 VGND.n28 9.0005
R157 VGND.n18 VGND.n17 6.77697
R158 VGND.n35 VGND.n34 6.77697
R159 VGND.n49 VGND.n48 3.76521
R160 VGND.n29 VGND.n25 1.4005
R161 VGND.n13 VGND.n11 1.02737
R162 VGND.n23 VGND.n22 0.753441
R163 VGND.n28 VGND.n7 0.2005
R164 VGND.n19 VGND.n11 0.120292
R165 VGND.n20 VGND.n19 0.120292
R166 VGND.n21 VGND.n20 0.120292
R167 VGND.n21 VGND.n8 0.120292
R168 VGND.n30 VGND.n8 0.120292
R169 VGND.n31 VGND.n30 0.120292
R170 VGND.n32 VGND.n31 0.120292
R171 VGND.n32 VGND.n5 0.120292
R172 VGND.n39 VGND.n5 0.120292
R173 VGND.n40 VGND.n39 0.120292
R174 VGND.n41 VGND.n40 0.120292
R175 VGND.n41 VGND.n3 0.120292
R176 VGND.n45 VGND.n3 0.120292
R177 VGND.n46 VGND.n45 0.120292
R178 VGND.n47 VGND.n46 0.120292
R179 VGND.n47 VGND.n0 0.120292
R180 VGND.n52 VGND.n0 0.120292
R181 VGND VGND.n52 0.0213333
R182 a_751_21.n17 a_751_21.n16 345.31
R183 a_751_21.n16 a_751_21.n15 300.885
R184 a_751_21.n3 a_751_21.t14 212.081
R185 a_751_21.n4 a_751_21.t15 212.081
R186 a_751_21.n1 a_751_21.t16 212.081
R187 a_751_21.n0 a_751_21.t17 212.081
R188 a_751_21.n6 a_751_21.n5 152
R189 a_751_21.n3 a_751_21.t19 139.78
R190 a_751_21.n4 a_751_21.t13 139.78
R191 a_751_21.n1 a_751_21.t12 139.78
R192 a_751_21.n0 a_751_21.t18 139.78
R193 a_751_21.n8 a_751_21.n7 98.982
R194 a_751_21.n10 a_751_21.n9 98.982
R195 a_751_21.n12 a_751_21.n11 98.982
R196 a_751_21.n14 a_751_21.n13 98.982
R197 a_751_21.n8 a_751_21.n6 98.0768
R198 a_751_21.n6 a_751_21.n2 96.7795
R199 a_751_21.n16 a_751_21.n14 72.4768
R200 a_751_21.n1 a_751_21.n0 61.346
R201 a_751_21.n5 a_751_21.n4 40.1672
R202 a_751_21.n10 a_751_21.n8 36.2672
R203 a_751_21.n12 a_751_21.n10 36.2672
R204 a_751_21.n14 a_751_21.n12 36.2672
R205 a_751_21.n4 a_751_21.n2 29.3979
R206 a_751_21.n15 a_751_21.t6 26.5955
R207 a_751_21.n15 a_751_21.t7 26.5955
R208 a_751_21.n17 a_751_21.t10 26.5955
R209 a_751_21.t0 a_751_21.n17 26.5955
R210 a_751_21.n2 a_751_21.n1 25.447
R211 a_751_21.n13 a_751_21.t5 24.9236
R212 a_751_21.n13 a_751_21.t11 24.9236
R213 a_751_21.n7 a_751_21.t4 24.9236
R214 a_751_21.n7 a_751_21.t3 24.9236
R215 a_751_21.n9 a_751_21.t1 24.9236
R216 a_751_21.n9 a_751_21.t2 24.9236
R217 a_751_21.n11 a_751_21.t8 24.9236
R218 a_751_21.n11 a_751_21.t9 24.9236
R219 a_751_21.n5 a_751_21.n3 21.1793
R220 A2_N.n2 A2_N.t2 212.081
R221 A2_N.n1 A2_N.t3 212.081
R222 A2_N.n7 A2_N.t6 212.081
R223 A2_N.n8 A2_N.t0 212.081
R224 A2_N.n4 A2_N.n3 173.761
R225 A2_N A2_N.n9 161.921
R226 A2_N.n5 A2_N.n4 152
R227 A2_N.n6 A2_N.n0 152
R228 A2_N.n2 A2_N.t1 139.78
R229 A2_N.n1 A2_N.t7 139.78
R230 A2_N.n7 A2_N.t4 139.78
R231 A2_N.n8 A2_N.t5 139.78
R232 A2_N.n6 A2_N.n5 49.6611
R233 A2_N.n3 A2_N.n1 44.549
R234 A2_N.n9 A2_N.n7 43.0884
R235 A2_N.n4 A2_N.n0 21.7605
R236 A2_N.n9 A2_N.n8 18.2581
R237 A2_N.n3 A2_N.n2 16.7975
R238 A2_N A2_N.n0 11.8405
R239 A2_N.n7 A2_N.n6 6.57323
R240 A2_N.n5 A2_N.n1 5.11262
R241 a_1139_297.n1 a_1139_297.n0 585
R242 a_1139_297.n1 a_1139_297.t2 374.668
R243 a_1139_297.n3 a_1139_297.t4 274.827
R244 a_1139_297.n3 a_1139_297.n2 209.06
R245 a_1139_297.n5 a_1139_297.n4 187.506
R246 a_1139_297.n4 a_1139_297.n1 67.8142
R247 a_1139_297.n4 a_1139_297.n3 65.8023
R248 a_1139_297.n2 a_1139_297.t6 26.5955
R249 a_1139_297.n2 a_1139_297.t7 26.5955
R250 a_1139_297.n0 a_1139_297.t1 26.5955
R251 a_1139_297.n0 a_1139_297.t0 26.5955
R252 a_1139_297.t3 a_1139_297.n5 26.5955
R253 a_1139_297.n5 a_1139_297.t5 26.5955
R254 VPB.t3 VPB.t12 556.386
R255 VPB.t5 VPB.t6 248.599
R256 VPB.t4 VPB.t5 248.599
R257 VPB.t7 VPB.t4 248.599
R258 VPB.t17 VPB.t7 248.599
R259 VPB.t18 VPB.t17 248.599
R260 VPB.t19 VPB.t18 248.599
R261 VPB.t12 VPB.t19 248.599
R262 VPB.t2 VPB.t3 248.599
R263 VPB.t1 VPB.t2 248.599
R264 VPB.t0 VPB.t1 248.599
R265 VPB.t9 VPB.t0 248.599
R266 VPB.t14 VPB.t9 248.599
R267 VPB.t13 VPB.t14 248.599
R268 VPB.t16 VPB.t13 248.599
R269 VPB.t15 VPB.t16 248.599
R270 VPB.t11 VPB.t15 248.599
R271 VPB.t10 VPB.t11 248.599
R272 VPB.t8 VPB.t10 248.599
R273 VPB VPB.t8 189.409
R274 A1_N.n3 A1_N.t0 212.081
R275 A1_N.n5 A1_N.t1 212.081
R276 A1_N.n7 A1_N.t2 212.081
R277 A1_N.n1 A1_N.t3 212.081
R278 A1_N.n4 A1_N.n0 173.761
R279 A1_N.n9 A1_N.n2 173.761
R280 A1_N.n6 A1_N.n0 152
R281 A1_N.n9 A1_N.n8 152
R282 A1_N.n3 A1_N.t6 139.78
R283 A1_N.n5 A1_N.t7 139.78
R284 A1_N.n7 A1_N.t5 139.78
R285 A1_N.n1 A1_N.t4 139.78
R286 A1_N.n8 A1_N.n6 49.6611
R287 A1_N.n7 A1_N.n2 46.0096
R288 A1_N.n5 A1_N.n4 41.6278
R289 A1_N.n4 A1_N.n3 19.7187
R290 A1_N.n2 A1_N.n1 15.3369
R291 A1_N A1_N.n0 13.1205
R292 A1_N A1_N.n9 8.6405
R293 A1_N.n6 A1_N.n5 8.03383
R294 A1_N.n8 A1_N.n7 3.65202
R295 VPWR.n30 VPWR.n3 606.505
R296 VPWR.n5 VPWR.n4 606.505
R297 VPWR.n24 VPWR.n7 606.505
R298 VPWR.n14 VPWR.n11 323.914
R299 VPWR.n13 VPWR.n12 323.192
R300 VPWR.n32 VPWR.n1 323.192
R301 VPWR.n26 VPWR.n25 34.6358
R302 VPWR.n17 VPWR.n10 34.6358
R303 VPWR.n18 VPWR.n17 34.6358
R304 VPWR.n19 VPWR.n18 34.6358
R305 VPWR.n19 VPWR.n8 34.6358
R306 VPWR.n23 VPWR.n8 34.6358
R307 VPWR.n30 VPWR.n29 32.0005
R308 VPWR.n13 VPWR.n10 30.4946
R309 VPWR.n1 VPWR.t2 26.5955
R310 VPWR.n1 VPWR.t0 26.5955
R311 VPWR.n3 VPWR.t10 26.5955
R312 VPWR.n3 VPWR.t3 26.5955
R313 VPWR.n4 VPWR.t8 26.5955
R314 VPWR.n4 VPWR.t11 26.5955
R315 VPWR.n7 VPWR.t1 26.5955
R316 VPWR.n7 VPWR.t9 26.5955
R317 VPWR.n12 VPWR.t5 26.5955
R318 VPWR.n12 VPWR.t4 26.5955
R319 VPWR.n11 VPWR.t7 26.5955
R320 VPWR.n11 VPWR.t6 26.5955
R321 VPWR.n32 VPWR.n31 25.977
R322 VPWR.n31 VPWR.n30 18.4476
R323 VPWR.n29 VPWR.n5 12.424
R324 VPWR.n24 VPWR.n23 9.41227
R325 VPWR.n15 VPWR.n10 9.3005
R326 VPWR.n17 VPWR.n16 9.3005
R327 VPWR.n18 VPWR.n9 9.3005
R328 VPWR.n20 VPWR.n19 9.3005
R329 VPWR.n21 VPWR.n8 9.3005
R330 VPWR.n23 VPWR.n22 9.3005
R331 VPWR.n25 VPWR.n6 9.3005
R332 VPWR.n27 VPWR.n26 9.3005
R333 VPWR.n29 VPWR.n28 9.3005
R334 VPWR.n30 VPWR.n2 9.3005
R335 VPWR.n31 VPWR.n0 9.3005
R336 VPWR.n33 VPWR.n32 7.4049
R337 VPWR.n14 VPWR.n13 6.64705
R338 VPWR.n25 VPWR.n24 6.4005
R339 VPWR.n26 VPWR.n5 3.38874
R340 VPWR.n15 VPWR.n14 0.581083
R341 VPWR.n33 VPWR.n0 0.144904
R342 VPWR.n16 VPWR.n15 0.120292
R343 VPWR.n16 VPWR.n9 0.120292
R344 VPWR.n20 VPWR.n9 0.120292
R345 VPWR.n21 VPWR.n20 0.120292
R346 VPWR.n22 VPWR.n21 0.120292
R347 VPWR.n22 VPWR.n6 0.120292
R348 VPWR.n27 VPWR.n6 0.120292
R349 VPWR.n28 VPWR.n27 0.120292
R350 VPWR.n28 VPWR.n2 0.120292
R351 VPWR.n2 VPWR.n0 0.120292
R352 VPWR VPWR.n33 0.117202
R353 a_27_297.n9 a_27_297.n8 301.233
R354 a_27_297.n3 a_27_297.n2 300.885
R355 a_27_297.n5 a_27_297.n4 300.885
R356 a_27_297.n7 a_27_297.n6 288.212
R357 a_27_297.n1 a_27_297.t4 287.399
R358 a_27_297.t3 a_27_297.n9 272.877
R359 a_27_297.n1 a_27_297.n0 195.78
R360 a_27_297.n9 a_27_297.n7 57.0969
R361 a_27_297.n7 a_27_297.n5 57.0969
R362 a_27_297.n3 a_27_297.n1 49.8182
R363 a_27_297.n5 a_27_297.n3 44.424
R364 a_27_297.n6 a_27_297.t0 26.5955
R365 a_27_297.n6 a_27_297.t5 26.5955
R366 a_27_297.n0 a_27_297.t7 26.5955
R367 a_27_297.n0 a_27_297.t6 26.5955
R368 a_27_297.n2 a_27_297.t11 26.5955
R369 a_27_297.n2 a_27_297.t10 26.5955
R370 a_27_297.n4 a_27_297.t9 26.5955
R371 a_27_297.n4 a_27_297.t8 26.5955
R372 a_27_297.n8 a_27_297.t2 26.5955
R373 a_27_297.n8 a_27_297.t1 26.5955
C0 VPB VPWR 0.183498f
C1 B1 VPWR 0.086497f
C2 VPB Y 0.008426f
C3 B2 VPWR 0.057634f
C4 VPB VGND 0.013584f
C5 B1 Y 0.091594f
C6 A1_N A2_N 0.063906f
C7 A1_N VPWR 0.083588f
C8 B1 VGND 0.083394f
C9 B2 Y 0.143852f
C10 A2_N VPWR 0.032262f
C11 A1_N Y 0.001125f
C12 B2 VGND 0.033595f
C13 A2_N Y 1.51e-19
C14 A1_N VGND 0.0612f
C15 VPWR Y 0.022096f
C16 A2_N VGND 0.050696f
C17 VPB B1 0.125636f
C18 VPWR VGND 0.188414f
C19 VPB B2 0.114821f
C20 Y VGND 0.273547f
C21 VPB A1_N 0.120638f
C22 B1 B2 0.293612f
C23 VPB A2_N 0.120825f
C24 VGND VNB 1.0804f
C25 Y VNB 0.019485f
C26 VPWR VNB 0.855614f
C27 A2_N VNB 0.379394f
C28 A1_N VNB 0.363338f
C29 B2 VNB 0.351341f
C30 B1 VNB 0.396552f
C31 VPB VNB 1.9337f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21bo_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_1 VNB VPB VGND VPWR X A2 A1 B1_N
X0 a_298_297.t1 a_27_413.t2 a_215_297.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297.t0 a_27_413.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297.t0 A2.t0 VPWR.t3 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X.t0 a_215_297.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR.t0 B1_N.t0 a_27_413.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X.t1 a_215_297.t4 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47.t0 A1.t0 a_215_297.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND.t3 B1_N.t1 a_27_413.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR.t2 A1.t1 a_298_297.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t2 A2.t1 a_382_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_27_413.t0 a_27_413.n1 695.548
R1 a_27_413.n1 a_27_413.n0 314.63
R2 a_27_413.n1 a_27_413.t1 275.144
R3 a_27_413.n0 a_27_413.t3 200.833
R4 a_27_413.n0 a_27_413.t2 192.8
R5 a_215_297.t1 a_215_297.n2 264.067
R6 a_215_297.n2 a_215_297.n0 244.399
R7 a_215_297.n0 a_215_297.t4 231.244
R8 a_215_297.n0 a_215_297.t3 158.945
R9 a_215_297.n2 a_215_297.n1 94.9644
R10 a_215_297.n1 a_215_297.t2 24.9236
R11 a_215_297.n1 a_215_297.t0 24.9236
R12 a_298_297.t0 a_298_297.n0 676.949
R13 a_298_297.n0 a_298_297.t2 26.5955
R14 a_298_297.n0 a_298_297.t1 26.5955
R15 VPB.t2 VPB.t1 559.346
R16 VPB.t0 VPB.t3 559.346
R17 VPB.t4 VPB.t2 254.518
R18 VPB.t3 VPB.t4 248.599
R19 VPB VPB.t0 192.369
R20 VGND.n3 VGND.n2 185
R21 VGND.n5 VGND.n4 185
R22 VGND.n11 VGND.n10 117.889
R23 VGND.n10 VGND.t3 68.1564
R24 VGND.n4 VGND.n3 64.6159
R25 VGND.n10 VGND.t1 41.6479
R26 VGND.n4 VGND.t0 41.539
R27 VGND.n3 VGND.t2 40.6159
R28 VGND.n9 VGND.n8 34.6358
R29 VGND.n11 VGND.n9 31.624
R30 VGND.n8 VGND.n1 26.3813
R31 VGND.n6 VGND.n5 9.50262
R32 VGND.n6 VGND.n1 9.3005
R33 VGND.n8 VGND.n7 9.3005
R34 VGND.n9 VGND.n0 9.3005
R35 VGND.n5 VGND.n2 8.2968
R36 VGND.n12 VGND.n11 6.88217
R37 VGND.n2 VGND.n1 0.711611
R38 VGND VGND.n12 0.226733
R39 VGND.n12 VGND.n0 0.15696
R40 VGND.n7 VGND.n6 0.120292
R41 VGND.n7 VGND.n0 0.120292
R42 VNB.t3 VNB.t0 2691.26
R43 VNB VNB.t4 1908.09
R44 VNB.t4 VNB.t1 1708.74
R45 VNB.t2 VNB.t3 1224.6
R46 VNB.t1 VNB.t2 1196.12
R47 A2.n0 A2.t0 231.017
R48 A2.n0 A2.t1 158.716
R49 A2.n1 A2.n0 152
R50 A2.n1 A2 14.0313
R51 A2 A2.n1 2.70819
R52 VPWR.n7 VPWR.t0 662.22
R53 VPWR.n2 VPWR.n1 603.619
R54 VPWR.n3 VPWR.t1 252.575
R55 VPWR.n6 VPWR.n5 34.6358
R56 VPWR.n1 VPWR.t3 27.5805
R57 VPWR.n1 VPWR.t2 27.5805
R58 VPWR.n7 VPWR.n6 21.4593
R59 VPWR.n5 VPWR.n2 20.7064
R60 VPWR.n5 VPWR.n4 9.3005
R61 VPWR.n6 VPWR.n0 9.3005
R62 VPWR.n8 VPWR.n7 7.12063
R63 VPWR.n3 VPWR.n2 6.71073
R64 VPWR.n4 VPWR.n3 0.560616
R65 VPWR.n8 VPWR.n0 0.148519
R66 VPWR.n4 VPWR.n0 0.120292
R67 VPWR VPWR.n8 0.114842
R68 X.n0 X.t1 353.317
R69 X.n1 X.t0 209.923
R70 X.n1 X 8.91479
R71 X X.n0 8.15228
R72 X.n0 X 7.23962
R73 X X.n1 6.62907
R74 B1_N.n1 B1_N.t1 299.911
R75 B1_N.n0 B1_N.t0 199.762
R76 B1_N.n0 B1_N 155.061
R77 B1_N.n2 B1_N.n1 152
R78 B1_N.n1 B1_N.n0 60.6968
R79 B1_N.n2 B1_N 15.8614
R80 B1_N B1_N.n2 3.06137
R81 A1.n0 A1.t1 241.536
R82 A1.n0 A1.t0 169.237
R83 A1.n1 A1.n0 152
R84 A1.n1 A1 8.58403
R85 A1 A1.n1 1.65697
R86 a_382_47.t0 a_382_47.t1 51.6928
C0 VPWR X 0.114913f
C1 A2 VGND 0.019667f
C2 VPWR VGND 0.07888f
C3 X VGND 0.057294f
C4 VPB B1_N 0.103238f
C5 VPB A1 0.027656f
C6 VPB A2 0.041742f
C7 B1_N A1 1.31e-20
C8 VPB VPWR 0.097622f
C9 B1_N A2 4.62e-21
C10 A1 A2 0.111772f
C11 B1_N VPWR 0.018972f
C12 VPB X 0.011733f
C13 A1 VPWR 0.021516f
C14 B1_N X 2.01e-19
C15 VPB VGND 0.011706f
C16 B1_N VGND 0.049226f
C17 A1 X 1.5e-19
C18 A2 VPWR 0.030697f
C19 A2 X 0.005686f
C20 A1 VGND 0.01436f
C21 VGND VNB 0.439582f
C22 X VNB 0.089001f
C23 VPWR VNB 0.36562f
C24 A2 VNB 0.107548f
C25 A1 VNB 0.089279f
C26 B1_N VNB 0.290462f
C27 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21bo_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_2 VNB VPB VGND VPWR B1_N A1 X A2
X0 VPWR.t0 A1.t0 a_485_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_485_297.t2 a_297_93.t2 a_79_21.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_297_93.t0 B1_N.t0 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.108375 ps=1.01 w=0.42 l=0.15
X3 a_581_47.t0 A1.t1 a_79_21.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 VGND.t2 a_79_21.t3 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.108375 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_79_21.t1 a_297_93.t3 VGND.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND.t4 A2.t0 a_581_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 VPWR.t2 a_79_21.t4 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1815 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X8 a_297_93.t1 B1_N.t1 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1815 ps=1.51 w=0.42 l=0.15
X9 X.t2 a_79_21.t5 VPWR.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 a_485_297.t1 A2.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 X.t0 a_79_21.t6 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t0 241.536
R1 A1.n0 A1.t1 169.237
R2 A1 A1.n0 160.791
R3 a_485_297.n0 a_485_297.t1 661.947
R4 a_485_297.t0 a_485_297.n0 26.5955
R5 a_485_297.n0 a_485_297.t2 26.5955
R6 VPWR.n6 VPWR.t3 868.5
R7 VPWR.n4 VPWR.n1 682.745
R8 VPWR.n3 VPWR.n2 613.097
R9 VPWR.n1 VPWR.t4 103.191
R10 VPWR.n1 VPWR.t2 27.2932
R11 VPWR.n2 VPWR.t1 26.5955
R12 VPWR.n2 VPWR.t0 26.5955
R13 VPWR.n5 VPWR.n4 26.3534
R14 VPWR.n6 VPWR.n5 19.9534
R15 VPWR.n5 VPWR.n0 9.3005
R16 VPWR.n7 VPWR.n6 9.3005
R17 VPWR.n4 VPWR.n3 6.78635
R18 VPWR.n3 VPWR.n0 0.172593
R19 VPWR.n7 VPWR.n0 0.120292
R20 VPWR VPWR.n7 0.0213333
R21 VPB.t5 VPB.t2 556.386
R22 VPB.t3 VPB.t5 301.87
R23 VPB.t4 VPB.t3 254.518
R24 VPB.t0 VPB.t1 248.599
R25 VPB.t2 VPB.t0 248.599
R26 VPB VPB.t4 189.409
R27 a_297_93.n1 a_297_93.t1 682.087
R28 a_297_93.t0 a_297_93.n1 252.819
R29 a_297_93.n0 a_297_93.t2 229.001
R30 a_297_93.n0 a_297_93.t3 155.607
R31 a_297_93.n1 a_297_93.n0 152
R32 a_79_21.t2 a_79_21.n4 316.846
R33 a_79_21.n4 a_79_21.n0 282.224
R34 a_79_21.n4 a_79_21.n3 262.772
R35 a_79_21.n1 a_79_21.t4 221.72
R36 a_79_21.n2 a_79_21.t5 221.72
R37 a_79_21.n1 a_79_21.t3 149.421
R38 a_79_21.n2 a_79_21.t6 149.421
R39 a_79_21.n3 a_79_21.n2 47.3079
R40 a_79_21.n0 a_79_21.t0 33.2313
R41 a_79_21.n3 a_79_21.n1 29.4561
R42 a_79_21.n0 a_79_21.t1 27.6928
R43 B1_N B1_N.n0 168.332
R44 B1_N.n0 B1_N.t1 148.35
R45 B1_N.n0 B1_N.t0 132.282
R46 VGND.n4 VGND.t4 303.769
R47 VGND.n9 VGND.t1 287.151
R48 VGND.n3 VGND.t3 282.817
R49 VGND.n7 VGND.n2 120.678
R50 VGND.n2 VGND.t0 62.8576
R51 VGND.n7 VGND.n1 29.3652
R52 VGND.n3 VGND.n1 27.4829
R53 VGND.n9 VGND.n8 25.977
R54 VGND.n2 VGND.t2 25.8467
R55 VGND.n8 VGND.n7 24.8476
R56 VGND.n10 VGND.n9 9.3005
R57 VGND.n8 VGND.n0 9.3005
R58 VGND.n5 VGND.n1 9.3005
R59 VGND.n7 VGND.n6 9.3005
R60 VGND.n4 VGND.n3 6.59816
R61 VGND.n5 VGND.n4 0.277343
R62 VGND.n6 VGND.n5 0.120292
R63 VGND.n6 VGND.n0 0.120292
R64 VGND.n10 VGND.n0 0.120292
R65 VGND VGND.n10 0.0213333
R66 VNB.t1 VNB.t4 2677.02
R67 VNB.t3 VNB.t1 1452.43
R68 VNB.t4 VNB.t0 1366.99
R69 VNB.t2 VNB.t3 1224.6
R70 VNB.t0 VNB.t5 1025.24
R71 VNB VNB.t2 911.327
R72 a_581_47.t0 a_581_47.t1 38.7697
R73 X X.n0 320.409
R74 X X.n1 163.37
R75 X.n0 X.t3 27.5805
R76 X.n0 X.t2 27.5805
R77 X.n1 X.t1 25.8467
R78 X.n1 X.t0 25.8467
R79 A2.n0 A2.t1 233.288
R80 A2.n0 A2.t0 160.988
R81 A2 A2.n0 154.429
C0 VPB B1_N 0.039976f
C1 A2 VPWR 0.015179f
C2 VPB VGND 0.009183f
C3 VPWR X 0.103084f
C4 A1 VGND 0.030331f
C5 VPWR B1_N 0.005133f
C6 A2 VGND 0.051376f
C7 VPWR VGND 0.075731f
C8 X B1_N 0.003766f
C9 X VGND 0.135311f
C10 B1_N VGND 0.035776f
C11 VPB A1 0.027109f
C12 VPB A2 0.037839f
C13 VPB VPWR 0.088877f
C14 A1 A2 0.120267f
C15 VPB X 0.009846f
C16 A1 VPWR 0.018599f
C17 VGND VNB 0.495515f
C18 B1_N VNB 0.107647f
C19 X VNB 0.06873f
C20 VPWR VNB 0.374383f
C21 A2 VNB 0.149031f
C22 A1 VNB 0.089425f
C23 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21bo_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_4 VNB VPB VGND VPWR B1_N A2 X A1
X0 a_1021_47.t1 A1.t0 a_205_21.t5 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X.t3 a_205_21.t6 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR.t3 a_205_21.t7 X.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X.t4 a_205_21.t8 VGND.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND.t0 A2.t0 a_1021_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND.t1 a_42_47.t2 a_205_21.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_861_47.t0 A2.t1 VGND.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X7 a_205_21.t4 A1.t1 a_861_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.07475 ps=0.88 w=0.65 l=0.15
X8 X.t1 a_205_21.t9 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_603_297.t3 A1.t2 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND.t3 B1_N.t0 a_42_47.t0 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.25025 ps=2.07 w=0.65 l=0.15
X11 VPWR.t5 A2.t2 a_603_297.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_603_297.t5 a_42_47.t3 a_205_21.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR.t1 a_205_21.t10 X.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X14 a_205_21.t2 a_42_47.t4 a_603_297.t4 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t6 a_205_21.t11 X.t7 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.26325 pd=1.46 as=0.091 ps=0.93 w=0.65 l=0.15
X16 VPWR.t0 B1_N.t1 a_42_47.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X17 VGND.t5 a_205_21.t12 X.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VPWR.t7 A1.t3 a_603_297.t2 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_603_297.t0 A2.t3 VPWR.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_205_21.t3 a_42_47.t5 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26325 ps=1.46 w=0.65 l=0.15
X21 X.t5 a_205_21.t13 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 A1.n0 A1.t3 212.081
R1 A1.n1 A1.t2 212.081
R2 A1 A1.n2 153.929
R3 A1.n0 A1.t0 139.78
R4 A1.n1 A1.t1 139.78
R5 A1.n2 A1.n0 35.055
R6 A1.n2 A1.n1 26.2914
R7 a_205_21.n12 a_205_21.n0 649.754
R8 a_205_21.n0 a_205_21.n2 271.764
R9 a_205_21.n9 a_205_21.t10 212.081
R10 a_205_21.n7 a_205_21.t9 212.081
R11 a_205_21.n5 a_205_21.t7 212.081
R12 a_205_21.n4 a_205_21.t6 212.081
R13 a_205_21.n11 a_205_21.n1 96.3742
R14 a_205_21.n0 a_205_21.n1 2.11365
R15 a_205_21.n6 a_205_21.n3 165.189
R16 a_205_21.n10 a_205_21.n9 160.034
R17 a_205_21.n8 a_205_21.n3 152
R18 a_205_21.n9 a_205_21.t11 139.78
R19 a_205_21.n7 a_205_21.t13 139.78
R20 a_205_21.n5 a_205_21.t12 139.78
R21 a_205_21.n4 a_205_21.t8 139.78
R22 a_205_21.n1 a_205_21.n10 88.2013
R23 a_205_21.n5 a_205_21.n4 62.8066
R24 a_205_21.n9 a_205_21.n8 41.6278
R25 a_205_21.n6 a_205_21.n5 34.3247
R26 a_205_21.n7 a_205_21.n6 28.4823
R27 a_205_21.t1 a_205_21.n12 26.5955
R28 a_205_21.n12 a_205_21.t2 26.5955
R29 a_205_21.n11 a_205_21.t0 24.9236
R30 a_205_21.n11 a_205_21.t3 24.9236
R31 a_205_21.n2 a_205_21.t5 24.9236
R32 a_205_21.n2 a_205_21.t4 24.9236
R33 a_205_21.n8 a_205_21.n7 21.1793
R34 a_205_21.n10 a_205_21.n3 13.1884
R35 a_1021_47.t0 a_1021_47.t1 49.8467
R36 VNB.t6 VNB.t2 2733.98
R37 VNB VNB.t3 1495.15
R38 VNB.t1 VNB.t8 1310.03
R39 VNB.t4 VNB.t6 1224.6
R40 VNB.t5 VNB.t4 1224.6
R41 VNB.t7 VNB.t5 1224.6
R42 VNB.t3 VNB.t7 1224.6
R43 VNB.t10 VNB.t0 1196.12
R44 VNB.t9 VNB.t10 1196.12
R45 VNB.t2 VNB.t1 1196.12
R46 VNB.t8 VNB.t9 1082.2
R47 VPWR.n4 VPWR.t1 862.595
R48 VPWR.n9 VPWR.n8 604.321
R49 VPWR.n20 VPWR.n1 598.965
R50 VPWR.n18 VPWR.n3 598.965
R51 VPWR.n7 VPWR.n6 598.965
R52 VPWR.n12 VPWR.n11 34.6358
R53 VPWR.n13 VPWR.n12 34.6358
R54 VPWR.n19 VPWR.n18 32.377
R55 VPWR.n1 VPWR.t4 27.5805
R56 VPWR.n1 VPWR.t0 27.5805
R57 VPWR.n3 VPWR.t2 27.5805
R58 VPWR.n3 VPWR.t3 27.5805
R59 VPWR.n17 VPWR.n4 27.4829
R60 VPWR.n6 VPWR.t8 26.5955
R61 VPWR.n6 VPWR.t5 26.5955
R62 VPWR.n8 VPWR.t6 26.5955
R63 VPWR.n8 VPWR.t7 26.5955
R64 VPWR.n11 VPWR.n7 24.4711
R65 VPWR.n13 VPWR.n4 16.5652
R66 VPWR.n18 VPWR.n17 12.0476
R67 VPWR.n21 VPWR.n20 9.91792
R68 VPWR.n11 VPWR.n10 9.3005
R69 VPWR.n12 VPWR.n5 9.3005
R70 VPWR.n14 VPWR.n13 9.3005
R71 VPWR.n15 VPWR.n4 9.3005
R72 VPWR.n17 VPWR.n16 9.3005
R73 VPWR.n18 VPWR.n2 9.3005
R74 VPWR.n19 VPWR.n0 9.3005
R75 VPWR.n20 VPWR.n19 7.52991
R76 VPWR.n9 VPWR.n7 6.37482
R77 VPWR.n10 VPWR.n9 0.658988
R78 VPWR.n21 VPWR.n0 0.141672
R79 VPWR VPWR.n21 0.121778
R80 VPWR.n10 VPWR.n5 0.120292
R81 VPWR.n14 VPWR.n5 0.120292
R82 VPWR.n15 VPWR.n14 0.120292
R83 VPWR.n16 VPWR.n15 0.120292
R84 VPWR.n16 VPWR.n2 0.120292
R85 VPWR.n2 VPWR.n0 0.120292
R86 X.n2 X.n0 649.754
R87 X.n2 X.n1 585
R88 X.n5 X.n3 249.754
R89 X.n5 X.n4 185
R90 X X.n5 46.6027
R91 X.n1 X.t2 27.5805
R92 X.n1 X.t3 27.5805
R93 X.n0 X.t0 27.5805
R94 X.n0 X.t1 27.5805
R95 X.n4 X.t6 25.8467
R96 X.n4 X.t4 25.8467
R97 X.n3 X.t7 25.8467
R98 X.n3 X.t5 25.8467
R99 X X.n2 18.824
R100 VPB.t3 VPB.t1 568.225
R101 VPB VPB.t2 310.748
R102 VPB.t4 VPB.t3 254.518
R103 VPB.t5 VPB.t4 254.518
R104 VPB.t6 VPB.t5 254.518
R105 VPB.t2 VPB.t6 254.518
R106 VPB.t9 VPB.t8 248.599
R107 VPB.t10 VPB.t9 248.599
R108 VPB.t7 VPB.t10 248.599
R109 VPB.t0 VPB.t7 248.599
R110 VPB.t1 VPB.t0 248.599
R111 VGND.n7 VGND.n6 198.964
R112 VGND.n19 VGND.n18 198.964
R113 VGND.n1 VGND.n0 198.554
R114 VGND.n12 VGND.n11 185
R115 VGND.n10 VGND.n9 185
R116 VGND.n5 VGND.t0 160.224
R117 VGND.n11 VGND.n10 74.7697
R118 VGND.n11 VGND.t6 46.1543
R119 VGND.n17 VGND.n3 33.8686
R120 VGND.n20 VGND.n19 32.377
R121 VGND.n6 VGND.t1 32.3082
R122 VGND.n8 VGND.n7 30.4946
R123 VGND.n10 VGND.t2 28.6159
R124 VGND.n18 VGND.t4 25.8467
R125 VGND.n18 VGND.t5 25.8467
R126 VGND.n0 VGND.t7 25.8467
R127 VGND.n0 VGND.t3 25.8467
R128 VGND.n6 VGND.t8 24.9236
R129 VGND.n9 VGND.n8 16.4089
R130 VGND.n19 VGND.n17 12.0476
R131 VGND.n21 VGND.n20 9.3005
R132 VGND.n19 VGND.n2 9.3005
R133 VGND.n17 VGND.n16 9.3005
R134 VGND.n15 VGND.n3 9.3005
R135 VGND.n14 VGND.n13 9.3005
R136 VGND.n8 VGND.n4 9.3005
R137 VGND.n22 VGND.n1 9.16498
R138 VGND.n20 VGND.n1 7.52991
R139 VGND.n13 VGND.n12 6.64201
R140 VGND.n7 VGND.n5 6.44231
R141 VGND.n12 VGND.n3 4.46842
R142 VGND.n13 VGND.n9 3.14012
R143 VGND.n5 VGND.n4 0.187327
R144 VGND.n22 VGND.n21 0.141672
R145 VGND VGND.n22 0.121778
R146 VGND.n14 VGND.n4 0.120292
R147 VGND.n15 VGND.n14 0.120292
R148 VGND.n16 VGND.n15 0.120292
R149 VGND.n16 VGND.n2 0.120292
R150 VGND.n21 VGND.n2 0.120292
R151 A2 A2.n1 248.62
R152 A2.n1 A2.t2 241.536
R153 A2.n0 A2.t3 241.536
R154 A2 A2.n0 174.838
R155 A2.n1 A2.t1 169.237
R156 A2.n0 A2.t0 169.237
R157 a_42_47.n2 a_42_47.n1 456.118
R158 a_42_47.t1 a_42_47.n2 322.793
R159 a_42_47.n0 a_42_47.t3 212.081
R160 a_42_47.n1 a_42_47.t4 212.081
R161 a_42_47.n2 a_42_47.t0 198.459
R162 a_42_47.n0 a_42_47.t2 139.78
R163 a_42_47.n1 a_42_47.t5 139.78
R164 a_42_47.n1 a_42_47.n0 61.346
R165 a_861_47.t0 a_861_47.t1 42.462
R166 a_603_297.n1 a_603_297.n0 585
R167 a_603_297.n2 a_603_297.t4 399.911
R168 a_603_297.n1 a_603_297.t0 380.762
R169 a_603_297.n3 a_603_297.n2 298.993
R170 a_603_297.n2 a_603_297.n1 58.1201
R171 a_603_297.n0 a_603_297.t2 26.5955
R172 a_603_297.n0 a_603_297.t3 26.5955
R173 a_603_297.t1 a_603_297.n3 26.5955
R174 a_603_297.n3 a_603_297.t5 26.5955
R175 B1_N.n0 B1_N.t1 241.536
R176 B1_N.n0 B1_N.t0 169.237
R177 B1_N B1_N.n0 153.25
C0 VPB VPWR 0.122978f
C1 VPB X 0.004885f
C2 B1_N VPWR 0.015105f
C3 A2 A1 0.21368f
C4 B1_N X 0.054645f
C5 VPB VGND 0.010715f
C6 A2 VPWR 0.046703f
C7 A1 VPWR 0.031007f
C8 B1_N VGND 0.024309f
C9 A2 VGND 0.067407f
C10 VPWR X 0.035832f
C11 A1 VGND 0.032382f
C12 VPWR VGND 0.120933f
C13 X VGND 0.11182f
C14 VPB B1_N 0.032827f
C15 VPB A2 0.063244f
C16 VPB A1 0.051661f
C17 VGND VNB 0.700609f
C18 X VNB 0.016464f
C19 VPWR VNB 0.563712f
C20 A1 VNB 0.168166f
C21 A2 VNB 0.223491f
C22 B1_N VNB 0.116163f
C23 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_0 VNB VPB VPWR VGND A1 A2 B1_N Y
X0 a_300_369.t0 A2.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.0896 ps=0.92 w=0.64 l=0.15
X1 a_400_47.t0 A1.t0 Y.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=0.95 w=0.42 l=0.15
X2 VGND.t0 A2.t1 a_400_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND.t1 B1_N.t0 a_27_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.04 as=0.1113 ps=1.37 w=0.42 l=0.15
X4 VPWR.t0 B1_N.t1 a_27_47.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 Y.t1 a_27_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=0.95 as=0.1302 ps=1.04 w=0.42 l=0.15
X6 a_300_369.t2 a_27_47.t3 Y.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0896 pd=0.92 as=0.1696 ps=1.81 w=0.64 l=0.15
X7 VPWR.t2 A1.t1 a_300_369.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
R0 A2.n0 A2.t0 277.577
R1 A2.n0 A2.t1 143.858
R2 A2 A2.n0 77.5035
R3 VPWR.n1 VPWR.t0 672.65
R4 VPWR.n1 VPWR.n0 616.984
R5 VPWR.n0 VPWR.t1 43.0943
R6 VPWR.n0 VPWR.t2 43.0943
R7 VPWR VPWR.n1 0.203625
R8 a_300_369.t0 a_300_369.n0 697.663
R9 a_300_369.n0 a_300_369.t1 43.0943
R10 a_300_369.n0 a_300_369.t2 43.0943
R11 VPB.t0 VPB.t3 562.306
R12 VPB.t2 VPB.t1 254.518
R13 VPB.t3 VPB.t2 254.518
R14 VPB VPB.t0 195.327
R15 A1.n0 A1.t1 288.577
R16 A1.n0 A1.t0 158.631
R17 A1 A1.n0 71.7279
R18 Y Y.t2 630.227
R19 Y Y.n0 253.512
R20 Y.n0 Y.t0 111.43
R21 Y.n0 Y.t1 40.0005
R22 a_400_47.t0 a_400_47.t1 60.0005
R23 VNB.t2 VNB.t3 2192.88
R24 VNB.t3 VNB.t0 1936.57
R25 VNB.t0 VNB.t1 1025.24
R26 VNB VNB.t2 939.807
R27 VGND.n4 VGND.t0 248.829
R28 VGND.n3 VGND.n2 185
R29 VGND.n1 VGND.n0 185
R30 VGND.n2 VGND.n1 97.1434
R31 VGND.n2 VGND.t2 40.0005
R32 VGND.n1 VGND.t1 40.0005
R33 VGND.n4 VGND.n3 10.0216
R34 VGND.n5 VGND.n0 7.37107
R35 VGND.n3 VGND.n0 6.26237
R36 VGND.n5 VGND.n4 0.245611
R37 VGND VGND.n5 0.118068
R38 B1_N.n0 B1_N.t0 303.125
R39 B1_N.n0 B1_N.t1 165.001
R40 B1_N B1_N.n0 69.656
R41 a_27_47.t0 a_27_47.n1 732.74
R42 a_27_47.n0 a_27_47.t2 291.233
R43 a_27_47.n1 a_27_47.t1 245.661
R44 a_27_47.n0 a_27_47.t3 229.623
R45 a_27_47.n1 a_27_47.n0 188.077
C0 VPWR Y 0.064114f
C1 A2 VGND 0.047201f
C2 VPWR VGND 0.053616f
C3 Y VGND 0.092994f
C4 VPB B1_N 0.101016f
C5 VPB A1 0.05114f
C6 VPB A2 0.06108f
C7 VPB VPWR 0.071207f
C8 A1 A2 0.166501f
C9 B1_N VPWR 0.051585f
C10 VPB Y 0.013402f
C11 A1 VPWR 0.016956f
C12 VPB VGND 0.009415f
C13 B1_N Y 0.065368f
C14 B1_N VGND 0.020527f
C15 A2 VPWR 0.016139f
C16 A1 Y 0.080527f
C17 A1 VGND 0.032972f
C18 A2 Y 0.002148f
C19 VGND VNB 0.364934f
C20 Y VNB 0.01781f
C21 VPWR VNB 0.288959f
C22 A2 VNB 0.184932f
C23 A1 VNB 0.112827f
C24 B1_N VNB 0.16219f
C25 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB B1_N Y A1 A2
X0 a_300_297.t0 a_27_413.t2 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND.t0 A2.t0 a_384_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR.t1 B1_N.t0 a_27_413.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y.t0 a_27_413.t3 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 VPWR.t2 A1.t0 a_300_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47.t1 A1.t1 Y.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND.t2 B1_N.t1 a_27_413.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297.t2 A2.t1 VPWR.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
R0 a_27_413.t0 a_27_413.n1 695.918
R1 a_27_413.n1 a_27_413.n0 276.07
R2 a_27_413.n1 a_27_413.t1 269.324
R3 a_27_413.n0 a_27_413.t2 233.77
R4 a_27_413.n0 a_27_413.t3 200.833
R5 Y.n4 Y 592.177
R6 Y.n4 Y.n0 585
R7 Y.n5 Y.n4 585
R8 Y.n2 Y.n1 185
R9 Y.n1 Y.t2 40.6159
R10 Y.n1 Y.t0 40.6159
R11 Y.n3 Y.n2 30.5104
R12 Y.n4 Y.t1 27.5805
R13 Y Y.n0 7.17626
R14 Y.n5 Y 7.17626
R15 Y.n3 Y 6.18717
R16 Y Y.n0 6.01262
R17 Y Y.n5 6.01262
R18 Y.n2 Y 4.0191
R19 Y Y.n3 3.87929
R20 a_300_297.n0 a_300_297.t2 711.6
R21 a_300_297.n0 a_300_297.t1 27.5805
R22 a_300_297.t0 a_300_297.n0 27.5805
R23 VPB.t1 VPB.t0 562.306
R24 VPB.t2 VPB.t3 254.518
R25 VPB.t0 VPB.t2 254.518
R26 VPB VPB.t1 195.327
R27 A2.n0 A2.t1 231.017
R28 A2.n0 A2.t0 158.716
R29 A2 A2.n0 154.429
R30 a_384_47.t0 a_384_47.t1 51.6928
R31 VGND.n1 VGND.t0 156.174
R32 VGND.n1 VGND.n0 123.02
R33 VGND.n0 VGND.t2 57.8164
R34 VGND.n0 VGND.t1 25.6749
R35 VGND VGND.n1 0.309116
R36 VNB VNB.t2 1765.7
R37 VNB.t1 VNB.t3 1680.26
R38 VNB.t2 VNB.t1 1395.47
R39 VNB.t3 VNB.t0 1224.6
R40 B1_N.n1 B1_N.t1 283.844
R41 B1_N.n0 B1_N.t0 201.369
R42 B1_N B1_N.n0 155.061
R43 B1_N.n2 B1_N.n1 152
R44 B1_N.n1 B1_N.n0 60.6968
R45 B1_N B1_N.n2 15.8614
R46 B1_N.n2 B1_N 3.06137
R47 VPWR.n1 VPWR.t1 671.092
R48 VPWR.n1 VPWR.n0 315.757
R49 VPWR.n0 VPWR.t0 27.5805
R50 VPWR.n0 VPWR.t2 27.5805
R51 VPWR VPWR.n1 0.209829
R52 A1.n0 A1.t0 241.536
R53 A1.n0 A1.t1 169.237
R54 A1 A1.n0 156.755
C0 VPB B1_N 0.102846f
C1 VPB A1 0.026219f
C2 B1_N A1 2.36e-19
C3 VPB A2 0.037549f
C4 VPB VPWR 0.068716f
C5 A1 A2 0.092312f
C6 B1_N VPWR 0.018411f
C7 VPB Y 0.010913f
C8 VPB VGND 0.01018f
C9 B1_N Y 0.003656f
C10 A1 VPWR 0.021177f
C11 A1 Y 0.083515f
C12 A2 VPWR 0.021185f
C13 B1_N VGND 0.027178f
C14 A2 Y 8.84e-19
C15 A1 VGND 0.077228f
C16 A2 VGND 0.049294f
C17 VPWR Y 0.069054f
C18 VPWR VGND 0.057442f
C19 Y VGND 0.125367f
C20 VGND VNB 0.375628f
C21 Y VNB 0.013292f
C22 VPWR VNB 0.290723f
C23 A2 VNB 0.144296f
C24 A1 VNB 0.100718f
C25 B1_N VNB 0.255296f
C26 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_2 VNB VPB VPWR VGND B1_N A2 Y A1
X0 Y.t4 a_61_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183125 ps=1.24 w=0.65 l=0.15
X1 VPWR.t1 A2.t0 a_217_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297.t5 a_61_47.t3 Y.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47.t0 A2.t1 VGND.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 a_217_297.t0 A2.t2 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y.t1 a_61_47.t4 a_217_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR.t3 A1.t0 a_217_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47.t0 B1_N.t0 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VGND.t3 A2.t3 a_637_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND.t1 a_61_47.t5 Y.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y.t5 A1.t1 a_479_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.06825 ps=0.86 w=0.65 l=0.15
X11 VGND.t0 B1_N.t1 a_61_47.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.183125 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297.t3 A1.t2 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47.t1 A1.t3 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R0 a_61_47.t0 a_61_47.n2 696.206
R1 a_61_47.n2 a_61_47.t1 292.594
R2 a_61_47.n0 a_61_47.t3 218.507
R3 a_61_47.n1 a_61_47.t4 218.507
R4 a_61_47.n2 a_61_47.n1 213.373
R5 a_61_47.n0 a_61_47.t5 146.208
R6 a_61_47.n1 a_61_47.t2 146.208
R7 a_61_47.n1 a_61_47.n0 69.8074
R8 VGND.n3 VGND.n2 198.964
R9 VGND.n1 VGND.t3 144.355
R10 VGND.n6 VGND.n5 117.09
R11 VGND.n5 VGND.t0 72.1983
R12 VGND.n5 VGND.t2 44.3082
R13 VGND.n2 VGND.t1 35.0774
R14 VGND.n6 VGND.n4 28.9887
R15 VGND.n2 VGND.t4 25.8467
R16 VGND.n4 VGND.n3 24.8476
R17 VGND.n4 VGND.n0 9.3005
R18 VGND.n7 VGND.n6 7.06748
R19 VGND.n3 VGND.n1 6.87979
R20 VGND VGND.n7 0.228243
R21 VGND.n1 VGND.n0 0.180349
R22 VGND.n7 VGND.n0 0.154189
R23 Y.n3 Y.n2 353.731
R24 Y Y.n4 185.321
R25 Y.n4 Y.n3 185
R26 Y.n1 Y.n0 171.732
R27 Y.n2 Y.t2 26.5955
R28 Y.n2 Y.t1 26.5955
R29 Y.n0 Y.t0 25.8467
R30 Y.n0 Y.t5 25.8467
R31 Y.n4 Y.t3 24.9236
R32 Y.n4 Y.t4 24.9236
R33 Y Y.n1 17.6005
R34 Y.n3 Y.n1 3.8405
R35 VNB.t0 VNB.t3 2107.44
R36 VNB VNB.t0 1509.39
R37 VNB.t2 VNB.t5 1366.99
R38 VNB.t1 VNB.t4 1224.6
R39 VNB.t6 VNB.t1 1224.6
R40 VNB.t3 VNB.t2 1196.12
R41 VNB.t5 VNB.t6 1025.24
R42 A2 A2.n0 243.185
R43 A2.n0 A2.t0 241.536
R44 A2.n1 A2.t2 239.685
R45 A2.n0 A2.t1 169.237
R46 A2.n1 A2.t3 167.386
R47 A2 A2.n1 164.579
R48 a_217_297.t4 a_217_297.n3 370.914
R49 a_217_297.n1 a_217_297.t0 363.389
R50 a_217_297.n1 a_217_297.n0 296.125
R51 a_217_297.n3 a_217_297.n2 289.24
R52 a_217_297.n3 a_217_297.n1 58.7765
R53 a_217_297.n0 a_217_297.t2 27.5805
R54 a_217_297.n0 a_217_297.t3 27.5805
R55 a_217_297.n2 a_217_297.t1 26.5955
R56 a_217_297.n2 a_217_297.t5 26.5955
R57 VPWR.n12 VPWR.t2 672.194
R58 VPWR.n5 VPWR.n4 605.707
R59 VPWR.n3 VPWR.n2 604.206
R60 VPWR.n6 VPWR.n1 34.6358
R61 VPWR.n10 VPWR.n1 34.6358
R62 VPWR.n11 VPWR.n10 34.6358
R63 VPWR.n6 VPWR.n5 30.1181
R64 VPWR.n2 VPWR.t0 27.5805
R65 VPWR.n2 VPWR.t3 27.5805
R66 VPWR.n4 VPWR.t4 26.5955
R67 VPWR.n4 VPWR.t1 26.5955
R68 VPWR.n12 VPWR.n11 19.9534
R69 VPWR.n5 VPWR.n3 11.6392
R70 VPWR.n7 VPWR.n6 9.3005
R71 VPWR.n8 VPWR.n1 9.3005
R72 VPWR.n10 VPWR.n9 9.3005
R73 VPWR.n11 VPWR.n0 9.3005
R74 VPWR.n13 VPWR.n12 9.3005
R75 VPWR.n7 VPWR.n3 0.585982
R76 VPWR.n8 VPWR.n7 0.120292
R77 VPWR.n9 VPWR.n8 0.120292
R78 VPWR.n9 VPWR.n0 0.120292
R79 VPWR.n13 VPWR.n0 0.120292
R80 VPWR VPWR.n13 0.0213333
R81 VPB.t2 VPB.t5 559.346
R82 VPB.t3 VPB.t0 254.518
R83 VPB.t4 VPB.t3 254.518
R84 VPB.t1 VPB.t4 248.599
R85 VPB.t6 VPB.t1 248.599
R86 VPB.t5 VPB.t6 248.599
R87 VPB VPB.t2 192.369
R88 a_479_47.t0 a_479_47.t1 38.7697
R89 A1.n0 A1.t0 212.081
R90 A1.n1 A1.t2 212.081
R91 A1.n0 A1.t3 139.78
R92 A1.n1 A1.t1 139.78
R93 A1 A1.n2 68.5618
R94 A1.n2 A1.n1 30.3387
R95 A1.n2 A1.n0 25.7468
R96 B1_N.n0 B1_N.t0 254.97
R97 B1_N.n0 B1_N.t1 167.773
R98 B1_N B1_N.n0 76.7459
R99 a_637_47.t0 a_637_47.t1 51.6928
C0 Y VGND 0.22564f
C1 VPB A2 0.069917f
C2 VPB A1 0.053858f
C3 VPB B1_N 0.096186f
C4 A2 A1 0.225255f
C5 VPB VPWR 0.102448f
C6 A2 B1_N 4.77e-19
C7 A2 VPWR 0.040335f
C8 VPB Y 0.006363f
C9 VPB VGND 0.011606f
C10 A2 Y 0.07129f
C11 A1 VPWR 0.027531f
C12 B1_N VPWR 0.039714f
C13 A1 Y 0.05697f
C14 A2 VGND 0.062392f
C15 A1 VGND 0.031942f
C16 B1_N Y 0.001426f
C17 VPWR Y 0.010202f
C18 B1_N VGND 0.021488f
C19 VPWR VGND 0.083594f
C20 VGND VNB 0.520551f
C21 Y VNB 0.019872f
C22 VPWR VNB 0.423864f
C23 B1_N VNB 0.244698f
C24 A1 VNB 0.173072f
C25 A2 VNB 0.235098f
C26 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_4 VNB VPB VGND VPWR Y A1 A2 B1_N
X0 a_223_297.t7 A2.t0 VPWR.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y.t3 A1.t0 a_658_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR.t8 B1_N.t0 a_27_47.t0 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3 a_223_297.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X4 Y.t10 a_27_47.t2 VGND.t8 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VGND.t4 A2.t1 a_658_47.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_223_297.t11 a_27_47.t3 Y.t11 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X7 Y.t4 a_27_47.t4 VGND.t7 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.1235 ps=1.03 w=0.65 l=0.15
X8 VPWR.t6 A2.t2 a_223_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_658_47.t6 A2.t3 VGND.t3 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2015 ps=1.27 w=0.65 l=0.15
X10 VPWR.t1 A1.t2 a_223_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_223_297.t2 A1.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_658_47.t5 A2.t4 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 Y.t5 a_27_47.t5 a_223_297.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_223_297.t5 A2.t5 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR.t4 A2.t6 a_223_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X16 VPWR.t3 A1.t4 a_223_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_658_47.t2 A1.t5 Y.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND.t0 B1_N.t1 a_27_47.t1 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.26975 ps=2.13 w=0.65 l=0.15
X19 a_223_297.t9 a_27_47.t6 Y.t6 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_658_47.t1 A1.t6 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 VGND.t1 A2.t7 a_658_47.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 VGND.t6 a_27_47.t7 Y.t7 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VGND.t5 a_27_47.t8 Y.t8 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 Y.t0 A1.t7 a_658_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X25 Y.t9 a_27_47.t9 a_223_297.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 A2.n2 A2.n1 280.188
R1 A2.n1 A2.t6 236.18
R2 A2.n0 A2.t5 212.081
R3 A2.n5 A2.t2 212.081
R4 A2.n3 A2.t0 212.081
R5 A2 A2.n0 164.014
R6 A2.n1 A2.t3 163.881
R7 A2.n4 A2.n2 152
R8 A2.n7 A2.n6 152
R9 A2.n0 A2.t1 139.78
R10 A2.n5 A2.t4 139.78
R11 A2.n3 A2.t7 139.78
R12 A2.n6 A2.n0 40.8975
R13 A2.n4 A2.n3 35.055
R14 A2.n5 A2.n4 27.752
R15 A2.n6 A2.n5 21.9096
R16 A2.n7 A2.n2 6.90844
R17 A2 A2.n7 3.65764
R18 VPWR.n24 VPWR.t8 867.614
R19 VPWR.n8 VPWR.n7 604.463
R20 VPWR.n16 VPWR.n4 598.965
R21 VPWR.n6 VPWR.n5 598.965
R22 VPWR.n10 VPWR.n9 598.965
R23 VPWR.n18 VPWR.n17 34.6358
R24 VPWR.n18 VPWR.n1 34.6358
R25 VPWR.n22 VPWR.n1 34.6358
R26 VPWR.n23 VPWR.n22 34.6358
R27 VPWR.n4 VPWR.t4 29.5505
R28 VPWR.n11 VPWR.n6 28.2358
R29 VPWR.n4 VPWR.t0 27.5805
R30 VPWR.n5 VPWR.t2 27.5805
R31 VPWR.n5 VPWR.t1 27.5805
R32 VPWR.n9 VPWR.t7 27.5805
R33 VPWR.n9 VPWR.t3 27.5805
R34 VPWR.n7 VPWR.t5 27.5805
R35 VPWR.n7 VPWR.t6 27.5805
R36 VPWR.n16 VPWR.n15 23.7181
R37 VPWR.n17 VPWR.n16 20.7064
R38 VPWR.n24 VPWR.n23 19.9534
R39 VPWR.n15 VPWR.n6 16.1887
R40 VPWR.n11 VPWR.n10 11.6711
R41 VPWR.n12 VPWR.n11 9.3005
R42 VPWR.n13 VPWR.n6 9.3005
R43 VPWR.n15 VPWR.n14 9.3005
R44 VPWR.n16 VPWR.n3 9.3005
R45 VPWR.n17 VPWR.n2 9.3005
R46 VPWR.n19 VPWR.n18 9.3005
R47 VPWR.n20 VPWR.n1 9.3005
R48 VPWR.n22 VPWR.n21 9.3005
R49 VPWR.n23 VPWR.n0 9.3005
R50 VPWR.n25 VPWR.n24 7.49328
R51 VPWR.n10 VPWR.n8 6.79
R52 VPWR.n12 VPWR.n8 0.839506
R53 VPWR.n25 VPWR.n0 0.143781
R54 VPWR.n13 VPWR.n12 0.120292
R55 VPWR.n14 VPWR.n13 0.120292
R56 VPWR.n14 VPWR.n3 0.120292
R57 VPWR.n3 VPWR.n2 0.120292
R58 VPWR.n19 VPWR.n2 0.120292
R59 VPWR.n20 VPWR.n19 0.120292
R60 VPWR.n21 VPWR.n20 0.120292
R61 VPWR.n21 VPWR.n0 0.120292
R62 VPWR VPWR.n25 0.119642
R63 a_223_297.n9 a_223_297.n8 598.867
R64 a_223_297.n4 a_223_297.n3 585
R65 a_223_297.n2 a_223_297.n1 585
R66 a_223_297.n6 a_223_297.n5 585
R67 a_223_297.n8 a_223_297.t5 367.079
R68 a_223_297.n2 a_223_297.t8 366.293
R69 a_223_297.n7 a_223_297.n0 295.748
R70 a_223_297.n6 a_223_297.n4 54.7858
R71 a_223_297.n7 a_223_297.n6 47.8614
R72 a_223_297.n8 a_223_297.n7 47.5831
R73 a_223_297.n4 a_223_297.n2 43.8159
R74 a_223_297.n3 a_223_297.t11 33.4905
R75 a_223_297.n5 a_223_297.t1 27.5805
R76 a_223_297.n5 a_223_297.t0 27.5805
R77 a_223_297.n0 a_223_297.t3 27.5805
R78 a_223_297.n0 a_223_297.t2 27.5805
R79 a_223_297.n1 a_223_297.t10 27.5805
R80 a_223_297.n1 a_223_297.t9 27.5805
R81 a_223_297.n3 a_223_297.t4 27.5805
R82 a_223_297.n9 a_223_297.t6 27.5805
R83 a_223_297.t7 a_223_297.n9 27.5805
R84 VPB.t11 VPB.t8 562.306
R85 VPB.t12 VPB.t4 272.274
R86 VPB.t4 VPB.t0 260.437
R87 VPB.t6 VPB.t5 254.518
R88 VPB.t7 VPB.t6 254.518
R89 VPB.t3 VPB.t7 254.518
R90 VPB.t2 VPB.t3 254.518
R91 VPB.t1 VPB.t2 254.518
R92 VPB.t0 VPB.t1 254.518
R93 VPB.t10 VPB.t12 254.518
R94 VPB.t9 VPB.t10 254.518
R95 VPB.t8 VPB.t9 254.518
R96 VPB VPB.t11 213.084
R97 A1.n0 A1.t4 221.72
R98 A1.n3 A1.t3 221.72
R99 A1.n6 A1.t2 221.72
R100 A1.n4 A1.t1 221.72
R101 A1.n5 A1.n2 169.763
R102 A1 A1.n1 154.613
R103 A1.n9 A1.n8 152
R104 A1.n7 A1.n2 152
R105 A1.n0 A1.t5 138.173
R106 A1.n3 A1.t7 138.173
R107 A1.n6 A1.t6 138.173
R108 A1.n4 A1.t0 138.173
R109 A1.n8 A1.n7 53.7316
R110 A1.n6 A1.n5 47.4103
R111 A1.n3 A1.n1 45.83
R112 A1.n1 A1.n0 22.1251
R113 A1.n5 A1.n4 20.5448
R114 A1.n9 A1.n2 17.7638
R115 A1 A1.n9 15.1515
R116 A1.n8 A1.n3 7.90214
R117 A1.n7 A1.n6 6.32181
R118 a_658_47.n4 a_658_47.n3 229.032
R119 a_658_47.n5 a_658_47.n4 185
R120 a_658_47.n2 a_658_47.n0 152.333
R121 a_658_47.n2 a_658_47.n1 88.9685
R122 a_658_47.n4 a_658_47.n2 46.7451
R123 a_658_47.n3 a_658_47.t3 25.8467
R124 a_658_47.n3 a_658_47.t6 25.8467
R125 a_658_47.n1 a_658_47.t4 25.8467
R126 a_658_47.n1 a_658_47.t2 25.8467
R127 a_658_47.n0 a_658_47.t7 25.8467
R128 a_658_47.n0 a_658_47.t5 25.8467
R129 a_658_47.t0 a_658_47.n5 25.8467
R130 a_658_47.n5 a_658_47.t1 25.8467
R131 Y Y.n9 607.044
R132 Y.n8 Y.n7 585
R133 Y.n2 Y.n0 235.036
R134 Y.n5 Y.n4 234.422
R135 Y.n2 Y.n1 185
R136 Y.n5 Y.n3 95.6721
R137 Y.n6 Y.n2 93.1916
R138 Y.n6 Y.n5 53.0406
R139 Y.n9 Y.t6 27.5805
R140 Y.n9 Y.t5 27.5805
R141 Y.n7 Y.t11 27.5805
R142 Y.n7 Y.t9 27.5805
R143 Y.n3 Y.t7 25.8467
R144 Y.n3 Y.t10 25.8467
R145 Y.n4 Y.t8 25.8467
R146 Y.n4 Y.t4 25.8467
R147 Y.n1 Y.t1 25.8467
R148 Y.n1 Y.t3 25.8467
R149 Y.n0 Y.t2 25.8467
R150 Y.n0 Y.t0 25.8467
R151 Y.n8 Y.n6 24.4818
R152 Y Y.n8 2.41828
R153 VNB.t9 VNB.t6 2192.88
R154 VNB.t11 VNB.t8 1509.39
R155 VNB VNB.t11 1366.99
R156 VNB.t5 VNB.t7 1224.6
R157 VNB.t4 VNB.t5 1224.6
R158 VNB.t2 VNB.t4 1224.6
R159 VNB.t0 VNB.t2 1224.6
R160 VNB.t1 VNB.t0 1224.6
R161 VNB.t3 VNB.t1 1224.6
R162 VNB.t6 VNB.t3 1224.6
R163 VNB.t12 VNB.t9 1224.6
R164 VNB.t10 VNB.t12 1224.6
R165 VNB.t8 VNB.t10 1224.6
R166 B1_N.n0 B1_N.t0 241.536
R167 B1_N.n0 B1_N.t1 169.237
R168 B1_N B1_N.n0 161.957
R169 a_27_47.t0 a_27_47.n13 388.997
R170 a_27_47.n2 a_27_47.t3 255.899
R171 a_27_47.n3 a_27_47.t9 212.081
R172 a_27_47.n7 a_27_47.t6 212.081
R173 a_27_47.n10 a_27_47.t5 212.081
R174 a_27_47.n13 a_27_47.t1 186.982
R175 a_27_47.n5 a_27_47.n4 166.04
R176 a_27_47.n12 a_27_47.n11 152
R177 a_27_47.n9 a_27_47.n0 152
R178 a_27_47.n6 a_27_47.n5 152
R179 a_27_47.n11 a_27_47.t4 148.544
R180 a_27_47.n8 a_27_47.t8 139.78
R181 a_27_47.n1 a_27_47.t2 139.78
R182 a_27_47.n2 a_27_47.t7 139.78
R183 a_27_47.n8 a_27_47.n7 43.8187
R184 a_27_47.n11 a_27_47.n10 35.055
R185 a_27_47.n4 a_27_47.n1 32.1338
R186 a_27_47.n3 a_27_47.n2 18.9884
R187 a_27_47.n6 a_27_47.n1 17.5278
R188 a_27_47.n10 a_27_47.n9 14.6066
R189 a_27_47.n5 a_27_47.n0 14.0392
R190 a_27_47.n12 a_27_47.n0 14.0392
R191 a_27_47.n4 a_27_47.n3 11.6853
R192 a_27_47.n13 a_27_47.n12 10.5295
R193 a_27_47.n9 a_27_47.n8 4.38232
R194 a_27_47.n7 a_27_47.n6 1.46111
R195 VGND.n9 VGND.n8 211.947
R196 VGND.n27 VGND.n26 198.964
R197 VGND.n20 VGND.n19 185
R198 VGND.n18 VGND.n17 185
R199 VGND.n1 VGND.n0 185
R200 VGND.n7 VGND.t4 161.159
R201 VGND.n19 VGND.n18 62.7697
R202 VGND.n0 VGND.t0 36.9236
R203 VGND.n11 VGND.n10 34.6358
R204 VGND.n11 VGND.n5 34.6358
R205 VGND.n15 VGND.n5 34.6358
R206 VGND.n16 VGND.n15 34.6358
R207 VGND.n29 VGND.n28 34.6358
R208 VGND.n0 VGND.t7 33.2313
R209 VGND.n25 VGND.n3 32.7349
R210 VGND.n17 VGND.n16 29.2665
R211 VGND.n18 VGND.t3 25.8467
R212 VGND.n19 VGND.t6 25.8467
R213 VGND.n8 VGND.t2 25.8467
R214 VGND.n8 VGND.t1 25.8467
R215 VGND.n26 VGND.t8 25.8467
R216 VGND.n26 VGND.t5 25.8467
R217 VGND.n10 VGND.n9 14.6829
R218 VGND.n31 VGND.n1 14.2651
R219 VGND.n9 VGND.n7 12.5018
R220 VGND.n30 VGND.n29 9.3005
R221 VGND.n28 VGND.n2 9.3005
R222 VGND.n25 VGND.n24 9.3005
R223 VGND.n23 VGND.n3 9.3005
R224 VGND.n22 VGND.n21 9.3005
R225 VGND.n16 VGND.n4 9.3005
R226 VGND.n15 VGND.n14 9.3005
R227 VGND.n13 VGND.n5 9.3005
R228 VGND.n12 VGND.n11 9.3005
R229 VGND.n10 VGND.n6 9.3005
R230 VGND.n29 VGND.n1 8.33968
R231 VGND.n27 VGND.n25 7.90638
R232 VGND.n21 VGND.n20 6.92509
R233 VGND.n20 VGND.n3 2.72837
R234 VGND.n28 VGND.n27 1.88285
R235 VGND.n7 VGND.n6 0.864349
R236 VGND.n21 VGND.n17 0.210336
R237 VGND.n31 VGND.n30 0.141672
R238 VGND VGND.n31 0.121778
R239 VGND.n12 VGND.n6 0.120292
R240 VGND.n13 VGND.n12 0.120292
R241 VGND.n14 VGND.n13 0.120292
R242 VGND.n14 VGND.n4 0.120292
R243 VGND.n22 VGND.n4 0.120292
R244 VGND.n23 VGND.n22 0.120292
R245 VGND.n24 VGND.n23 0.120292
R246 VGND.n24 VGND.n2 0.120292
R247 VGND.n30 VGND.n2 0.120292
C0 A2 Y 0.101573f
C1 A1 VPWR 0.058505f
C2 B1_N VGND 0.015117f
C3 A1 Y 0.143328f
C4 A2 VGND 0.080206f
C5 VPWR Y 0.027628f
C6 A1 VGND 0.035311f
C7 VPWR VGND 0.13556f
C8 Y VGND 0.260291f
C9 VPB B1_N 0.039664f
C10 VPB A2 0.143723f
C11 VPB A1 0.118826f
C12 VPB VPWR 0.140339f
C13 A2 A1 0.29479f
C14 B1_N VPWR 0.01899f
C15 VPB Y 0.007808f
C16 VPB VGND 0.012735f
C17 B1_N Y 6.37e-19
C18 A2 VPWR 0.086093f
C19 VGND VNB 0.788785f
C20 Y VNB 0.019101f
C21 VPWR VNB 0.633685f
C22 A1 VNB 0.356038f
C23 A2 VNB 0.425068f
C24 B1_N VNB 0.145752f
C25 VPB VNB 1.40213f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21.t2 B1.t0 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297.t2 B1.t1 a_81_21.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR.t2 a_81_21.t3 X.t0 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR.t0 A1.t0 a_299_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND.t0 a_81_21.t4 X.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND.t1 A2.t0 a_384_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297.t1 A2.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47.t1 A1.t1 a_81_21.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
R0 B1.n0 B1.t1 230.793
R1 B1.n0 B1.t0 158.494
R2 B1 B1.n0 157.781
R3 VGND.n4 VGND.t1 241.518
R4 VGND.n3 VGND.n2 185
R5 VGND.n1 VGND.n0 185
R6 VGND.n2 VGND.n1 62.7697
R7 VGND.n2 VGND.t2 41.539
R8 VGND.n1 VGND.t0 41.539
R9 VGND.n5 VGND.n0 9.66405
R10 VGND.n3 VGND.n0 8.05976
R11 VGND.n4 VGND.n3 7.96699
R12 VGND.n5 VGND.n4 0.254179
R13 VGND VGND.n5 0.120124
R14 a_81_21.t1 a_81_21.n2 408.337
R15 a_81_21.n2 a_81_21.n0 251.718
R16 a_81_21.n1 a_81_21.t3 230.793
R17 a_81_21.n1 a_81_21.t4 158.494
R18 a_81_21.n2 a_81_21.n1 152
R19 a_81_21.n0 a_81_21.t0 25.8467
R20 a_81_21.n0 a_81_21.t2 24.9236
R21 VNB.t3 VNB.t2 2677.02
R22 VNB.t0 VNB.t1 1224.6
R23 VNB.t2 VNB.t0 1210.36
R24 VNB VNB.t3 954.045
R25 a_299_297.n0 a_299_297.t1 719.394
R26 a_299_297.t0 a_299_297.n0 27.5805
R27 a_299_297.n0 a_299_297.t2 26.5955
R28 VPB.t3 VPB.t2 556.386
R29 VPB.t0 VPB.t1 254.518
R30 VPB.t2 VPB.t0 251.559
R31 VPB VPB.t3 198.287
R32 X.t0 X 759.665
R33 X.n0 X.t0 747.904
R34 X.n1 X.t1 209.923
R35 X X.n0 16.0005
R36 X X.n1 10.0928
R37 X.n1 X 6.64665
R38 X.n0 X 0.738962
R39 VPWR.n1 VPWR.t2 342.221
R40 VPWR.n1 VPWR.n0 315.748
R41 VPWR.n0 VPWR.t1 27.5805
R42 VPWR.n0 VPWR.t0 27.5805
R43 VPWR VPWR.n1 0.213345
R44 A1.n0 A1.t0 241.536
R45 A1.n0 A1.t1 169.237
R46 A1 A1.n0 157.781
R47 A2.n0 A2.t1 231.017
R48 A2.n0 A2.t0 158.716
R49 A2 A2.n0 154.347
R50 a_384_47.t0 a_384_47.t1 51.6928
C0 VPB VGND 0.007132f
C1 B1 VPWR 0.019602f
C2 B1 VGND 0.018138f
C3 A1 VPWR 0.020947f
C4 A2 VPWR 0.020087f
C5 A1 VGND 0.078569f
C6 X VPWR 0.084724f
C7 A2 VGND 0.049499f
C8 X VGND 0.05115f
C9 VPWR VGND 0.057888f
C10 VPB B1 0.038719f
C11 VPB A1 0.026428f
C12 B1 A1 0.081725f
C13 VPB A2 0.03733f
C14 VPB X 0.010847f
C15 A1 A2 0.092059f
C16 VPB VPWR 0.068018f
C17 B1 X 3.04e-20
C18 VGND VNB 0.364132f
C19 VPWR VNB 0.285747f
C20 X VNB 0.094473f
C21 A2 VNB 0.144001f
C22 A1 VNB 0.099647f
C23 B1 VNB 0.108793f
C24 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR.t3 a_80_199.t3 X.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X.t2 a_80_199.t4 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND.t3 a_80_199.t5 X.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X.t0 a_80_199.t6 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199.t0 B1.t0 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297.t1 B1.t1 a_80_199.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47.t1 A1.t0 a_80_199.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR.t1 A1.t1 a_386_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND.t0 A2.t1 a_458_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
R0 a_80_199.t1 a_80_199.n4 361.635
R1 a_80_199.n1 a_80_199.t4 324.548
R2 a_80_199.n4 a_80_199.n0 260.582
R3 a_80_199.n3 a_80_199.t3 231.017
R4 a_80_199.n4 a_80_199.n3 152
R5 a_80_199.n2 a_80_199.t5 148.387
R6 a_80_199.n1 a_80_199.t6 139.78
R7 a_80_199.n0 a_80_199.t2 66.462
R8 a_80_199.n2 a_80_199.n1 59.4472
R9 a_80_199.n0 a_80_199.t0 25.8467
R10 a_80_199.n3 a_80_199.n2 10.3291
R11 X X.n0 594.74
R12 X.n2 X.n0 585
R13 X.n2 X.n1 267.937
R14 X.n0 X.t3 27.5805
R15 X.n0 X.t2 27.5805
R16 X.n1 X.t1 25.8467
R17 X.n1 X.t0 25.8467
R18 X X.n2 16.6962
R19 VPWR.n3 VPWR.t3 863.645
R20 VPWR.n2 VPWR.n1 605.73
R21 VPWR.n5 VPWR.t2 342.214
R22 VPWR.n1 VPWR.t1 31.5205
R23 VPWR.n1 VPWR.t0 30.5355
R24 VPWR.n5 VPWR.n4 22.9652
R25 VPWR.n4 VPWR.n3 19.9534
R26 VPWR.n4 VPWR.n0 9.3005
R27 VPWR.n6 VPWR.n5 9.3005
R28 VPWR.n3 VPWR.n2 7.11182
R29 VPWR.n2 VPWR.n0 0.225794
R30 VPWR.n6 VPWR.n0 0.120292
R31 VPWR VPWR.n6 0.0213333
R32 VPB.t4 VPB.t1 562.306
R33 VPB.t2 VPB.t0 275.235
R34 VPB.t1 VPB.t2 254.518
R35 VPB.t3 VPB.t4 254.518
R36 VPB VPB.t3 192.369
R37 VGND.n1 VGND.t0 288.596
R38 VGND.n5 VGND.t2 281.25
R39 VGND.n3 VGND.n2 198.964
R40 VGND.n2 VGND.t1 36.9236
R41 VGND.n4 VGND.n3 32.7534
R42 VGND.n2 VGND.t3 25.8467
R43 VGND.n6 VGND.n5 11.9358
R44 VGND.n4 VGND.n0 9.3005
R45 VGND.n5 VGND.n4 7.15344
R46 VGND.n3 VGND.n1 6.21844
R47 VGND.n1 VGND.n0 0.191579
R48 VGND.n6 VGND.n0 0.120292
R49 VGND VGND.n6 0.0213333
R50 VNB.t1 VNB.t2 1851.13
R51 VNB.t2 VNB.t0 1509.39
R52 VNB VNB.t3 1409.71
R53 VNB.t4 VNB.t1 1395.47
R54 VNB.t3 VNB.t4 1224.6
R55 A2.n0 A2.t0 236.661
R56 A2.n0 A2.t1 183.829
R57 A2 A2.n0 154.236
R58 a_386_297.t0 a_386_297.n0 664.957
R59 a_386_297.n0 a_386_297.t2 27.5805
R60 a_386_297.n0 a_386_297.t1 27.5805
R61 B1.n0 B1.t1 230.155
R62 B1.n0 B1.t0 157.856
R63 B1 B1.n0 155.856
R64 A1.n0 A1.t1 236.934
R65 A1 A1.n0 165.305
R66 A1.n0 A1.t0 164.633
R67 a_458_47.t0 a_458_47.t1 70.1543
C0 X VGND 0.080574f
C1 VPB B1 0.041674f
C2 VPB A1 0.029009f
C3 VPB A2 0.036695f
C4 B1 A1 0.066922f
C5 B1 A2 1.86e-19
C6 VPB VPWR 0.081424f
C7 B1 VPWR 0.016706f
C8 VPB X 0.006439f
C9 A1 A2 0.104392f
C10 VPB VGND 0.008332f
C11 A1 VPWR 0.020369f
C12 B1 X 8.47e-19
C13 A2 VPWR 0.018943f
C14 B1 VGND 0.015566f
C15 A1 VGND 0.068348f
C16 VPWR X 0.127834f
C17 A2 VGND 0.051922f
C18 VPWR VGND 0.074512f
C19 VGND VNB 0.428053f
C20 X VNB 0.044067f
C21 VPWR VNB 0.356209f
C22 A2 VNB 0.15339f
C23 A1 VNB 0.107801f
C24 B1 VNB 0.110336f
C25 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR.t2 A2.t0 a_109_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297.t1 B1.t0 a_109_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND.t2 A2.t1 a_373_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X.t1 a_27_297.t4 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297.t0 B1.t1 a_109_297.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297.t1 A1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47.t0 A1.t1 a_27_297.t3 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X.t0 a_27_297.t5 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297.t0 B2.t0 a_27_297.t2 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47.t1 B2.t1 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t0 722.096
R1 A2.n0 A2.t1 162.963
R2 A2 A2.n0 162.282
R3 a_109_297.n1 a_109_297.n0 960.074
R4 a_109_297.n0 a_109_297.t3 34.4755
R5 a_109_297.n0 a_109_297.t1 28.5655
R6 a_109_297.n1 a_109_297.t2 26.5955
R7 a_109_297.t0 a_109_297.n1 26.5955
R8 VPWR.n1 VPWR.t0 795.005
R9 VPWR.n1 VPWR.n0 321.094
R10 VPWR.n0 VPWR.t2 34.4755
R11 VPWR.n0 VPWR.t1 26.5955
R12 VPWR VPWR.n1 0.666646
R13 VPB.t3 VPB.t1 550.467
R14 VPB.t1 VPB.t4 278.193
R15 VPB.t4 VPB.t2 272.274
R16 VPB.t0 VPB.t3 248.599
R17 VPB VPB.t0 192.369
R18 B1.n0 B1.t1 239.505
R19 B1.n0 B1.t0 167.204
R20 B1 B1.n0 161.85
R21 a_109_47.t0 a_109_47.t1 42.462
R22 a_27_297.t0 a_27_297.n3 774.126
R23 a_27_297.n0 a_27_297.t1 299.772
R24 a_27_297.n3 a_27_297.t2 289.397
R25 a_27_297.n0 a_27_297.t3 268.077
R26 a_27_297.n1 a_27_297.t4 233.576
R27 a_27_297.n1 a_27_297.t5 161.275
R28 a_27_297.n2 a_27_297.n1 152.892
R29 a_27_297.n3 a_27_297.n2 139.825
R30 a_27_297.n4 a_27_297.t0 110.32
R31 a_27_297.n2 a_27_297.n0 106.153
R32 VNB.t0 VNB.t2 2677.02
R33 VNB.t2 VNB.t4 1423.95
R34 VNB.t4 VNB.t3 1310.03
R35 VNB.t1 VNB.t0 1082.2
R36 VNB VNB.t1 925.567
R37 a_373_47.t0 a_373_47.t1 64.6159
R38 VGND.n1 VGND.n0 205.256
R39 VGND.n1 VGND.t0 151.368
R40 VGND.n0 VGND.t2 32.3082
R41 VGND.n0 VGND.t1 24.9236
R42 VGND VGND.n1 0.0752166
R43 X.n0 X 593.615
R44 X.n1 X.n0 585
R45 X X.t0 348.091
R46 X.n0 X.t1 26.5955
R47 X X.n1 8.61589
R48 X.n1 X 8.12358
R49 A1.n0 A1.t0 256.716
R50 A1.n0 A1.t1 161.275
R51 A1.n1 A1.n0 155.657
R52 A1 A1.n1 18.8957
R53 A1.n1 A1 3.9624
R54 B2.n0 B2.t0 241.536
R55 B2.n0 B2.t1 169.237
R56 B2 B2.n0 168.641
C0 VPWR X 0.09141f
C1 A2 VGND 0.016221f
C2 VPB B2 0.029852f
C3 VPWR VGND 0.064099f
C4 VPB B1 0.03168f
C5 X VGND 0.054267f
C6 B2 B1 0.073857f
C7 VPB A1 0.038674f
C8 VPB A2 0.028389f
C9 B1 A1 0.065706f
C10 VPB VPWR 0.07143f
C11 B2 A2 8.94e-20
C12 B1 A2 1.81e-19
C13 VPB X 0.011018f
C14 B2 VPWR 0.012568f
C15 B2 X 3.26e-20
C16 VPB VGND 0.007463f
C17 A1 A2 0.073773f
C18 B1 VPWR 0.013891f
C19 A1 VPWR 0.016808f
C20 B2 VGND 0.053784f
C21 B1 X 8.38e-20
C22 A2 VPWR 0.017794f
C23 B1 VGND 0.026654f
C24 A1 X 2.98e-19
C25 A1 VGND 0.013674f
C26 A2 X 0.001099f
C27 VGND VNB 0.421193f
C28 X VNB 0.091659f
C29 VPWR VNB 0.328062f
C30 A2 VNB 0.092694f
C31 A1 VNB 0.111912f
C32 B1 VNB 0.111541f
C33 B2 VNB 0.126407f
C34 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_4 VNB VPB VGND VPWR A2 B1 Y A1
X0 a_28_297.t4 B1.t0 Y.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47.t5 A1.t0 Y.t8 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y.t2 B1.t1 a_28_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y.t5 B1.t2 VGND.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47.t4 A1.t1 Y.t9 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297.t6 A2.t0 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47.t7 A2.t1 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y.t1 B1.t3 a_28_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND.t3 B1.t4 Y.t4 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND.t2 B1.t5 Y.t7 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y.t10 A1.t2 a_462_47.t3 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297.t8 A1.t3 VPWR.t7 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR.t2 A2.t2 a_28_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y.t6 B1.t6 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X14 VGND.t5 A2.t3 a_462_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297.t1 B1.t7 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR.t6 A1.t4 a_28_297.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297.t10 A1.t5 VPWR.t5 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND.t0 A2.t4 a_462_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR.t1 A2.t5 a_28_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297.t7 A2.t6 VPWR.t0 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y.t11 A1.t6 a_462_47.t2 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47.t6 A2.t7 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR.t4 A1.t7 a_28_297.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 B1.n0 B1.t7 212.081
R1 B1.n1 B1.t3 212.081
R2 B1.n5 B1.t0 212.081
R3 B1.n3 B1.t1 212.081
R4 B1 B1.n2 158.569
R5 B1.n7 B1.n6 152
R6 B1.n0 B1.t4 139.78
R7 B1.n1 B1.t2 139.78
R8 B1.n5 B1.t5 139.78
R9 B1.n3 B1.t6 139.78
R10 B1.n7 B1.n4 93.4859
R11 B1.n1 B1.n0 62.8066
R12 B1.n5 B1.n4 53.4291
R13 B1.n6 B1.n2 49.6611
R14 B1.n2 B1.n1 10.2247
R15 B1.n4 B1.n3 8.67196
R16 B1 B1.n7 4.88471
R17 B1.n6 B1.n5 2.92171
R18 Y Y.n12 608.894
R19 Y.n11 Y.n10 585
R20 Y.n2 Y.n0 235.036
R21 Y.n5 Y.n4 233.142
R22 Y.n7 Y.n6 186.325
R23 Y.n2 Y.n1 185
R24 Y.n6 Y.n3 185
R25 Y.n9 Y.n2 93.1916
R26 Y.n8 Y.n7 62.5783
R27 Y.n9 Y.n8 31.7798
R28 Y.n12 Y.t3 27.5805
R29 Y.n12 Y.t2 27.5805
R30 Y.n10 Y.t0 27.5805
R31 Y.n10 Y.t1 27.5805
R32 Y.n1 Y.t9 25.8467
R33 Y.n1 Y.t10 25.8467
R34 Y.n0 Y.t8 25.8467
R35 Y.n0 Y.t11 25.8467
R36 Y.n4 Y.t7 25.8467
R37 Y.n4 Y.t6 25.8467
R38 Y.n6 Y.t4 25.8467
R39 Y.n6 Y.t5 25.8467
R40 Y.n11 Y.n9 25.4168
R41 Y.n7 Y.n5 15.8902
R42 Y.n8 Y.n3 2.5605
R43 Y.n5 Y.n3 1.2805
R44 Y Y.n11 0.569389
R45 a_28_297.n3 a_28_297.n2 598.867
R46 a_28_297.n7 a_28_297.n6 585
R47 a_28_297.n9 a_28_297.n8 585
R48 a_28_297.n3 a_28_297.t7 367.079
R49 a_28_297.n8 a_28_297.t3 366.293
R50 a_28_297.n5 a_28_297.n0 295.748
R51 a_28_297.n4 a_28_297.n1 295.748
R52 a_28_297.n7 a_28_297.n5 54.7858
R53 a_28_297.n5 a_28_297.n4 47.8614
R54 a_28_297.n4 a_28_297.n3 47.5831
R55 a_28_297.n8 a_28_297.n7 43.8159
R56 a_28_297.n6 a_28_297.t1 33.4905
R57 a_28_297.n6 a_28_297.t0 27.5805
R58 a_28_297.n0 a_28_297.t9 27.5805
R59 a_28_297.n0 a_28_297.t8 27.5805
R60 a_28_297.n1 a_28_297.t11 27.5805
R61 a_28_297.n1 a_28_297.t10 27.5805
R62 a_28_297.n2 a_28_297.t5 27.5805
R63 a_28_297.n2 a_28_297.t6 27.5805
R64 a_28_297.n9 a_28_297.t2 27.5805
R65 a_28_297.t4 a_28_297.n9 27.5805
R66 VPB.t1 VPB.t0 272.274
R67 VPB.t0 VPB.t8 260.437
R68 VPB.t5 VPB.t7 254.518
R69 VPB.t6 VPB.t5 254.518
R70 VPB.t11 VPB.t6 254.518
R71 VPB.t10 VPB.t11 254.518
R72 VPB.t9 VPB.t10 254.518
R73 VPB.t8 VPB.t9 254.518
R74 VPB.t2 VPB.t1 254.518
R75 VPB.t4 VPB.t2 254.518
R76 VPB.t3 VPB.t4 254.518
R77 VPB VPB.t3 192.369
R78 A1.n1 A1.t7 221.72
R79 A1.n8 A1.t5 221.72
R80 A1.n2 A1.t4 221.72
R81 A1.n3 A1.t3 221.72
R82 A1.n5 A1.n4 169.763
R83 A1.n10 A1.n9 152
R84 A1.n7 A1.n0 152
R85 A1.n6 A1.n5 152
R86 A1.n1 A1.t0 138.173
R87 A1.n8 A1.t6 138.173
R88 A1.n2 A1.t1 138.173
R89 A1.n3 A1.t2 138.173
R90 A1.n7 A1.n6 53.7316
R91 A1.n4 A1.n2 47.4103
R92 A1.n9 A1.n8 45.83
R93 A1.n9 A1.n1 22.1251
R94 A1.n4 A1.n3 20.5448
R95 A1.n10 A1.n0 17.7638
R96 A1.n5 A1.n0 17.7638
R97 A1.n8 A1.n7 7.90214
R98 A1.n6 A1.n2 6.32181
R99 A1 A1.n10 0.784173
R100 a_462_47.n3 a_462_47.n1 229.032
R101 a_462_47.n3 a_462_47.n2 185
R102 a_462_47.n4 a_462_47.n0 152.333
R103 a_462_47.n5 a_462_47.n4 88.9685
R104 a_462_47.n4 a_462_47.n3 46.7451
R105 a_462_47.n1 a_462_47.t3 25.8467
R106 a_462_47.n1 a_462_47.t7 25.8467
R107 a_462_47.n2 a_462_47.t2 25.8467
R108 a_462_47.n2 a_462_47.t4 25.8467
R109 a_462_47.n0 a_462_47.t1 25.8467
R110 a_462_47.n0 a_462_47.t6 25.8467
R111 a_462_47.n5 a_462_47.t0 25.8467
R112 a_462_47.t5 a_462_47.n5 25.8467
R113 VNB.t3 VNB.t11 1338.51
R114 VNB.t10 VNB.t5 1224.6
R115 VNB.t0 VNB.t10 1224.6
R116 VNB.t9 VNB.t0 1224.6
R117 VNB.t6 VNB.t9 1224.6
R118 VNB.t8 VNB.t6 1224.6
R119 VNB.t7 VNB.t8 1224.6
R120 VNB.t11 VNB.t7 1224.6
R121 VNB.t4 VNB.t3 1224.6
R122 VNB.t2 VNB.t4 1224.6
R123 VNB.t1 VNB.t2 1224.6
R124 VNB VNB.t1 925.567
R125 VGND.n8 VGND.n7 211.947
R126 VGND.n17 VGND.n16 201.458
R127 VGND.n21 VGND.n2 198.964
R128 VGND.n6 VGND.t5 160.786
R129 VGND.n23 VGND.t1 148.752
R130 VGND.n10 VGND.n9 34.6358
R131 VGND.n10 VGND.n4 34.6358
R132 VGND.n14 VGND.n4 34.6358
R133 VGND.n15 VGND.n14 34.6358
R134 VGND.n16 VGND.t3 33.2313
R135 VGND.n17 VGND.n15 31.2476
R136 VGND.n7 VGND.t6 25.8467
R137 VGND.n7 VGND.t0 25.8467
R138 VGND.n16 VGND.t7 25.8467
R139 VGND.n2 VGND.t4 25.8467
R140 VGND.n2 VGND.t2 25.8467
R141 VGND.n21 VGND.n1 24.4711
R142 VGND.n22 VGND.n21 19.9534
R143 VGND.n23 VGND.n22 19.9534
R144 VGND.n17 VGND.n1 16.9417
R145 VGND.n8 VGND.n6 16.7917
R146 VGND.n9 VGND.n8 10.1652
R147 VGND.n24 VGND.n23 9.3005
R148 VGND.n22 VGND.n0 9.3005
R149 VGND.n21 VGND.n20 9.3005
R150 VGND.n19 VGND.n1 9.3005
R151 VGND.n18 VGND.n17 9.3005
R152 VGND.n15 VGND.n3 9.3005
R153 VGND.n14 VGND.n13 9.3005
R154 VGND.n12 VGND.n4 9.3005
R155 VGND.n11 VGND.n10 9.3005
R156 VGND.n9 VGND.n5 9.3005
R157 VGND.n6 VGND.n5 1.09207
R158 VGND.n11 VGND.n5 0.120292
R159 VGND.n12 VGND.n11 0.120292
R160 VGND.n13 VGND.n12 0.120292
R161 VGND.n13 VGND.n3 0.120292
R162 VGND.n18 VGND.n3 0.120292
R163 VGND.n19 VGND.n18 0.120292
R164 VGND.n20 VGND.n19 0.120292
R165 VGND.n20 VGND.n0 0.120292
R166 VGND.n24 VGND.n0 0.120292
R167 VGND VGND.n24 0.0213333
R168 A2.n2 A2.n1 280.188
R169 A2.n1 A2.t5 236.18
R170 A2.n0 A2.t6 212.081
R171 A2.n5 A2.t2 212.081
R172 A2.n3 A2.t0 212.081
R173 A2.n1 A2.t1 163.881
R174 A2 A2.n0 162.695
R175 A2.n4 A2.n2 152
R176 A2.n7 A2.n6 152
R177 A2.n0 A2.t3 139.78
R178 A2.n5 A2.t7 139.78
R179 A2.n3 A2.t4 139.78
R180 A2.n6 A2.n0 40.8975
R181 A2.n4 A2.n3 35.055
R182 A2.n5 A2.n4 27.752
R183 A2.n6 A2.n5 21.9096
R184 A2.n7 A2.n2 6.90844
R185 A2 A2.n7 4.97828
R186 VPWR.n7 VPWR.n6 604.183
R187 VPWR.n12 VPWR.n1 598.965
R188 VPWR.n10 VPWR.n3 598.965
R189 VPWR.n5 VPWR.n4 598.965
R190 VPWR.n10 VPWR.n9 32.7534
R191 VPWR.n1 VPWR.t1 29.5505
R192 VPWR.n12 VPWR.n11 28.2358
R193 VPWR.n1 VPWR.t7 27.5805
R194 VPWR.n3 VPWR.t5 27.5805
R195 VPWR.n3 VPWR.t6 27.5805
R196 VPWR.n4 VPWR.t3 27.5805
R197 VPWR.n4 VPWR.t4 27.5805
R198 VPWR.n6 VPWR.t0 27.5805
R199 VPWR.n6 VPWR.t2 27.5805
R200 VPWR.n11 VPWR.n10 11.6711
R201 VPWR.n9 VPWR.n8 9.3005
R202 VPWR.n10 VPWR.n2 9.3005
R203 VPWR.n11 VPWR.n0 9.3005
R204 VPWR.n7 VPWR.n5 9.22973
R205 VPWR.n9 VPWR.n5 7.15344
R206 VPWR.n13 VPWR.n12 6.65763
R207 VPWR.n8 VPWR.n7 1.10236
R208 VPWR VPWR.n13 0.581628
R209 VPWR.n13 VPWR.n0 0.161829
R210 VPWR.n8 VPWR.n2 0.120292
R211 VPWR.n2 VPWR.n0 0.120292
C0 VPB VPWR 0.116188f
C1 B1 Y 0.284714f
C2 A2 A1 0.29568f
C3 B1 VPWR 0.034918f
C4 VPB VGND 0.011278f
C5 A2 Y 0.10137f
C6 B1 VGND 0.106094f
C7 A1 Y 0.143519f
C8 A2 VPWR 0.084484f
C9 A2 VGND 0.079244f
C10 A1 VPWR 0.052519f
C11 Y VPWR 0.027138f
C12 A1 VGND 0.033537f
C13 Y VGND 0.254192f
C14 VPWR VGND 0.118007f
C15 VPB B1 0.139525f
C16 VPB A2 0.144443f
C17 B1 A2 0.052499f
C18 VPB A1 0.118826f
C19 VPB Y 0.007137f
C20 VGND VNB 0.723386f
C21 VPWR VNB 0.557809f
C22 Y VNB 0.031524f
C23 A1 VNB 0.356041f
C24 A2 VNB 0.421609f
C25 B1 VNB 0.426869f
C26 VPB VNB 1.22494f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_2 VNB VPB VGND VPWR A2 A1 Y B1
X0 VGND.t2 A2.t0 a_285_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND.t3 B1.t0 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t4 A1.t0 a_114_47.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47.t1 A2.t1 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297.t3 B1.t1 Y.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297.t0 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y.t0 B1.t2 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR.t3 A2.t2 a_27_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297.t4 A2.t3 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR.t0 A1.t2 a_27_297.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47.t1 A1.t3 Y.t5 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y.t2 B1.t3 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
R0 A2.n1 A2.t2 671.731
R1 A2.n2 A2.n0 241.905
R2 A2.n0 A2.t3 241.536
R3 A2.n0 A2.t0 169.237
R4 A2.n1 A2.t1 167.07
R5 A2.n2 A2.n1 152
R6 A2 A2.n2 5.1005
R7 a_285_47.t0 a_285_47.t1 38.7697
R8 VGND.n3 VGND.n2 198.964
R9 VGND.n4 VGND.t3 168.058
R10 VGND.n9 VGND.t1 137.514
R11 VGND.n2 VGND.t0 35.0774
R12 VGND.n7 VGND.n1 34.6358
R13 VGND.n8 VGND.n7 34.6358
R14 VGND.n2 VGND.t2 25.8467
R15 VGND.n9 VGND.n8 22.2123
R16 VGND.n3 VGND.n1 11.2946
R17 VGND.n10 VGND.n9 9.3005
R18 VGND.n5 VGND.n1 9.3005
R19 VGND.n7 VGND.n6 9.3005
R20 VGND.n8 VGND.n0 9.3005
R21 VGND.n4 VGND.n3 7.11056
R22 VGND.n5 VGND.n4 0.56796
R23 VGND.n6 VGND.n5 0.120292
R24 VGND.n6 VGND.n0 0.120292
R25 VGND.n10 VGND.n0 0.120292
R26 VGND VGND.n10 0.0226354
R27 VNB.t2 VNB.t0 1366.99
R28 VNB.t4 VNB.t5 1224.6
R29 VNB.t1 VNB.t4 1210.36
R30 VNB.t0 VNB.t3 1196.12
R31 VNB.t5 VNB.t2 1025.24
R32 VNB VNB.t1 996.764
R33 B1.n1 B1.t1 218.507
R34 B1.n0 B1.t2 218.507
R35 B1.n2 B1.n1 208.511
R36 B1.n1 B1.t0 146.208
R37 B1.n0 B1.t3 146.208
R38 B1.n1 B1.n0 69.8074
R39 B1.n2 B1 13.266
R40 B1 B1.n2 2.5605
R41 Y.n3 Y.n2 332.284
R42 Y Y.n4 185.201
R43 Y.n4 Y.n3 185
R44 Y.n1 Y.n0 170.469
R45 Y.n2 Y.t1 26.5955
R46 Y.n2 Y.t0 26.5955
R47 Y.n0 Y.t5 25.8467
R48 Y.n0 Y.t4 25.8467
R49 Y.n4 Y.t3 24.9236
R50 Y.n4 Y.t2 24.9236
R51 Y Y.n1 11.0005
R52 Y.n3 Y.n1 2.4005
R53 A1.n0 A1.t2 212.081
R54 A1.n1 A1.t1 212.081
R55 A1.n0 A1.t3 139.78
R56 A1.n1 A1.t0 139.78
R57 A1 A1.n2 68.5511
R58 A1.n2 A1.n0 30.5224
R59 A1.n2 A1.n1 25.563
R60 a_114_47.t0 a_114_47.t1 50.7697
R61 a_27_297.t3 a_27_297.n3 398.082
R62 a_27_297.n1 a_27_297.t5 363.389
R63 a_27_297.n1 a_27_297.n0 296.125
R64 a_27_297.n3 a_27_297.n2 289.24
R65 a_27_297.n3 a_27_297.n1 58.7765
R66 a_27_297.n0 a_27_297.t1 27.5805
R67 a_27_297.n0 a_27_297.t0 27.5805
R68 a_27_297.n2 a_27_297.t2 26.5955
R69 a_27_297.n2 a_27_297.t4 26.5955
R70 VPB.t1 VPB.t0 254.518
R71 VPB.t5 VPB.t1 254.518
R72 VPB.t2 VPB.t3 248.599
R73 VPB.t4 VPB.t2 248.599
R74 VPB.t0 VPB.t4 248.599
R75 VPB VPB.t5 204.207
R76 VPWR.n2 VPWR.n0 614.221
R77 VPWR.n2 VPWR.n1 604.294
R78 VPWR.n1 VPWR.t1 27.5805
R79 VPWR.n1 VPWR.t3 27.5805
R80 VPWR.n0 VPWR.t2 26.5955
R81 VPWR.n0 VPWR.t0 26.5955
R82 VPWR VPWR.n2 0.560285
C0 VPB Y 0.005049f
C1 A1 B1 2.94e-19
C2 A2 VPWR 0.042572f
C3 VPB VGND 0.007263f
C4 A1 VPWR 0.028734f
C5 A2 Y 0.071413f
C6 B1 VPWR 0.017987f
C7 A2 VGND 0.071822f
C8 A1 Y 0.058671f
C9 B1 Y 0.117296f
C10 A1 VGND 0.031725f
C11 B1 VGND 0.059494f
C12 VPWR Y 0.01257f
C13 VPWR VGND 0.064971f
C14 Y VGND 0.251472f
C15 VPB A2 0.069044f
C16 VPB A1 0.053858f
C17 VPB B1 0.07973f
C18 A2 A1 0.22587f
C19 A2 B1 0.059508f
C20 VPB VPWR 0.066122f
C21 VGND VNB 0.443841f
C22 Y VNB 0.029544f
C23 VPWR VNB 0.326032f
C24 B1 VNB 0.258529f
C25 A1 VNB 0.172911f
C26 A2 VNB 0.23941f
C27 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22oi_2 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 a_109_297.t1 A2.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47.t3 A1.t0 Y.t3 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t0 A2.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47.t1 A2.t2 VGND.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y.t0 B1.t0 a_109_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y.t4 A1.t1 a_467_47.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297.t7 B1.t1 Y.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t0 A2.t3 a_467_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t1 B2.t0 a_109_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47.t1 B2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47.t3 B1.t2 Y.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297.t5 A1.t2 VPWR.t2 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR.t3 A1.t3 a_109_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y.t5 B1.t3 a_27_47.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_297.t4 B2.t2 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t3 B2.t3 a_27_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t0 212.081
R1 A2.n1 A2.t1 212.081
R2 A2.n3 A2.n2 152
R3 A2.n0 A2.t2 139.78
R4 A2.n1 A2.t3 139.78
R5 A2.n2 A2.n0 48.2005
R6 A2 A2.n3 16.0005
R7 A2.n3 A2 13.4405
R8 A2.n2 A2.n1 13.146
R9 VPWR.n5 VPWR.n4 332.697
R10 VPWR.n6 VPWR.n3 320.976
R11 VPWR.n14 VPWR 37.9123
R12 VPWR.n8 VPWR.n7 34.6358
R13 VPWR.n8 VPWR.n1 34.6358
R14 VPWR.n12 VPWR.n1 34.6358
R15 VPWR.n13 VPWR.n12 34.6358
R16 VPWR.n3 VPWR.t2 26.5955
R17 VPWR.n3 VPWR.t3 26.5955
R18 VPWR.n4 VPWR.t1 26.5955
R19 VPWR.n4 VPWR.t0 26.5955
R20 VPWR.n7 VPWR.n6 26.3534
R21 VPWR.n6 VPWR.n5 15.1733
R22 VPWR.n7 VPWR.n2 9.3005
R23 VPWR.n9 VPWR.n8 9.3005
R24 VPWR.n10 VPWR.n1 9.3005
R25 VPWR.n12 VPWR.n11 9.3005
R26 VPWR.n13 VPWR.n0 9.3005
R27 VPWR VPWR.n13 6.02403
R28 VPWR.n5 VPWR.n2 0.857451
R29 VPWR.n9 VPWR.n2 0.120292
R30 VPWR.n10 VPWR.n9 0.120292
R31 VPWR.n11 VPWR.n10 0.120292
R32 VPWR.n11 VPWR.n0 0.120292
R33 VPWR.n14 VPWR.n0 0.120292
R34 VPWR VPWR.n14 0.0213333
R35 a_109_297.n2 a_109_297.n1 355.683
R36 a_109_297.n2 a_109_297.n0 297.95
R37 a_109_297.t1 a_109_297.n5 270.663
R38 a_109_297.n3 a_109_297.t6 214.101
R39 a_109_297.n5 a_109_297.n4 205.668
R40 a_109_297.n3 a_109_297.n2 83.3307
R41 a_109_297.n5 a_109_297.n3 59.9146
R42 a_109_297.n0 a_109_297.t2 26.5955
R43 a_109_297.n0 a_109_297.t7 26.5955
R44 a_109_297.n1 a_109_297.t3 26.5955
R45 a_109_297.n1 a_109_297.t4 26.5955
R46 a_109_297.n4 a_109_297.t0 26.5955
R47 a_109_297.n4 a_109_297.t5 26.5955
R48 VPB.t2 VPB.t6 556.386
R49 VPB.t0 VPB.t1 248.599
R50 VPB.t5 VPB.t0 248.599
R51 VPB.t6 VPB.t5 248.599
R52 VPB.t7 VPB.t2 248.599
R53 VPB.t3 VPB.t7 248.599
R54 VPB.t4 VPB.t3 248.599
R55 VPB VPB.t4 189.409
R56 A1.n0 A1.t2 212.081
R57 A1.n1 A1.t3 212.081
R58 A1.n2 A1.n1 160.764
R59 A1.n0 A1.t0 139.78
R60 A1.n1 A1.t1 139.78
R61 A1.n1 A1.n0 61.346
R62 A1 A1.n2 20.4805
R63 A1.n2 A1 8.9605
R64 Y.n4 Y.t2 417.452
R65 Y.n5 Y.t0 319.837
R66 Y.n4 Y.n3 299.252
R67 Y.n2 Y.n1 239.213
R68 Y.n2 Y.n0 211.353
R69 Y.n6 Y.n4 38.4005
R70 Y.n3 Y.t6 26.5955
R71 Y.n3 Y.t1 26.5955
R72 Y.n1 Y.t3 24.9236
R73 Y.n1 Y.t4 24.9236
R74 Y.n0 Y.t7 24.9236
R75 Y.n0 Y.t5 24.9236
R76 Y.n6 Y.n5 5.05125
R77 Y.n7 Y.n6 2.82647
R78 Y.n5 Y 2.08419
R79 Y.n7 Y 1.76602
R80 Y Y.n7 1.33037
R81 Y Y.n2 0.22119
R82 a_467_47.t2 a_467_47.n1 297.517
R83 a_467_47.n1 a_467_47.t1 282.853
R84 a_467_47.n1 a_467_47.n0 185
R85 a_467_47.n0 a_467_47.t0 24.9236
R86 a_467_47.n0 a_467_47.t3 24.9236
R87 VNB.t7 VNB.t3 2677.02
R88 VNB.t0 VNB.t1 1196.12
R89 VNB.t4 VNB.t0 1196.12
R90 VNB.t3 VNB.t4 1196.12
R91 VNB.t5 VNB.t7 1196.12
R92 VNB.t2 VNB.t5 1196.12
R93 VNB.t6 VNB.t2 1196.12
R94 VNB VNB.t6 911.327
R95 VGND.n3 VGND.n0 207.178
R96 VGND.n2 VGND.n1 200.516
R97 VGND.n1 VGND.t2 24.9236
R98 VGND.n1 VGND.t3 24.9236
R99 VGND.n0 VGND.t1 24.9236
R100 VGND.n0 VGND.t0 24.9236
R101 VGND.n3 VGND.n2 5.74908
R102 VGND.n2 VGND 3.29747
R103 VGND VGND.n3 0.146863
R104 B1.n0 B1.t0 212.081
R105 B1.n1 B1.t1 212.081
R106 B1.n3 B1.n2 152
R107 B1.n0 B1.t2 139.78
R108 B1.n1 B1.t3 139.78
R109 B1.n2 B1.n0 48.2005
R110 B1 B1.n3 21.1205
R111 B1.n2 B1.n1 13.146
R112 B1.n3 B1 8.3205
R113 B2.n0 B2.t0 212.081
R114 B2.n1 B2.t2 212.081
R115 B2.n2 B2.n1 160.764
R116 B2.n0 B2.t1 139.78
R117 B2.n1 B2.t3 139.78
R118 B2.n1 B2.n0 61.346
R119 B2 B2.n2 16.6405
R120 B2.n2 B2 12.8005
R121 a_27_47.n0 a_27_47.t3 297.517
R122 a_27_47.n0 a_27_47.t0 285.036
R123 a_27_47.n1 a_27_47.n0 185
R124 a_27_47.n1 a_27_47.t2 24.9236
R125 a_27_47.t1 a_27_47.n1 24.9236
C0 A2 VPWR 0.029794f
C1 A1 VGND 0.01849f
C2 Y VPWR 0.061068f
C3 A2 VGND 0.031595f
C4 VPB B2 0.061652f
C5 Y VGND 0.030561f
C6 VPB B1 0.057421f
C7 VPWR VGND 0.087423f
C8 B2 B1 0.065715f
C9 VPB A1 0.062991f
C10 VPB A2 0.06193f
C11 VPB Y 0.02733f
C12 B1 A1 0.018686f
C13 B2 Y 0.080261f
C14 VPB VPWR 0.094878f
C15 A1 A2 0.0637f
C16 VPB VGND 0.011121f
C17 B1 Y 0.141728f
C18 B2 VPWR 0.020367f
C19 B2 VGND 0.033658f
C20 A1 Y 0.072036f
C21 B1 VPWR 0.016371f
C22 B1 VGND 0.01814f
C23 A2 Y 0.001108f
C24 A1 VPWR 0.030763f
C25 VGND VNB 0.533379f
C26 VPWR VNB 0.449025f
C27 Y VNB 0.07338f
C28 A2 VNB 0.2108f
C29 A1 VNB 0.191157f
C30 B1 VNB 0.179572f
C31 B2 VNB 0.217478f
C32 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 Y.t2 B1.t0 a_109_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1 Y.t1 B1.t1 a_109_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t1 A2.t0 a_109_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297.t2 A1.t0 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47.t0 A1.t1 Y.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297.t0 B2.t0 Y.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47.t1 B2.t1 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND.t1 A2.t1 a_381_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
R0 B1.n0 B1.t1 239.505
R1 B1.n0 B1.t0 167.204
R2 B1 B1.n0 159.424
R3 a_109_47.t0 a_109_47.t1 42.462
R4 Y.n2 Y.t1 916.889
R5 Y.n0 Y.t2 278.288
R6 Y.n0 Y.t3 249.615
R7 Y.n2 Y.t0 215.875
R8 Y.n1 Y.n0 192.98
R9 Y Y.n3 78.5783
R10 Y.n3 Y.n2 17.7469
R11 Y Y.n1 6.04494
R12 Y.n1 Y 4.94595
R13 Y.n3 Y 3.49141
R14 VNB.t0 VNB.t3 2790.94
R15 VNB.t2 VNB.t0 1082.2
R16 VNB.t3 VNB.t1 1025.24
R17 VNB VNB.t2 911.327
R18 a_109_297.n1 a_109_297.n0 1243.69
R19 a_109_297.n0 a_109_297.t3 26.5955
R20 a_109_297.n0 a_109_297.t2 26.5955
R21 a_109_297.n1 a_109_297.t1 26.5955
R22 a_109_297.t0 a_109_297.n1 26.5955
R23 VPB.t1 VPB.t2 556.386
R24 VPB.t2 VPB.t3 248.599
R25 VPB.t0 VPB.t1 248.599
R26 VPB VPB.t0 189.409
R27 A2.n0 A2.t0 241.536
R28 A2.n0 A2.t1 169.237
R29 A2 A2.n0 161.31
R30 VPWR.n0 VPWR.t0 872.039
R31 VPWR.n0 VPWR.t1 347.286
R32 VPWR VPWR.n0 0.826376
R33 A1.n0 A1.t0 232.738
R34 A1.n0 A1.t1 160.438
R35 A1 A1.n0 155.352
R36 a_381_47.t0 a_381_47.t1 38.7697
R37 B2.n0 B2.t0 241.536
R38 B2.n0 B2.t1 169.237
R39 B2 B2.n0 158.525
R40 VGND.n0 VGND.t1 245.642
R41 VGND.n0 VGND.t0 230.584
R42 VGND VGND.n0 0.0752964
C0 VPB VPWR 0.068173f
C1 B2 Y 0.06212f
C2 B1 A2 1.75e-19
C3 B2 VPWR 0.008709f
C4 A1 A2 0.08596f
C5 B1 Y 0.093024f
C6 VPB VGND 0.007244f
C7 B2 VGND 0.057276f
C8 B1 VPWR 0.009634f
C9 A1 Y 0.094336f
C10 A2 Y 0.110184f
C11 B1 VGND 0.01766f
C12 A1 VPWR 0.017432f
C13 A2 VPWR 0.022438f
C14 A1 VGND 0.013245f
C15 Y VPWR 0.200418f
C16 A2 VGND 0.015611f
C17 VPB B2 0.029596f
C18 Y VGND 0.244976f
C19 VPB B1 0.032023f
C20 VPWR VGND 0.054941f
C21 VPB A1 0.036289f
C22 B2 B1 0.089809f
C23 VPB A2 0.030148f
C24 B2 A2 8.37e-20
C25 B1 A1 0.063097f
C26 VPB Y 0.030249f
C27 VGND VNB 0.375267f
C28 VPWR VNB 0.30925f
C29 Y VNB 0.112408f
C30 A2 VNB 0.117076f
C31 A1 VNB 0.110245f
C32 B1 VNB 0.107307f
C33 B2 VNB 0.139677f
C34 VPB VNB 0.604764f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_4 VNB VPB VGND VPWR X B2 A1 A2 B1
X0 a_484_297.t3 B2.t0 a_96_21.t5 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t2 B2.t1 a_566_47.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X.t7 a_96_21.t8 VGND.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t6 a_96_21.t9 X.t3 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 X.t2 a_96_21.t10 VPWR.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_96_21.t7 B1.t0 a_484_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR.t4 a_96_21.t11 X.t1 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t6 a_96_21.t12 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND.t4 a_96_21.t13 X.t5 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_484_297.t1 B1.t1 a_96_21.t3 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_484_297.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND.t7 A2.t1 a_918_47.t3 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_96_21.t4 B2.t2 a_484_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_96_21.t0 B1.t2 a_566_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_484_297.t4 A1.t0 VPWR.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR.t2 A1.t1 a_484_297.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_96_21.t6 A1.t2 a_918_47.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR.t7 A2.t2 a_484_297.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_566_47.t2 B2.t3 VGND.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X19 a_918_47.t0 A1.t3 a_96_21.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_566_47.t1 B1.t3 a_96_21.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_918_47.t2 A2.t3 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X22 X.t0 a_96_21.t14 VPWR.t3 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND.t3 a_96_21.t15 X.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 B2.n1 B2.t2 241.536
R1 B2.n0 B2.t0 241.536
R2 B2.n2 B2.n0 238.481
R3 B2.n1 B2.t3 169.237
R4 B2.n0 B2.t1 169.237
R5 B2.n2 B2.n1 152
R6 B2 B2.n2 6.87457
R7 a_96_21.n16 a_96_21.n0 638.836
R8 a_96_21.n17 a_96_21.n16 585
R9 a_96_21.n14 a_96_21.n12 306.31
R10 a_96_21.n2 a_96_21.t9 212.081
R11 a_96_21.n9 a_96_21.t10 212.081
R12 a_96_21.n3 a_96_21.t11 212.081
R13 a_96_21.n4 a_96_21.t14 212.081
R14 a_96_21.n14 a_96_21.n13 185
R15 a_96_21.n6 a_96_21.n5 173.761
R16 a_96_21.n7 a_96_21.n6 152
R17 a_96_21.n8 a_96_21.n1 152
R18 a_96_21.n11 a_96_21.n10 152
R19 a_96_21.n2 a_96_21.t13 139.78
R20 a_96_21.n9 a_96_21.t8 139.78
R21 a_96_21.n3 a_96_21.t15 139.78
R22 a_96_21.n4 a_96_21.t12 139.78
R23 a_96_21.n15 a_96_21.n14 96.4955
R24 a_96_21.n16 a_96_21.n15 77.5934
R25 a_96_21.n8 a_96_21.n7 49.6611
R26 a_96_21.n10 a_96_21.n9 48.2005
R27 a_96_21.n5 a_96_21.n3 39.4369
R28 a_96_21.n0 a_96_21.t5 26.5955
R29 a_96_21.n0 a_96_21.t7 26.5955
R30 a_96_21.t3 a_96_21.n17 26.5955
R31 a_96_21.n17 a_96_21.t4 26.5955
R32 a_96_21.n13 a_96_21.t1 24.9236
R33 a_96_21.n13 a_96_21.t0 24.9236
R34 a_96_21.n12 a_96_21.t2 24.9236
R35 a_96_21.n12 a_96_21.t6 24.9236
R36 a_96_21.n5 a_96_21.n4 21.9096
R37 a_96_21.n11 a_96_21.n1 21.7605
R38 a_96_21.n6 a_96_21.n1 21.7605
R39 a_96_21.n10 a_96_21.n2 13.146
R40 a_96_21.n15 a_96_21.n11 11.2005
R41 a_96_21.n7 a_96_21.n3 10.2247
R42 a_96_21.n9 a_96_21.n8 1.46111
R43 a_484_297.n3 a_484_297.t2 877.509
R44 a_484_297.n3 a_484_297.n2 585
R45 a_484_297.n1 a_484_297.n0 301.397
R46 a_484_297.n5 a_484_297.n4 289.24
R47 a_484_297.n1 a_484_297.t0 276.938
R48 a_484_297.n4 a_484_297.n3 58.7539
R49 a_484_297.n4 a_484_297.n1 54.4359
R50 a_484_297.n5 a_484_297.t7 35.4605
R51 a_484_297.t3 a_484_297.n5 33.4905
R52 a_484_297.n2 a_484_297.t5 26.5955
R53 a_484_297.n2 a_484_297.t1 26.5955
R54 a_484_297.n0 a_484_297.t6 26.5955
R55 a_484_297.n0 a_484_297.t4 26.5955
R56 VPB.t10 VPB.t2 556.386
R57 VPB.t3 VPB.t11 295.95
R58 VPB.t6 VPB.t0 248.599
R59 VPB.t4 VPB.t6 248.599
R60 VPB.t11 VPB.t4 248.599
R61 VPB.t5 VPB.t3 248.599
R62 VPB.t1 VPB.t5 248.599
R63 VPB.t2 VPB.t1 248.599
R64 VPB.t9 VPB.t10 248.599
R65 VPB.t8 VPB.t9 248.599
R66 VPB.t7 VPB.t8 248.599
R67 VPB VPB.t7 242.679
R68 a_566_47.n1 a_566_47.n0 418.873
R69 a_566_47.n0 a_566_47.t3 24.9236
R70 a_566_47.n0 a_566_47.t1 24.9236
R71 a_566_47.t0 a_566_47.n1 24.9236
R72 a_566_47.n1 a_566_47.t2 24.9236
R73 VGND.n25 VGND.t5 280.822
R74 VGND.n9 VGND.n7 207.965
R75 VGND.n2 VGND.n1 207.965
R76 VGND.n19 VGND.n18 185
R77 VGND.n17 VGND.n16 185
R78 VGND.n8 VGND.t7 173.998
R79 VGND.n18 VGND.n17 96.0005
R80 VGND.n11 VGND.n10 34.6358
R81 VGND.n11 VGND.n5 34.6358
R82 VGND.n24 VGND.n23 34.6358
R83 VGND.n7 VGND.t2 33.2313
R84 VGND.n20 VGND.n2 32.0005
R85 VGND.n7 VGND.t0 31.3851
R86 VGND.n16 VGND.n5 28.8064
R87 VGND.n10 VGND.n9 27.1064
R88 VGND.n20 VGND.n19 26.5476
R89 VGND.n25 VGND.n24 25.977
R90 VGND.n17 VGND.t1 24.9236
R91 VGND.n18 VGND.t4 24.9236
R92 VGND.n1 VGND.t6 24.9236
R93 VGND.n1 VGND.t3 24.9236
R94 VGND.n26 VGND.n25 17.9593
R95 VGND.n9 VGND.n8 15.1039
R96 VGND.n24 VGND.n0 9.3005
R97 VGND.n23 VGND.n22 9.3005
R98 VGND.n21 VGND.n20 9.3005
R99 VGND.n4 VGND.n3 9.3005
R100 VGND.n15 VGND.n14 9.3005
R101 VGND.n10 VGND.n6 9.3005
R102 VGND.n12 VGND.n11 9.3005
R103 VGND.n13 VGND.n5 9.3005
R104 VGND.n15 VGND.n4 9.2005
R105 VGND.n23 VGND.n2 2.63579
R106 VGND.n19 VGND.n4 0.9005
R107 VGND.n16 VGND.n15 0.3005
R108 VGND.n8 VGND.n6 0.173777
R109 VGND.n12 VGND.n6 0.120292
R110 VGND.n13 VGND.n12 0.120292
R111 VGND.n14 VGND.n13 0.120292
R112 VGND.n14 VGND.n3 0.120292
R113 VGND.n21 VGND.n3 0.120292
R114 VGND.n22 VGND.n21 0.120292
R115 VGND.n22 VGND.n0 0.120292
R116 VGND.n26 VGND.n0 0.120292
R117 VGND VGND.n26 0.0226354
R118 VNB.t8 VNB.t4 2677.02
R119 VNB.t5 VNB.t2 1423.95
R120 VNB.t3 VNB.t11 1196.12
R121 VNB.t6 VNB.t3 1196.12
R122 VNB.t2 VNB.t6 1196.12
R123 VNB.t1 VNB.t5 1196.12
R124 VNB.t0 VNB.t1 1196.12
R125 VNB.t4 VNB.t0 1196.12
R126 VNB.t10 VNB.t8 1196.12
R127 VNB.t7 VNB.t10 1196.12
R128 VNB.t9 VNB.t7 1196.12
R129 VNB VNB.t9 1167.64
R130 X.n2 X.n0 253.444
R131 X.n2 X.n1 209.02
R132 X.n5 X.n3 135.249
R133 X.n5 X.n4 98.982
R134 X X.n2 39.4176
R135 X X.n5 29.3806
R136 X.n0 X.t3 26.5955
R137 X.n0 X.t2 26.5955
R138 X.n1 X.t1 26.5955
R139 X.n1 X.t0 26.5955
R140 X.n3 X.t5 24.9236
R141 X.n3 X.t7 24.9236
R142 X.n4 X.t4 24.9236
R143 X.n4 X.t6 24.9236
R144 VPWR.n3 VPWR.t6 845.178
R145 VPWR.n7 VPWR.n6 613.389
R146 VPWR.n9 VPWR.n8 606.505
R147 VPWR.n23 VPWR.t3 343.351
R148 VPWR.n21 VPWR.n2 316.757
R149 VPWR.n10 VPWR.n5 34.6358
R150 VPWR.n14 VPWR.n5 34.6358
R151 VPWR.n15 VPWR.n14 34.6358
R152 VPWR.n16 VPWR.n15 34.6358
R153 VPWR.n16 VPWR.n3 28.6123
R154 VPWR.n22 VPWR.n21 27.8593
R155 VPWR.n2 VPWR.t5 26.5955
R156 VPWR.n2 VPWR.t4 26.5955
R157 VPWR.n8 VPWR.t1 26.5955
R158 VPWR.n8 VPWR.t7 26.5955
R159 VPWR.n6 VPWR.t0 26.5955
R160 VPWR.n6 VPWR.t2 26.5955
R161 VPWR.n21 VPWR.n20 22.5887
R162 VPWR.n20 VPWR.n3 21.8358
R163 VPWR.n10 VPWR.n9 17.3181
R164 VPWR.n23 VPWR.n22 16.5652
R165 VPWR.n11 VPWR.n10 9.3005
R166 VPWR.n12 VPWR.n5 9.3005
R167 VPWR.n14 VPWR.n13 9.3005
R168 VPWR.n15 VPWR.n4 9.3005
R169 VPWR.n17 VPWR.n16 9.3005
R170 VPWR.n18 VPWR.n3 9.3005
R171 VPWR.n20 VPWR.n19 9.3005
R172 VPWR.n21 VPWR.n1 9.3005
R173 VPWR.n22 VPWR.n0 9.3005
R174 VPWR.n24 VPWR.n23 9.3005
R175 VPWR.n9 VPWR.n7 6.86355
R176 VPWR.n11 VPWR.n7 0.801108
R177 VPWR.n12 VPWR.n11 0.120292
R178 VPWR.n13 VPWR.n12 0.120292
R179 VPWR.n13 VPWR.n4 0.120292
R180 VPWR.n17 VPWR.n4 0.120292
R181 VPWR.n18 VPWR.n17 0.120292
R182 VPWR.n19 VPWR.n18 0.120292
R183 VPWR.n19 VPWR.n1 0.120292
R184 VPWR.n1 VPWR.n0 0.120292
R185 VPWR.n24 VPWR.n0 0.120292
R186 VPWR VPWR.n24 0.0226354
R187 B1.n0 B1.t0 212.081
R188 B1.n1 B1.t1 212.081
R189 B1 B1.n2 153.268
R190 B1.n0 B1.t3 139.78
R191 B1.n1 B1.t2 139.78
R192 B1.n2 B1.n0 30.6732
R193 B1.n2 B1.n1 30.6732
R194 A2.n2 A2.n0 260.188
R195 A2.n1 A2.t0 241.536
R196 A2.n0 A2.t2 241.536
R197 A2.n1 A2.t1 169.237
R198 A2.n0 A2.t3 169.237
R199 A2.n2 A2.n1 152
R200 A2 A2.n2 22.4005
R201 a_918_47.n1 a_918_47.n0 326.865
R202 a_918_47.n0 a_918_47.t3 24.9236
R203 a_918_47.n0 a_918_47.t0 24.9236
R204 a_918_47.n1 a_918_47.t1 24.9236
R205 a_918_47.t2 a_918_47.n1 24.9236
R206 A1.n0 A1.t1 212.081
R207 A1.n1 A1.t0 212.081
R208 A1 A1.n2 157.12
R209 A1.n0 A1.t3 139.78
R210 A1.n1 A1.t2 139.78
R211 A1.n2 A1.n0 30.6732
R212 A1.n2 A1.n1 30.6732
C0 A2 VPWR 0.045362f
C1 B2 VGND 0.032502f
C2 B1 X 2.22e-19
C3 B1 VGND 0.018255f
C4 A1 VPWR 0.029506f
C5 A2 X 3.03e-20
C6 A2 VGND 0.056173f
C7 A1 X 4.1e-20
C8 A1 VGND 0.01734f
C9 VPWR X 0.335103f
C10 VPB B2 0.066686f
C11 VPWR VGND 0.12676f
C12 VPB B1 0.050999f
C13 X VGND 0.265017f
C14 B2 B1 0.212706f
C15 VPB A2 0.070993f
C16 B2 A2 0.092645f
C17 VPB A1 0.050973f
C18 VPB VPWR 0.138504f
C19 B2 VPWR 0.023285f
C20 VPB X 0.015145f
C21 A2 A1 0.207246f
C22 VPB VGND 0.01099f
C23 B1 VPWR 0.015596f
C24 B2 X 7.6e-19
C25 VGND VNB 0.758061f
C26 X VNB 0.060097f
C27 VPWR VNB 0.613178f
C28 A1 VNB 0.166288f
C29 A2 VNB 0.230172f
C30 B1 VNB 0.166404f
C31 B2 VNB 0.193215f
C32 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_2 VPWR VGND VPB VNB B2 B1 A1 A2 X
X0 VPWR.t3 a_27_297.t4 X.t1 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND.t0 A2.t0 a_381_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X.t3 a_27_297.t5 VGND.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X3 X.t0 a_27_297.t6 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X4 a_27_297.t1 B1.t0 a_109_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5 a_27_297.t3 B1.t1 a_109_297.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND.t2 a_27_297.t7 X.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_109_297.t3 A1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR.t0 A2.t1 a_109_297.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9 a_381_47.t1 A1.t1 a_27_297.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_109_297.t0 B2.t0 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_109_47.t1 B2.t1 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
R0 a_27_297.n4 a_27_297.t3 916.889
R1 a_27_297.n0 a_27_297.t1 278.288
R2 a_27_297.n0 a_27_297.t2 249.615
R3 a_27_297.t0 a_27_297.n4 215.875
R4 a_27_297.n4 a_27_297.n3 213.317
R5 a_27_297.n1 a_27_297.t4 212.081
R6 a_27_297.n2 a_27_297.t6 212.081
R7 a_27_297.n3 a_27_297.n2 158.573
R8 a_27_297.n1 a_27_297.t7 139.78
R9 a_27_297.n2 a_27_297.t5 139.78
R10 a_27_297.n3 a_27_297.n0 109.493
R11 a_27_297.n2 a_27_297.n1 61.346
R12 X.n1 X 593.615
R13 X.n2 X.n1 585
R14 X X.n0 283.476
R15 X.n1 X.t1 26.5955
R16 X.n1 X.t0 26.5955
R17 X.n0 X.t2 24.9236
R18 X.n0 X.t3 24.9236
R19 X X.n2 8.61589
R20 X.n2 X 8.12358
R21 VPWR.n5 VPWR.t1 838.817
R22 VPWR.n3 VPWR.n1 312.053
R23 VPWR.n2 VPWR.t3 270.457
R24 VPWR.n1 VPWR.t0 35.4605
R25 VPWR.n1 VPWR.t2 26.5955
R26 VPWR.n4 VPWR.n3 24.8476
R27 VPWR.n5 VPWR.n4 19.577
R28 VPWR.n4 VPWR.n0 9.3005
R29 VPWR.n6 VPWR.n5 7.10563
R30 VPWR.n3 VPWR.n2 6.37948
R31 VPWR.n2 VPWR.n0 0.684108
R32 VPWR VPWR.n6 0.348167
R33 VPWR.n6 VPWR.n0 0.154648
R34 VPB.t2 VPB.t3 556.386
R35 VPB.t3 VPB.t1 284.113
R36 VPB.t1 VPB.t4 275.235
R37 VPB.t4 VPB.t5 248.599
R38 VPB.t0 VPB.t2 248.599
R39 VPB VPB.t0 189.409
R40 A2.n0 A2.t1 241.536
R41 A2.n0 A2.t0 169.237
R42 A2 A2.n0 167.361
R43 a_381_47.t0 a_381_47.t1 60.9236
R44 VGND.n4 VGND.n3 200.516
R45 VGND.n2 VGND.t2 168.667
R46 VGND.n11 VGND.t1 145.362
R47 VGND.n5 VGND.n1 34.6358
R48 VGND.n9 VGND.n1 34.6358
R49 VGND.n10 VGND.n9 34.6358
R50 VGND.n3 VGND.t3 33.2313
R51 VGND.n3 VGND.t0 24.9236
R52 VGND.n5 VGND.n4 21.4593
R53 VGND.n11 VGND.n10 10.9181
R54 VGND.n12 VGND.n11 9.3005
R55 VGND.n6 VGND.n5 9.3005
R56 VGND.n7 VGND.n1 9.3005
R57 VGND.n9 VGND.n8 9.3005
R58 VGND.n10 VGND.n0 9.3005
R59 VGND.n4 VGND.n2 6.62655
R60 VGND.n6 VGND.n2 0.636469
R61 VGND.n7 VGND.n6 0.120292
R62 VGND.n8 VGND.n7 0.120292
R63 VGND.n8 VGND.n0 0.120292
R64 VGND.n12 VGND.n0 0.120292
R65 VGND VGND.n12 0.0213333
R66 VNB.t1 VNB.t2 2790.94
R67 VNB.t2 VNB.t0 1366.99
R68 VNB.t0 VNB.t5 1324.27
R69 VNB.t5 VNB.t4 1196.12
R70 VNB.t3 VNB.t1 1082.2
R71 VNB VNB.t3 911.327
R72 B1.n0 B1.t1 239.505
R73 B1.n0 B1.t0 167.204
R74 B1 B1.n0 161.85
R75 a_109_47.t0 a_109_47.t1 42.462
R76 a_109_297.n1 a_109_297.n0 953.038
R77 a_109_297.n0 a_109_297.t2 33.4905
R78 a_109_297.n0 a_109_297.t3 31.5205
R79 a_109_297.n1 a_109_297.t1 26.5955
R80 a_109_297.t0 a_109_297.n1 26.5955
R81 A1.n0 A1.t0 233.869
R82 A1.n0 A1.t1 161.57
R83 A1.n1 A1.n0 155.657
R84 A1 A1.n1 18.8957
R85 A1.n1 A1 3.9624
R86 B2.n0 B2.t0 241.536
R87 B2.n0 B2.t1 169.237
R88 B2 B2.n0 168.641
C0 VPB VPWR 0.085341f
C1 VPB A1 0.036285f
C2 B2 B1 0.073857f
C3 B2 VPWR 0.008225f
C4 VPB X 0.004164f
C5 VPB A2 0.027075f
C6 VPB VGND 0.009426f
C7 B2 X 5.48e-20
C8 B1 VPWR 0.009814f
C9 B1 A1 0.061274f
C10 B2 VGND 0.053141f
C11 B1 X 9.58e-20
C12 A1 VPWR 0.016511f
C13 VPWR X 0.176244f
C14 A2 VPWR 0.020999f
C15 B1 VGND 0.026201f
C16 A1 X 2.78e-19
C17 VPWR VGND 0.085699f
C18 A1 A2 0.069791f
C19 A2 X 0.00156f
C20 A1 VGND 0.012952f
C21 X VGND 0.12295f
C22 A2 VGND 0.016888f
C23 VPB B2 0.029838f
C24 VPB B1 0.032101f
C25 VGND VNB 0.501765f
C26 X VNB 0.019986f
C27 VPWR VNB 0.404843f
C28 A2 VNB 0.089869f
C29 A1 VNB 0.110582f
C30 B1 VNB 0.112455f
C31 B2 VNB 0.126345f
C32 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22oi_4 VNB VPB VGND VPWR A1 A2 B2 Y B1
X0 a_27_47.t7 B1.t0 Y.t8 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47.t6 B1.t1 Y.t7 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297.t14 A2.t0 VPWR.t6 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 Y.t12 B1.t2 a_27_297.t10 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297.t4 B2.t0 Y.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t5 A2.t1 a_27_297.t13 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297.t12 A2.t2 VPWR.t4 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y.t13 A1.t0 a_803_47.t3 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y.t3 B2.t1 a_27_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR.t3 A2.t3 a_27_297.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y.t1 A1.t1 a_803_47.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND.t7 A2.t4 a_803_47.t7 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_297.t6 B2.t2 Y.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47.t0 B2.t3 VGND.t3 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_27_47.t1 B2.t4 VGND.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_803_47.t1 A1.t2 Y.t14 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_297.t9 B1.t3 Y.t11 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47.t0 A1.t3 Y.t15 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_803_47.t6 A2.t5 VGND.t6 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_803_47.t5 A2.t6 VGND.t5 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND.t1 B2.t5 a_27_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y.t6 B1.t4 a_27_47.t5 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t10 B1.t5 a_27_297.t8 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297.t15 A1.t4 VPWR.t7 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y.t5 B1.t6 a_27_47.t4 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_27_297.t7 B1.t7 Y.t9 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR.t0 A1.t5 a_27_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_27_297.t1 A1.t6 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND.t4 A2.t7 a_803_47.t4 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y.t0 B2.t6 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR.t2 A1.t7 a_27_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND.t0 B2.t7 a_27_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n0 B1.t3 212.081
R1 B1.n2 B1.t5 212.081
R2 B1.n4 B1.t7 212.081
R3 B1.n3 B1.t2 212.081
R4 B1 B1.n5 158.081
R5 B1.n0 B1.t1 139.78
R6 B1.n2 B1.t6 139.78
R7 B1.n4 B1.t0 139.78
R8 B1.n3 B1.t4 139.78
R9 B1 B1.n1 91.0594
R10 B1.n4 B1.n3 61.346
R11 B1.n2 B1.n1 39.1809
R12 B1.n5 B1.n4 35.7853
R13 B1.n5 B1.n2 25.5611
R14 B1.n1 B1.n0 18.4714
R15 Y.n9 Y.n8 351.986
R16 Y.n14 Y.n13 302.774
R17 Y.n12 Y.n11 301.14
R18 Y.n9 Y.n7 296.726
R19 Y.n2 Y.n0 229.8
R20 Y.n6 Y.n5 186.792
R21 Y.n2 Y.n1 185
R22 Y.n4 Y.n3 185
R23 Y.n4 Y.n2 72.5338
R24 Y.n12 Y.n10 48.0005
R25 Y.n14 Y.n12 41.9561
R26 Y.n6 Y.n4 40.2672
R27 Y.n10 Y.n6 34.8165
R28 Y.n13 Y.t4 26.5955
R29 Y.n13 Y.t0 26.5955
R30 Y.n7 Y.t9 26.5955
R31 Y.n7 Y.t12 26.5955
R32 Y.n8 Y.t11 26.5955
R33 Y.n8 Y.t10 26.5955
R34 Y.n11 Y.t2 26.5955
R35 Y.n11 Y.t3 26.5955
R36 Y.n5 Y.t8 24.9236
R37 Y.n5 Y.t6 24.9236
R38 Y.n3 Y.t7 24.9236
R39 Y.n3 Y.t5 24.9236
R40 Y.n1 Y.t15 24.9236
R41 Y.n1 Y.t1 24.9236
R42 Y.n0 Y.t14 24.9236
R43 Y.n0 Y.t13 24.9236
R44 Y Y.n14 5.48621
R45 Y.n10 Y.n9 2.84494
R46 a_27_47.t6 a_27_47.n5 312.334
R47 a_27_47.n5 a_27_47.n4 185
R48 a_27_47.n1 a_27_47.t3 174.512
R49 a_27_47.n1 a_27_47.n0 98.982
R50 a_27_47.n3 a_27_47.n2 88.3446
R51 a_27_47.n5 a_27_47.n3 53.5212
R52 a_27_47.n3 a_27_47.n1 48.9326
R53 a_27_47.n4 a_27_47.t4 24.9236
R54 a_27_47.n4 a_27_47.t7 24.9236
R55 a_27_47.n2 a_27_47.t5 24.9236
R56 a_27_47.n2 a_27_47.t1 24.9236
R57 a_27_47.n0 a_27_47.t2 24.9236
R58 a_27_47.n0 a_27_47.t0 24.9236
R59 VNB.t7 VNB.t4 2677.02
R60 VNB.t10 VNB.t12 1196.12
R61 VNB.t11 VNB.t10 1196.12
R62 VNB.t15 VNB.t11 1196.12
R63 VNB.t13 VNB.t15 1196.12
R64 VNB.t9 VNB.t13 1196.12
R65 VNB.t14 VNB.t9 1196.12
R66 VNB.t4 VNB.t14 1196.12
R67 VNB.t5 VNB.t7 1196.12
R68 VNB.t8 VNB.t5 1196.12
R69 VNB.t6 VNB.t8 1196.12
R70 VNB.t1 VNB.t6 1196.12
R71 VNB.t2 VNB.t1 1196.12
R72 VNB.t0 VNB.t2 1196.12
R73 VNB.t3 VNB.t0 1196.12
R74 VNB VNB.t3 911.327
R75 A2.n3 A2.t0 212.081
R76 A2.n5 A2.t1 212.081
R77 A2.n7 A2.t2 212.081
R78 A2.n1 A2.t3 212.081
R79 A2.n4 A2.n0 172.725
R80 A2.n9 A2.n2 172.725
R81 A2.n6 A2.n0 152
R82 A2.n9 A2.n8 152
R83 A2.n3 A2.t6 139.78
R84 A2.n5 A2.t7 139.78
R85 A2.n7 A2.t5 139.78
R86 A2.n1 A2.t4 139.78
R87 A2.n8 A2.n6 49.6611
R88 A2.n7 A2.n2 48.2005
R89 A2.n5 A2.n4 39.4369
R90 A2.n4 A2.n3 21.9096
R91 A2.n2 A2.n1 13.146
R92 A2 A2.n0 11.5815
R93 A2.n6 A2.n5 10.2247
R94 A2 A2.n9 9.14336
R95 A2.n8 A2.n7 1.46111
R96 VPWR.n7 VPWR.n6 323.952
R97 VPWR.n10 VPWR.n3 318.293
R98 VPWR.n5 VPWR.n4 318.293
R99 VPWR.n12 VPWR.n1 318.293
R100 VPWR.n11 VPWR.n10 33.5064
R101 VPWR.n9 VPWR.n5 27.4829
R102 VPWR.n1 VPWR.t1 26.5955
R103 VPWR.n1 VPWR.t2 26.5955
R104 VPWR.n3 VPWR.t7 26.5955
R105 VPWR.n3 VPWR.t0 26.5955
R106 VPWR.n4 VPWR.t4 26.5955
R107 VPWR.n4 VPWR.t3 26.5955
R108 VPWR.n6 VPWR.t6 26.5955
R109 VPWR.n6 VPWR.t5 26.5955
R110 VPWR.n10 VPWR.n9 16.9417
R111 VPWR.n13 VPWR.n12 12.4952
R112 VPWR.n12 VPWR.n11 10.9181
R113 VPWR.n9 VPWR.n8 9.3005
R114 VPWR.n10 VPWR.n2 9.3005
R115 VPWR.n11 VPWR.n0 9.3005
R116 VPWR.n7 VPWR.n5 6.64428
R117 VPWR VPWR.n13 1.078
R118 VPWR.n8 VPWR.n7 0.584064
R119 VPWR.n13 VPWR.n0 0.147187
R120 VPWR.n8 VPWR.n2 0.120292
R121 VPWR.n2 VPWR.n0 0.120292
R122 a_27_297.n14 a_27_297.n13 585
R123 a_27_297.n13 a_27_297.n3 585
R124 a_27_297.n16 a_27_297.n15 300.885
R125 a_27_297.n1 a_27_297.n0 300.885
R126 a_27_297.n18 a_27_297.n17 300.885
R127 a_27_297.n11 a_27_297.n2 291.094
R128 a_27_297.n5 a_27_297.t14 279.526
R129 a_27_297.n1 a_27_297.t3 272.372
R130 a_27_297.n12 a_27_297.n10 268.952
R131 a_27_297.n5 a_27_297.n4 208.507
R132 a_27_297.n7 a_27_297.n6 208.507
R133 a_27_297.n9 a_27_297.n8 208.507
R134 a_27_297.n12 a_27_297.n11 47.0974
R135 a_27_297.n13 a_27_297.n12 47.0974
R136 a_27_297.n10 a_27_297.n9 45.7539
R137 a_27_297.n16 a_27_297.n14 45.7539
R138 a_27_297.n7 a_27_297.n5 44.424
R139 a_27_297.n9 a_27_297.n7 44.424
R140 a_27_297.n17 a_27_297.n1 44.424
R141 a_27_297.n17 a_27_297.n16 44.424
R142 a_27_297.n13 a_27_297.t2 26.5955
R143 a_27_297.n11 a_27_297.t9 26.5955
R144 a_27_297.n4 a_27_297.t13 26.5955
R145 a_27_297.n4 a_27_297.t12 26.5955
R146 a_27_297.n6 a_27_297.t11 26.5955
R147 a_27_297.n6 a_27_297.t15 26.5955
R148 a_27_297.n8 a_27_297.t0 26.5955
R149 a_27_297.n8 a_27_297.t1 26.5955
R150 a_27_297.n15 a_27_297.t8 26.5955
R151 a_27_297.n15 a_27_297.t7 26.5955
R152 a_27_297.n0 a_27_297.t5 26.5955
R153 a_27_297.n0 a_27_297.t6 26.5955
R154 a_27_297.t10 a_27_297.n18 26.5955
R155 a_27_297.n18 a_27_297.t4 26.5955
R156 a_27_297.n10 a_27_297.n3 5.65245
R157 a_27_297.n3 a_27_297.n2 2.81339
R158 a_27_297.n14 a_27_297.n2 2.81339
R159 VPB.t9 VPB.t2 556.386
R160 VPB.t13 VPB.t14 248.599
R161 VPB.t12 VPB.t13 248.599
R162 VPB.t11 VPB.t12 248.599
R163 VPB.t15 VPB.t11 248.599
R164 VPB.t0 VPB.t15 248.599
R165 VPB.t1 VPB.t0 248.599
R166 VPB.t2 VPB.t1 248.599
R167 VPB.t8 VPB.t9 248.599
R168 VPB.t7 VPB.t8 248.599
R169 VPB.t10 VPB.t7 248.599
R170 VPB.t4 VPB.t10 248.599
R171 VPB.t5 VPB.t4 248.599
R172 VPB.t6 VPB.t5 248.599
R173 VPB.t3 VPB.t6 248.599
R174 VPB VPB.t3 189.409
R175 B2.n3 B2.t0 212.081
R176 B2.n5 B2.t1 212.081
R177 B2.n7 B2.t2 212.081
R178 B2.n1 B2.t6 212.081
R179 B2.n4 B2.n0 173.761
R180 B2.n9 B2.n2 173.761
R181 B2.n6 B2.n0 152
R182 B2.n9 B2.n8 152
R183 B2.n3 B2.t4 139.78
R184 B2.n5 B2.t5 139.78
R185 B2.n7 B2.t3 139.78
R186 B2.n1 B2.t7 139.78
R187 B2.n8 B2.n6 49.6611
R188 B2.n5 B2.n4 48.2005
R189 B2.n7 B2.n2 39.4369
R190 B2.n2 B2.n1 21.9096
R191 B2 B2.n0 14.7205
R192 B2.n4 B2.n3 13.146
R193 B2.n8 B2.n7 10.2247
R194 B2 B2.n9 7.0405
R195 B2.n6 B2.n5 1.46111
R196 A1.n2 A1.t4 212.081
R197 A1.n1 A1.t5 212.081
R198 A1.n7 A1.t6 212.081
R199 A1.n8 A1.t7 212.081
R200 A1.n4 A1.n3 172.725
R201 A1 A1.n9 172.114
R202 A1.n5 A1.n4 152
R203 A1.n6 A1.n0 152
R204 A1.n2 A1.t2 139.78
R205 A1.n1 A1.t0 139.78
R206 A1.n7 A1.t3 139.78
R207 A1.n8 A1.t1 139.78
R208 A1.n6 A1.n5 49.6611
R209 A1.n9 A1.n7 48.2005
R210 A1.n3 A1.n1 39.4369
R211 A1.n3 A1.n2 21.9096
R212 A1.n4 A1.n0 20.7243
R213 A1.n9 A1.n8 13.146
R214 A1.n5 A1.n1 10.2247
R215 A1.n7 A1.n6 1.46111
R216 A1 A1.n0 0.610024
R217 a_803_47.n4 a_803_47.t2 312.334
R218 a_803_47.n5 a_803_47.n4 185
R219 a_803_47.n1 a_803_47.t5 174.512
R220 a_803_47.n1 a_803_47.n0 98.982
R221 a_803_47.n3 a_803_47.n2 88.3446
R222 a_803_47.n4 a_803_47.n3 53.5212
R223 a_803_47.n3 a_803_47.n1 48.9326
R224 a_803_47.n2 a_803_47.t7 24.9236
R225 a_803_47.n2 a_803_47.t1 24.9236
R226 a_803_47.n0 a_803_47.t4 24.9236
R227 a_803_47.n0 a_803_47.t6 24.9236
R228 a_803_47.t3 a_803_47.n5 24.9236
R229 a_803_47.n5 a_803_47.t0 24.9236
R230 VGND.n12 VGND.n11 214.865
R231 VGND.n10 VGND.n9 207.965
R232 VGND.n3 VGND.n2 207.965
R233 VGND.n33 VGND.n1 207.965
R234 VGND.n34 VGND.n33 43.1829
R235 VGND.n12 VGND.n10 37.9269
R236 VGND.n15 VGND.n14 34.6358
R237 VGND.n16 VGND.n15 34.6358
R238 VGND.n16 VGND.n7 34.6358
R239 VGND.n20 VGND.n7 34.6358
R240 VGND.n21 VGND.n20 34.6358
R241 VGND.n22 VGND.n21 34.6358
R242 VGND.n22 VGND.n5 34.6358
R243 VGND.n26 VGND.n5 34.6358
R244 VGND.n27 VGND.n26 34.6358
R245 VGND.n28 VGND.n27 34.6358
R246 VGND.n32 VGND.n31 34.6358
R247 VGND.n31 VGND.n3 27.8593
R248 VGND.n11 VGND.t5 24.9236
R249 VGND.n11 VGND.t4 24.9236
R250 VGND.n9 VGND.t6 24.9236
R251 VGND.n9 VGND.t7 24.9236
R252 VGND.n2 VGND.t2 24.9236
R253 VGND.n2 VGND.t1 24.9236
R254 VGND.n1 VGND.t3 24.9236
R255 VGND.n1 VGND.t0 24.9236
R256 VGND.n14 VGND.n13 9.3005
R257 VGND.n15 VGND.n8 9.3005
R258 VGND.n17 VGND.n16 9.3005
R259 VGND.n18 VGND.n7 9.3005
R260 VGND.n20 VGND.n19 9.3005
R261 VGND.n21 VGND.n6 9.3005
R262 VGND.n23 VGND.n22 9.3005
R263 VGND.n24 VGND.n5 9.3005
R264 VGND.n26 VGND.n25 9.3005
R265 VGND.n27 VGND.n4 9.3005
R266 VGND.n29 VGND.n28 9.3005
R267 VGND.n31 VGND.n30 9.3005
R268 VGND.n32 VGND.n0 9.3005
R269 VGND.n28 VGND.n3 6.77697
R270 VGND.n14 VGND.n10 2.25932
R271 VGND.n13 VGND.n12 2.19951
R272 VGND.n33 VGND.n32 0.753441
R273 VGND.n13 VGND.n8 0.120292
R274 VGND.n17 VGND.n8 0.120292
R275 VGND.n18 VGND.n17 0.120292
R276 VGND.n19 VGND.n18 0.120292
R277 VGND.n19 VGND.n6 0.120292
R278 VGND.n23 VGND.n6 0.120292
R279 VGND.n24 VGND.n23 0.120292
R280 VGND.n25 VGND.n24 0.120292
R281 VGND.n25 VGND.n4 0.120292
R282 VGND.n29 VGND.n4 0.120292
R283 VGND.n30 VGND.n29 0.120292
R284 VGND.n30 VGND.n0 0.120292
R285 VGND.n34 VGND.n0 0.120292
R286 VGND VGND.n34 0.0213333
C0 VPB B2 0.120076f
C1 Y VGND 0.052741f
C2 VPB B1 0.129554f
C3 VPWR VGND 0.148029f
C4 VPB A1 0.12053f
C5 B2 B1 0.05266f
C6 VPB A2 0.122062f
C7 VPB Y 0.013831f
C8 B1 A1 0.034476f
C9 VPB VPWR 0.141473f
C10 B2 Y 0.179587f
C11 VPB VGND 0.010415f
C12 B2 VPWR 0.033971f
C13 B1 Y 0.311549f
C14 A1 A2 0.065868f
C15 A1 Y 0.13232f
C16 B2 VGND 0.059432f
C17 B1 VPWR 0.031189f
C18 A1 VPWR 0.078224f
C19 B1 VGND 0.033279f
C20 A2 Y 3.06e-19
C21 A2 VPWR 0.092162f
C22 A1 VGND 0.033779f
C23 A2 VGND 0.062836f
C24 Y VPWR 0.034964f
C25 VGND VNB 0.85071f
C26 VPWR VNB 0.701484f
C27 Y VNB 0.030159f
C28 A2 VNB 0.393622f
C29 A1 VNB 0.362302f
C30 B1 VNB 0.381938f
C31 B2 VNB 0.392365f
C32 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47.t1 A1.t0 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y.t2 B1.t0 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR.t1 A1.t1 a_113_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297.t1 B1.t1 Y.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND.t1 A2.t1 a_199_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
R0 A1.n0 A1.t1 241.536
R1 A1.n0 A1.t0 169.237
R2 A1 A1.n0 156.655
R3 Y.n0 Y.t0 358.224
R4 Y Y.n1 270.289
R5 Y.n1 Y.t1 25.8467
R6 Y.n1 Y.t2 25.8467
R7 Y Y.n0 8.33467
R8 Y.n0 Y 7.34578
R9 a_199_47.t0 a_199_47.t1 54.462
R10 VNB.t1 VNB.t0 1267.31
R11 VNB.t2 VNB.t1 1224.6
R12 VNB VNB.t2 982.524
R13 A2.n0 A2.t0 231.017
R14 A2.n0 A2.t1 158.716
R15 A2 A2.n0 154.387
R16 VPWR VPWR.n0 614.966
R17 VPWR.n0 VPWR.t0 30.5355
R18 VPWR.n0 VPWR.t1 27.5805
R19 a_113_297.t0 a_113_297.n0 538.659
R20 a_113_297.n0 a_113_297.t2 27.5805
R21 a_113_297.n0 a_113_297.t1 27.5805
R22 VPB.t2 VPB.t0 263.397
R23 VPB.t1 VPB.t2 254.518
R24 VPB VPB.t1 204.207
R25 B1.n0 B1.t1 229.369
R26 B1.n0 B1.t0 157.07
R27 B1 B1.n0 154.934
R28 VGND.n0 VGND.t0 288
R29 VGND.n0 VGND.t1 240.708
R30 VGND VGND.n0 0.160744
C0 Y VPB 0.014642f
C1 VPWR VGND 0.036961f
C2 Y B1 0.112603f
C3 VPWR VPB 0.042396f
C4 VGND VPB 0.005478f
C5 VPWR B1 0.01343f
C6 VGND B1 0.043596f
C7 VPB B1 0.038865f
C8 A1 A2 0.091231f
C9 A1 Y 0.081255f
C10 A1 VPWR 0.015389f
C11 A2 Y 0.001218f
C12 A1 VGND 0.077964f
C13 A2 VPWR 0.014703f
C14 A1 VPB 0.026387f
C15 A2 VGND 0.049477f
C16 Y VPWR 0.044654f
C17 A2 VPB 0.037282f
C18 A1 B1 0.051837f
C19 Y VGND 0.065351f
C20 VGND VNB 0.285624f
C21 VPWR VNB 0.210674f
C22 Y VNB 0.054434f
C23 A2 VNB 0.143834f
C24 A1 VNB 0.098086f
C25 B1 VNB 0.161998f
C26 VPB VNB 0.427572f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_4 VNB VPB VGND VPWR X B1 A1 A2
X0 VGND.t3 B1.t0 a_84_21.t4 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_741_47.t0 A2.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_84_21.t5 A1.t0 a_741_47.t1 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.07475 ps=0.88 w=0.65 l=0.15
X3 VGND.t1 A2.t1 a_901_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t7 a_84_21.t6 X.t7 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR.t1 A2.t2 a_483_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_483_297.t1 B1.t1 a_84_21.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X.t3 a_84_21.t7 VGND.t5 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X8 a_84_21.t1 B1.t2 a_483_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND.t4 a_84_21.t8 X.t2 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.264875 pd=1.465 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VPWR.t6 a_84_21.t9 X.t6 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_483_297.t2 A2.t3 VPWR.t0 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=2.79 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR.t3 A1.t1 a_483_297.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND.t7 a_84_21.t10 X.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 X.t5 a_84_21.t11 VPWR.t5 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X15 a_84_21.t3 B1.t3 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.264875 ps=1.465 w=0.65 l=0.15
X16 a_483_297.t4 A1.t2 VPWR.t2 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X.t0 a_84_21.t12 VGND.t6 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_901_47.t1 A1.t3 a_84_21.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X.t4 a_84_21.t13 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 B1.n0 B1.t1 212.081
R1 B1.n1 B1.t2 212.081
R2 B1 B1.n1 174.732
R3 B1.n0 B1.t0 139.78
R4 B1.n1 B1.t3 139.78
R5 B1.n1 B1.n0 61.346
R6 a_84_21.n12 a_84_21.n0 363.517
R7 a_84_21.n0 a_84_21.n2 271.764
R8 a_84_21.n9 a_84_21.t6 212.081
R9 a_84_21.n7 a_84_21.t13 212.081
R10 a_84_21.n5 a_84_21.t9 212.081
R11 a_84_21.n4 a_84_21.t11 212.081
R12 a_84_21.n11 a_84_21.n1 96.3742
R13 a_84_21.n0 a_84_21.n1 2.11365
R14 a_84_21.n6 a_84_21.n3 165.189
R15 a_84_21.n10 a_84_21.n9 160.034
R16 a_84_21.n8 a_84_21.n3 152
R17 a_84_21.n9 a_84_21.t8 139.78
R18 a_84_21.n7 a_84_21.t12 139.78
R19 a_84_21.n5 a_84_21.t10 139.78
R20 a_84_21.n4 a_84_21.t7 139.78
R21 a_84_21.n1 a_84_21.n10 85.8738
R22 a_84_21.n5 a_84_21.n4 62.8066
R23 a_84_21.n9 a_84_21.n8 41.6278
R24 a_84_21.n6 a_84_21.n5 34.3247
R25 a_84_21.n7 a_84_21.n6 28.4823
R26 a_84_21.n12 a_84_21.t2 26.5955
R27 a_84_21.t1 a_84_21.n12 26.5955
R28 a_84_21.n11 a_84_21.t4 24.9236
R29 a_84_21.n11 a_84_21.t3 24.9236
R30 a_84_21.n2 a_84_21.t0 24.9236
R31 a_84_21.n2 a_84_21.t5 24.9236
R32 a_84_21.n8 a_84_21.n7 21.1793
R33 a_84_21.n10 a_84_21.n3 13.1884
R34 VGND.n20 VGND.t5 282.764
R35 VGND.n5 VGND.n4 198.964
R36 VGND.n18 VGND.n2 198.964
R37 VGND.n13 VGND.n12 185
R38 VGND.n11 VGND.n10 185
R39 VGND.n6 VGND.t1 160.863
R40 VGND.n12 VGND.n11 75.6928
R41 VGND.n12 VGND.t4 46.1543
R42 VGND.n4 VGND.t3 32.3082
R43 VGND.n11 VGND.t2 28.6159
R44 VGND.n9 VGND.n8 26.7086
R45 VGND.n14 VGND.n1 26.4529
R46 VGND.n2 VGND.t6 25.8467
R47 VGND.n2 VGND.t7 25.8467
R48 VGND.n4 VGND.t0 24.9236
R49 VGND.n18 VGND.n1 22.9652
R50 VGND.n19 VGND.n18 21.4593
R51 VGND.n8 VGND.n5 19.9534
R52 VGND.n20 VGND.n19 18.4476
R53 VGND.n13 VGND.n10 9.90239
R54 VGND.n21 VGND.n20 9.3005
R55 VGND.n19 VGND.n0 9.3005
R56 VGND.n18 VGND.n17 9.3005
R57 VGND.n16 VGND.n1 9.3005
R58 VGND.n15 VGND.n14 9.3005
R59 VGND.n9 VGND.n3 9.3005
R60 VGND.n8 VGND.n7 9.3005
R61 VGND.n6 VGND.n5 7.15453
R62 VGND.n14 VGND.n13 0.966538
R63 VGND.n10 VGND.n9 0.242009
R64 VGND.n7 VGND.n6 0.184012
R65 VGND.n7 VGND.n3 0.120292
R66 VGND.n15 VGND.n3 0.120292
R67 VGND.n16 VGND.n15 0.120292
R68 VGND.n17 VGND.n16 0.120292
R69 VGND.n17 VGND.n0 0.120292
R70 VGND.n21 VGND.n0 0.120292
R71 VGND VGND.n21 0.0226354
R72 VNB.t8 VNB.t3 2748.22
R73 VNB.t4 VNB.t0 1310.03
R74 VNB.t6 VNB.t8 1224.6
R75 VNB.t7 VNB.t6 1224.6
R76 VNB.t9 VNB.t7 1224.6
R77 VNB.t2 VNB.t1 1196.12
R78 VNB.t5 VNB.t2 1196.12
R79 VNB.t3 VNB.t4 1196.12
R80 VNB.t0 VNB.t5 1082.2
R81 VNB VNB.t9 996.764
R82 A2 A2.n0 254.977
R83 A2.n1 A2.t3 241.536
R84 A2.n0 A2.t2 241.536
R85 A2.n1 A2.t1 169.237
R86 A2.n0 A2.t0 169.237
R87 A2 A2.n1 166.593
R88 a_741_47.t0 a_741_47.t1 42.462
R89 A1.n0 A1.t1 212.081
R90 A1.n1 A1.t2 212.081
R91 A1 A1.n2 157.555
R92 A1.n0 A1.t3 139.78
R93 A1.n1 A1.t0 139.78
R94 A1.n2 A1.n0 35.055
R95 A1.n2 A1.n1 26.2914
R96 a_901_47.t0 a_901_47.t1 49.8467
R97 X.n2 X.n1 355.265
R98 X.n2 X.n0 297.406
R99 X.n5 X.n3 249.754
R100 X.n5 X.n4 185
R101 X.n0 X.t6 27.5805
R102 X.n0 X.t5 27.5805
R103 X.n1 X.t7 27.5805
R104 X.n1 X.t4 27.5805
R105 X.n4 X.t1 25.8467
R106 X.n4 X.t3 25.8467
R107 X.n3 X.t2 25.8467
R108 X.n3 X.t0 25.8467
R109 X X.n5 25.6859
R110 X.n6 X.n2 24.4711
R111 X X.n6 18.0711
R112 X.n6 X 3.69535
R113 VPWR.n8 VPWR.n7 604.317
R114 VPWR.n6 VPWR.n5 598.965
R115 VPWR.n19 VPWR.t5 337.305
R116 VPWR.n17 VPWR.n2 309.726
R117 VPWR.n3 VPWR.t7 250.424
R118 VPWR.n11 VPWR.n10 34.6358
R119 VPWR.n12 VPWR.n11 34.6358
R120 VPWR.n2 VPWR.t4 27.5805
R121 VPWR.n2 VPWR.t6 27.5805
R122 VPWR.n12 VPWR.n3 27.4829
R123 VPWR.n5 VPWR.t2 26.5955
R124 VPWR.n5 VPWR.t1 26.5955
R125 VPWR.n7 VPWR.t0 26.5955
R126 VPWR.n7 VPWR.t3 26.5955
R127 VPWR.n16 VPWR.n3 22.9652
R128 VPWR.n17 VPWR.n16 22.9652
R129 VPWR.n18 VPWR.n17 21.4593
R130 VPWR.n19 VPWR.n18 18.4476
R131 VPWR.n10 VPWR.n6 13.9299
R132 VPWR.n10 VPWR.n9 9.3005
R133 VPWR.n11 VPWR.n4 9.3005
R134 VPWR.n13 VPWR.n12 9.3005
R135 VPWR.n14 VPWR.n3 9.3005
R136 VPWR.n16 VPWR.n15 9.3005
R137 VPWR.n17 VPWR.n1 9.3005
R138 VPWR.n18 VPWR.n0 9.3005
R139 VPWR.n20 VPWR.n19 9.3005
R140 VPWR.n8 VPWR.n6 6.71935
R141 VPWR.n9 VPWR.n8 0.822144
R142 VPWR.n9 VPWR.n4 0.120292
R143 VPWR.n13 VPWR.n4 0.120292
R144 VPWR.n14 VPWR.n13 0.120292
R145 VPWR.n15 VPWR.n14 0.120292
R146 VPWR.n15 VPWR.n1 0.120292
R147 VPWR.n1 VPWR.n0 0.120292
R148 VPWR.n20 VPWR.n0 0.120292
R149 VPWR VPWR.n20 0.0226354
R150 VPB.t9 VPB.t0 571.184
R151 VPB.t6 VPB.t9 254.518
R152 VPB.t8 VPB.t6 254.518
R153 VPB.t7 VPB.t8 254.518
R154 VPB.t5 VPB.t2 248.599
R155 VPB.t4 VPB.t5 248.599
R156 VPB.t3 VPB.t4 248.599
R157 VPB.t1 VPB.t3 248.599
R158 VPB.t0 VPB.t1 248.599
R159 VPB VPB.t7 207.166
R160 a_483_297.n2 a_483_297.t0 415.298
R161 a_483_297.n1 a_483_297.t2 312.822
R162 a_483_297.n1 a_483_297.n0 297.678
R163 a_483_297.n3 a_483_297.n2 296.05
R164 a_483_297.n2 a_483_297.n1 61.1665
R165 a_483_297.n0 a_483_297.t5 26.5955
R166 a_483_297.n0 a_483_297.t4 26.5955
R167 a_483_297.n3 a_483_297.t3 26.5955
R168 a_483_297.t1 a_483_297.n3 26.5955
C0 A1 VGND 0.030546f
C1 VPWR X 0.24746f
C2 VPWR VGND 0.113278f
C3 X VGND 0.139527f
C4 VPB B1 0.070497f
C5 VPB A2 0.065645f
C6 VPB A1 0.051281f
C7 B1 A2 0.058455f
C8 VPB VPWR 0.127685f
C9 B1 VPWR 0.024437f
C10 VPB X 0.011541f
C11 A2 A1 0.210667f
C12 B1 X 0.002734f
C13 VPB VGND 0.011955f
C14 A2 VPWR 0.039898f
C15 B1 VGND 0.036448f
C16 A1 VPWR 0.026688f
C17 A2 VGND 0.059931f
C18 VGND VNB 0.661897f
C19 X VNB 0.067151f
C20 VPWR VNB 0.541237f
C21 A1 VNB 0.168575f
C22 A2 VNB 0.222527f
C23 B1 VNB 0.195735f
C24 VPB VNB 1.13634f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR.t2 a_80_21.t3 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297.t2 A3.t0 VPWR.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47.t0 A2.t0 a_209_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47.t1 A3.t1 VGND.t2 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND.t0 a_80_21.t4 X.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND.t1 B1.t0 a_80_21.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21.t2 A1.t0 a_303_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR.t3 A2.t1 a_209_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21.t0 B1.t1 a_209_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297.t1 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
R0 a_80_21.t0 a_80_21.n2 467.872
R1 a_80_21.n2 a_80_21.n0 269.12
R2 a_80_21.n0 a_80_21.t3 241
R3 a_80_21.n0 a_80_21.t4 168.701
R4 a_80_21.n2 a_80_21.n1 95.685
R5 a_80_21.n1 a_80_21.t1 34.1543
R6 a_80_21.n1 a_80_21.t2 26.7697
R7 X X.n0 593.34
R8 X.n3 X.n0 585
R9 X.n2 X.n0 585
R10 X.n1 X.t0 128.517
R11 X.n2 X.n1 63.7581
R12 X.n0 X.t1 27.5805
R13 X.n3 X 8.33989
R14 X.n1 X 5.759
R15 X X.n3 4.84898
R16 X X.n2 4.84898
R17 VPWR.n2 VPWR.n0 608.785
R18 VPWR.n2 VPWR.n1 229.508
R19 VPWR.n1 VPWR.t0 34.4755
R20 VPWR.n1 VPWR.t2 33.4905
R21 VPWR.n0 VPWR.t1 32.5055
R22 VPWR.n0 VPWR.t3 32.5055
R23 VPWR VPWR.n2 0.432488
R24 VPB.t3 VPB.t1 292.991
R25 VPB.t2 VPB.t0 284.113
R26 VPB.t4 VPB.t2 284.113
R27 VPB.t1 VPB.t4 278.193
R28 VPB VPB.t3 192.369
R29 A3.n0 A3.t0 241.536
R30 A3.n0 A3.t1 169.237
R31 A3.n1 A3.n0 152
R32 A3.n1 A3 14.0693
R33 A3 A3.n1 2.3087
R34 a_209_297.n1 a_209_297.n0 653.061
R35 a_209_297.n0 a_209_297.t3 32.5055
R36 a_209_297.t0 a_209_297.n1 32.5055
R37 a_209_297.n1 a_209_297.t1 32.5055
R38 a_209_297.n0 a_209_297.t2 30.5355
R39 A2.n0 A2.t1 241.536
R40 A2.n0 A2.t0 169.237
R41 A2.n1 A2.n0 152
R42 A2.n1 A2 12.8005
R43 A2 A2.n1 2.47068
R44 a_209_47.t0 a_209_47.t1 59.0774
R45 a_303_47.t0 a_303_47.t1 60.9236
R46 VNB.t1 VNB.t3 1409.71
R47 VNB.t4 VNB.t2 1366.99
R48 VNB.t0 VNB.t4 1366.99
R49 VNB.t3 VNB.t0 1338.51
R50 VNB VNB.t1 925.567
R51 VGND.n1 VGND.t1 237.055
R52 VGND.n1 VGND.n0 206.165
R53 VGND.n0 VGND.t0 38.7697
R54 VGND.n0 VGND.t2 24.9236
R55 VGND VGND.n1 0.167132
R56 B1.n0 B1.t1 241.536
R57 B1.n0 B1.t0 169.237
R58 B1.n1 B1.n0 152
R59 B1.n1 B1 14.8903
R60 B1 B1.n1 2.87397
R61 A1.n0 A1.t1 241.536
R62 A1.n0 A1.t0 169.237
R63 A1.n1 A1.n0 152
R64 A1.n1 A1 13.7665
R65 A1 A1.n1 2.6571
C0 VPB VPWR 0.071542f
C1 A3 X 0.00625f
C2 VPB VGND 0.007686f
C3 A3 VPWR 0.040256f
C4 A1 B1 0.101116f
C5 A2 X 3.42e-19
C6 A1 X 1.56e-19
C7 A3 VGND 0.016898f
C8 A2 VPWR 0.022678f
C9 A2 VGND 0.014804f
C10 A1 VPWR 0.018013f
C11 B1 VPWR 0.01773f
C12 A1 VGND 0.013522f
C13 B1 VGND 0.017205f
C14 X VPWR 0.117035f
C15 VPB A3 0.02968f
C16 X VGND 0.057244f
C17 VPB A2 0.028537f
C18 VPWR VGND 0.06622f
C19 A3 A2 0.108535f
C20 VPB A1 0.028686f
C21 VPB B1 0.034195f
C22 A2 A1 0.104261f
C23 VPB X 0.010822f
C24 VGND VNB 0.410332f
C25 VPWR VNB 0.331823f
C26 X VNB 0.08952f
C27 B1 VNB 0.11534f
C28 A1 VNB 0.089669f
C29 A2 VNB 0.089585f
C30 A3 VNB 0.089866f
C31 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31o_2 VNB VPB VGND VPWR B1 A1 A2 A3 X
X0 VPWR.t0 A2.t0 a_277_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297.t3 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_79_21.t0 B1.t0 a_277_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 a_277_297.t1 A3.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t3 a_79_21.t3 X.t1 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t3 a_79_21.t4 X.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_361_47.t0 A2.t1 a_277_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_277_47.t1 A3.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND.t0 B1.t1 a_79_21.t1 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X9 a_79_21.t2 A1.t1 a_361_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 X.t0 a_79_21.t5 VPWR.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 X.t2 a_79_21.t6 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n0 A2.t0 241.536
R1 A2 A2.n0 199.649
R2 A2.n0 A2.t1 169.237
R3 a_277_297.n1 a_277_297.n0 648.543
R4 a_277_297.n0 a_277_297.t3 38.4155
R5 a_277_297.n0 a_277_297.t2 26.5955
R6 a_277_297.t0 a_277_297.n1 26.5955
R7 a_277_297.n1 a_277_297.t1 26.5955
R8 VPWR.n6 VPWR.t4 873.438
R9 VPWR.n2 VPWR.n1 608.192
R10 VPWR.n4 VPWR.n3 316.245
R11 VPWR.n1 VPWR.t0 34.4755
R12 VPWR.n1 VPWR.t2 30.5355
R13 VPWR.n3 VPWR.t1 26.5955
R14 VPWR.n3 VPWR.t3 26.5955
R15 VPWR.n6 VPWR.n5 22.9652
R16 VPWR.n5 VPWR.n4 18.4476
R17 VPWR.n5 VPWR.n0 9.3005
R18 VPWR.n7 VPWR.n6 9.3005
R19 VPWR.n4 VPWR.n2 7.05667
R20 VPWR.n2 VPWR.n0 0.564795
R21 VPWR.n7 VPWR.n0 0.120292
R22 VPWR VPWR.n7 0.0213333
R23 VPB.t3 VPB.t2 284.113
R24 VPB.t0 VPB.t3 284.113
R25 VPB.t1 VPB.t0 248.599
R26 VPB.t4 VPB.t1 248.599
R27 VPB.t5 VPB.t4 248.599
R28 VPB VPB.t5 189.409
R29 A1.n0 A1.t0 241.536
R30 A1 A1.n0 202.931
R31 A1.n0 A1.t1 169.237
R32 B1.n0 B1.t0 227.987
R33 B1.n0 B1.t1 155.686
R34 B1 B1.n0 155.611
R35 a_79_21.t0 a_79_21.n4 384.991
R36 a_79_21.n4 a_79_21.n3 323.204
R37 a_79_21.n4 a_79_21.n0 263.637
R38 a_79_21.n1 a_79_21.t3 212.081
R39 a_79_21.n2 a_79_21.t5 212.081
R40 a_79_21.n1 a_79_21.t4 139.78
R41 a_79_21.n2 a_79_21.t6 139.78
R42 a_79_21.n0 a_79_21.t2 47.0774
R43 a_79_21.n3 a_79_21.n2 36.5157
R44 a_79_21.n0 a_79_21.t1 24.9236
R45 a_79_21.n3 a_79_21.n1 24.8308
R46 A3.n0 A3.t0 241.536
R47 A3.n0 A3.t1 169.237
R48 A3.n1 A3.n0 157.625
R49 A3.n1 A3 14.3615
R50 A3 A3.n1 3.68535
R51 X X.n1 639.212
R52 X.n2 X.n0 232.435
R53 X.n1 X.t1 26.5955
R54 X.n1 X.t0 26.5955
R55 X.n0 X.t3 24.9236
R56 X.n0 X.t2 24.9236
R57 X.n2 X 15.3103
R58 X X.n2 1.75736
R59 VGND.n5 VGND.t2 287.151
R60 VGND.n1 VGND.t0 286.2
R61 VGND.n3 VGND.n2 199.739
R62 VGND.n5 VGND.n4 25.977
R63 VGND.n2 VGND.t1 24.9236
R64 VGND.n2 VGND.t3 24.9236
R65 VGND.n4 VGND.n3 19.9534
R66 VGND.n6 VGND.n5 9.3005
R67 VGND.n4 VGND.n0 9.3005
R68 VGND.n3 VGND.n1 7.17083
R69 VGND.n1 VGND.n0 0.167755
R70 VGND.n6 VGND.n0 0.120292
R71 VGND VGND.n6 0.0213333
R72 VNB.t3 VNB.t0 1537.86
R73 VNB.t1 VNB.t3 1366.99
R74 VNB.t2 VNB.t1 1196.12
R75 VNB.t5 VNB.t2 1196.12
R76 VNB.t4 VNB.t5 1196.12
R77 VNB VNB.t4 911.327
R78 a_277_47.t0 a_277_47.t1 49.8467
R79 a_361_47.t0 a_361_47.t1 60.9236
C0 A1 VPWR 0.016019f
C1 A2 X 0.006462f
C2 A3 VGND 0.039164f
C3 A1 X 1.19e-19
C4 B1 VPWR 0.015249f
C5 A2 VGND 0.045029f
C6 A1 VGND 0.037217f
C7 B1 X 7.74e-20
C8 B1 VGND 0.037926f
C9 VPWR X 0.148098f
C10 VPB A3 0.025579f
C11 VPWR VGND 0.065156f
C12 VPB A2 0.026329f
C13 X VGND 0.11041f
C14 A3 A2 0.093978f
C15 VPB A1 0.027532f
C16 A3 A1 0.001914f
C17 VPB B1 0.041784f
C18 A2 A1 0.109286f
C19 VPB VPWR 0.069285f
C20 A3 VPWR 0.017034f
C21 VPB X 0.008894f
C22 A2 VPWR 0.016221f
C23 A3 X 0.014406f
C24 VPB VGND 0.007704f
C25 A1 B1 0.04921f
C26 VGND VNB 0.419014f
C27 X VNB 0.069146f
C28 VPWR VNB 0.334845f
C29 B1 VNB 0.162453f
C30 A1 VNB 0.093223f
C31 A2 VNB 0.092951f
C32 A3 VNB 0.09066f
C33 VPB VNB 0.69336f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31o_4 VNB VPB VGND VPWR X B1 A2 A1 A3
X0 VPWR.t3 a_277_47.t6 X.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X.t2 a_277_47.t7 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X.t1 a_277_47.t8 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR.t5 A2.t0 a_27_297.t1 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297.t2 A3.t0 VPWR.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47.t0 B1.t0 a_27_297.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297.t6 A1.t0 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND.t3 a_277_47.t9 X.t7 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR.t9 A1.t1 a_27_297.t7 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND.t2 a_277_47.t10 X.t6 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297.t0 A2.t1 VPWR.t6 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47.t0 A2.t2 a_109_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_361_47.t1 A1.t2 a_277_47.t4 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 X.t5 a_277_47.t11 VGND.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND.t5 A3.t1 a_445_47.t1 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X15 X.t4 a_277_47.t12 VGND.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X16 a_277_47.t5 A1.t3 a_193_47.t1 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_445_47.t0 A2.t3 a_361_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND.t7 B1.t1 a_277_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297.t4 B1.t2 a_277_47.t2 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR.t7 A3.t2 a_27_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR.t0 a_277_47.t13 X.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47.t1 A3.t3 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47.t3 B1.t3 VGND.t6 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
R0 a_277_47.n13 a_277_47.n11 318.272
R1 a_277_47.n15 a_277_47.n14 299.82
R2 a_277_47.n2 a_277_47.t13 212.081
R3 a_277_47.n1 a_277_47.t7 212.081
R4 a_277_47.n6 a_277_47.t6 212.081
R5 a_277_47.n8 a_277_47.t8 212.081
R6 a_277_47.n10 a_277_47.n9 152
R7 a_277_47.n7 a_277_47.n0 152
R8 a_277_47.n5 a_277_47.n4 152
R9 a_277_47.n2 a_277_47.t9 139.78
R10 a_277_47.n1 a_277_47.t11 139.78
R11 a_277_47.n6 a_277_47.t10 139.78
R12 a_277_47.n8 a_277_47.t12 139.78
R13 a_277_47.n13 a_277_47.n12 102.272
R14 a_277_47.n4 a_277_47.n3 88.8951
R15 a_277_47.n14 a_277_47.n10 78.8882
R16 a_277_47.n9 a_277_47.n7 49.6611
R17 a_277_47.n14 a_277_47.n13 48.4343
R18 a_277_47.n3 a_277_47.n1 42.5272
R19 a_277_47.n6 a_277_47.n5 40.8975
R20 a_277_47.n15 a_277_47.t2 26.5955
R21 a_277_47.t0 a_277_47.n15 26.5955
R22 a_277_47.n12 a_277_47.t1 24.9236
R23 a_277_47.n12 a_277_47.t3 24.9236
R24 a_277_47.n11 a_277_47.t4 24.9236
R25 a_277_47.n11 a_277_47.t5 24.9236
R26 a_277_47.n5 a_277_47.n1 20.449
R27 a_277_47.n3 a_277_47.n2 16.0056
R28 a_277_47.n4 a_277_47.n0 13.1884
R29 a_277_47.n10 a_277_47.n0 13.1884
R30 a_277_47.n7 a_277_47.n6 8.76414
R31 a_277_47.n9 a_277_47.n8 2.92171
R32 X.n2 X.n1 362.101
R33 X.n2 X.n0 298.853
R34 X.n5 X.n3 248.248
R35 X.n5 X.n4 185
R36 X X.n2 45.5534
R37 X X.n5 45.5534
R38 X.n1 X.t3 26.5955
R39 X.n1 X.t1 26.5955
R40 X.n0 X.t0 26.5955
R41 X.n0 X.t2 26.5955
R42 X.n3 X.t6 24.9236
R43 X.n3 X.t4 24.9236
R44 X.n4 X.t7 24.9236
R45 X.n4 X.t5 24.9236
R46 X X.n6 21.0829
R47 X.n6 X 6.4005
R48 X.n6 X 4.51815
R49 VPWR.n13 VPWR.t1 775.264
R50 VPWR.n10 VPWR.t0 698.62
R51 VPWR.n25 VPWR.n1 604.783
R52 VPWR.n23 VPWR.n3 604.783
R53 VPWR.n5 VPWR.n4 604.783
R54 VPWR.n11 VPWR.n9 604.783
R55 VPWR.n4 VPWR.t4 38.4155
R56 VPWR.n17 VPWR.n7 34.6358
R57 VPWR.n18 VPWR.n17 34.6358
R58 VPWR.n19 VPWR.n18 34.6358
R59 VPWR.n13 VPWR.n12 30.4946
R60 VPWR.n23 VPWR.n22 28.9887
R61 VPWR.n1 VPWR.t6 26.5955
R62 VPWR.n1 VPWR.t7 26.5955
R63 VPWR.n3 VPWR.t8 26.5955
R64 VPWR.n3 VPWR.t9 26.5955
R65 VPWR.n4 VPWR.t5 26.5955
R66 VPWR.n9 VPWR.t2 26.5955
R67 VPWR.n9 VPWR.t3 26.5955
R68 VPWR.n25 VPWR.n24 22.9652
R69 VPWR.n24 VPWR.n23 15.4358
R70 VPWR.n13 VPWR.n7 13.9299
R71 VPWR.n22 VPWR.n5 9.41227
R72 VPWR.n12 VPWR.n8 9.3005
R73 VPWR.n14 VPWR.n13 9.3005
R74 VPWR.n15 VPWR.n7 9.3005
R75 VPWR.n17 VPWR.n16 9.3005
R76 VPWR.n18 VPWR.n6 9.3005
R77 VPWR.n20 VPWR.n19 9.3005
R78 VPWR.n22 VPWR.n21 9.3005
R79 VPWR.n23 VPWR.n2 9.3005
R80 VPWR.n24 VPWR.n0 9.3005
R81 VPWR.n11 VPWR.n10 8.39785
R82 VPWR.n12 VPWR.n11 7.90638
R83 VPWR.n26 VPWR.n25 7.12063
R84 VPWR.n10 VPWR.n8 1.18757
R85 VPWR.n19 VPWR.n5 0.376971
R86 VPWR.n26 VPWR.n0 0.148519
R87 VPWR.n14 VPWR.n8 0.120292
R88 VPWR.n15 VPWR.n14 0.120292
R89 VPWR.n16 VPWR.n15 0.120292
R90 VPWR.n16 VPWR.n6 0.120292
R91 VPWR.n20 VPWR.n6 0.120292
R92 VPWR.n21 VPWR.n20 0.120292
R93 VPWR.n21 VPWR.n2 0.120292
R94 VPWR.n2 VPWR.n0 0.120292
R95 VPWR VPWR.n26 0.11354
R96 VPB.t8 VPB.t1 556.386
R97 VPB.t4 VPB.t5 284.113
R98 VPB.t6 VPB.t4 284.113
R99 VPB.t2 VPB.t0 248.599
R100 VPB.t3 VPB.t2 248.599
R101 VPB.t1 VPB.t3 248.599
R102 VPB.t5 VPB.t8 248.599
R103 VPB.t10 VPB.t6 248.599
R104 VPB.t11 VPB.t10 248.599
R105 VPB.t7 VPB.t11 248.599
R106 VPB.t9 VPB.t7 248.599
R107 VPB VPB.t9 189.409
R108 A2.n2 A2.n1 250.544
R109 A2.n1 A2.t1 241.536
R110 A2.n0 A2.t0 241.536
R111 A2.n1 A2.t2 169.237
R112 A2.n0 A2.t3 169.237
R113 A2.n3 A2.n0 156.8
R114 A2.n3 A2.n2 17.6437
R115 A2 A2.n3 5.4405
R116 A2.n2 A2 3.80591
R117 a_27_297.n1 a_27_297.t4 401.041
R118 a_27_297.n3 a_27_297.t5 388.695
R119 a_27_297.n3 a_27_297.n2 298.853
R120 a_27_297.n5 a_27_297.n4 298.853
R121 a_27_297.n1 a_27_297.n0 286.238
R122 a_27_297.n4 a_27_297.n1 84.8093
R123 a_27_297.n4 a_27_297.n3 63.2476
R124 a_27_297.n0 a_27_297.t2 38.4155
R125 a_27_297.n2 a_27_297.t7 26.5955
R126 a_27_297.n2 a_27_297.t0 26.5955
R127 a_27_297.n0 a_27_297.t3 26.5955
R128 a_27_297.t1 a_27_297.n5 26.5955
R129 a_27_297.n5 a_27_297.t6 26.5955
R130 A3 A3.n0 319.841
R131 A3.n0 A3.t0 241.536
R132 A3.n1 A3.t2 236.934
R133 A3.n0 A3.t1 169.237
R134 A3.n1 A3.t3 164.633
R135 A3.n2 A3.n1 152
R136 A3.n2 A3 9.7285
R137 A3 A3.n2 1.87783
R138 B1.n1 B1.t2 212.081
R139 B1.n0 B1.t0 212.081
R140 B1 B1.n1 196.091
R141 B1.n1 B1.t1 139.78
R142 B1.n0 B1.t3 139.78
R143 B1.n1 B1.n0 61.346
R144 A1.n0 A1.t0 221.72
R145 A1.n1 A1.t1 221.72
R146 A1 A1.n2 154.012
R147 A1.n0 A1.t2 149.421
R148 A1.n1 A1.t3 149.421
R149 A1.n2 A1.n0 37.4894
R150 A1.n2 A1.n1 37.4894
R151 VGND.n7 VGND.t3 279.55
R152 VGND.n21 VGND.n20 201.393
R153 VGND.n6 VGND.n5 200.516
R154 VGND.n14 VGND.n13 185
R155 VGND.n12 VGND.n11 185
R156 VGND.n29 VGND.t4 161.302
R157 VGND.n13 VGND.n12 66.462
R158 VGND.n12 VGND.t0 39.6928
R159 VGND.n13 VGND.t7 39.6928
R160 VGND.n10 VGND.n9 34.6358
R161 VGND.n19 VGND.n3 34.6358
R162 VGND.n23 VGND.n22 34.6358
R163 VGND.n23 VGND.n1 34.6358
R164 VGND.n27 VGND.n1 34.6358
R165 VGND.n28 VGND.n27 34.6358
R166 VGND.n29 VGND.n28 32.377
R167 VGND.n20 VGND.t5 32.3082
R168 VGND.n20 VGND.t6 28.6159
R169 VGND.n5 VGND.t1 24.9236
R170 VGND.n5 VGND.t2 24.9236
R171 VGND.n14 VGND.n3 23.1332
R172 VGND.n22 VGND.n21 12.8005
R173 VGND.n30 VGND.n29 11.5593
R174 VGND.n11 VGND.n10 9.58023
R175 VGND.n28 VGND.n0 9.3005
R176 VGND.n27 VGND.n26 9.3005
R177 VGND.n25 VGND.n1 9.3005
R178 VGND.n24 VGND.n23 9.3005
R179 VGND.n22 VGND.n2 9.3005
R180 VGND.n9 VGND.n8 9.3005
R181 VGND.n10 VGND.n4 9.3005
R182 VGND.n16 VGND.n15 9.3005
R183 VGND.n17 VGND.n3 9.3005
R184 VGND.n19 VGND.n18 9.3005
R185 VGND.n7 VGND.n6 8.39785
R186 VGND.n9 VGND.n6 7.90638
R187 VGND.n15 VGND.n11 5.31742
R188 VGND.n15 VGND.n14 1.77281
R189 VGND.n8 VGND.n7 1.18757
R190 VGND.n21 VGND.n19 0.376971
R191 VGND.n8 VGND.n4 0.120292
R192 VGND.n16 VGND.n4 0.120292
R193 VGND.n17 VGND.n16 0.120292
R194 VGND.n18 VGND.n17 0.120292
R195 VGND.n18 VGND.n2 0.120292
R196 VGND.n24 VGND.n2 0.120292
R197 VGND.n25 VGND.n24 0.120292
R198 VGND.n26 VGND.n25 0.120292
R199 VGND.n26 VGND.n0 0.120292
R200 VGND.n30 VGND.n0 0.120292
R201 VGND VGND.n30 0.0213333
R202 VNB.t9 VNB.t2 2677.02
R203 VNB.t7 VNB.t8 1366.99
R204 VNB.t0 VNB.t7 1366.99
R205 VNB.t3 VNB.t5 1196.12
R206 VNB.t4 VNB.t3 1196.12
R207 VNB.t2 VNB.t4 1196.12
R208 VNB.t8 VNB.t9 1196.12
R209 VNB.t11 VNB.t0 1196.12
R210 VNB.t10 VNB.t11 1196.12
R211 VNB.t1 VNB.t10 1196.12
R212 VNB.t6 VNB.t1 1196.12
R213 VNB VNB.t6 911.327
R214 a_109_47.t0 a_109_47.t1 49.8467
R215 a_193_47.t0 a_193_47.t1 49.8467
R216 a_361_47.t0 a_361_47.t1 49.8467
R217 a_445_47.t0 a_445_47.t1 60.9236
C0 A2 A1 0.190561f
C1 VPB VPWR 0.134195f
C2 A3 B1 0.054967f
C3 A3 VPWR 0.050448f
C4 A2 B1 3.8e-19
C5 VPB X 0.015356f
C6 A2 VPWR 0.032461f
C7 VPB VGND 0.012116f
C8 A3 VGND 0.063405f
C9 A1 VPWR 0.033174f
C10 A2 VGND 0.060083f
C11 B1 VPWR 0.019072f
C12 B1 X 0.005949f
C13 A1 VGND 0.021609f
C14 VPWR X 0.287347f
C15 B1 VGND 0.063769f
C16 VPB A3 0.073455f
C17 VPWR VGND 0.132425f
C18 VPB A2 0.052208f
C19 X VGND 0.145505f
C20 VPB A1 0.051082f
C21 A3 A2 0.225382f
C22 VPB B1 0.071503f
C23 A3 A1 0.048434f
C24 VGND VNB 0.771663f
C25 X VNB 0.077665f
C26 VPWR VNB 0.608678f
C27 B1 VNB 0.210582f
C28 A1 VNB 0.167132f
C29 A2 VNB 0.194857f
C30 A3 VNB 0.240522f
C31 VPB VNB 1.31353f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR VPB VNB A3 A2 A1 Y B1
X0 Y.t2 A1.t0 a_181_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 a_181_47.t0 A2.t0 a_109_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 VGND.t1 B1.t0 Y.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.105625 ps=0.975 w=0.65 l=0.15
X3 VPWR.t0 A2.t1 a_109_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 Y.t0 B1.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_109_297.t3 A1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X6 a_109_297.t2 A3.t0 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47.t0 A3.t1 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A1.n0 A1.t1 241.536
R1 A1 A1.n0 188.593
R2 A1.n0 A1.t0 169.237
R3 a_181_47.t0 a_181_47.t1 67.3851
R4 Y.n2 Y 593.216
R5 Y.n2 Y.n0 585
R6 Y.n3 Y.n2 585
R7 Y.n3 Y.n1 176.892
R8 Y.n1 Y.t1 35.0774
R9 Y.n2 Y.t0 28.5655
R10 Y.n1 Y.t2 24.9236
R11 Y Y.n0 8.21543
R12 Y Y.n0 4.77662
R13 Y Y.n3 4.77662
R14 VNB.t2 VNB.t3 1466.67
R15 VNB.t3 VNB.t1 1352.75
R16 VNB.t0 VNB.t2 1025.24
R17 VNB VNB.t0 911.327
R18 A2.n0 A2.t1 241.536
R19 A2.n0 A2.t0 169.237
R20 A2 A2.n0 153.583
R21 a_109_47.t0 a_109_47.t1 38.7697
R22 B1.n0 B1.t1 229.754
R23 B1.n0 B1.t0 157.453
R24 B1 B1.n0 154.91
R25 VGND.n0 VGND.t1 283.457
R26 VGND.n0 VGND.t0 156.424
R27 VGND VGND.n0 0.075072
R28 a_109_297.n1 a_109_297.n0 1265.99
R29 a_109_297.t0 a_109_297.n1 37.4305
R30 a_109_297.n0 a_109_297.t1 26.5955
R31 a_109_297.n0 a_109_297.t2 26.5955
R32 a_109_297.n1 a_109_297.t3 26.5955
R33 VPWR.n1 VPWR.n0 605.063
R34 VPWR.n1 VPWR.t1 249.919
R35 VPWR.n0 VPWR.t2 33.4905
R36 VPWR.n0 VPWR.t0 26.5955
R37 VPWR VPWR.n1 0.550712
R38 VPB.t3 VPB.t0 281.154
R39 VPB.t1 VPB.t3 269.315
R40 VPB.t2 VPB.t1 248.599
R41 VPB VPB.t2 189.409
R42 A3.n0 A3.t0 230.155
R43 A3.n0 A3.t1 157.856
R44 A3 A3.n0 155.685
C0 B1 Y 0.088202f
C1 A1 VGND 0.020244f
C2 VPWR Y 0.054494f
C3 B1 VGND 0.030992f
C4 VPB A3 0.037896f
C5 VPWR VGND 0.05116f
C6 VPB A2 0.02628f
C7 Y VGND 0.079497f
C8 A3 A2 0.088858f
C9 VPB A1 0.030533f
C10 A3 A1 0.002561f
C11 VPB B1 0.039111f
C12 A2 A1 0.079352f
C13 VPB VPWR 0.057476f
C14 A3 VPWR 0.054344f
C15 VPB Y 0.012212f
C16 A3 Y 2.43e-19
C17 A1 B1 0.048219f
C18 A2 VPWR 0.020535f
C19 VPB VGND 0.005776f
C20 A2 Y 0.033818f
C21 A3 VGND 0.049571f
C22 A1 VPWR 0.026688f
C23 A1 Y 0.074326f
C24 A2 VGND 0.095109f
C25 B1 VPWR 0.013695f
C26 VGND VNB 0.34044f
C27 Y VNB 0.059409f
C28 VPWR VNB 0.28219f
C29 B1 VNB 0.147606f
C30 A1 VNB 0.094864f
C31 A2 VNB 0.098148f
C32 A3 VNB 0.145026f
C33 VPB VNB 0.516168f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_2 VNB VPB VPWR VGND B1 Y A1 A2 A3
X0 VGND.t3 B1.t0 Y.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR.t3 A1.t0 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297.t5 B1.t1 Y.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47.t3 A1.t1 Y.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR.t1 A2.t1 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297.t6 A3.t0 VPWR.t4 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47.t3 A3.t1 VGND.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47.t1 A2.t2 a_277_47.t0 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297.t2 A1.t2 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y.t4 B1.t2 a_27_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47.t1 A2.t3 a_27_47.t0 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y.t2 B1.t3 VGND.t2 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X13 Y.t0 A1.t3 a_277_47.t2 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR.t5 A3.t2 a_27_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND.t0 A3.t3 a_27_47.t2 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 B1.n4 B1.t1 212.081
R1 B1.n1 B1.t2 212.081
R2 B1.n5 B1.n4 180.482
R3 B1.n3 B1.n2 152
R4 B1.n4 B1.t3 139.78
R5 B1.n1 B1.t0 139.78
R6 B1.n3 B1.n1 51.852
R7 B1.n4 B1.n3 21.1793
R8 B1.n2 B1.n0 17.9205
R9 B1.n0 B1 15.3605
R10 B1.n2 B1 10.5605
R11 B1 B1.n5 3.12939
R12 B1.n5 B1.n0 0.853833
R13 Y.n1 Y.t1 327.937
R14 Y Y.n0 317.591
R15 Y.n1 Y.t2 182.994
R16 Y.n3 Y.n2 97.3
R17 Y.n0 Y.t4 42.3555
R18 Y.n2 Y.t3 39.6928
R19 Y.n2 Y.t0 26.7697
R20 Y.n0 Y.t5 26.5955
R21 Y Y.n3 0.587757
R22 Y.n3 Y.n1 0.428431
R23 VGND.n2 VGND.n0 206.22
R24 VGND.n2 VGND.n1 205.488
R25 VGND.n0 VGND.t2 39.6928
R26 VGND.n0 VGND.t3 24.9236
R27 VGND.n1 VGND.t1 24.9236
R28 VGND.n1 VGND.t0 24.9236
R29 VGND VGND.n2 0.147009
R30 VNB.t6 VNB.t3 2677.02
R31 VNB.t1 VNB.t5 1452.43
R32 VNB.t5 VNB.t4 1423.95
R33 VNB.t3 VNB.t1 1281.55
R34 VNB.t7 VNB.t6 1196.12
R35 VNB.t2 VNB.t7 1196.12
R36 VNB.t0 VNB.t2 1196.12
R37 VNB VNB.t0 911.327
R38 A1.n3 A1.t0 212.081
R39 A1.n0 A1.t2 212.081
R40 A1 A1.n2 154.272
R41 A1.n4 A1.n3 152
R42 A1.n0 A1.t3 139.78
R43 A1.n1 A1.t1 139.78
R44 A1.n1 A1.n0 65.7278
R45 A1.n3 A1.n2 62.8066
R46 A1.n2 A1.n1 13.146
R47 A1 A1.n4 6.60695
R48 A1.n4 A1 3.30373
R49 a_27_297.t5 a_27_297.n5 407.067
R50 a_27_297.n2 a_27_297.t7 388.695
R51 a_27_297.n2 a_27_297.n1 298.853
R52 a_27_297.n3 a_27_297.n0 298.853
R53 a_27_297.n5 a_27_297.n4 286.238
R54 a_27_297.n5 a_27_297.n3 123.963
R55 a_27_297.n3 a_27_297.n2 63.2476
R56 a_27_297.n4 a_27_297.t2 44.3255
R57 a_27_297.n1 a_27_297.t1 26.5955
R58 a_27_297.n1 a_27_297.t6 26.5955
R59 a_27_297.n0 a_27_297.t3 26.5955
R60 a_27_297.n0 a_27_297.t0 26.5955
R61 a_27_297.n4 a_27_297.t4 26.5955
R62 VPWR.n12 VPWR.n1 604.783
R63 VPWR.n10 VPWR.n3 604.783
R64 VPWR.n7 VPWR.n6 587.37
R65 VPWR.n5 VPWR.n4 585
R66 VPWR.n6 VPWR.n5 66.9805
R67 VPWR.n5 VPWR.t3 49.2505
R68 VPWR.n6 VPWR.t2 45.3105
R69 VPWR.n10 VPWR.n9 28.9887
R70 VPWR.n1 VPWR.t4 26.5955
R71 VPWR.n1 VPWR.t5 26.5955
R72 VPWR.n3 VPWR.t0 26.5955
R73 VPWR.n3 VPWR.t1 26.5955
R74 VPWR.n12 VPWR.n11 22.9652
R75 VPWR.n9 VPWR.n4 21.177
R76 VPWR.n11 VPWR.n10 15.4358
R77 VPWR.n9 VPWR.n8 9.3005
R78 VPWR.n10 VPWR.n2 9.3005
R79 VPWR.n11 VPWR.n0 9.3005
R80 VPWR.n13 VPWR.n12 7.12063
R81 VPWR.n8 VPWR.n7 4.22922
R82 VPWR.n7 VPWR.n4 2.9355
R83 VPWR.n13 VPWR.n0 0.148519
R84 VPWR.n8 VPWR.n2 0.120292
R85 VPWR.n2 VPWR.n0 0.120292
R86 VPWR VPWR.n13 0.11354
R87 VPB.t3 VPB.t2 574.144
R88 VPB.t2 VPB.t4 301.87
R89 VPB.t4 VPB.t5 295.95
R90 VPB.t0 VPB.t3 248.599
R91 VPB.t1 VPB.t0 248.599
R92 VPB.t6 VPB.t1 248.599
R93 VPB.t7 VPB.t6 248.599
R94 VPB VPB.t7 189.409
R95 A2.n2 A2.t1 212.081
R96 A2.n0 A2.t0 212.081
R97 A2 A2.n1 154.891
R98 A2.n3 A2.n2 152
R99 A2.n2 A2.t3 139.78
R100 A2.n0 A2.t2 139.78
R101 A2.n2 A2.n1 52.5823
R102 A2.n1 A2.n0 8.76414
R103 A2.n3 A2 4.95534
R104 A2 A2.n3 4.54244
R105 a_277_47.n1 a_277_47.n0 474.659
R106 a_277_47.n1 a_277_47.t3 30.462
R107 a_277_47.n0 a_277_47.t0 24.9236
R108 a_277_47.n0 a_277_47.t1 24.9236
R109 a_277_47.t2 a_277_47.n1 24.9236
R110 A3.n1 A3.t0 212.081
R111 A3.n2 A3.t2 212.081
R112 A3.n2 A3.n0 184.864
R113 A3.n4 A3.n3 152
R114 A3.n1 A3.t1 139.78
R115 A3.n2 A3.t3 139.78
R116 A3.n3 A3.n1 41.6278
R117 A3.n3 A3.n2 19.7187
R118 A3.n4 A3.n0 7.43276
R119 A3.n0 A3 1.96179
R120 A3 A3.n4 0.103726
R121 a_27_47.n1 a_27_47.t2 331.325
R122 a_27_47.t1 a_27_47.n1 331.325
R123 a_27_47.n1 a_27_47.n0 185
R124 a_27_47.n0 a_27_47.t0 24.9236
R125 a_27_47.n0 a_27_47.t3 24.9236
C0 A1 Y 0.118427f
C1 A2 VGND 0.024575f
C2 B1 VPWR 0.021777f
C3 B1 Y 0.176713f
C4 A1 VGND 0.028066f
C5 VPWR Y 0.019647f
C6 B1 VGND 0.034395f
C7 VPB A3 0.073055f
C8 VPWR VGND 0.091425f
C9 VPB A2 0.056781f
C10 Y VGND 0.168059f
C11 A3 A2 0.106345f
C12 VPB A1 0.097086f
C13 VPB B1 0.080838f
C14 A2 A1 0.096461f
C15 VPB VPWR 0.088451f
C16 A3 VPWR 0.041498f
C17 VPB Y 0.007792f
C18 A3 Y 3.4e-19
C19 A1 B1 0.038222f
C20 A2 VPWR 0.039623f
C21 VPB VGND 0.005754f
C22 A3 VGND 0.035547f
C23 A2 Y 7.37e-19
C24 A1 VPWR 0.047505f
C25 VGND VNB 0.538381f
C26 Y VNB 0.060039f
C27 VPWR VNB 0.43614f
C28 B1 VNB 0.257598f
C29 A1 VNB 0.240167f
C30 A2 VNB 0.178539f
C31 A3 VNB 0.246114f
C32 VPB VNB 0.959148f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_4 VNB VPB VPWR VGND Y B1 A1 A2 A3
X0 a_27_47.t3 A2.t0 a_445_47.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47.t2 A2.t1 a_445_47.t2 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR.t7 A1.t0 a_27_297.t7 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297.t6 A1.t1 VPWR.t6 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297.t8 B1.t0 Y.t3 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t3 A2.t2 a_27_297.t3 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297.t5 A1.t2 VPWR.t5 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_297.t10 A3.t0 VPWR.t8 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR.t4 A1.t3 a_27_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X9 Y.t2 B1.t1 a_27_297.t9 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_297.t14 B1.t2 Y.t1 VPB.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_445_47.t4 A1.t4 Y.t11 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t9 A3.t1 a_27_297.t11 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y.t0 B1.t3 a_27_297.t12 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X14 a_445_47.t5 A1.t5 Y.t10 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VGND.t3 B1.t4 Y.t7 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_297.t13 A3.t2 VPWR.t10 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_47.t4 A3.t3 VGND.t7 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_47.t5 A3.t4 VGND.t6 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y.t9 A1.t6 a_445_47.t6 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_27_297.t2 A2.t3 VPWR.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X21 Y.t8 A1.t7 a_445_47.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y.t6 B1.t5 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y.t5 B1.t6 VGND.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VGND.t5 A3.t5 a_27_47.t6 VNB.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_445_47.t1 A2.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR.t1 A2.t5 a_27_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_445_47.t0 A2.t6 a_27_47.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_27_297.t0 A2.t7 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND.t0 B1.t7 Y.t4 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR.t11 A3.t6 a_27_297.t15 VPB.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 VGND.t4 A3.t7 a_27_47.t7 VNB.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A2.n1 A2.t3 212.081
R1 A2.n9 A2.t5 212.081
R2 A2.n2 A2.t7 212.081
R3 A2.n3 A2.t2 212.081
R4 A2.n11 A2.n10 152
R5 A2.n8 A2.n0 152
R6 A2.n7 A2.n6 152
R7 A2.n5 A2.n4 152
R8 A2.n1 A2.t1 139.78
R9 A2.n9 A2.t6 139.78
R10 A2.n2 A2.t0 139.78
R11 A2.n3 A2.t4 139.78
R12 A2.n8 A2.n7 54.0429
R13 A2.n4 A2.n2 52.5823
R14 A2.n10 A2.n9 48.2005
R15 A2.n11 A2.n0 14.352
R16 A2.n10 A2.n1 13.146
R17 A2.n6 A2 12.8005
R18 A2 A2.n5 9.30959
R19 A2.n4 A2.n3 8.76414
R20 A2.n5 A2 8.53383
R21 A2.n9 A2.n8 5.84292
R22 A2.n6 A2 5.04292
R23 A2 A2.n11 1.93989
R24 A2 A2.n0 1.55202
R25 A2.n7 A2.n2 1.46111
R26 a_445_47.n2 a_445_47.n0 248.248
R27 a_445_47.n4 a_445_47.n3 248.248
R28 a_445_47.n2 a_445_47.n1 185
R29 a_445_47.n5 a_445_47.n4 185
R30 a_445_47.n4 a_445_47.n2 102.4
R31 a_445_47.n3 a_445_47.t3 24.9236
R32 a_445_47.n3 a_445_47.t1 24.9236
R33 a_445_47.n1 a_445_47.t7 24.9236
R34 a_445_47.n1 a_445_47.t5 24.9236
R35 a_445_47.n0 a_445_47.t6 24.9236
R36 a_445_47.n0 a_445_47.t4 24.9236
R37 a_445_47.n5 a_445_47.t2 24.9236
R38 a_445_47.t0 a_445_47.n5 24.9236
R39 a_27_47.n2 a_27_47.t7 329.051
R40 a_27_47.n4 a_27_47.t2 322.094
R41 a_27_47.n2 a_27_47.n1 201.189
R42 a_27_47.n3 a_27_47.n0 201.189
R43 a_27_47.n5 a_27_47.n4 185
R44 a_27_47.n4 a_27_47.n3 63.2476
R45 a_27_47.n3 a_27_47.n2 63.2476
R46 a_27_47.n1 a_27_47.t6 24.9236
R47 a_27_47.n1 a_27_47.t4 24.9236
R48 a_27_47.n0 a_27_47.t1 24.9236
R49 a_27_47.n0 a_27_47.t5 24.9236
R50 a_27_47.n5 a_27_47.t0 24.9236
R51 a_27_47.t3 a_27_47.n5 24.9236
R52 VNB.t2 VNB.t9 2677.02
R53 VNB.t7 VNB.t6 1196.12
R54 VNB.t5 VNB.t7 1196.12
R55 VNB.t4 VNB.t5 1196.12
R56 VNB.t10 VNB.t4 1196.12
R57 VNB.t8 VNB.t10 1196.12
R58 VNB.t11 VNB.t8 1196.12
R59 VNB.t9 VNB.t11 1196.12
R60 VNB.t0 VNB.t2 1196.12
R61 VNB.t3 VNB.t0 1196.12
R62 VNB.t1 VNB.t3 1196.12
R63 VNB.t13 VNB.t1 1196.12
R64 VNB.t14 VNB.t13 1196.12
R65 VNB.t12 VNB.t14 1196.12
R66 VNB.t15 VNB.t12 1196.12
R67 VNB VNB.t15 911.327
R68 A1.n10 A1.t3 213.917
R69 A1.n3 A1.t1 205.654
R70 A1.n7 A1.t0 205.654
R71 A1.n11 A1.t2 205.654
R72 A1.n2 A1.t6 204.049
R73 A1.n5 A1.n4 152
R74 A1.n8 A1.n0 152
R75 A1.n13 A1.n12 152
R76 A1.n10 A1.n1 152
R77 A1.n2 A1.t4 150.754
R78 A1.n9 A1.t5 139.78
R79 A1.n6 A1.t7 139.78
R80 A1.n11 A1.n10 49.5776
R81 A1.n9 A1.n8 41.3148
R82 A1.n6 A1.n5 34.4291
R83 A1.n13 A1.n1 14.352
R84 A1 A1.n0 13.1884
R85 A1.n5 A1.n3 12.3948
R86 A1.n7 A1.n6 11.0176
R87 A1.n4 A1 9.69747
R88 A1.n12 A1.n9 9.6405
R89 A1.n4 A1 8.14595
R90 A1.n3 A1.n2 6.55122
R91 A1.n8 A1.n7 5.50907
R92 A1 A1.n0 4.65505
R93 A1.n1 A1 2.32777
R94 A1.n12 A1.n11 1.37764
R95 A1 A1.n13 1.16414
R96 a_27_297.n3 a_27_297.n2 585
R97 a_27_297.n10 a_27_297.t15 410.818
R98 a_27_297.n6 a_27_297.n1 320.976
R99 a_27_297.n7 a_27_297.n0 320.976
R100 a_27_297.n11 a_27_297.n8 320.976
R101 a_27_297.n10 a_27_297.n9 320.976
R102 a_27_297.n13 a_27_297.n12 320.976
R103 a_27_297.n3 a_27_297.t8 287.853
R104 a_27_297.n5 a_27_297.n4 284.18
R105 a_27_297.n4 a_27_297.t12 125.096
R106 a_27_297.n5 a_27_297.n3 117.537
R107 a_27_297.n6 a_27_297.n5 90.0549
R108 a_27_297.n7 a_27_297.n6 64.7534
R109 a_27_297.n12 a_27_297.n7 63.2476
R110 a_27_297.n12 a_27_297.n11 63.2476
R111 a_27_297.n11 a_27_297.n10 63.2476
R112 a_27_297.n0 a_27_297.t4 30.5355
R113 a_27_297.n4 a_27_297.t6 26.5955
R114 a_27_297.n2 a_27_297.t9 26.5955
R115 a_27_297.n2 a_27_297.t14 26.5955
R116 a_27_297.n1 a_27_297.t7 26.5955
R117 a_27_297.n1 a_27_297.t5 26.5955
R118 a_27_297.n0 a_27_297.t2 26.5955
R119 a_27_297.n8 a_27_297.t3 26.5955
R120 a_27_297.n8 a_27_297.t10 26.5955
R121 a_27_297.n9 a_27_297.t11 26.5955
R122 a_27_297.n9 a_27_297.t13 26.5955
R123 a_27_297.n13 a_27_297.t1 26.5955
R124 a_27_297.t0 a_27_297.n13 26.5955
R125 VPWR.n11 VPWR.n10 605.029
R126 VPWR.n20 VPWR.n3 310.502
R127 VPWR.n5 VPWR.n4 310.502
R128 VPWR.n14 VPWR.n7 310.502
R129 VPWR.n9 VPWR.n8 310.502
R130 VPWR.n22 VPWR.n1 310.5
R131 VPWR.n16 VPWR.n15 34.6358
R132 VPWR.n13 VPWR.n9 33.5064
R133 VPWR.n20 VPWR.n19 28.9887
R134 VPWR.n1 VPWR.t10 26.5955
R135 VPWR.n1 VPWR.t11 26.5955
R136 VPWR.n3 VPWR.t8 26.5955
R137 VPWR.n3 VPWR.t9 26.5955
R138 VPWR.n4 VPWR.t0 26.5955
R139 VPWR.n4 VPWR.t3 26.5955
R140 VPWR.n7 VPWR.t2 26.5955
R141 VPWR.n7 VPWR.t1 26.5955
R142 VPWR.n8 VPWR.t5 26.5955
R143 VPWR.n8 VPWR.t4 26.5955
R144 VPWR.n10 VPWR.t6 26.5955
R145 VPWR.n10 VPWR.t7 26.5955
R146 VPWR.n22 VPWR.n21 22.9652
R147 VPWR.n21 VPWR.n20 15.4358
R148 VPWR.n19 VPWR.n5 9.41227
R149 VPWR.n13 VPWR.n12 9.3005
R150 VPWR.n15 VPWR.n6 9.3005
R151 VPWR.n17 VPWR.n16 9.3005
R152 VPWR.n19 VPWR.n18 9.3005
R153 VPWR.n20 VPWR.n2 9.3005
R154 VPWR.n21 VPWR.n0 9.3005
R155 VPWR.n23 VPWR.n22 7.12063
R156 VPWR.n14 VPWR.n13 6.4005
R157 VPWR.n11 VPWR.n9 5.64089
R158 VPWR.n15 VPWR.n14 3.38874
R159 VPWR.n12 VPWR.n11 0.653702
R160 VPWR.n16 VPWR.n5 0.376971
R161 VPWR.n23 VPWR.n0 0.148519
R162 VPWR.n12 VPWR.n6 0.120292
R163 VPWR.n17 VPWR.n6 0.120292
R164 VPWR.n18 VPWR.n17 0.120292
R165 VPWR.n18 VPWR.n2 0.120292
R166 VPWR.n2 VPWR.n0 0.120292
R167 VPWR VPWR.n23 0.11354
R168 VPB.t6 VPB.t12 544.548
R169 VPB.t2 VPB.t4 260.437
R170 VPB.t9 VPB.t8 248.599
R171 VPB.t14 VPB.t9 248.599
R172 VPB.t12 VPB.t14 248.599
R173 VPB.t7 VPB.t6 248.599
R174 VPB.t5 VPB.t7 248.599
R175 VPB.t4 VPB.t5 248.599
R176 VPB.t1 VPB.t2 248.599
R177 VPB.t0 VPB.t1 248.599
R178 VPB.t3 VPB.t0 248.599
R179 VPB.t10 VPB.t3 248.599
R180 VPB.t11 VPB.t10 248.599
R181 VPB.t13 VPB.t11 248.599
R182 VPB.t15 VPB.t13 248.599
R183 VPB VPB.t15 189.409
R184 B1.n6 B1.t3 212.081
R185 B1.n1 B1.t0 212.081
R186 B1.n2 B1.t1 212.081
R187 B1.n0 B1.t2 212.081
R188 B1 B1.n3 155.226
R189 B1.n5 B1.n4 152
R190 B1.n7 B1.n6 152
R191 B1.n6 B1.t4 139.78
R192 B1.n1 B1.t6 139.78
R193 B1.n2 B1.t7 139.78
R194 B1.n0 B1.t5 139.78
R195 B1.n2 B1.n1 61.346
R196 B1.n6 B1.n5 54.0429
R197 B1.n3 B1.n0 46.7399
R198 B1.n3 B1.n2 14.6066
R199 B1.n5 B1.n0 7.30353
R200 B1 B1.n7 6.85404
R201 B1.n4 B1 5.03987
R202 B1.n4 B1 4.23357
R203 B1.n7 B1 2.4194
R204 Y.n2 Y.n0 645.612
R205 Y.n2 Y.n1 585
R206 Y.n5 Y.t10 322.094
R207 Y.n9 Y.t5 272.889
R208 Y.n8 Y.n3 201.189
R209 Y.n7 Y.n6 185
R210 Y.n5 Y.n4 185
R211 Y.n8 Y.n7 63.2476
R212 Y.n7 Y.n5 63.2476
R213 Y.n9 Y.n8 28.9887
R214 Y.n1 Y.t3 26.5955
R215 Y.n1 Y.t2 26.5955
R216 Y.n0 Y.t1 26.5955
R217 Y.n0 Y.t0 26.5955
R218 Y.n4 Y.t11 24.9236
R219 Y.n4 Y.t8 24.9236
R220 Y.n6 Y.t7 24.9236
R221 Y.n6 Y.t9 24.9236
R222 Y.n3 Y.t4 24.9236
R223 Y.n3 Y.t6 24.9236
R224 Y Y.n2 13.7605
R225 Y Y.n9 2.8805
R226 A3.n1 A3.t0 212.081
R227 A3.n4 A3.t1 212.081
R228 A3.n0 A3.t2 212.081
R229 A3.n9 A3.t6 212.081
R230 A3.n10 A3.n9 179.022
R231 A3.n3 A3.n2 152
R232 A3.n6 A3.n5 152
R233 A3.n8 A3.n7 152
R234 A3.n1 A3.t4 139.78
R235 A3.n4 A3.t5 139.78
R236 A3.n0 A3.t3 139.78
R237 A3.n9 A3.t7 139.78
R238 A3.n3 A3.n1 48.9308
R239 A3.n5 A3.n4 41.6278
R240 A3.n8 A3.n0 34.3247
R241 A3.n9 A3.n8 27.0217
R242 A3.n5 A3.n0 19.7187
R243 A3.n7 A3.n6 14.352
R244 A3.n2 A3 12.6066
R245 A3.n10 A3 12.6066
R246 A3.n4 A3.n3 12.4157
R247 A3.n2 A3 5.23686
R248 A3 A3.n10 5.23686
R249 A3.n6 A3 1.74595
R250 A3.n7 A3 1.74595
R251 VGND.n10 VGND.n7 205.096
R252 VGND.n9 VGND.n8 199.739
R253 VGND.n25 VGND.n2 199.739
R254 VGND.n28 VGND.n27 199.739
R255 VGND.n13 VGND.n6 34.6358
R256 VGND.n14 VGND.n13 34.6358
R257 VGND.n15 VGND.n14 34.6358
R258 VGND.n15 VGND.n4 34.6358
R259 VGND.n19 VGND.n4 34.6358
R260 VGND.n20 VGND.n19 34.6358
R261 VGND.n21 VGND.n20 34.6358
R262 VGND.n21 VGND.n1 34.6358
R263 VGND.n25 VGND.n1 28.9887
R264 VGND.n7 VGND.t1 24.9236
R265 VGND.n7 VGND.t0 24.9236
R266 VGND.n8 VGND.t2 24.9236
R267 VGND.n8 VGND.t3 24.9236
R268 VGND.n2 VGND.t6 24.9236
R269 VGND.n2 VGND.t5 24.9236
R270 VGND.n27 VGND.t7 24.9236
R271 VGND.n27 VGND.t4 24.9236
R272 VGND.n9 VGND.n6 24.4711
R273 VGND.n28 VGND.n26 22.9652
R274 VGND.n26 VGND.n25 15.4358
R275 VGND.n11 VGND.n6 9.3005
R276 VGND.n13 VGND.n12 9.3005
R277 VGND.n14 VGND.n5 9.3005
R278 VGND.n16 VGND.n15 9.3005
R279 VGND.n17 VGND.n4 9.3005
R280 VGND.n19 VGND.n18 9.3005
R281 VGND.n20 VGND.n3 9.3005
R282 VGND.n22 VGND.n21 9.3005
R283 VGND.n23 VGND.n1 9.3005
R284 VGND.n25 VGND.n24 9.3005
R285 VGND.n26 VGND.n0 9.3005
R286 VGND.n29 VGND.n28 7.12063
R287 VGND.n10 VGND.n9 6.37482
R288 VGND.n11 VGND.n10 0.658988
R289 VGND.n29 VGND.n0 0.148519
R290 VGND.n12 VGND.n11 0.120292
R291 VGND.n12 VGND.n5 0.120292
R292 VGND.n16 VGND.n5 0.120292
R293 VGND.n17 VGND.n16 0.120292
R294 VGND.n18 VGND.n17 0.120292
R295 VGND.n18 VGND.n3 0.120292
R296 VGND.n22 VGND.n3 0.120292
R297 VGND.n23 VGND.n22 0.120292
R298 VGND.n24 VGND.n23 0.120292
R299 VGND.n24 VGND.n0 0.120292
R300 VGND VGND.n29 0.11354
C0 A3 VGND 0.070001f
C1 A2 Y 2.1e-19
C2 A1 VPWR 0.074227f
C3 A1 Y 0.146396f
C4 B1 VPWR 0.040174f
C5 A2 VGND 0.035952f
C6 A1 VGND 0.042759f
C7 B1 Y 0.297699f
C8 B1 VGND 0.068854f
C9 VPWR Y 0.022237f
C10 VPB A3 0.134098f
C11 VPWR VGND 0.152442f
C12 VPB A2 0.116743f
C13 Y VGND 0.245405f
C14 A3 A2 0.078238f
C15 VPB A1 0.144401f
C16 VPB B1 0.134627f
C17 VPB VPWR 0.14435f
C18 A3 B1 8.72e-20
C19 A2 A1 0.060707f
C20 A3 VPWR 0.084451f
C21 VPB Y 0.005021f
C22 A2 B1 2.23e-19
C23 VPB VGND 0.011279f
C24 A3 Y 5.71e-20
C25 A2 VPWR 0.069156f
C26 A1 B1 0.076635f
C27 VGND VNB 0.849013f
C28 Y VNB 0.0689f
C29 VPWR VNB 0.709165f
C30 B1 VNB 0.386112f
C31 A1 VNB 0.406506f
C32 A2 VNB 0.359599f
C33 A3 VNB 0.420909f
C34 VPB VNB 1.57932f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21.t2 A1.t0 a_346_47.t1 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21.t1 B1.t0 a_250_297.t3 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47.t1 B1.t1 a_93_21.t3 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR.t2 a_93_21.t4 X.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND.t1 B2.t0 a_584_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47.t1 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297.t1 B2.t1 a_93_21.t0 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND.t2 a_93_21.t5 X.t0 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297.t0 A3.t1 VPWR.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR.t3 A2.t0 a_250_297.t4 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297.t2 A1.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47.t0 A2.t1 a_256_47.t0 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
R0 A1.n0 A1.t1 241.536
R1 A1.n0 A1.t0 169.237
R2 A1 A1.n0 154.429
R3 a_346_47.t0 a_346_47.t1 83.0774
R4 a_93_21.n3 a_93_21.n2 792.583
R5 a_93_21.n2 a_93_21.n0 349.666
R6 a_93_21.n1 a_93_21.t4 236.552
R7 a_93_21.n1 a_93_21.t5 164.251
R8 a_93_21.n2 a_93_21.n1 152
R9 a_93_21.n0 a_93_21.t3 41.539
R10 a_93_21.n0 a_93_21.t2 39.6928
R11 a_93_21.t0 a_93_21.n3 27.5805
R12 a_93_21.n3 a_93_21.t1 27.5805
R13 VNB.t4 VNB.t0 1893.85
R14 VNB.t2 VNB.t3 1708.74
R15 VNB.t3 VNB.t5 1680.26
R16 VNB.t0 VNB.t2 1281.55
R17 VNB VNB.t4 1110.68
R18 VNB.t5 VNB.t1 1025.24
R19 B1.n0 B1.t0 241.536
R20 B1.n0 B1.t1 169.237
R21 B1 B1.n0 153.677
R22 a_250_297.n1 a_250_297.t1 390.42
R23 a_250_297.n2 a_250_297.n1 365.33
R24 a_250_297.n1 a_250_297.n0 289.24
R25 a_250_297.n0 a_250_297.t3 37.4305
R26 a_250_297.n0 a_250_297.t2 35.4605
R27 a_250_297.n2 a_250_297.t4 32.5055
R28 a_250_297.t0 a_250_297.n2 32.5055
R29 VPB.t3 VPB.t0 375.858
R30 VPB.t5 VPB.t2 355.14
R31 VPB.t2 VPB.t4 307.788
R32 VPB.t0 VPB.t5 284.113
R33 VPB.t4 VPB.t1 254.518
R34 VPB VPB.t3 230.841
R35 a_584_47.t0 a_584_47.t1 38.7697
R36 X.n4 X 593.216
R37 X.n4 X.n3 585
R38 X.n5 X.n4 585
R39 X.n1 X 186.529
R40 X.n2 X.n1 185
R41 X.n4 X.t1 40.3855
R42 X.n1 X.t0 37.8467
R43 X.n3 X 10.7927
R44 X.n2 X.n0 8.28285
R45 X.n0 X 6.77697
R46 X.n6 X 6.52599
R47 X.n3 X 6.27501
R48 X X.n0 5.15871
R49 X X.n6 4.96766
R50 X.n5 X 4.77662
R51 X.n6 X.n5 3.24826
R52 X X.n2 2.00834
R53 VPWR.n2 VPWR.n0 605.413
R54 VPWR.n2 VPWR.n1 315.74
R55 VPWR.n1 VPWR.t0 51.2205
R56 VPWR.n1 VPWR.t2 44.3255
R57 VPWR.n0 VPWR.t1 44.3255
R58 VPWR.n0 VPWR.t3 44.3255
R59 VPWR VPWR.n2 0.292128
R60 B2.n0 B2.t1 241.536
R61 B2.n0 B2.t0 169.237
R62 B2.n1 B2.n0 152
R63 B2 B2.n1 13.5275
R64 B2.n1 B2 2.01193
R65 VGND.n1 VGND.n0 206.173
R66 VGND.n1 VGND.t1 156.615
R67 VGND.n0 VGND.t0 68.3082
R68 VGND.n0 VGND.t2 26.7697
R69 VGND VGND.n1 0.157741
R70 A3.n0 A3.t1 241.536
R71 A3.n0 A3.t0 169.237
R72 A3 A3.n0 158.4
R73 a_256_47.t0 a_256_47.t1 55.3851
R74 A2.n0 A2.t0 241.536
R75 A2.n0 A2.t1 169.237
R76 A2 A2.n0 154.607
C0 B1 B2 0.082331f
C1 A1 X 6.03e-20
C2 A2 VPWR 0.013294f
C3 A3 VGND 0.009742f
C4 A1 VPWR 0.015992f
C5 B1 X 3.83e-20
C6 A2 VGND 0.011437f
C7 A1 VGND 0.01333f
C8 B1 VPWR 0.010035f
C9 VPB A3 0.029118f
C10 B2 VPWR 0.010807f
C11 B1 VGND 0.034397f
C12 VPB A2 0.028677f
C13 X VPWR 0.084928f
C14 B2 VGND 0.046938f
C15 A3 A2 0.078809f
C16 VPB A1 0.029574f
C17 X VGND 0.059994f
C18 VPB B1 0.027632f
C19 VPWR VGND 0.075955f
C20 VPB B2 0.035517f
C21 A2 A1 0.09713f
C22 A3 B1 7.88e-22
C23 VPB X 0.010825f
C24 A3 B2 9.12e-20
C25 A2 B1 1.44e-20
C26 A3 X 2.45e-19
C27 VPB VPWR 0.075576f
C28 A1 B1 0.096524f
C29 A2 B2 1.46e-19
C30 A2 X 1.19e-19
C31 A3 VPWR 0.015799f
C32 A1 B2 3.14e-19
C33 VPB VGND 0.007881f
C34 VGND VNB 0.465075f
C35 VPWR VNB 0.364756f
C36 X VNB 0.093662f
C37 B2 VNB 0.140129f
C38 B1 VNB 0.100974f
C39 A1 VNB 0.095135f
C40 A2 VNB 0.092101f
C41 A3 VNB 0.092873f
C42 VPB VNB 0.781956f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_2 VNB VPB VGND VPWR X A3 A2 B2 B1 A1
X0 VPWR.t0 A3.t0 a_299_297.t0 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_299_297.t3 A2.t0 VPWR.t1 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_352_47.t0 B2.t0 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.209625 ps=1.295 w=0.65 l=0.15
X3 a_549_47.t0 A1.t0 a_21_199.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 X.t3 a_21_199.t4 VPWR.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND.t3 a_21_199.t5 X.t1 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.209625 pd=1.295 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47.t1 A2.t1 a_549_47.t1 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 VPWR.t2 A1.t1 a_299_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 a_299_297.t1 B1.t0 a_21_199.t2 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_21_199.t0 B2.t1 a_299_297.t2 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND.t1 A3.t1 a_665_47.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR.t4 a_21_199.t6 X.t2 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X.t0 a_21_199.t7 VGND.t2 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_21_199.t1 B1.t1 a_352_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
R0 A3.n0 A3.t0 230.155
R1 A3.n0 A3.t1 157.856
R2 A3.n1 A3.n0 152
R3 A3.n1 A3 15.2005
R4 A3 A3.n1 2.93383
R5 a_299_297.n1 a_299_297.t2 400.861
R6 a_299_297.n2 a_299_297.n1 386.134
R7 a_299_297.n1 a_299_297.n0 286.418
R8 a_299_297.n0 a_299_297.t4 26.5955
R9 a_299_297.n0 a_299_297.t1 26.5955
R10 a_299_297.t0 a_299_297.n2 26.5955
R11 a_299_297.n2 a_299_297.t3 26.5955
R12 VPWR.n12 VPWR.n1 604.783
R13 VPWR.n5 VPWR.n4 604.201
R14 VPWR.n3 VPWR.t0 343.481
R15 VPWR.n4 VPWR.t1 58.1155
R16 VPWR.n6 VPWR.n2 34.6358
R17 VPWR.n10 VPWR.n2 34.6358
R18 VPWR.n11 VPWR.n10 34.6358
R19 VPWR.n1 VPWR.t3 26.5955
R20 VPWR.n1 VPWR.t4 26.5955
R21 VPWR.n4 VPWR.t2 26.5955
R22 VPWR.n12 VPWR.n11 22.9652
R23 VPWR.n6 VPWR.n5 13.9299
R24 VPWR.n7 VPWR.n6 9.3005
R25 VPWR.n8 VPWR.n2 9.3005
R26 VPWR.n10 VPWR.n9 9.3005
R27 VPWR.n11 VPWR.n0 9.3005
R28 VPWR.n13 VPWR.n12 7.12063
R29 VPWR.n5 VPWR.n3 6.98769
R30 VPWR.n7 VPWR.n3 0.593044
R31 VPWR.n13 VPWR.n0 0.148519
R32 VPWR.n8 VPWR.n7 0.120292
R33 VPWR.n9 VPWR.n8 0.120292
R34 VPWR.n9 VPWR.n0 0.120292
R35 VPWR VPWR.n13 0.11354
R36 VPB.t5 VPB.t2 556.386
R37 VPB.t4 VPB.t3 343.303
R38 VPB.t3 VPB.t0 248.599
R39 VPB.t1 VPB.t4 248.599
R40 VPB.t2 VPB.t1 248.599
R41 VPB.t6 VPB.t5 248.599
R42 VPB VPB.t6 189.409
R43 A2.n0 A2.t0 241.536
R44 A2.n0 A2.t1 169.237
R45 A2.n1 A2.n0 152
R46 A2.n1 A2 11.9584
R47 A2 A2.n1 1.85313
R48 B2.n0 B2.t1 233.26
R49 B2 B2.n0 200.436
R50 B2.n0 B2.t0 139.78
R51 VGND.n9 VGND.t2 282.596
R52 VGND.n7 VGND.n6 185
R53 VGND.n5 VGND.n4 185
R54 VGND.n3 VGND.t1 156.953
R55 VGND.n6 VGND.n5 69.2313
R56 VGND.n5 VGND.t0 24.9236
R57 VGND.n6 VGND.t3 24.9236
R58 VGND.n8 VGND.n7 22.4325
R59 VGND.n9 VGND.n8 19.9534
R60 VGND.n4 VGND.n3 10.807
R61 VGND.n10 VGND.n9 9.3005
R62 VGND.n8 VGND.n0 9.3005
R63 VGND.n2 VGND.n1 9.3005
R64 VGND.n4 VGND.n1 7.84956
R65 VGND.n7 VGND.n1 1.20805
R66 VGND.n3 VGND.n2 0.150444
R67 VGND.n2 VGND.n0 0.120292
R68 VGND.n10 VGND.n0 0.120292
R69 VGND VGND.n10 0.0213333
R70 a_352_47.t0 a_352_47.t1 65.539
R71 VNB.t6 VNB.t0 2264.08
R72 VNB.t3 VNB.t4 1651.78
R73 VNB.t0 VNB.t2 1438.19
R74 VNB.t2 VNB.t3 1366.99
R75 VNB.t4 VNB.t1 1196.12
R76 VNB.t5 VNB.t6 1196.12
R77 VNB VNB.t5 911.327
R78 A1.n0 A1.t1 237.736
R79 A1.n1 A1.n0 185.512
R80 A1.n0 A1.t0 165.435
R81 A1 A1.n1 9.06717
R82 A1.n1 A1 4.73093
R83 a_21_199.n5 a_21_199.n4 313.736
R84 a_21_199.n4 a_21_199.n3 261.93
R85 a_21_199.n1 a_21_199.t4 212.081
R86 a_21_199.n2 a_21_199.t6 212.081
R87 a_21_199.n4 a_21_199.n0 173.357
R88 a_21_199.n1 a_21_199.t5 139.78
R89 a_21_199.n2 a_21_199.t7 139.78
R90 a_21_199.n3 a_21_199.n1 39.4369
R91 a_21_199.n0 a_21_199.t3 32.3082
R92 a_21_199.n0 a_21_199.t1 28.6159
R93 a_21_199.n5 a_21_199.t2 26.5955
R94 a_21_199.t0 a_21_199.n5 26.5955
R95 a_21_199.n3 a_21_199.n2 21.9096
R96 a_549_47.t0 a_549_47.t1 79.3851
R97 X.n0 X 595.668
R98 X.n1 X.n0 585
R99 X.n2 X.t3 382.296
R100 X X.n3 211.748
R101 X.n0 X.t2 26.5955
R102 X.n3 X.t1 24.9236
R103 X.n3 X.t0 24.9236
R104 X.n1 X 10.6672
R105 X X.n2 5.18145
R106 X.n2 X.n1 4.87669
R107 a_665_47.t0 a_665_47.t1 49.8467
R108 B1.n0 B1.t0 241.536
R109 B1 B1.n0 186.26
R110 B1.n0 B1.t1 169.237
C0 A2 VPWR 0.021079f
C1 A1 VGND 0.045479f
C2 VPB B2 0.050179f
C3 A2 VGND 0.071858f
C4 A3 VPWR 0.0436f
C5 VPB B1 0.028468f
C6 X VPWR 0.163132f
C7 A3 VGND 0.046816f
C8 VPB A1 0.030074f
C9 B2 B1 0.05353f
C10 X VGND 0.062548f
C11 B2 A1 2.33e-20
C12 VPB A2 0.030283f
C13 VPWR VGND 0.088767f
C14 B1 A1 0.081828f
C15 VPB A3 0.040792f
C16 VPB X 0.012534f
C17 B1 A2 0.009005f
C18 B1 A3 4.82e-21
C19 B2 X 0.010447f
C20 VPB VPWR 0.094904f
C21 A1 A2 0.113791f
C22 VPB VGND 0.009082f
C23 A1 A3 4.43e-20
C24 B2 VPWR 0.011087f
C25 B1 VPWR 0.011885f
C26 B2 VGND 0.054077f
C27 A2 A3 0.109993f
C28 A1 VPWR 0.020137f
C29 B1 VGND 0.013119f
C30 VGND VNB 0.519497f
C31 VPWR VNB 0.422561f
C32 X VNB 0.076859f
C33 A3 VNB 0.157082f
C34 A2 VNB 0.098913f
C35 A1 VNB 0.099001f
C36 B1 VNB 0.094195f
C37 B2 VNB 0.135553f
C38 VPB VNB 0.870552f
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_4 VNB VPB VGND VPWR X A3 A2 A1 B1 B2
X0 VGND.t1 A3.t0 a_445_47.t1 VNB.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_445_297.t6 A2.t0 VPWR.t7 VPB.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR.t6 A2.t1 a_445_297.t5 VPB.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_635_47.t2 A2.t2 a_445_47.t2 VNB.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_445_297.t2 A3.t1 VPWR.t1 VPB.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR.t2 a_79_21.t8 X.t3 VPB.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_297.t0 B2.t0 a_79_21.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_79_21.t6 B1.t0 a_1142_47.t1 VNB.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_79_21.t7 B2.t1 a_445_297.t9 VPB.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X.t2 a_79_21.t9 VPWR.t3 VPB.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_445_47.t3 A2.t3 a_635_47.t1 VNB.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_79_21.t5 A1.t0 a_635_47.t3 VNB.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR.t4 a_79_21.t10 X.t1 VPB.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_445_297.t3 B1.t1 a_79_21.t2 VPB.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND.t2 a_79_21.t11 X.t7 VNB.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND.t3 a_79_21.t12 X.t6 VNB.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_1142_47.t0 B1.t2 a_79_21.t3 VNB.t3 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND.t6 B2.t2 a_1142_47.t3 VNB.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X18 a_635_47.t0 A1.t1 a_79_21.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X.t5 a_79_21.t13 VGND.t4 VNB.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_445_47.t0 A3.t2 VGND.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_79_21.t4 B1.t3 a_445_297.t4 VPB.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.585 ps=2.17 w=1 l=0.15
X22 a_1142_47.t2 B2.t3 VGND.t7 VNB.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VPWR.t0 A3.t3 a_445_297.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 a_445_297.t7 A1.t2 VPWR.t8 VPB.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.585 pd=2.17 as=0.135 ps=1.27 w=1 l=0.15
X25 X.t0 a_79_21.t14 VPWR.t5 VPB.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 VPWR.t9 A1.t3 a_445_297.t8 VPB.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 X.t4 a_79_21.t15 VGND.t5 VNB.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 A3.n2 A3.t3 212.081
R1 A3.n0 A3.t1 212.081
R2 A3.n3 A3.n2 173.28
R3 A3.n1 A3 156.364
R4 A3.n2 A3.t0 139.78
R5 A3.n0 A3.t2 139.78
R6 A3.n1 A3.n0 32.8641
R7 A3.n2 A3.n1 28.4823
R8 A3.n3 A3 15.4187
R9 A3 A3.n3 11.346
R10 a_445_47.n1 a_445_47.n0 490.094
R11 a_445_47.n0 a_445_47.t2 24.9236
R12 a_445_47.n0 a_445_47.t3 24.9236
R13 a_445_47.n1 a_445_47.t1 24.9236
R14 a_445_47.t0 a_445_47.n1 24.9236
R15 VGND.n6 VGND.t1 282.817
R16 VGND.n15 VGND.t5 282.817
R17 VGND.n5 VGND.n4 206.54
R18 VGND.n9 VGND.n8 199.739
R19 VGND.n13 VGND.n2 199.739
R20 VGND.n9 VGND.n7 32.0005
R21 VGND.n13 VGND.n1 25.977
R22 VGND.n4 VGND.t7 24.9236
R23 VGND.n4 VGND.t6 24.9236
R24 VGND.n8 VGND.t0 24.9236
R25 VGND.n8 VGND.t3 24.9236
R26 VGND.n2 VGND.t4 24.9236
R27 VGND.n2 VGND.t2 24.9236
R28 VGND.n15 VGND.n14 19.9534
R29 VGND.n14 VGND.n13 18.4476
R30 VGND.n9 VGND.n1 12.424
R31 VGND.n6 VGND.n5 10.9894
R32 VGND.n16 VGND.n15 9.3005
R33 VGND.n7 VGND.n3 9.3005
R34 VGND.n10 VGND.n9 9.3005
R35 VGND.n11 VGND.n1 9.3005
R36 VGND.n13 VGND.n12 9.3005
R37 VGND.n14 VGND.n0 9.3005
R38 VGND.n7 VGND.n6 6.4005
R39 VGND.n5 VGND.n3 0.147189
R40 VGND.n10 VGND.n3 0.120292
R41 VGND.n11 VGND.n10 0.120292
R42 VGND.n12 VGND.n11 0.120292
R43 VGND.n12 VGND.n0 0.120292
R44 VGND.n16 VGND.n0 0.120292
R45 VGND VGND.n16 0.0213333
R46 VNB.t0 VNB.t9 3631.07
R47 VNB.t2 VNB.t13 2677.02
R48 VNB.t3 VNB.t10 1324.27
R49 VNB.t10 VNB.t11 1196.12
R50 VNB.t9 VNB.t3 1196.12
R51 VNB.t8 VNB.t0 1196.12
R52 VNB.t12 VNB.t8 1196.12
R53 VNB.t13 VNB.t12 1196.12
R54 VNB.t1 VNB.t2 1196.12
R55 VNB.t5 VNB.t1 1196.12
R56 VNB.t6 VNB.t5 1196.12
R57 VNB.t4 VNB.t6 1196.12
R58 VNB.t7 VNB.t4 1196.12
R59 VNB VNB.t7 911.327
R60 A2.n1 A2.t0 205.654
R61 A2.n2 A2.t1 205.654
R62 A2.n2 A2.n0 153.377
R63 A2.n4 A2.n3 152
R64 A2.n1 A2.t2 139.78
R65 A2.n2 A2.t3 139.78
R66 A2.n3 A2.n2 45.4462
R67 A2.n4 A2.n0 17.4085
R68 A2.n3 A2.n1 12.3948
R69 A2.n0 A2 5.6325
R70 A2 A2.n4 0.5125
R71 VPWR.n13 VPWR.t0 868.721
R72 VPWR.n9 VPWR.n8 604.741
R73 VPWR.n7 VPWR.n6 599.74
R74 VPWR.n21 VPWR.t5 337.096
R75 VPWR.n19 VPWR.n2 310.502
R76 VPWR.n4 VPWR.n3 310.502
R77 VPWR.n12 VPWR.n11 34.6358
R78 VPWR.n14 VPWR.n4 32.0005
R79 VPWR.n2 VPWR.t3 26.5955
R80 VPWR.n2 VPWR.t4 26.5955
R81 VPWR.n3 VPWR.t1 26.5955
R82 VPWR.n3 VPWR.t2 26.5955
R83 VPWR.n6 VPWR.t7 26.5955
R84 VPWR.n6 VPWR.t6 26.5955
R85 VPWR.n8 VPWR.t8 26.5955
R86 VPWR.n8 VPWR.t9 26.5955
R87 VPWR.n19 VPWR.n18 25.977
R88 VPWR.n21 VPWR.n20 19.9534
R89 VPWR.n20 VPWR.n19 18.4476
R90 VPWR.n18 VPWR.n4 12.424
R91 VPWR.n11 VPWR.n10 9.3005
R92 VPWR.n12 VPWR.n5 9.3005
R93 VPWR.n15 VPWR.n14 9.3005
R94 VPWR.n16 VPWR.n4 9.3005
R95 VPWR.n18 VPWR.n17 9.3005
R96 VPWR.n19 VPWR.n1 9.3005
R97 VPWR.n20 VPWR.n0 9.3005
R98 VPWR.n22 VPWR.n21 9.3005
R99 VPWR.n9 VPWR.n7 8.42954
R100 VPWR.n11 VPWR.n7 7.90638
R101 VPWR.n14 VPWR.n13 6.4005
R102 VPWR.n13 VPWR.n12 3.38874
R103 VPWR.n10 VPWR.n9 1.1494
R104 VPWR.n10 VPWR.n5 0.120292
R105 VPWR.n15 VPWR.n5 0.120292
R106 VPWR.n16 VPWR.n15 0.120292
R107 VPWR.n17 VPWR.n16 0.120292
R108 VPWR.n17 VPWR.n1 0.120292
R109 VPWR.n1 VPWR.n0 0.120292
R110 VPWR.n22 VPWR.n0 0.120292
R111 VPWR VPWR.n22 0.0213333
R112 a_445_297.n6 a_445_297.t5 839.861
R113 a_445_297.n7 a_445_297.n6 671.966
R114 a_445_297.n5 a_445_297.n0 601.188
R115 a_445_297.n2 a_445_297.n1 585
R116 a_445_297.n4 a_445_297.n3 585
R117 a_445_297.n2 a_445_297.t0 381.223
R118 a_445_297.n3 a_445_297.t7 203.895
R119 a_445_297.n5 a_445_297.n4 143.812
R120 a_445_297.n4 a_445_297.n2 63.2476
R121 a_445_297.n6 a_445_297.n5 63.2476
R122 a_445_297.n3 a_445_297.t4 26.5955
R123 a_445_297.n1 a_445_297.t9 26.5955
R124 a_445_297.n1 a_445_297.t3 26.5955
R125 a_445_297.n0 a_445_297.t8 26.5955
R126 a_445_297.n0 a_445_297.t6 26.5955
R127 a_445_297.n7 a_445_297.t1 26.5955
R128 a_445_297.t2 a_445_297.n7 26.5955
R129 VPB.t11 VPB.t4 781.308
R130 VPB.t1 VPB.t9 556.386
R131 VPB.t13 VPB.t0 248.599
R132 VPB.t3 VPB.t13 248.599
R133 VPB.t4 VPB.t3 248.599
R134 VPB.t12 VPB.t11 248.599
R135 VPB.t10 VPB.t12 248.599
R136 VPB.t9 VPB.t10 248.599
R137 VPB.t2 VPB.t1 248.599
R138 VPB.t5 VPB.t2 248.599
R139 VPB.t6 VPB.t5 248.599
R140 VPB.t7 VPB.t6 248.599
R141 VPB.t8 VPB.t7 248.599
R142 VPB VPB.t8 189.409
R143 a_635_47.n0 a_635_47.t1 331.325
R144 a_635_47.n0 a_635_47.t0 331.325
R145 a_635_47.n1 a_635_47.n0 185
R146 a_635_47.n1 a_635_47.t3 24.9236
R147 a_635_47.t2 a_635_47.n1 24.9236
R148 a_79_21.n15 a_79_21.n14 648.247
R149 a_79_21.n14 a_79_21.n13 585
R150 a_79_21.n12 a_79_21.n11 293.83
R151 a_79_21.n2 a_79_21.n0 252.012
R152 a_79_21.n2 a_79_21.n1 245.613
R153 a_79_21.n4 a_79_21.t8 212.081
R154 a_79_21.n9 a_79_21.t9 212.081
R155 a_79_21.n7 a_79_21.t10 212.081
R156 a_79_21.n5 a_79_21.t14 212.081
R157 a_79_21.n6 a_79_21.n3 166.352
R158 a_79_21.n8 a_79_21.n3 152
R159 a_79_21.n11 a_79_21.n10 152
R160 a_79_21.n4 a_79_21.t12 139.78
R161 a_79_21.n9 a_79_21.t13 139.78
R162 a_79_21.n7 a_79_21.t11 139.78
R163 a_79_21.n5 a_79_21.t15 139.78
R164 a_79_21.n14 a_79_21.n12 88.1992
R165 a_79_21.n12 a_79_21.n2 51.9534
R166 a_79_21.n10 a_79_21.n4 48.9308
R167 a_79_21.n9 a_79_21.n8 41.6278
R168 a_79_21.n7 a_79_21.n6 34.3247
R169 a_79_21.n6 a_79_21.n5 27.0217
R170 a_79_21.n13 a_79_21.t2 26.5955
R171 a_79_21.n13 a_79_21.t4 26.5955
R172 a_79_21.t1 a_79_21.n15 26.5955
R173 a_79_21.n15 a_79_21.t7 26.5955
R174 a_79_21.n1 a_79_21.t0 24.9236
R175 a_79_21.n1 a_79_21.t5 24.9236
R176 a_79_21.n0 a_79_21.t3 24.9236
R177 a_79_21.n0 a_79_21.t6 24.9236
R178 a_79_21.n8 a_79_21.n7 19.7187
R179 a_79_21.n11 a_79_21.n3 14.352
R180 a_79_21.n10 a_79_21.n9 12.4157
R181 X.n2 X.n1 384.223
R182 X.n2 X.n0 320.976
R183 X.n5 X.n4 264.435
R184 X.n5 X.n3 201.189
R185 X X.n2 33.455
R186 X X.n5 28.2187
R187 X.n1 X.t3 26.5955
R188 X.n1 X.t2 26.5955
R189 X.n0 X.t1 26.5955
R190 X.n0 X.t0 26.5955
R191 X.n3 X.t7 24.9236
R192 X.n3 X.t4 24.9236
R193 X.n4 X.t6 24.9236
R194 X.n4 X.t5 24.9236
R195 B2.n1 B2.t0 260.281
R196 B2.n2 B2.t1 212.081
R197 B2.n0 B2.t3 192.8
R198 B2.n0 B2 174.564
R199 B2.n4 B2.n3 152
R200 B2.n2 B2.t2 149.421
R201 B2.n3 B2.n2 44.1838
R202 B2.n4 B2 17.1641
R203 B2.n3 B2.n1 11.2472
R204 B2.n5 B2 9.84665
R205 B2 B2.n5 4.94595
R206 B2.n1 B2.n0 4.8205
R207 B2.n5 B2.n4 4.65505
R208 B1.n1 B1.t1 219.31
R209 B1.n3 B1.t3 212.081
R210 B1.n4 B1.t0 155.742
R211 B1.n2 B1.n0 152
R212 B1.n5 B1.n4 152
R213 B1.n1 B1.t2 149.421
R214 B1.n3 B1.n2 53.0205
R215 B1.n5 B1 9.77505
R216 B1.n2 B1.n1 7.2305
R217 B1 B1.n0 6.98232
R218 B1.n0 B1 3.72414
R219 B1.n4 B1.n3 1.60717
R220 B1 B1.n5 0.931409
R221 a_1142_47.n1 a_1142_47.t2 343.358
R222 a_1142_47.t1 a_1142_47.n1 334.712
R223 a_1142_47.n1 a_1142_47.n0 185
R224 a_1142_47.n0 a_1142_47.t0 33.2313
R225 a_1142_47.n0 a_1142_47.t3 24.9236
R226 A1.n1 A1.t2 257.067
R227 A1.n2 A1.t3 205.654
R228 A1.n0 A1.t1 192.8
R229 A1 A1.n0 169.971
R230 A1.n4 A1.n3 152
R231 A1.n2 A1.t0 149.421
R232 A1.n3 A1.n2 33.138
R233 A1.n3 A1.n1 18.8286
R234 A1.n4 A1 13.3125
R235 A1 A1.n4 10.2405
R236 A1.n1 A1.n0 8.03383
C0 VPB B1 0.068644f
C1 X VGND 0.220326f
C2 A2 A1 0.067525f
C3 VPB B2 0.072875f
C4 VPB VPWR 0.152894f
C5 VPB X 0.011488f
C6 A1 B1 0.014686f
C7 A3 VPWR 0.032628f
C8 A3 X 0.003006f
C9 A2 VPWR 0.0259f
C10 VPB VGND 0.011649f
C11 A3 VGND 0.034595f
C12 A2 X 3.16e-19
C13 A1 VPWR 0.025908f
C14 B1 B2 0.091927f
C15 A2 VGND 0.017666f
C16 B1 VPWR 0.02213f
C17 A1 X 1.74e-19
C18 B2 VPWR 0.019443f
C19 A1 VGND 0.017612f
C20 VPB A3 0.069231f
C21 B1 VGND 0.024353f
C22 VPB A2 0.061857f
C23 VPWR X 0.313446f
C24 B2 VGND 0.03545f
C25 VPB A1 0.069753f
C26 A3 A2 0.038299f
C27 VPWR VGND 0.15219f
C28 VGND VNB 0.874478f
C29 X VNB 0.07253f
C30 VPWR VNB 0.730185f
C31 B2 VNB 0.2437f
C32 B1 VNB 0.198464f
C33 A1 VNB 0.204622f
C34 A2 VNB 0.188224f
C35 A3 VNB 0.202988f
C36 VPB VNB 1.57932f
.ends

