


.subckt sky130_fd_sc_hs__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_93_264# a_257_126# a_530_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_530_392# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND A1_N a_257_126# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 VPWR A1_N a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_93_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_257_126# a_93_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_257_126# A2_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 a_258_392# A2_N a_257_126# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR B1 a_530_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_605_126# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 X a_93_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_93_264# B2 a_605_126# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_221_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_293_333# A2_N a_546_378# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_149_74# B2 a_221_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR B2 a_61_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND A2_N a_293_333# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 a_61_392# a_293_333# a_221_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 X a_221_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_293_333# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 X a_221_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND B1 a_149_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_221_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_61_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_546_378# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_221_74# a_293_333# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_586_94# A2_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND a_162_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_162_48# a_586_94# a_820_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_162_48# B2 a_1009_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_820_392# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_1009_74# B2 a_162_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_820_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_162_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND a_586_94# a_162_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_1009_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 X a_162_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_820_392# a_586_94# a_162_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VGND B1 a_1009_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VPWR A1_N a_583_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR B2 a_820_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VPWR a_162_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND A1_N a_586_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 X a_162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR B1 a_820_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 VPWR a_162_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_583_368# A2_N a_586_94# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND a_162_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A1_N a_117_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR B1 a_399_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_399_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B2 a_488_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_117_392# A2_N a_126_112# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND A1_N a_126_112# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 VGND a_126_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_126_112# A2_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 Y a_126_112# a_399_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_488_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_615_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_212_102# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y a_212_102# a_424_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B2 a_615_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR B2 a_424_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR B1 a_424_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A1_N a_209_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND B1 a_615_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y a_212_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_615_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_209_392# A2_N a_212_102# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_212_102# A2_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_424_368# a_212_102# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_424_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_424_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND A1_N a_212_102# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_914_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_539_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B2 a_914_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND B1 a_914_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_114_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_539_368# a_114_392# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR B1 a_539_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y B2 a_914_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND B1 a_914_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y a_114_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_539_368# a_114_392# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_914_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_114_392# A2_N a_29_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_539_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR A1_N a_29_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 Y a_114_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VPWR B2 a_539_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_914_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_914_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR B2 a_539_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR B1 a_539_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VGND a_114_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_539_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VGND A2_N a_114_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_29_392# A2_N a_114_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 Y a_114_392# a_539_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 Y a_114_392# a_539_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_29_392# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X28 a_114_392# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_539_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR a_194_136# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_34_392# a_272_110# a_194_136# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND a_194_136# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_194_136# a_272_110# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_122_136# A1 a_194_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_34_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_272_110# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 VPWR A1 a_34_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND A2 a_122_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_272_110# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR A2 a_504_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_187_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_187_244# A1 a_587_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_32_368# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 X a_187_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND a_32_368# a_187_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_504_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_187_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_187_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_32_368# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_587_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_187_244# a_32_368# a_504_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_864_123# A1 a_187_338# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND a_187_338# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR a_187_338# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 X a_187_338# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_187_338# a_29_392# a_596_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR a_187_338# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A1 a_596_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_596_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_596_392# a_29_392# a_187_338# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 X a_187_338# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_596_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_29_392# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 X a_187_338# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_187_338# a_29_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_187_338# A1 a_864_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VGND a_29_392# a_187_338# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 VPWR A2 a_596_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 VGND a_187_338# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 X a_187_338# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND A2 a_864_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_29_392# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_864_123# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VPWR A2 a_348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_29_424# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_348_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y A1 a_437_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_29_424# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y a_29_424# a_348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_29_424# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 a_437_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VPWR B1_N a_62_94# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_241_368# a_62_94# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_241_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_241_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_62_94# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_436_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_62_94# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VPWR A2 a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y A1 a_436_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y a_62_94# a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR A1 a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A2 a_436_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y a_62_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_436_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_31_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_31_368# a_803_323# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_46_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y a_803_323# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y a_803_323# a_31_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_46_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_31_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_31_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_31_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_46_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_803_323# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_31_368# a_803_323# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND A2 a_46_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR B1_N a_803_323# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 Y a_803_323# a_31_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Y a_803_323# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VPWR A1 a_31_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Y A1 a_46_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR A1 a_31_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR A2 a_31_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Y A1 a_46_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR A2 a_31_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND a_803_323# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND B1_N a_803_323# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_46_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VGND A2 a_46_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_803_323# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_264# B1 a_364_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_81_264# A1 a_452_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 X a_81_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A2 a_364_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_364_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_81_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_452_136# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VGND B1 a_81_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VGND a_84_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_484_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_84_244# B1 a_401_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VPWR A2 a_401_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_84_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND B1 a_84_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_84_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_401_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 X a_84_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_84_244# A1 a_484_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR a_91_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_503_392# B1 a_91_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_91_48# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_503_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND A2 a_700_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR a_91_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_503_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_91_48# A1 a_700_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR A2 a_503_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 X a_91_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_91_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_700_74# A1 a_91_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 X a_91_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_700_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VGND a_91_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_91_48# B1 a_503_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 X a_91_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR A1 a_503_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 X a_91_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND B1 a_91_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_29_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A2 a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_29_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_117_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A1 a_280_107# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_280_107# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A2 a_131_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A1 a_131_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_131_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_131_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_280_107# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_131_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y B1 a_131_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A2 a_280_107# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_69_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_84_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR A2 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A2 a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_84_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_69_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_69_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND A2 a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y A1 a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_69_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_84_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y A1 a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y B1 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_84_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_69_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_69_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR A2 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR A1 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VPWR A1 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_132_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_132_392# B2 a_222_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_52_123# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VPWR a_222_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_222_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_222_392# B1 a_132_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_132_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND B2 a_230_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_222_392# A1 a_52_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_230_79# B1 a_222_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_491_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR a_81_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_81_48# B2 a_388_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_388_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_81_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A1 a_388_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND a_81_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_81_48# B1 a_491_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_304_74# A1 a_81_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 X a_81_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A2 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_388_368# B1 a_81_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_95_306# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A2 a_1064_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_1064_123# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_555_392# B2 a_95_306# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_95_306# B2 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_95_306# B1 a_645_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 VPWR a_95_306# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_1064_123# A1 a_95_306# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_95_306# A1 a_1064_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 VPWR A1 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_555_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND a_95_306# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_95_306# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND B2 a_645_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_95_306# B1 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VGND a_95_306# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_555_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 X a_95_306# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_645_120# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_555_392# B1 a_95_306# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 a_645_120# B1 a_95_306# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 X a_95_306# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 X a_95_306# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR A2 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A2 a_71_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_71_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y A1 a_339_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_339_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_159_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_71_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y B1 a_71_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND B2 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_66_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y B1 a_558_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_558_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_148_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_66_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_66_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_558_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND B2 a_558_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y B2 a_66_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR A1 a_66_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y B1 a_66_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR A2 a_66_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_148_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Y A1 a_148_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VGND A2 a_148_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_66_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B1 a_48_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_840_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_45_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B2 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_45_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y A1 a_840_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND A2 a_840_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y B1 a_48_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_840_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y B2 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_45_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y B1 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y A1 a_840_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND A2 a_840_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR A2 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Y B1 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_840_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND B2 a_48_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR A1 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_45_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VGND B2 a_48_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR A1 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_48_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_45_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR A2 a_45_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_45_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_48_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_45_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_48_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_45_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_840_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_48_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VGND A3 a_265_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_265_120# A2 a_337_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_81_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 X a_81_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_250_392# B1 a_81_270# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_81_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_250_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_337_120# A1 a_81_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR A1 a_250_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR A3 a_250_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_97_296# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_97_296# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_371_74# A2 a_449_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 X a_97_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A3 a_362_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR A1 a_362_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_362_368# B1 a_97_296# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_97_296# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND A3 a_371_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_362_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_449_74# A1 a_97_296# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 X a_97_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_83_274# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND a_83_274# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A1 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_83_274# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A3 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_83_274# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_529_392# B1 a_83_274# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_83_274# A1 a_775_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_83_274# B1 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_529_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_529_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND a_83_274# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_83_274# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_1000_74# A2 a_775_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 X a_83_274# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 X a_83_274# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR A2 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_1000_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 X a_83_274# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_775_74# A2 a_1000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_529_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VGND B1 a_83_274# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_775_74# A1 a_83_274# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 VGND A3 a_1000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_136_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_136_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A3 a_145_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_223_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A3 a_136_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_145_74# A2 a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_136_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_200_74# A2 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y A1 a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_114_74# A2 a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_114_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_200_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND A3 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_475_74# A2 a_30_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y A1 a_475_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND A3 a_30_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_30_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_30_74# A2 a_475_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_475_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_475_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_30_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_30_74# A2 a_475_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_475_74# A2 a_30_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VGND A3 a_30_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 Y A1 a_475_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_84_48# B2 a_244_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_601_94# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VPWR A3 a_244_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_244_368# B1 a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_84_48# B1 a_601_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 X a_84_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A1 a_244_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_244_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_259_94# A2 a_337_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 X a_84_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND A3 a_259_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_337_94# A1 a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_45_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A3 a_346_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR A1 a_346_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_661_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_433_74# A1 a_45_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_45_264# B2 a_346_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_346_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_45_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_346_368# B1 a_45_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VGND a_45_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 X a_45_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_45_264# B1 a_661_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_355_74# A2 a_433_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND A3 a_355_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_83_283# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND a_83_283# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_83_283# B1 a_587_110# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND A3 a_992_122# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VPWR A1 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND a_83_283# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_587_110# B1 a_83_283# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_1079_122# A2 a_992_122# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_509_392# B1 a_83_283# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_509_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 X a_83_283# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_992_122# A2 a_1079_122# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_587_110# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 X a_83_283# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_83_283# B2 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VPWR A3 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_509_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_1079_122# A1 a_83_283# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 a_992_122# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 X a_83_283# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR A2 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 a_509_392# B2 a_83_283# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_83_283# A1 a_1079_122# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 VGND B2 a_587_110# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 VPWR a_83_283# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_509_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X26 X a_83_283# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_83_283# B1 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_391_74# A2 a_469_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_119_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND B2 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y A1 a_391_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_469_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 Y A1 a_507_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND A3 a_771_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_771_74# A2 a_507_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_507_74# A2 a_771_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_771_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_507_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_1313_74# A2 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_868_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 Y A1 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_1313_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Y A1 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_1313_74# A2 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_1313_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_868_74# A2 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_868_74# A2 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 VGND A3 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 a_868_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X39 VGND A3 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 X a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_83_244# A1 a_449_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND B1 a_83_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_83_244# B1 a_354_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_354_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_354_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VPWR A4 a_354_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_657_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_449_74# A2 a_543_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A2 a_354_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_543_74# A3 a_657_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_121_74# A3 a_199_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_313_74# A1 a_441_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_27_392# B1 a_441_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VPWR a_441_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_441_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A3 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_27_392# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND A4 a_121_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_199_74# A2 a_313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 X a_441_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 X a_441_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_27_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_441_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VGND a_113_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A2 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_1205_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_113_98# A1 a_751_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 X a_113_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_751_74# A1 a_113_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR A1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_27_392# B1 a_113_98# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR a_113_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR a_113_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_392# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND a_113_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR A3 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_751_74# A2 a_1010_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_113_98# B1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_113_98# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 X a_113_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_27_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VGND B1 a_113_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_27_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 a_1010_74# A2 a_751_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_1010_74# A3 a_1205_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 X a_113_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR A4 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_1205_74# A3 a_1010_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 X a_113_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND A4 a_1205_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A3 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_355_74# A2 a_469_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_116_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_116_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_469_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_277_74# A3 a_355_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND A4 a_277_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_709_74# A3 a_512_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_709_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_512_74# A2 a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_512_74# A3 a_709_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_239_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_239_74# A2 a_512_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 Y A1 a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND A4 a_709_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_1235_74# A3 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_325_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_325_74# A2 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_852_74# A2 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_325_74# A2 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_1235_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Y A1 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_852_74# A3 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y A1 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_1235_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_27_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VGND A4 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_27_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_325_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_852_74# A3 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 a_852_74# A2 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 VGND A4 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X36 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 a_1235_74# A3 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 X a_81_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A1 a_279_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_279_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND C1 a_81_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 X a_81_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_279_392# B1 a_550_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_550_392# C1 a_81_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_81_264# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VGND A2 a_366_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_366_136# A1 a_81_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_600_392# C1 a_85_270# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_85_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND C1 a_85_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_317_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_85_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_399_74# A1 a_85_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR A1 a_317_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND A2 a_399_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_85_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 X a_85_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_85_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_317_392# B1 a_600_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_105_280# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND A2 a_1064_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_1064_123# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_105_280# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_105_280# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 X a_105_280# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_517_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_105_280# C1 a_602_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_1064_123# A1 a_105_280# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_105_280# A1 a_1064_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR A1 a_517_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 X a_105_280# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_517_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_105_280# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VPWR a_105_280# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_517_392# B1 a_602_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 X a_105_280# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND B1 a_105_280# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 X a_105_280# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_602_392# C1 a_105_280# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 VGND C1 a_105_280# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_602_392# B1 a_517_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 VPWR A2 a_517_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VGND a_105_280# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_354_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_71_368# B1 a_354_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_71_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A1 a_71_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_159_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A2 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_114_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_114_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_497_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_497_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y A1 a_38_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_38_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A2 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_38_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_114_368# B1 a_497_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y C1 a_497_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND A2 a_38_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_77_368# B1 a_901_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_77_368# B1 a_901_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A2 a_77_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y C1 a_901_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_901_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A2 a_77_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_77_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_77_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_92_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_92_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_901_368# B1 a_77_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_92_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_77_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_901_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VGND A2 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Y A1 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_77_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 Y C1 a_901_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 Y A1 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND A2 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 VPWR A1 a_77_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_92_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VPWR A1 a_77_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_901_368# B1 a_77_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_509_392# C1 a_148_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VGND A2 a_417_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_310_392# B2 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_417_79# A1 a_148_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 X a_148_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_148_260# B1 a_597_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_310_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_509_392# B1 a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND C1 a_148_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 X a_148_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_597_79# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VPWR A2 a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_515_392# C1 a_89_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 X a_89_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR a_89_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_603_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_316_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND C1 a_89_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_316_392# B2 a_515_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND A2 a_337_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_337_74# A1 a_89_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_89_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A2 a_316_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 X a_89_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_515_392# B1 a_316_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_89_260# B1 a_603_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 X a_154_135# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_154_135# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_1102_392# C1 a_154_135# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_154_135# A1 a_71_135# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_1346_123# B1 a_154_135# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_1102_392# B2 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND A2 a_71_135# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_157_376# B1 a_1102_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 X a_154_135# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND B2 a_1346_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_157_376# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 X a_154_135# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_154_135# B1 a_1346_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VGND C1 a_154_135# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_71_135# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_157_376# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_1346_123# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_154_135# C1 a_1102_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_1102_392# B1 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 a_154_135# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_157_376# B2 a_1102_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VPWR a_154_135# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR A2 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VPWR a_154_135# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 X a_154_135# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR A1 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X26 a_71_135# A1 a_154_135# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 VGND a_154_135# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_263_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_118_368# B1 a_263_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y A1 a_567_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR A2 a_263_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND B2 a_351_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_351_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_567_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y C1 a_118_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_263_368# B2 a_118_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y C1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_29_368# B2 a_294_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_293_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_294_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_675_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y A1 a_675_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_29_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_294_368# B2 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_29_368# B1 a_294_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y B1 a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_294_368# B1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR A1 a_294_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR A2 a_294_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_294_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_293_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND B2 a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_675_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND A2 a_675_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_114_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_114_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_534_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B1 a_1326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_531_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_531_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_531_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_1326_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_531_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y A1 a_534_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_1326_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND B2 a_1326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_531_368# B2 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_531_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_1326_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y C1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR A1 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Y A1 a_534_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_114_368# B2 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND B2 a_1326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_534_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Y C1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VPWR A1 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_534_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_534_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_114_368# B1 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VPWR A2 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_114_368# B1 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 VGND A2 a_534_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_1326_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 VPWR A2 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_114_368# B2 a_531_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 VGND A2 a_534_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_531_368# B2 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 a_531_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 Y B1 a_1326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
X0 a_651_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_119_74# C2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_32_74# C2 a_27_390# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_32_74# C1 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_27_390# C1 a_32_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_337_390# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_337_390# B1 a_27_390# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VPWR a_32_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_390# B2 a_337_390# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_32_74# A1 a_651_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VGND a_32_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_386_74# B1 a_32_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 VPWR A1 a_337_390# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VGND B2 a_386_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a222o_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
X0 a_639_368# B1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_27_82# C1 a_114_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_775_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_27_82# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_82# B1 a_775_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 X a_27_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 X a_27_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A2 a_557_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_27_82# C1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR A1 a_639_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_639_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_116_392# B2 a_639_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VPWR a_27_82# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_557_74# A1 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_116_392# C2 a_27_82# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_114_82# C2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
X0 a_116_392# B1 a_369_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_697_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 Y A1 a_697_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND B2 a_461_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_369_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_119_74# C2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 Y C1 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 Y C1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_116_392# C2 Y VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR A2 a_369_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_461_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_369_392# B2 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a222oi_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
X0 VPWR A2 a_515_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VGND C2 a_137_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VGND A2 a_981_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_515_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VPWR A1 a_515_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_137_74# C2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_515_392# B1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 Y A1 a_981_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_981_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_515_392# B2 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 Y C2 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_981_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_116_392# C2 Y VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_116_392# B1 a_515_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_515_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_116_392# B2 a_515_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VGND B2 a_593_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_593_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 Y C1 a_137_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 Y B1 a_593_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 Y C1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 a_137_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_593_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_116_392# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VGND A3 a_264_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_89_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_359_123# A1 a_89_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VPWR A1 a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_264_120# A2 a_359_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 X a_89_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A3 a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_89_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_546_392# C1 a_89_270# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VGND C1 a_89_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_258_392# B1 a_546_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_258_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VGND A3 a_351_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_330_392# B1 a_660_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR A1 a_330_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_351_74# A2 a_423_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_660_392# C1 a_21_270# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_21_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND C1 a_21_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_330_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 X a_21_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR A3 a_330_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VGND a_21_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_423_74# A1 a_21_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_21_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 X a_21_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_334_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_154_392# A1 a_1081_39# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_69_392# B1 a_334_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_334_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_154_392# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_334_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND a_154_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_334_392# B1 a_69_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_888_105# A2 a_1081_39# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_1081_39# A2 a_888_105# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VGND C1 a_154_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_888_105# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 X a_154_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND B1 a_154_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 X a_154_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_154_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 X a_154_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 X a_154_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_154_392# C1 a_69_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VPWR A2 a_334_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 VPWR A1 a_334_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 a_1081_39# A1 a_154_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_154_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR a_154_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR A3 a_334_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_154_392# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 VGND A3 a_888_105# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 a_69_392# C1 a_154_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A3 a_156_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_231_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_156_368# B1 a_462_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_159_74# A2 a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_462_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A1 a_156_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_156_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND A3 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_45_74# A2 a_300_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y A1 a_300_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_127_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A1 a_127_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_127_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_127_368# B1 a_692_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_45_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A3 a_127_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR A2 a_127_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_127_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_692_368# B1 a_127_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_692_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND A3 a_45_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y C1 a_692_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_300_74# A2 a_45_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_300_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_114_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_114_368# B1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_114_368# B1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_114_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y C1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_114_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_114_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y A1 a_465_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND A3 a_34_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR A3 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR A1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_34_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_114_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_1213_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND A3 a_34_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 Y A1 a_465_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_1213_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR A3 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_34_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_1213_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR A2 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VPWR A2 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_1213_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_34_74# A2 a_465_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 Y C1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_465_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VPWR A1 a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_465_74# A2 a_34_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 a_114_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_34_74# A2 a_465_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_465_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_465_74# A2 a_34_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR A2 a_80_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_431_392# D1 a_85_136# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR a_85_136# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_80_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND B1 a_85_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_80_392# B1 a_353_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_85_136# A1 a_168_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VGND D1 a_85_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_85_136# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_353_392# C1 a_431_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_168_136# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VGND a_85_136# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR a_91_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A1 a_630_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_522_368# B1 a_630_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_444_368# C1 a_522_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_91_244# D1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_91_244# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_91_244# D1 a_444_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND A2 a_771_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND a_91_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 X a_91_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_630_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 X a_91_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND C1 a_91_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_771_74# A1 a_91_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 X a_137_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A2 a_1013_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_137_260# D1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND A2 a_1210_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_137_260# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 X a_137_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_549_392# C1 a_814_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_137_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_1013_392# B1 a_814_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_1013_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_1013_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 X a_137_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND a_137_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_137_260# A1 a_1210_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VGND C1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_549_392# D1 a_137_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_1210_74# A1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 VPWR a_137_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_137_260# D1 a_549_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VGND a_137_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND D1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VPWR a_137_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_814_392# C1 a_549_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_1210_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 VGND B1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 a_814_392# B1 a_1013_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X26 a_137_260# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 VPWR A1 a_1013_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_342_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y A1 a_461_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y D1 a_156_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_461_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_156_368# C1 a_234_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A2 a_342_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_234_368# B1 a_342_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR A2 a_533_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y D1 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_722_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_334_368# B1 a_533_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR A1 a_533_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_722_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y A1 a_722_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_69_368# D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_69_368# C1 a_334_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A2 a_722_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_334_368# C1 a_69_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_533_368# B1 a_334_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_533_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_533_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y D1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_853_368# B1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A2 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A2 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y D1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_474_368# B1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_474_368# C1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_853_368# B1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_474_368# C1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_853_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_1228_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_853_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_29_368# D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_853_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_853_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_1228_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_29_368# D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Y D1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_29_368# C1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_1228_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_29_368# C1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_474_368# B1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 Y A1 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR A1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_1228_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VPWR A1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 VGND A2 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 Y A1 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 VPWR A2 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR A a_56_136# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_56_136# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_143_136# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_56_136# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_56_136# A a_143_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR a_56_136# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X
X0 a_31_74# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_118_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_31_74# A a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A a_31_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X
X0 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and2b_1 A_N B VGND VNB VPB VPWR X
X0 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_266_98# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VGND a_266_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_353_98# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_266_98# a_27_74# a_353_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR a_27_74# a_266_98# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR a_266_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__and2b_2 A_N B VGND VNB VPB VPWR X
X0 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND a_198_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR B a_198_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_198_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 X a_198_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_505_74# a_27_74# a_198_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_198_48# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND B a_505_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_198_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__and2b_4 A_N B VGND VNB VPB VPWR X
X0 X a_218_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_233_74# a_27_392# a_218_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 X a_218_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 X a_218_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_218_424# a_27_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VPWR B a_218_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND B a_233_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_233_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR a_218_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_392# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 X a_218_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR a_218_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND a_218_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_218_424# a_27_392# a_233_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_27_392# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VPWR a_27_392# a_218_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_218_424# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 VGND a_218_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and3_1 A B C VGND VNB VPB VPWR X
X0 a_27_398# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR B a_27_398# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_121_136# B a_233_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_27_398# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_27_398# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_398# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_27_398# A a_121_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_233_136# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__and3_2 A B C VGND VNB VPB VPWR X
X0 a_41_384# A a_133_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND a_41_384# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_133_136# B a_247_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_41_384# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_247_136# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 X a_41_384# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 X a_41_384# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_41_384# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VPWR B a_41_384# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VPWR a_41_384# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__and3_4 A B C VGND VNB VPB VPWR X
X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR B a_83_260# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_83_260# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VGND C a_489_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_686_74# B a_489_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_83_260# A a_686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_489_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_489_74# B a_686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_83_260# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR C a_83_260# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_686_74# A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_431_94# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_266_94# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR a_266_94# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_353_94# B a_431_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_266_94# a_114_74# a_353_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR A_N a_114_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND a_266_94# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_266_94# a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VPWR B a_266_94# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VGND A_N a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__and3b_2 A_N B C VGND VNB VPB VPWR X
X0 a_454_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_284_368# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 X a_284_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR a_284_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_284_368# a_27_88# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_284_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR B a_284_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_284_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_376_74# B a_454_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_27_88# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_27_88# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X11 a_284_368# a_27_88# a_376_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and3b_4 A_N B C VGND VNB VPB VPWR X
X0 a_298_368# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_239_98# B a_498_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 X a_298_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 X a_298_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_298_368# a_27_74# a_239_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR B a_298_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_298_368# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND C a_498_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR C a_298_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR a_298_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR a_298_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_498_98# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 VGND a_298_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_298_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VPWR a_27_74# a_298_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VGND a_298_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_498_98# B a_239_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_239_98# a_27_74# a_298_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 X a_298_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 X a_298_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_96_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_335_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VPWR a_96_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A a_96_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_96_74# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VPWR C a_96_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_257_74# C a_335_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_179_74# B a_257_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_96_74# A a_179_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 VGND a_96_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4_2 A B C D VGND VNB VPB VPWR X
X0 VPWR C a_56_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_335_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 X a_56_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_143_74# B a_221_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_56_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_56_74# A a_143_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_56_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A a_56_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 X a_56_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_56_74# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VGND a_56_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_221_74# C a_335_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4_4 A B C D VGND VNB VPB VPWR X
X0 X a_116_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_116_392# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_463_119# C a_32_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 X a_116_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_463_119# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_32_119# C a_463_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 VGND a_116_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_116_392# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR a_116_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR B a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 X a_116_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 X a_116_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_116_392# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VPWR A a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_32_119# B a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VPWR a_116_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_116_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_119_119# A a_116_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 VPWR C a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VGND D a_463_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 VPWR D a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 a_119_119# B a_32_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_116_392# A a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_116_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_526_139# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_353_124# B a_448_139# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VPWR C a_226_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VGND a_226_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_448_139# C a_526_139# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_226_424# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR a_226_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_226_424# a_27_74# a_353_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR a_27_74# a_226_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_226_424# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4b_2 A_N B C D VGND VNB VPB VPWR X
X0 a_27_112# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR D a_186_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_459_74# C a_537_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_186_48# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VPWR a_186_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND D a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_537_74# B a_645_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_645_74# a_27_112# a_186_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND a_186_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_186_48# a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_27_112# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X11 X a_186_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 X a_186_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR B a_186_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4b_4 A_N B C D VGND VNB VPB VPWR X
X0 a_27_368# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_27_368# a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR C a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_751_125# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_199_294# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND a_199_294# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_199_294# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_199_294# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_664_125# C a_751_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_1136_125# a_27_368# a_199_294# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_199_294# a_27_368# a_1136_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VPWR B a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_1136_125# B a_664_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VPWR D a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_199_294# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_199_294# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_27_368# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 X a_199_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_199_294# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 a_664_125# B a_1136_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_751_125# C a_664_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VGND D a_751_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_199_294# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 X a_199_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 X a_199_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 X a_199_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND a_179_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_179_48# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VPWR B_N a_503_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_647_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VGND B_N a_503_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 VPWR a_27_74# a_179_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 VPWR a_179_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR C a_179_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_455_74# a_503_48# a_533_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_179_48# a_503_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_179_48# a_27_74# a_455_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_533_74# C a_647_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR a_225_82# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR C a_225_82# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_225_82# a_354_252# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_498_82# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND B_N a_354_252# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR B_N a_354_252# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 X a_225_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_390_82# C a_498_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_27_74# a_225_82# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_225_82# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND a_225_82# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_312_82# a_354_252# a_390_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_225_82# a_27_74# a_312_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 X a_225_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
X0 a_472_388# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VGND a_472_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_685_140# a_27_74# a_412_140# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_685_140# C a_882_137# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VGND A_N a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_472_388# a_200_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND a_472_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A_N a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_27_74# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VGND D a_882_137# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 X a_472_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR D a_472_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VPWR a_200_74# a_472_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_472_388# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 X a_472_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 X a_472_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_882_137# C a_685_140# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_882_137# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 VPWR a_27_74# a_472_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 a_472_388# a_200_74# a_412_140# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_412_140# a_200_74# a_472_388# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VPWR a_472_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR C a_472_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VPWR a_472_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_27_74# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 a_412_140# a_27_74# a_685_140# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 X a_472_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_472_388# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__buf_1 A VGND VNB VPB VPWR X
X0 VGND a_27_164# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_164# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 a_27_164# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VPWR a_27_164# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__buf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_21_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 X a_21_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND A a_21_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_21_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_21_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 X a_21_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__buf_4 A VGND VNB VPB VPWR X
X0 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_86_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A a_86_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR A a_86_260# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__buf_8 A VGND VNB VPB VPWR X
X0 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X
X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X41 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends

.subckt sky130_fd_sc_hs__bufbuf_1 A VGND VNB VPB VPWR X
X0 a_27_112# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_27_112# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15

X2 VGND a_27_112# a_221_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_27_112# a_221_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15

X4 a_334_368# a_221_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_221_368# a_334_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15

X6 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends

.subckt sky130_fd_sc_hs__bufbuf_8 A VGND VNB VPB VPWR X
X0 a_27_112# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_334_368# a_221_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND a_221_368# a_334_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_334_368# a_221_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR a_221_368# a_334_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_112# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X20 VGND a_27_112# a_221_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_334_368# a_221_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VPWR a_27_112# a_221_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_334_368# a_221_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__bufbuf_16 A VGND VNB VPB VPWR X
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_203_74# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VPWR a_27_368# a_203_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 VPWR a_27_368# a_203_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X36 a_203_74# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X41 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X42 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X43 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X44 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X45 VGND a_27_368# a_203_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X46 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X47 VGND a_27_368# a_203_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X48 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X49 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X50 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X51 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends


.subckt sky130_fd_sc_hs__bufinv_1 A VGND VNB VPB VPWR Y
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15

X2 VPWR a_27_368# a_183_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_27_368# a_183_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15

X4 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends

.subckt sky130_fd_sc_hs__bufinv_8 A VGND VNB VPB VPWR Y
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR a_27_368# a_183_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_183_48# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_27_368# a_183_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND a_27_368# a_183_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND a_27_368# a_183_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_183_48# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__bufinv_16 A VGND VNB VPB VPWR Y
X0 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X39 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X41 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X42 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X43 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X44 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X45 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X46 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X47 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X48 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X49 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__clkbuf_1 A VGND VNB VPB VPWR X
X0 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__clkbuf_2 A VGND VNB VPB VPWR X
X0 X a_43_192# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A a_43_192# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 X a_43_192# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 VPWR a_43_192# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A a_43_192# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_43_192# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR a_83_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR a_83_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND A a_83_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 X a_83_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VGND a_83_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 X a_83_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 X a_83_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_83_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 X a_83_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR A a_83_270# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__clkbuf_8 A VGND VNB VPB VPWR X
X0 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_125_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A a_125_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 a_125_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 VPWR A a_125_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__clkbuf_16 A VGND VNB VPB VPWR X
X0 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__clkdlyinv3sd1_1 A VGND VNB VPB VPWR Y
X0 VPWR a_28_74# a_285_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_285_392# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_285_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 VGND a_28_74# a_285_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__clkdlyinv3sd2_1 A VGND VNB VPB VPWR Y
X0 VPWR a_288_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_288_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X5 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.25
.ends



.subckt sky130_fd_sc_hs__clkdlyinv3sd3_1 A VGND VNB VPB VPWR Y
X0 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X1 VPWR a_288_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_288_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
.ends



.subckt sky130_fd_sc_hs__clkdlyinv5sd1_1 A VGND VNB VPB VPWR Y
X0 a_682_74# a_549_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_288_74# a_549_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_682_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR a_682_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_682_74# a_549_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VGND a_288_74# a_549_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__clkdlyinv5sd2_1 A VGND VNB VPB VPWR Y
X0 a_682_74# a_549_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.25
X1 VGND a_682_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_288_74# a_549_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.25
X5 VPWR a_682_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X7 VGND a_288_74# a_549_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X8 a_682_74# a_549_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X9 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.25
.ends



.subckt sky130_fd_sc_hs__clkdlyinv5sd3_1 A VGND VNB VPB VPWR Y
X0 VPWR a_288_74# a_549_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X1 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X2 VGND a_682_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR a_682_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X7 VGND a_288_74# a_549_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X8 a_682_74# a_549_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X9 a_682_74# a_549_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
.ends



.subckt sky130_fd_sc_hs__clkinv_0 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hs__clkinv_1 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hs__clkinv_2 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__clkinv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__clkinv_8 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__clkinv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X30 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X36 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__conb_1 VGND VNB VPB VPWR HI LO
XR0 HI VPWR sky130_fd_pr__res_generic_po w=0.51 l=0.045
XR1 VGND LO sky130_fd_pr__res_generic_po w=0.51 l=0.045
.ends



.subckt sky130_fd_sc_hs__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=1.0
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=1.0
.ends



.subckt sky130_fd_sc_hs__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=1.0
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=1.0
X2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=1.0
X3 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=1.0
.ends



.subckt sky130_fd_sc_hs__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR a_27_74# a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_595_119# a_200_74# a_311_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_1534_446# a_1349_114# a_1818_76# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_311_119# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 a_1349_114# a_27_74# a_1483_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 VGND a_1534_446# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_474_405# a_537_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 VPWR a_1534_446# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_1611_140# a_1534_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_595_119# a_27_74# a_311_119# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 a_1483_508# a_1534_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 VGND a_27_74# a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_1917_392# a_1349_114# a_1534_446# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_537_503# a_200_74# a_595_119# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_978_357# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X15 a_27_74# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR a_2412_410# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR a_474_405# a_1297_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_311_119# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 a_474_405# a_978_357# a_867_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X20 a_867_119# a_595_119# a_474_405# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 VPWR a_978_357# a_1917_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_1254_119# a_27_74# a_1349_114# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X23 VGND SET_B a_1818_76# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_978_357# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_1297_424# a_200_74# a_1349_114# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 a_2412_410# a_1534_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X27 a_867_119# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X28 a_933_424# a_978_357# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X29 VGND a_2412_410# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VGND a_474_405# a_523_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_523_119# a_27_74# a_595_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_1534_446# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X33 a_1349_114# a_200_74# a_1611_140# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 VPWR SET_B a_474_405# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X35 a_1818_76# a_978_357# a_1534_446# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_2412_410# a_1534_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 a_27_74# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 VGND a_474_405# a_1254_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X39 a_474_405# a_595_119# a_933_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR a_27_74# a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1240_125# a_27_74# a_1335_112# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 Q a_2516_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_473_405# a_529_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VPWR a_1555_410# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Q_N a_1555_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_311_119# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 VGND a_2516_368# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_1931_392# a_1335_112# a_1555_410# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VGND SET_B a_1832_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_930_424# a_975_322# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_867_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X12 VPWR a_2516_368# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_1640_138# a_1555_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 VGND a_27_74# a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_1335_112# a_27_74# a_1504_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X16 VPWR a_473_405# a_536_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 a_1555_410# a_1335_112# a_1832_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_601_119# a_27_74# a_311_119# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_601_119# a_200_74# a_311_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_27_74# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_1504_508# a_1555_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_529_119# a_27_74# a_601_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VGND a_473_405# a_1240_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X24 a_1335_112# a_200_74# a_1640_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_311_119# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_975_322# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 a_536_503# a_200_74# a_601_119# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 a_473_405# a_601_119# a_930_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X29 VPWR a_975_322# a_1931_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X30 VPWR SET_B a_473_405# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X31 Q_N a_1555_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 VGND a_1555_410# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 a_2516_368# a_1555_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X34 a_1555_410# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X35 VPWR a_473_405# a_1312_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X36 a_2516_368# a_1555_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X37 Q a_2516_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 a_1832_74# a_975_322# a_1555_410# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 a_975_322# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X40 a_1312_424# a_200_74# a_1335_112# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X41 a_27_74# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X42 a_473_405# a_975_322# a_867_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X43 a_867_125# a_601_119# a_473_405# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_671_93# a_520_87# a_1017_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_1318_119# a_214_74# a_1311_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 a_1474_446# a_1062_93# a_1708_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_671_93# a_1203_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_520_87# a_27_74# a_713_379# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 VGND SET_B a_1708_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_422_125# a_214_74# a_520_87# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 a_1814_392# a_1062_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_1017_379# a_1062_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VPWR SET_B a_1474_446# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_713_379# a_671_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_2320_410# a_1474_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VPWR a_2320_410# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_671_93# a_1062_93# a_872_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 a_872_119# a_520_87# a_671_93# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 a_1062_93# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_1062_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X18 a_1311_424# a_27_74# a_1498_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VPWR a_27_74# a_214_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_606_87# a_671_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VGND a_1474_446# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VPWR D a_422_125# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 a_520_87# a_214_74# a_606_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_1498_74# a_1474_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_1418_508# a_1474_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 a_422_125# a_27_74# a_520_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VGND a_27_74# a_214_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR SET_B a_671_93# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X29 VGND SET_B a_872_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X30 VGND a_671_93# a_1318_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X31 VPWR a_1474_446# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 VGND a_2320_410# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 a_2320_410# a_1474_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X34 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_1203_379# a_27_74# a_1311_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X36 VGND D a_422_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 a_1474_446# a_1311_424# a_1814_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X38 a_1708_74# a_1311_424# a_1474_446# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 a_1311_424# a_214_74# a_1418_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 VGND RESET_B a_1624_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_125_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VPWR a_1224_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_38_78# D a_125_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VGND a_319_360# a_498_360# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_910_118# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 VPWR a_319_360# a_498_360# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_1224_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_706_463# a_841_401# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_841_401# a_319_360# a_1224_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_1434_74# a_1482_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_1224_74# a_498_360# a_1465_471# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 VPWR a_2026_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_706_463# a_319_360# a_796_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VPWR RESET_B a_706_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_1482_48# a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X16 a_38_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 a_1465_471# a_1482_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 VGND a_2026_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_319_360# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_2026_424# a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 a_38_78# a_319_360# a_706_463# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 a_796_463# a_841_401# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 VGND a_706_463# a_841_401# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_319_360# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_1224_74# a_319_360# a_1434_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_2026_424# a_1224_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X27 a_706_463# a_498_360# a_832_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 a_841_401# a_498_360# a_1224_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 a_1624_74# a_1224_74# a_1482_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X30 VPWR D a_38_78# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X31 a_38_78# a_498_360# a_706_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 VPWR RESET_B a_1482_48# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X33 a_832_118# a_841_401# a_910_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X16 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X27 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X32 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X36 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
X0 VGND CLK_N a_300_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR a_300_74# a_507_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR D a_33_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_120_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_714_127# a_300_74# a_850_127# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_1550_119# a_1598_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 VPWR RESET_B a_1598_93# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 a_1598_93# a_1266_119# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_714_127# a_507_368# a_817_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 VPWR RESET_B a_714_127# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 a_1266_119# a_507_368# a_1550_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VGND a_714_127# a_856_304# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_33_74# D a_120_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_1547_508# a_1598_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_33_74# a_507_368# a_714_127# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_817_508# a_856_304# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X16 VGND RESET_B a_1736_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_850_127# a_856_304# a_922_127# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_922_127# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 a_1934_94# a_1266_119# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 VPWR a_1934_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_1736_119# a_1266_119# a_1598_93# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 a_33_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 a_33_74# a_300_74# a_714_127# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_856_304# a_300_74# a_1266_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR CLK_N a_300_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_856_304# a_507_368# a_1266_119# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_1934_94# a_1266_119# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X28 VGND a_1934_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VGND a_300_74# a_507_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VPWR a_714_127# a_856_304# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X31 a_1266_119# a_300_74# a_1547_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1468_493# a_1518_203# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 VGND a_1266_74# a_1864_409# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 VGND a_306_74# a_490_366# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_30_78# a_306_74# a_695_457# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_830_359# a_490_366# a_1266_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND a_695_457# a_830_359# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_1266_74# a_1864_409# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_306_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_695_457# a_306_74# a_785_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 VPWR RESET_B a_695_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 Q a_1864_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR D a_30_78# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_306_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_1266_74# a_490_366# a_1468_493# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_695_457# a_490_366# a_816_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 Q a_1864_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND RESET_B a_1656_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_785_457# a_830_359# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_1518_203# a_1266_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_1656_81# a_1266_74# a_1518_203# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_894_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VPWR a_695_457# a_830_359# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_30_78# a_490_366# a_695_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 VPWR a_306_74# a_490_366# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_117_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_30_78# D a_117_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_830_359# a_306_74# a_1266_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_1476_81# a_1518_203# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 a_816_138# a_830_359# a_894_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_30_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 VPWR RESET_B a_1518_203# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X31 a_1266_74# a_306_74# a_1476_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_817_138# a_837_359# a_895_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_696_457# a_306_74# a_786_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 a_1271_74# a_490_362# a_1478_493# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_30_78# a_306_74# a_696_457# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_1481_81# a_1525_212# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_306_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND a_1271_74# a_1921_409# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR D a_30_78# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_306_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_696_457# a_490_362# a_817_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_1525_212# a_1271_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 VGND a_696_457# a_837_359# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Q a_1921_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_30_78# a_490_362# a_696_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VPWR RESET_B a_696_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 Q a_1921_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_895_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 VGND a_1921_409# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR a_696_457# a_837_359# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VGND a_306_74# a_490_362# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_1271_74# a_306_74# a_1481_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_786_457# a_837_359# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_1478_493# a_1525_212# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 a_837_359# a_306_74# a_1271_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X24 a_117_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 VPWR a_1271_74# a_1921_409# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 a_1663_81# a_1271_74# a_1525_212# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VPWR a_306_74# a_490_362# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_30_78# D a_117_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_837_359# a_490_362# a_1271_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VGND RESET_B a_1663_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 VPWR RESET_B a_1525_212# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 VPWR a_1921_409# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_30_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 VPWR a_313_74# a_494_366# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_890_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_313_74# a_494_366# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_2010_409# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR D a_37_78# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_699_463# a_494_366# a_812_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 VPWR RESET_B a_1678_395# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 Q a_2010_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_124_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 Q a_2010_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_37_78# D a_124_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_1350_392# a_313_74# a_1647_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_699_463# a_313_74# a_789_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 VPWR a_699_463# a_834_355# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_1827_81# a_1350_392# a_1678_395# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_834_355# a_494_366# a_1350_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND RESET_B a_1827_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_313_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_1627_493# a_1678_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_789_463# a_834_355# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X20 Q a_2010_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VPWR a_1350_392# a_2010_409# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 VPWR a_2010_409# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR RESET_B a_699_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_1678_395# a_1350_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 a_37_78# a_494_366# a_699_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 a_812_138# a_834_355# a_890_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VGND a_2010_409# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_37_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X29 a_313_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_834_355# a_313_74# a_1350_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X31 a_1350_392# a_494_366# a_1627_493# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 a_2010_409# a_1350_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X33 VGND a_699_463# a_834_355# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_1647_81# a_1678_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 Q a_2010_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_37_78# a_313_74# a_699_463# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 VGND a_1350_392# a_2010_409# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 VGND a_2010_409# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1517_508# a_1510_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_1462_74# a_1510_48# a_1540_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_1355_377# a_225_74# a_1462_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_779_380# a_596_81# a_1061_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_2113_74# a_1355_377# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VGND a_1355_377# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_80# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1355_377# a_398_74# a_1517_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_748_81# a_779_380# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VPWR a_2113_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_1540_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 VPWR a_596_81# a_779_380# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 a_1510_48# a_1355_377# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VPWR SET_B a_1355_377# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_2113_74# a_1355_377# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 VPWR a_1355_377# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_728_463# a_779_380# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 VGND a_2113_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR a_596_81# a_1254_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 VGND a_596_81# a_1262_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_1262_74# a_398_74# a_1355_377# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_27_80# a_398_74# a_596_81# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_27_80# a_225_74# a_596_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_1254_341# a_225_74# a_1355_377# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X26 a_596_81# a_398_74# a_748_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_1061_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_779_380# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_596_81# a_225_74# a_728_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 VGND a_1355_377# a_1510_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_27_80# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1001_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 VPWR a_1339_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND a_1339_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_1258_341# a_225_74# a_1339_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_1453_118# a_1501_92# a_1531_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_1339_74# a_398_74# a_1521_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 a_595_97# a_398_74# a_731_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1501_92# a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_2221_74# a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_731_97# a_757_401# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VPWR a_2221_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_1521_508# a_1501_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_757_401# a_595_97# a_1001_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_2221_74# a_1339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 Q_N a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_1261_74# a_398_74# a_1339_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_27_74# a_225_74# a_595_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_27_74# a_398_74# a_595_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_1339_74# a_225_74# a_1453_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_706_463# a_757_401# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VGND a_1339_74# a_1501_92# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VPWR a_595_97# a_757_401# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 Q a_2221_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND a_595_97# a_1261_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VPWR SET_B a_1339_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 Q_N a_1339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 Q a_2221_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VPWR a_595_97# a_1258_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X31 a_1531_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 VGND a_2221_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X36 a_595_97# a_225_74# a_706_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X37 a_757_401# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_1457_508# a_1470_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_1027_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_709_463# a_760_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 VGND a_1902_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# a_398_74# a_604_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_1215_74# a_398_74# a_1298_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_1500_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1902_74# a_1298_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 a_760_395# a_604_74# a_1027_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_1902_74# a_1298_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_1298_392# a_398_74# a_1457_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 VPWR a_224_350# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_604_74# a_224_350# a_709_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VPWR SET_B a_1298_392# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 VPWR a_604_74# a_1197_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_604_74# a_398_74# a_740_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_1422_74# a_1470_48# a_1500_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 VGND a_224_350# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR a_1902_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_1298_392# a_224_350# a_1422_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VGND a_604_74# a_1215_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_1197_341# a_224_350# a_1298_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_224_350# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_27_74# a_224_350# a_604_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 VGND a_1298_392# a_1470_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_224_350# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VPWR a_604_74# a_760_395# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 VPWR a_1298_392# a_1470_48# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X29 a_740_74# a_760_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X30 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_760_395# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_1489_118# a_1566_92# a_1596_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_716_456# a_767_384# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 VGND a_2022_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_74# a_225_74# a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_27_74# a_398_74# a_612_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_1266_341# a_225_74# a_1356_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_1356_74# a_398_74# a_1521_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 a_1356_74# a_225_74# a_1489_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 VPWR a_612_74# a_767_384# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 a_781_74# a_767_384# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 Q a_2022_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_1521_508# a_1566_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_767_384# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 a_612_74# a_225_74# a_716_456# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_1057_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_2022_94# a_1356_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 Q a_2022_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_1596_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VPWR SET_B a_1356_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X20 VPWR a_1356_74# a_1566_92# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 a_612_74# a_398_74# a_781_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_767_384# a_612_74# a_1057_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 VPWR a_2022_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_1278_74# a_398_74# a_1356_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 VPWR a_612_74# a_1266_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X30 VGND a_612_74# a_1278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X31 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 VGND a_1356_74# a_1566_92# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_2022_94# a_1356_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_1225_74# a_398_74# a_1321_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_1514_88# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 VPWR a_612_74# a_767_402# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 a_1220_347# a_225_74# a_1321_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR a_1321_392# a_1484_62# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 a_27_74# a_225_74# a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1436_88# a_1484_62# a_1514_88# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_767_402# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 VGND a_1940_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_767_402# a_612_74# a_1035_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_1035_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_612_74# a_398_74# a_732_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 VPWR a_1321_392# a_1940_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 VPWR a_1940_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_716_463# a_767_402# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 VPWR SET_B a_1321_392# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 Q a_1940_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Q a_1940_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_1940_74# a_1321_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Q a_1940_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_27_74# a_398_74# a_612_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 a_1321_392# a_225_74# a_1436_88# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_612_74# a_225_74# a_716_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 a_1321_392# a_398_74# a_1480_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 Q a_1940_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_1480_508# a_1484_62# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 VGND a_612_74# a_1225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X31 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 VPWR a_612_74# a_1220_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X33 a_1940_74# a_1321_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X34 VGND a_1321_392# a_1484_62# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 VPWR a_1940_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X36 a_732_74# a_767_402# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 VGND a_1940_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
X0 VGND D a_420_503# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 VPWR a_543_447# a_701_463# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VGND a_1644_94# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR D a_420_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 a_1158_482# a_1191_120# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_543_447# a_205_368# a_713_102# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_713_102# a_701_463# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_1644_94# a_1191_120# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VPWR a_1644_94# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_543_447# a_27_74# a_650_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_1191_120# a_1005_120# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VPWR a_1191_120# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND a_27_74# a_205_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_701_463# a_27_74# a_1005_120# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_420_503# a_27_74# a_543_447# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_1005_120# a_27_74# a_1143_146# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_650_508# a_701_463# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_1143_146# a_1191_120# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VGND a_1191_120# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_420_503# a_205_368# a_543_447# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 a_1191_120# a_1005_120# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_27_74# a_205_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_1005_120# a_205_368# a_1158_482# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_701_463# a_205_368# a_1005_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X25 a_1644_94# a_1191_120# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 VGND a_543_447# a_701_463# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X27 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
X0 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1248_128# a_1290_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND D a_451_503# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_753_284# a_206_368# a_1000_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VPWR a_1835_368# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_558_445# a_27_74# a_702_445# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VPWR a_1000_424# a_1290_102# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_1000_424# a_27_74# a_1248_128# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_753_284# a_27_74# a_1000_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_1290_102# a_1000_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 Q_N a_1835_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_558_445# a_206_368# a_717_102# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 VGND a_558_445# a_753_284# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X13 a_1835_368# a_1290_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_702_445# a_753_284# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_1208_479# a_1290_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 a_451_503# a_27_74# a_558_445# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 VPWR D a_451_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 VPWR a_1290_102# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Q_N a_1835_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Q a_1290_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND a_1835_368# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_451_503# a_206_368# a_558_445# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_1835_368# a_1290_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 VGND a_1290_102# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VPWR a_558_445# a_753_284# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X28 a_1290_102# a_1000_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_1000_424# a_206_368# a_1208_479# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 Q a_1290_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_717_102# a_753_284# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_454_503# a_206_368# a_561_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 a_1118_508# a_1210_314# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 VPWR a_561_463# a_713_458# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_1210_314# a_1011_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VPWR a_1210_314# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND a_1210_314# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_561_463# a_27_74# a_668_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_1210_314# a_1011_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_561_463# a_206_368# a_731_101# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VGND D a_454_503# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_1011_424# a_27_74# a_1168_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_1011_424# a_206_368# a_1118_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 a_668_503# a_713_458# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_1168_124# a_1210_314# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND a_561_463# a_713_458# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X18 a_713_458# a_27_74# a_1011_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 a_731_101# a_713_458# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_713_458# a_206_368# a_1011_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 VPWR D a_454_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_454_503# a_27_74# a_561_463# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_538_429# a_27_74# a_644_504# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 Q a_1217_314# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_695_459# a_206_368# a_1019_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VGND a_1217_314# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_695_459# a_27_74# a_1019_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_1125_508# a_1217_314# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 a_431_508# a_27_74# a_538_429# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_708_101# a_695_459# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_1217_314# a_1019_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_1172_124# a_1217_314# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Q a_1217_314# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR D a_431_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VGND a_538_429# a_695_459# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 a_1217_314# a_1019_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VPWR a_1217_314# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_1019_424# a_206_368# a_1125_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_431_508# a_206_368# a_538_429# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 VPWR a_538_429# a_695_459# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_644_504# a_695_459# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_538_429# a_206_368# a_708_101# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_1019_424# a_27_74# a_1172_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VGND D a_431_508# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
X0 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_651_503# a_696_458# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 VGND a_1226_296# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_544_485# a_696_458# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 a_1034_424# a_27_74# a_1178_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 VGND a_1226_296# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_1034_424# a_206_368# a_1141_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 a_1226_296# a_1034_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_544_485# a_206_368# a_735_102# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 Q a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_1226_296# a_1034_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Q a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Q a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Q a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_437_503# a_206_368# a_544_485# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X16 a_696_458# a_27_74# a_1034_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VPWR a_1034_424# a_1226_296# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 VGND D a_437_503# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_735_102# a_696_458# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_1141_508# a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_544_485# a_27_74# a_651_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 VPWR a_1226_296# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_696_458# a_206_368# a_1034_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X25 VPWR a_544_485# a_696_458# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 VPWR D a_437_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X27 a_437_503# a_27_74# a_544_485# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 VPWR a_1226_296# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_1178_124# a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



*
* Updated May 2, 2024 with subcircuit compatible with continuous models

.subckt sky130_fd_sc_hs__diode_2 DIODE VGND VNB VPB VPWR
XD0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=7.32e+06 area=6.417e+11
.ends



.subckt sky130_fd_sc_hs__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_27_74# a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_258_392# a_309_338# a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_83_260# a_315_54# a_484_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_267_80# a_315_54# a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VGND CLK a_984_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_987_393# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_477_124# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_315_54# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VGND GATE a_267_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_484_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 VPWR GATE a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND a_315_54# a_309_338# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR CLK a_987_393# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 a_984_125# a_27_74# a_987_393# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VPWR a_315_54# a_309_338# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_83_260# a_309_338# a_477_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 VPWR a_987_393# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_27_74# a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VGND a_987_393# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_315_54# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_27_74# a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR a_1041_387# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_1044_119# a_27_74# a_1041_387# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_315_48# a_315_338# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_508_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_494_118# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_1041_387# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_1041_387# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 GCLK a_1041_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_83_244# a_315_338# a_494_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VGND CLK a_1044_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_315_48# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR GATE a_264_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_83_244# a_315_48# a_508_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_267_74# a_315_48# a_83_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VGND a_315_48# a_315_338# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_315_48# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 GCLK a_1041_387# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VGND GATE a_267_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_27_74# a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_264_392# a_315_338# a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VPWR CLK a_1041_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_1047_74# a_27_74# a_1044_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_524_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 GCLK a_1044_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_334_54# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# a_84_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_1044_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_1044_368# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR GATE a_283_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND CLK a_1047_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 GCLK a_1044_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR CLK a_1044_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 GCLK a_1044_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND a_1044_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_283_392# a_334_338# a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_286_80# a_334_54# a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VPWR a_1044_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_334_54# a_334_338# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND GATE a_286_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 VPWR a_334_54# a_334_338# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 GCLK a_1044_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR a_1044_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_334_54# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 a_491_124# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_84_48# a_334_54# a_524_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_27_74# a_84_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_84_48# a_334_338# a_491_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_802_508# a_889_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 VGND a_889_92# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_373_74# a_231_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VPWR a_1437_112# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_889_92# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_608_74# a_231_74# a_686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_1133_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND a_27_424# a_608_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_1437_112# a_889_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_373_74# a_231_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_841_118# a_889_92# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VPWR a_27_424# a_611_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VPWR a_686_74# a_889_92# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_611_392# a_373_74# a_686_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VGND GATE_N a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_1437_112# a_889_92# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 VPWR GATE_N a_231_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_686_74# a_231_74# a_802_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_889_92# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_686_74# a_373_74# a_841_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_27_424# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 a_889_92# a_686_74# a_1133_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_424# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X23 VGND a_1437_112# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR GATE_N a_230_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND a_27_112# a_592_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_670_74# a_230_74# a_783_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_838_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_1446_368# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR a_27_112# a_595_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_363_74# a_230_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_838_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND a_838_48# a_1446_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_790_74# a_838_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 Q_N a_1446_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_363_74# a_230_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_1066_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_595_392# a_363_74# a_670_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 Q a_838_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_27_112# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 a_838_48# a_670_74# a_1066_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND a_838_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_783_508# a_838_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 VGND GATE_N a_230_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 Q_N a_1446_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_27_112# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 a_670_74# a_363_74# a_790_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 Q a_838_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR a_838_48# a_1446_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 VPWR a_1446_368# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_592_74# a_230_74# a_670_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 VPWR a_670_74# a_838_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR a_823_98# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_642_392# a_353_98# a_753_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 a_753_508# a_823_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 VPWR a_1342_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR GATE a_226_104# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_823_98# a_642_392# a_1051_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_142# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_353_98# a_226_104# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_642_392# a_226_104# a_775_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VGND a_27_142# a_571_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR a_27_142# a_564_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND GATE a_226_104# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_1051_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_353_98# a_226_104# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_142# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 VPWR a_642_392# a_823_98# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_823_98# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_564_392# a_226_104# a_642_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_823_98# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_1342_74# a_823_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X20 a_571_80# a_353_98# a_642_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_1342_74# a_823_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 a_775_124# a_823_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VGND a_1342_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 Q a_821_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1449_368# a_821_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_569_80# a_363_82# a_641_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 Q a_821_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_27_112# a_566_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_821_98# a_641_80# a_1049_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_821_98# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_641_80# a_821_98# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_641_80# a_230_74# a_773_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR GATE a_230_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_641_80# a_363_82# a_757_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_27_112# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_757_508# a_821_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 a_363_82# a_230_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_821_98# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_27_112# a_569_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 VGND a_1449_368# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR a_821_98# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 Q_N a_1449_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_1449_368# a_821_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_27_112# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 VGND GATE a_230_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Q_N a_1449_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_1049_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_566_392# a_230_74# a_641_80# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_773_124# a_821_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 VPWR a_1449_368# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_363_82# a_230_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_570_392# a_357_392# a_654_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 VPWR a_654_392# a_897_406# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_357_392# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_681_74# a_232_98# a_654_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_1139_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_357_392# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_897_406# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_793_508# a_897_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 VPWR a_897_406# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_654_392# a_232_98# a_793_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_897_406# a_654_392# a_1139_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND a_27_136# a_681_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_654_392# a_357_392# a_854_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 VPWR a_27_136# a_570_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_854_74# a_897_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VGND a_897_406# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_697_74# a_232_98# a_670_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_586_392# a_373_82# a_670_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_27_136# a_697_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 VPWR a_913_406# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_778_504# a_913_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 VPWR a_27_136# a_586_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_670_392# a_373_82# a_870_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_670_392# a_232_98# a_778_504# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 a_870_74# a_913_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 VGND a_913_406# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR a_670_392# a_913_406# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_373_82# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_1153_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_913_406# a_670_392# a_1153_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_373_82# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_913_406# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 Q a_913_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 Q a_913_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR a_27_136# a_561_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_666_74# a_232_98# a_639_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_888_406# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VPWR a_888_406# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_27_136# a_666_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_639_392# a_348_392# a_839_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X9 a_839_74# a_888_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VGND a_888_406# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_888_406# a_639_392# a_1035_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 VPWR a_888_406# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_747_504# a_888_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_1035_74# a_639_392# a_888_406# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_888_406# a_639_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 Q a_888_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_1035_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 Q a_888_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR RESET_B a_888_406# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_348_392# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 a_639_392# a_232_98# a_747_504# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X23 VGND a_888_406# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_561_392# a_348_392# a_639_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_348_392# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VGND RESET_B a_1035_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 Q a_888_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 VPWR a_639_392# a_888_406# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X29 Q a_888_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 VPWR GATE a_216_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR a_643_74# a_817_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_1045_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_817_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_568_392# a_216_424# a_643_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_565_74# a_363_74# a_643_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_769_74# a_817_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VGND GATE a_216_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND a_27_424# a_565_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_643_74# a_216_424# a_769_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_759_508# a_817_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_27_424# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X12 a_817_48# a_643_74# a_1045_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR a_27_424# a_568_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VPWR a_817_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_817_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_424# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_643_74# a_363_74# a_759_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_363_74# a_216_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 a_363_74# a_216_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
X0 VGND GATE a_235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_568_74# a_347_98# a_646_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VGND a_27_392# a_568_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VPWR a_646_74# a_832_55# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND a_832_55# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Q a_832_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR GATE a_235_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_347_98# a_235_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VPWR a_27_392# a_565_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_27_392# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_832_55# a_646_74# a_1060_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_565_392# a_235_74# a_646_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_784_81# a_832_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_646_74# a_347_98# a_756_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VPWR a_832_55# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Q a_832_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_646_74# a_235_74# a_784_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_832_55# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_27_392# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X19 a_347_98# a_235_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_756_508# a_832_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 a_1060_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
X0 Q a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_755_74# a_797_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_562_392# a_240_394# a_640_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VPWR RESET_B a_797_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 Q a_797_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR GATE a_240_394# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_938_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_27_126# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VGND GATE a_240_394# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_797_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Q a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_797_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_797_48# a_640_74# a_938_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VGND a_797_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_126# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 VGND RESET_B a_938_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 VPWR a_797_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_640_74# a_364_120# a_747_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 Q a_797_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_364_120# a_240_394# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_747_508# a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 a_559_74# a_364_120# a_640_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_797_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR a_640_74# a_797_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X24 VPWR a_27_126# a_562_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_364_120# a_240_394# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_938_74# a_640_74# a_797_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 VGND a_27_126# a_559_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 a_797_48# a_640_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X29 a_640_74# a_240_394# a_755_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 a_653_79# a_343_80# a_852_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 VPWR a_1347_424# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_805_392# a_863_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_27_120# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VPWR a_653_79# a_863_294# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR a_863_294# a_1347_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND a_863_294# a_1347_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 VPWR GATE_N a_232_82# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_653_79# a_232_82# a_805_392# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 Q a_863_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND GATE_N a_232_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_575_79# a_232_82# a_653_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_343_80# a_232_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND a_27_120# a_575_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_27_120# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 a_852_123# a_863_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_343_80# a_232_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 Q a_863_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR a_27_120# a_571_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VGND a_653_79# a_863_294# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_571_392# a_343_80# a_653_79# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VGND a_1347_424# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_27_136# a_569_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VGND a_647_79# a_887_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VPWR a_887_270# a_1442_94# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_647_79# a_232_98# a_814_392# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 VPWR a_647_79# a_887_270# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR a_27_136# a_565_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR a_887_270# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_565_392# a_343_74# a_647_79# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 Q a_887_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND a_1442_94# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Q_N a_1442_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VGND a_887_270# a_1442_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_343_74# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_839_123# a_887_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 Q_N a_1442_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND a_887_270# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_343_74# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 a_647_79# a_343_74# a_839_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 Q a_887_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_814_392# a_887_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 VPWR a_1442_94# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_569_79# a_232_98# a_647_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
X0 a_770_508# a_863_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 VGND a_1347_424# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Q a_863_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_664_392# a_863_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_863_98# a_1347_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_373_82# a_231_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_664_392# a_863_98# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_664_392# a_231_74# a_815_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_589_80# a_373_82# a_664_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_373_82# a_231_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 VPWR a_27_413# a_586_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 Q a_863_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND a_27_413# a_589_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VPWR GATE a_231_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 VGND GATE a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND a_863_98# a_1347_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 a_27_413# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X17 a_586_392# a_231_74# a_664_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_27_413# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 VPWR a_1347_424# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_664_392# a_373_82# a_770_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 a_815_124# a_863_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
X0 a_27_115# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 VPWR a_669_392# a_863_441# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_669_392# a_369_392# a_871_139# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_655_79# a_217_419# a_669_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_27_115# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_669_392# a_217_419# a_812_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VGND GATE_N a_217_419# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND a_27_115# a_655_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_871_139# a_863_441# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_812_508# a_863_441# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 VGND a_669_392# a_863_441# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VPWR GATE_N a_217_419# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 VPWR a_27_115# a_585_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_369_392# a_217_419# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VGND a_863_441# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_585_392# a_369_392# a_669_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VPWR a_863_441# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_369_392# a_217_419# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
X0 VPWR GATE_N a_232_82# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_669_392# a_369_392# a_875_139# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VPWR a_842_405# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_120# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VGND GATE_N a_232_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND a_669_392# a_842_405# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_842_405# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Q a_842_405# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_120# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X9 VPWR a_27_120# a_585_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_369_392# a_232_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_669_392# a_232_82# a_791_503# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 Q a_842_405# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_585_392# a_369_392# a_669_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_791_503# a_842_405# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_658_79# a_232_82# a_669_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_369_392# a_232_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_875_139# a_842_405# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 VPWR a_669_392# a_842_405# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND a_27_120# a_658_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
X0 a_27_115# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 Q a_840_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR GATE_N a_230_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VPWR a_27_115# a_591_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 Q a_840_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_591_392# a_369_392# a_675_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND GATE_N a_230_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_675_392# a_369_392# a_895_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_895_123# a_840_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VGND a_675_392# a_840_395# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VGND a_840_395# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Q a_840_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_840_395# a_675_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_840_395# a_675_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 VPWR a_840_395# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_27_115# D VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_789_508# a_840_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 a_369_392# a_230_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR a_840_395# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Q a_840_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_658_79# a_230_424# a_675_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_369_392# a_230_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 VGND a_840_395# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND a_27_115# a_658_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_675_392# a_230_424# a_789_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 VPWR a_675_392# a_840_395# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlxtp_1 D GATE VGND VNB VPB VPWR Q
X0 a_592_149# a_685_59# a_239_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_386_326# a_514_149# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_229_392# a_562_123# a_592_149# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND D a_116_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VGND a_386_326# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_562_123# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_239_85# a_116_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_386_326# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_386_326# a_592_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_229_392# a_116_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VPWR a_386_326# a_419_392# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_592_149# a_685_59# a_419_392# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_386_326# a_592_149# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_514_149# a_562_123# a_592_149# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 a_562_123# GATE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 VPWR D a_116_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 VGND a_562_123# a_685_59# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR a_562_123# a_685_59# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlygate4sd1_1 A VGND VNB VPB VPWR X
X0 a_405_138# a_288_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.18
X1 VGND a_405_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_405_138# a_288_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.18
X5 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VPWR a_405_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__dlygate4sd2_1 A VGND VNB VPB VPWR X
X0 a_405_138# a_288_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X1 VGND a_405_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_405_138# a_288_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.25
X4 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 VGND a_28_74# a_288_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X6 VPWR a_28_74# a_288_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.25
X7 VPWR a_405_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 a_405_138# a_289_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X1 VPWR a_28_74# a_289_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X2 VGND a_405_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VGND a_28_74# a_289_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.18
X5 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 a_405_138# a_289_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.50
X7 VPWR a_405_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 VGND a_28_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_316_138# X VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_604_138# a_785_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_28_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_316_138# a_497_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_604_138# a_497_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VPWR a_604_138# a_785_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_28_138# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 VGND a_316_138# a_497_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_28_138# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_316_138# X VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_604_138# a_497_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlymetal6s4s_1 A VGND VNB VPB VPWR X
X0 VGND a_28_138# a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_316_138# a_209_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_604_138# a_785_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_28_138# a_209_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_316_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_604_138# X VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VPWR a_604_138# a_785_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_28_138# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 VGND a_316_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_28_138# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_316_138# a_209_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_604_138# X VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__dlymetal6s6s_1 A VGND VNB VPB VPWR X
X0 VGND a_28_138# a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_316_138# a_209_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_604_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_28_138# a_209_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_316_138# a_497_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_604_138# a_497_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VPWR a_604_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_28_138# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 VGND a_316_138# a_497_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_28_138# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_316_138# a_209_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_604_138# a_497_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__ebufn_1 A TE_B VGND VNB VPB VPWR Z
X0 VGND A a_229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 VPWR A a_229_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_27_404# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_566_368# a_229_74# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_27_404# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 VPWR TE_B a_566_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_569_74# a_229_74# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND a_27_404# a_569_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__ebufn_2 A TE_B VGND VNB VPB VPWR Z
X0 VPWR TE_B a_33_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_283_48# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND A a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_33_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR A a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_27_74# a_283_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_283_48# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 Z a_84_48# a_33_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND a_283_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_33_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__ebufn_4 A TE_B VGND VNB VPB VPWR Z
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_378_74# a_208_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_348_368# a_27_368# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Z a_27_368# a_378_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_208_74# a_378_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_348_368# a_27_368# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Z a_27_368# a_348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND TE_B a_208_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR TE_B a_208_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_378_74# a_27_368# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_348_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR TE_B a_348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Z a_27_368# a_378_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR TE_B a_348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Z a_27_368# a_348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_378_74# a_208_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_378_74# a_27_368# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VGND a_208_74# a_378_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_348_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__ebufn_8 A TE_B VGND VNB VPB VPWR Z
X0 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_833_48# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR A a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_84_48# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_84_48# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_833_48# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
X0 a_1334_97# a_1419_71# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_27_74# a_818_74# a_1198_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_1419_71# a_1807_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR DE a_556_504# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 VPWR a_818_74# a_1008_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_2227_118# a_575_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_161_446# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VPWR a_1879_74# a_575_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_116_508# a_161_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 VPWR a_575_48# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_74# D a_145_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_2008_392# a_818_74# a_1879_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_161_446# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X13 a_556_504# a_575_48# a_27_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 VGND a_818_74# a_1008_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR CLK a_818_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_1423_508# a_1419_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 a_1807_74# a_1008_74# a_1879_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_27_74# a_1008_74# a_1198_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 VPWR a_1198_97# a_1419_71# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_1879_74# a_818_74# a_2227_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_1198_97# a_818_74# a_1423_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 VGND a_575_48# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_527_74# a_575_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 VGND a_1198_97# a_1419_71# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 Q a_1879_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 VGND a_161_446# a_527_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VGND a_1879_74# a_575_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 a_1198_97# a_1008_74# a_1334_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 VGND CLK a_818_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 Q a_1879_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_145_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 VPWR a_1419_71# a_2008_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X33 a_2206_443# a_575_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X34 a_27_74# D a_116_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X35 a_1879_74# a_1008_74# a_2206_443# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
X0 VPWR DE a_554_436# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_1997_74# a_533_61# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VPWR a_1156_90# a_1409_64# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VGND a_1409_64# a_1797_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_131_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_1797_74# a_958_74# a_1895_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_1156_90# a_763_74# a_1382_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 a_1382_508# a_1409_64# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 VGND a_763_74# a_958_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_763_74# a_958_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_554_436# a_533_61# a_27_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_159_446# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_1349_90# a_1409_64# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VGND CLK a_763_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_1895_74# a_958_74# a_2088_502# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 Q a_1895_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_508# D a_114_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 VPWR a_1895_74# a_533_61# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X18 VPWR CLK a_763_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Q a_1895_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_27_508# a_763_74# a_1156_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VGND a_159_446# a_491_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 a_27_508# a_958_74# a_1156_90# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 a_1156_90# a_958_74# a_1349_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 VGND a_1895_74# a_533_61# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_1895_74# a_763_74# a_1997_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 VPWR a_1409_64# a_1794_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_114_508# a_159_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 VGND a_1156_90# a_1409_64# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 a_27_508# D a_131_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X30 a_491_87# a_533_61# a_27_508# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_159_446# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X32 a_1794_392# a_763_74# a_1895_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X33 a_2088_502# a_533_61# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvn_1 A TE_B VGND VNB VPB VPWR Z
X0 a_22_46# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 a_278_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND a_22_46# a_281_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR TE_B a_278_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_281_100# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_22_46# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvn_2 A TE_B VGND VNB VPB VPWR Z
X0 a_231_74# a_115_464# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR TE_B a_227_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Z A a_227_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_115_464# a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Z A a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_231_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_227_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND TE_B a_115_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_227_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR TE_B a_115_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvn_4 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_281_74# a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_241_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR TE_B a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR TE_B a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Z A a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Z A a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_241_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR TE_B a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_281_74# a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_114_74# a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND a_114_74# a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Z A a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_281_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_241_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_241_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_281_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND TE_B a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvn_8 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VPWR TE_B a_126_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND TE_B a_126_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__einvp_1 A TE VGND VNB VPB VPWR Z
X0 VGND TE a_318_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_310_392# A Z VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_44_549# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_44_549# TE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 VPWR a_44_549# a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_318_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvp_2 A TE VGND VNB VPB VPWR Z
X0 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Z A a_36_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_36_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_368# a_263_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_36_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND TE a_36_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR a_263_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_263_323# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_263_323# TE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvp_4 A TE VGND VNB VPB VPWR Z
X0 a_27_368# a_473_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_473_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_27_368# a_473_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_473_323# TE VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_473_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_473_323# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__einvp_8 A TE VGND VNB VPB VPWR Z
X0 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_802_323# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_802_323# TE VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VGND a_465_249# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_217_368# B a_318_389# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR A a_217_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND A a_936_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_315_75# CIN a_69_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_318_389# CIN a_69_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_237_75# B a_315_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_69_260# a_465_249# a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VGND B a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 SUM a_69_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_465_249# CIN a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_509_347# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VGND A a_237_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VPWR A a_509_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_509_347# CIN VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_1107_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VPWR a_465_249# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR B a_1107_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_1100_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_69_260# a_465_249# a_509_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 a_501_75# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_936_75# B a_465_249# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_501_75# CIN VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 VPWR A a_916_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X24 a_916_347# B a_465_249# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 VGND A a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 a_465_249# CIN a_1107_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 SUM a_69_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_27_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_1094_347# B a_1202_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND CIN a_701_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND A a_701_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_992_347# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_1202_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND a_336_347# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_336_347# B a_484_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_701_79# a_336_347# a_992_347# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_27_378# CIN a_336_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 COUT a_336_347# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND B a_27_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_484_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_683_347# a_336_347# a_992_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 COUT a_336_347# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND a_992_347# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_992_347# CIN a_1119_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_487_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_336_347# B a_487_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_683_347# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 SUM a_992_347# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_1205_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_378# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_1119_79# B a_1205_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 SUM a_992_347# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_992_347# CIN a_1094_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X26 VPWR B a_27_378# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 VPWR a_336_347# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_27_79# CIN a_336_347# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VPWR A a_683_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X30 VPWR CIN a_683_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X31 a_701_79# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_418_74# B a_535_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_1141_347# B a_1235_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND CIN a_734_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_734_74# a_418_74# a_1024_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR CIN a_737_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_737_347# a_418_74# a_1024_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND A a_734_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_1024_74# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR a_418_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 COUT a_418_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_737_347# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_1024_74# CIN a_1160_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_1024_74# CIN a_1141_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VPWR A a_737_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_1235_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VPWR a_1024_74# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_27_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 COUT a_418_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_392# CIN a_418_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 VGND a_1024_74# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 COUT a_418_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VGND a_418_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 SUM a_1024_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_1238_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 SUM a_1024_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 SUM a_1024_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_418_74# B a_532_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_1160_74# B a_1238_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_535_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X30 VPWR a_418_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_27_74# CIN a_418_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 a_532_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 VGND a_1024_74# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 VGND a_418_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 VPWR B a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X36 SUM a_1024_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 COUT a_418_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 a_734_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
X0 SUM a_83_21# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 COUT a_410_58# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_1849_374# a_879_55# a_811_379# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_879_55# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_231_132# a_811_379# a_83_21# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_1660_374# a_879_55# a_1023_379# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_1023_379# B a_1849_374# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_1849_374# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_410_58# a_1023_379# a_231_132# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_1849_374# a_879_55# a_1023_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_644_104# a_811_379# a_83_21# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 VGND a_231_132# a_644_104# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 VGND A a_2342_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_879_55# a_811_379# a_410_58# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_1849_374# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_410_58# a_1023_379# a_879_55# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_83_21# a_1023_379# a_231_132# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 SUM a_83_21# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_811_379# B a_1660_374# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_231_132# a_811_379# a_410_58# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_83_21# a_1023_379# a_644_104# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VPWR a_231_132# a_644_104# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 VPWR A a_2342_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_1023_379# B a_1660_374# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X24 a_1660_374# a_2342_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_1660_374# a_879_55# a_811_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 a_1660_374# a_2342_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VPWR CI a_231_132# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X28 a_879_55# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VGND CI a_231_132# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X30 COUT a_410_58# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_811_379# B a_1849_374# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
X0 a_1689_424# a_849_424# a_1895_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_849_424# a_481_379# a_413_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_1689_424# a_514_424# a_1895_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VPWR a_1451_424# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_413_392# a_481_379# a_514_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_1895_424# a_849_424# a_2052_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR a_1895_424# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND CI a_1689_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_1451_424# a_849_424# a_1689_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_114_368# B a_849_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_114_368# a_481_379# a_849_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_481_379# a_514_424# a_1451_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 SUM a_1895_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR a_81_260# a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VGND A a_413_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VGND B a_481_379# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 SUM a_1895_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_81_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 VGND a_1895_424# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_1895_424# a_514_424# a_2052_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_481_379# a_849_424# a_1451_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_2052_424# a_1689_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 VPWR A a_413_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_413_392# B a_514_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 VPWR CI a_1689_424# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 COUT a_1451_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 COUT a_1451_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_514_424# B a_114_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X28 VGND a_81_260# a_114_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_849_424# B a_413_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X30 VPWR B a_481_379# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 VGND a_1451_424# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 a_1451_424# a_514_424# a_1689_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X33 a_2052_424# a_1689_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X34 a_81_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X35 a_514_424# a_481_379# a_114_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
X0 a_1183_102# a_1378_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_536_114# a_586_257# a_427_362# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_1378_125# CI VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_427_362# B a_536_114# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 SUM a_1278_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_586_257# a_528_362# a_1265_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 COUT a_1265_379# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 SUM a_1278_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 COUT a_1265_379# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_1265_379# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND a_1265_379# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_1378_125# CI VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VPWR a_27_74# a_427_362# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_200_74# B a_528_362# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_1183_102# a_528_362# a_1278_102# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_427_362# B a_528_362# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_1278_102# a_536_114# a_1378_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_1183_102# a_1378_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_1278_102# a_536_114# a_1183_102# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 VGND a_27_74# a_427_362# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VPWR a_1278_102# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VGND B a_586_257# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 COUT a_1265_379# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_200_74# B a_536_114# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 VPWR B a_586_257# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VPWR a_1265_379# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_1378_125# a_528_362# a_1265_379# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 SUM a_1278_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_528_362# a_586_257# a_200_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X31 a_1378_125# a_528_362# a_1278_102# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X32 VPWR a_1265_379# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 VPWR a_1278_102# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 a_1265_379# a_536_114# a_586_257# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X35 VGND a_1278_102# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 COUT a_1265_379# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 a_536_114# a_586_257# a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X38 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X39 VGND a_1278_102# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 VPWR A a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X41 a_1265_379# a_536_114# a_1378_125# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X42 a_528_362# a_586_257# a_427_362# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X43 SUM a_1278_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 COUT a_430_418# a_1595_400# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_492_48# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_1967_384# a_608_74# a_2004_136# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_1197_368# a_430_418# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_28_74# B a_608_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_1854_368# a_608_74# a_2004_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_608_74# a_492_48# a_256_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_256_368# B a_608_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VGND a_28_74# a_256_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_430_418# a_492_48# a_28_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR a_492_48# a_1197_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VPWR a_28_74# a_256_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_1967_384# a_1854_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_608_74# a_492_48# a_28_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 VGND a_2004_136# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_1595_400# CIN VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND a_492_48# a_1197_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 a_1595_400# CIN VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_2004_136# a_430_418# a_1854_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_1967_384# a_1854_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VPWR CIN a_1854_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR a_2004_136# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_2004_136# a_430_418# a_1967_384# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_430_418# a_492_48# a_256_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X25 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_492_48# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 COUT a_608_74# a_1595_400# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 a_28_74# B a_430_418# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X29 a_1197_368# a_608_74# COUT VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X30 a_256_368# B a_430_418# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X31 VGND CIN a_1854_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
X0 a_369_365# B a_27_100# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_27_100# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_1023_389# a_374_120# COUT_N VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_369_365# B a_241_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 COUT_N a_369_365# a_1261_421# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_241_368# a_336_263# a_374_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_1719_368# a_369_365# a_1744_94# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 VPWR CI a_1606_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND B a_1023_389# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_1261_421# CI VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR B a_1023_389# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_27_100# a_336_263# a_369_365# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_27_100# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_1744_94# a_374_120# a_1719_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_241_368# a_336_263# a_369_365# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_336_263# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_336_263# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_1261_421# CI VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 VPWR a_1744_94# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_1606_368# a_369_365# a_1744_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_27_100# a_336_263# a_374_120# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 a_1744_94# a_374_120# a_1606_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 VGND CI a_1606_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND a_1744_94# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 VPWR a_27_100# a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_374_120# B a_241_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 a_1719_368# a_1606_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_1719_368# a_1606_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 VGND a_27_100# a_241_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 a_1023_389# a_369_365# COUT_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X30 a_374_120# B a_27_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X31 COUT_N a_374_120# a_1261_421# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__fill_1 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__fill_2 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__fill_4 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__fill_8 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__fill_diode_2 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__fill_diode_4 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__fill_diode_8 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__ha_1 A B VGND VNB VPB VPWR COUT SUM
X0 SUM a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR a_239_294# a_83_260# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR B a_239_294# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VGND A a_305_130# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_239_294# B a_695_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_83_260# B a_386_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_695_119# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_305_130# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_239_294# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VPWR a_239_294# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_386_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_83_260# a_239_294# a_305_130# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 SUM a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND a_239_294# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__ha_2 A B VGND VNB VPB VPWR COUT SUM
X0 a_391_388# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_278_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_391_388# a_27_74# a_278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_27_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR A a_307_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR a_391_388# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR a_27_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 COUT a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 COUT a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR B a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 SUM a_391_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_307_388# B a_391_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 SUM a_391_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VGND A a_278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND a_391_388# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_74# B a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__ha_4 A B VGND VNB VPB VPWR COUT SUM
X0 SUM a_294_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR B a_435_99# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VGND B a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_435_99# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 COUT a_435_99# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_707_119# B a_435_99# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 SUM a_294_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_294_392# a_435_99# a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VGND a_435_99# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_294_392# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_435_99# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 VGND a_294_392# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_294_392# B a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 SUM a_294_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_435_99# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_294_392# a_435_99# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_435_99# B a_707_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 COUT a_435_99# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 SUM a_294_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 COUT a_435_99# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_27_125# a_435_99# a_294_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VGND A a_707_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_27_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 VPWR a_435_99# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_27_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X26 a_707_119# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 COUT a_435_99# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR a_294_392# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_27_125# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X30 VPWR a_294_392# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_27_392# B a_294_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X32 VPWR A a_435_99# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X33 VGND A a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X34 VPWR a_435_99# a_294_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X35 VPWR a_435_99# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__inv_1 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__inv_8 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__maj3_1 A B C VGND VNB VPB VPWR X
X0 a_223_120# B a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_226_384# B a_84_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_406_384# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_84_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND A a_223_120# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_403_136# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 VPWR A a_226_384# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_595_136# C a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_84_74# B a_406_384# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_598_384# C a_84_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VGND A a_595_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 X a_84_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_84_74# B a_403_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VPWR A a_598_384# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__maj3_2 A B C VGND VNB VPB VPWR X
X0 a_393_368# B a_87_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_87_264# B a_577_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A a_790_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_413_74# B a_87_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_793_74# C a_87_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 X a_87_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND a_87_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A a_413_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND A a_793_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_790_368# C a_87_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_87_264# B a_584_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_577_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_584_347# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 X a_87_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR a_87_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A a_393_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__maj3_4 A B C VGND VNB VPB VPWR X
X0 X a_219_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_119_392# B a_219_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_501_392# B a_219_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_219_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A a_906_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_119_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_905_392# C a_219_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_219_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_219_392# B a_114_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_219_392# C a_905_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_219_392# B a_501_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_504_125# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 X a_219_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_114_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VPWR a_219_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_501_392# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 X a_219_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR C a_501_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 VPWR a_219_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_219_392# B a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 a_906_78# C a_219_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_219_392# C a_906_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR A a_905_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VGND a_219_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 VGND A a_114_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 VGND C a_504_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 a_114_125# B a_219_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 VPWR A a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X28 a_905_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X29 a_219_392# B a_504_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X30 a_504_125# B a_219_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X31 a_906_78# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 a_27_112# S VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_304_74# A1 a_524_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_443_74# a_27_112# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_226_74# A1 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR S a_223_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND S a_226_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_524_368# a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_27_112# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 VGND a_304_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_223_368# A0 a_304_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_304_74# A0 a_443_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR a_304_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 a_27_368# A0 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 X a_116_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_116_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_459_48# a_38_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_459_48# S VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 X a_116_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_270_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_459_48# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X9 a_116_368# A1 a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VPWR a_116_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR a_459_48# a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_38_74# A0 a_116_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_116_368# A1 a_270_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X
X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
X0 a_426_74# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_114_74# a_426_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR S a_114_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_223_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_223_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y A1 a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y A1 a_399_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR a_114_74# a_399_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_225_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND S a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
X0 VPWR a_922_72# a_340_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_115_74# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y A1 a_340_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_340_368# a_922_72# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_340_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_118_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR S a_922_72# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_337_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND S a_337_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_922_72# a_115_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y A1 a_337_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y A0 a_118_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND S a_922_72# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_337_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR S a_118_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Y A0 a_115_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_115_74# a_922_72# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_118_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
X0 Y A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_114_85# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND a_1030_268# a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_1030_268# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_475_85# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_114_85# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_116_368# a_1030_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_475_85# a_1030_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y A0 a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_478_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR S a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_475_85# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_1030_268# S VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 Y A1 a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y A0 a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_478_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_116_368# a_1030_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_116_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Y A1 a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 Y A0 a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_116_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_114_85# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_475_85# a_1030_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 VPWR S a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND S a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VGND S a_1030_268# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VGND a_1030_268# a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_478_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR S a_1030_268# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X30 VGND S a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 Y A0 a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_478_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 VPWR a_1030_268# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 a_114_85# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 VPWR a_1338_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_846_74# S0 a_979_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_1338_125# a_1396_99# a_342_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_1396_99# S1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_255_341# S0 a_342_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_264_74# a_27_74# a_342_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_846_74# S1 a_1338_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VGND A0 a_264_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_342_74# S0 a_450_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_979_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_27_74# S0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_537_341# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_768_74# a_27_74# a_846_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_846_74# a_27_74# a_1065_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_342_74# S1 a_1338_125# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VGND a_1338_125# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND A2 a_768_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_1065_387# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_342_74# a_27_74# a_537_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 a_450_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_763_341# S0 a_846_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VPWR A0 a_255_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_1338_125# a_1396_99# a_846_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_1396_99# S1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X24 VPWR A2 a_763_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 a_27_74# S0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_909_74# S0 a_1152_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_255_74# S0 a_333_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR a_1429_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_1429_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_333_74# S0 a_618_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_1152_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND A1 a_255_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_1429_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A3 a_831_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_1429_74# a_1500_94# a_333_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_31_94# S0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_1429_74# a_1500_94# a_909_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_909_74# a_31_94# a_1047_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_1047_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_1500_94# S1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_831_74# S0 a_909_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VPWR A3 a_840_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_1500_94# S1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 a_333_74# a_31_94# a_507_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_507_74# A0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_840_392# a_31_94# a_909_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 a_618_392# A0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_333_74# S1 a_1429_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 a_31_94# S0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_909_74# S1 a_1429_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 X a_1429_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VPWR A1 a_264_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_264_392# a_31_94# a_333_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_509_392# S1 a_2199_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_2199_74# a_2489_347# a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_116_392# a_758_306# a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_1285_377# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_1450_121# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_1278_121# a_758_306# a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_1285_377# a_758_306# a_1191_121# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND A2 a_1278_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_1465_377# S0 a_1191_121# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_2199_74# a_2489_347# a_1191_121# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VPWR A2 a_1465_377# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_509_392# a_2489_347# a_2199_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_509_392# a_758_306# a_299_126# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_758_306# S0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_114_126# S0 a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VPWR A1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_296_392# S0 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_509_392# S0 a_114_126# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 a_1450_121# S0 a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 VGND A3 a_1450_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_1191_121# S0 a_1450_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_1191_121# a_2489_347# a_2199_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 VPWR a_2199_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_1278_121# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_758_306# S0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_2199_74# S1 a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 VPWR A0 a_296_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_509_392# a_758_306# a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X28 VGND A1 a_114_126# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 X a_2199_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 X a_2199_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VGND A0 a_299_126# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X32 a_299_126# a_758_306# a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X33 a_2489_347# S1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_1191_121# a_758_306# a_1285_377# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X35 a_1191_121# S1 a_2199_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X36 a_114_126# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X37 X a_2199_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_1191_121# S0 a_1465_377# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X39 a_296_392# A0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X40 a_509_392# S0 a_296_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X41 VPWR A3 a_1285_377# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X42 X a_2199_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X43 VGND a_2199_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X44 VGND a_2199_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X45 a_1465_377# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X46 a_2199_74# S1 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X47 a_299_126# A0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X48 a_2489_347# S1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X49 a_1191_121# a_758_306# a_1278_121# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X50 a_116_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X51 VPWR a_2199_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2_1 A B VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_117_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND B a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2_2 A B VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y
X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 a_27_112# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_112# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 a_269_74# a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND B a_269_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2b_2 A_N B VGND VNB VPB VPWR Y
X0 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 Y a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y a_27_74# a_242_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND B a_242_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_242_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_27_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_242_74# a_27_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand2b_4 A_N B VGND VNB VPB VPWR Y
X0 Y a_31_74# a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR a_31_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A_N a_31_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_243_74# a_31_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND B a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_31_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_243_74# a_31_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_243_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y a_31_74# a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND B a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_31_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 Y a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_243_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand3_1 A B C VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_155_74# B a_233_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND C a_155_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_233_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand3_2 A B C VGND VNB VPB VPWR Y
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND C a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_27_74# B a_283_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_283_74# B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_283_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y A a_283_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand3_4 A B C VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y A a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_27_82# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_82# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_82# B a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_456_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND C a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_27_82# B a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND C a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y A a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_456_82# B a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_456_82# B a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_456_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand3b_1 A_N B C VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_116# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_116# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 a_269_78# B a_347_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND C a_269_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_347_78# a_27_116# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_27_116# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand3b_2 A_N B C VGND VNB VPB VPWR Y
X0 Y a_27_94# a_403_54# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_403_54# B a_206_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_27_94# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_206_74# B a_403_54# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND C a_206_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_94# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_206_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_403_54# a_27_94# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y a_27_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_94# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand3b_4 A_N B C VGND VNB VPB VPWR Y
X0 Y a_89_172# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_297_82# B a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR a_89_172# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND C a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_297_82# B a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_744_74# a_89_172# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y a_89_172# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR A_N a_89_172# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_297_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_89_172# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_744_74# a_89_172# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_297_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y a_89_172# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND C a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_744_74# B a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_89_172# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_744_74# B a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 VGND D a_181_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_259_74# B a_373_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_373_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_181_74# C a_259_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4_2 A B C D VGND VNB VPB VPWR Y
X0 a_515_74# B a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_515_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND D a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_74# C a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_304_74# C a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y A a_515_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_304_74# B a_515_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4_4 A B C D VGND VNB VPB VPWR Y
X0 a_923_74# B a_554_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_923_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y A a_923_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# C a_554_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y A a_923_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_923_74# B a_554_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_74# C a_554_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_554_74# C a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_554_74# B a_923_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND D a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND D a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_554_74# C a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_554_74# B a_923_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_923_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
X0 a_27_112# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 a_27_112# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_263_74# C a_341_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND D a_263_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_341_74# B a_443_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_443_74# a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
X0 a_490_74# C a_719_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND D a_719_123# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y a_27_74# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_490_74# B a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_225_74# B a_490_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR a_27_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_719_123# C a_490_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_225_74# a_27_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_719_123# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
X0 VPWR A_N a_27_158# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR a_27_158# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y a_27_158# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_225_74# B a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y a_27_158# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_656_74# B a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_656_74# C a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_1025_158# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_656_74# B a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_656_74# C a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_1025_158# C a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_1025_158# C a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND D a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_158# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Y a_27_158# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND D a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_1025_158# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_225_74# a_27_158# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_27_158# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_225_74# a_27_158# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_225_74# B a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_27_398# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_398# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR B_N a_226_398# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_435_74# a_226_398# a_513_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_226_398# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_627_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND B_N a_226_398# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_513_74# C a_627_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y a_27_398# a_435_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_398# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 a_27_368# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_27_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_678_74# C a_886_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y a_27_368# a_373_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_678_74# a_231_74# a_373_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_373_74# a_27_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_231_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND B_N a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_27_368# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VGND D a_886_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_886_74# C a_678_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_373_74# a_231_74# a_678_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR B_N a_231_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_886_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Y a_231_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 a_1229_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y a_232_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y a_27_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y a_27_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_374_74# a_27_114# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_27_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_1229_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_828_74# a_232_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_27_114# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_374_74# a_27_114# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR a_232_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND B_N a_232_114# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Y a_27_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_1229_74# C a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_374_74# a_232_114# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_27_114# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_232_114# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 VPWR a_232_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_1229_74# C a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_828_74# a_232_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_828_74# C a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 Y a_27_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 Y a_232_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_828_74# C a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VPWR A_N a_27_114# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X32 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 VPWR a_27_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 VGND D a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 VGND D a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_374_74# a_232_114# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 VPWR B_N a_232_114# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_116_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2_2 A B VGND VNB VPB VPWR Y
X0 a_35_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_35_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B a_35_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A a_35_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2_8 A B VGND VNB VPB VPWR Y
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2b_1 A B_N VGND VNB VPB VPWR Y
X0 a_278_368# a_27_112# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_112# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_27_112# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 VPWR A a_278_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y a_27_112# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2b_2 A B_N VGND VNB VPB VPWR Y
X0 a_228_368# a_27_392# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_392# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_228_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_392# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 Y a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND a_27_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y a_27_392# a_228_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR A a_228_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor2b_4 A B_N VGND VNB VPB VPWR Y
X0 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_353_323# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 Y a_353_323# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y a_353_323# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y a_353_323# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND B_N a_353_323# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR B_N a_353_323# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_116_368# a_353_323# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_116_368# a_353_323# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VGND a_353_323# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_114_368# B a_198_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_198_368# C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor3_2 A B C VGND VNB VPB VPWR Y
X0 a_27_368# C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_306_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A a_306_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_306_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_368# B a_306_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor3_4 A B C VGND VNB VPB VPWR Y
X0 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_295_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_368# B a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y C a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_295_368# C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y C a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_368# B a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_295_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_295_368# C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 a_27_112# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 VPWR A a_260_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_260_368# B a_344_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_344_368# a_27_112# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_112# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor3b_2 A B C_N VGND VNB VPB VPWR Y
X0 Y a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND a_27_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y a_27_392# a_227_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_495_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_495_368# B a_227_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_392# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_227_368# a_27_392# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR A a_495_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_227_368# B a_495_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_27_392# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor3b_4 A B C_N VGND VNB VPB VPWR Y
X0 Y a_468_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_126_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND a_468_264# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_468_264# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR C_N a_468_264# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_27_368# a_468_264# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_368# a_468_264# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_126_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y a_468_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND C_N a_468_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR A a_126_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_126_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_27_368# B a_126_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_468_264# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 Y a_468_264# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Y a_468_264# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_27_368# B a_126_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR A a_126_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_126_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_144_368# B a_228_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_228_368# C a_342_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_342_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A a_144_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4_2 A B C D VGND VNB VPB VPWR Y
X0 a_27_368# C a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_116_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND D Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y D a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_490_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_490_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_368# B a_490_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_116_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR A a_490_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4_4 A B C D VGND VNB VPB VPWR Y
X0 Y D a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_496_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND D Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_879_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_496_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_496_368# B a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_879_368# B a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y D a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_496_368# B a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_368# C a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_27_368# C a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_27_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_879_368# B a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_879_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Y D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_27_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
X0 a_344_368# C a_446_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A a_260_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_260_368# B a_344_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_57_368# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_57_368# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 a_446_368# a_57_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y a_57_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
X0 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_27_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_229_368# a_27_392# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR A a_701_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_229_368# C a_498_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_392# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_701_368# B a_498_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_701_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y a_27_392# a_229_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_498_368# C a_229_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_392# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_498_368# B a_701_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Y a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y a_47_88# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y a_47_88# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y a_47_88# a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_778_368# B a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_1191_368# B a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR A a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR A a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_47_88# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 a_319_368# a_47_88# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_319_368# C a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_778_368# B a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_319_368# C a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND a_47_88# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_319_368# a_47_88# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_778_368# C a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_778_368# C a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_1191_368# B a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_1191_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_47_88# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VPWR D_N a_47_88# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X31 a_1191_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 VGND a_47_88# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 Y a_47_88# a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
X0 a_27_112# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_530_368# a_611_244# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR A a_313_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_313_368# B a_397_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR D_N a_611_244# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND D_N a_611_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y a_611_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_397_368# a_27_112# a_530_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_112# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
X0 VGND D_N a_311_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND a_27_392# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_392# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VPWR D_N a_311_124# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_985_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_392# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y a_311_124# a_493_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_985_368# B a_772_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_493_368# a_27_392# a_772_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR A a_985_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Y a_311_124# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_772_368# a_27_392# a_493_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_311_124# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_493_368# a_311_124# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_772_368# B a_985_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
X0 a_27_368# B a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_897_349# a_864_48# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND a_864_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y a_1162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_864_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_116_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_897_349# a_1162_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_368# a_864_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_116_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_1162_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND D_N a_1162_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 Y a_1162_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_864_48# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VGND a_1162_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_27_368# a_864_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VGND C_N a_864_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_897_349# a_864_48# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 Y a_1162_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 Y a_1162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VPWR D_N a_1162_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X30 a_1162_48# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X31 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 Y a_864_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 a_27_368# B a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_897_349# a_1162_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X36 VPWR C_N a_864_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X37 Y a_864_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_83_260# B2 a_693_384# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_83_260# a_233_384# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VPWR A1_N a_233_384# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_693_384# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_233_384# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR a_233_384# a_83_260# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_588_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_253_94# A2_N a_233_384# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND A1_N a_253_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VGND B1 a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_27_74# a_270_48# a_201_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A2_N a_270_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 VPWR B1 a_117_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_500_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_270_48# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 X a_201_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_270_48# A2_N a_500_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_201_392# a_270_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 X a_201_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_117_392# B2 a_201_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_27_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND a_201_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR a_201_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_476_48# A2_N a_835_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND a_310_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_310_392# a_476_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_310_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR a_476_48# a_310_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 X a_310_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 X a_310_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 X a_310_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_41_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VPWR a_310_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR B1 a_41_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_310_392# B2 a_41_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VPWR a_310_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A2_N a_476_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_476_48# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_835_94# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_310_392# a_476_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_27_74# a_476_48# a_310_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 X a_310_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_27_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_41_392# B2 a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_131_383# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_490_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR a_131_383# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_397_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y B2 a_490_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y a_131_383# a_397_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND B1 a_397_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A1_N a_131_383# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VGND A1_N a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_114_74# A2_N a_131_383# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR a_133_387# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_518_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND B2 a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR B1 a_796_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y B2 a_796_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_134_74# A2_N a_133_387# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 VGND B1 a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_796_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A1_N a_134_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_518_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A1_N a_133_387# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_133_387# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_518_74# a_133_387# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_796_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VPWR A2_N a_133_387# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_134_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_133_387# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 Y a_133_387# a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 Y a_133_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_133_387# A2_N a_134_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_114_368# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_857_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_857_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR B1 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_114_368# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y a_114_368# a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND A1_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_114_368# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_857_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_114_368# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y a_114_368# a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_1215_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND A1_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_114_368# A2_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_1215_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR A1_N a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR a_114_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_27_74# A2_N a_114_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_1215_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Y a_114_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_1215_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VPWR A1_N a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_857_74# a_114_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VPWR A2_N a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR A2_N a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_27_74# A2_N a_114_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VGND B2 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VPWR a_114_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 Y B2 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VGND B2 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_114_368# A2_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 Y a_114_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_857_74# a_114_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 Y B2 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 a_27_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 VGND B1 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 VGND B1 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 VPWR B1 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 a_27_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 a_857_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 X a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR B1 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_320_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_83_244# A2 a_376_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_83_244# B1 a_320_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VGND A1 a_320_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_376_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_160_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 X a_244_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_160_368# A2 a_244_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_244_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_244_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_54_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_54_74# B1 a_244_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_244_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_244_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND A2 a_54_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_116_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_116_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND a_216_387# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VPWR a_216_387# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_116_387# A2 a_216_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR B1 a_216_387# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 X a_216_387# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_216_387# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND A1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VGND a_216_387# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR a_216_387# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_216_387# B1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_27_125# B1 a_216_387# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_27_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 X a_216_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 X a_216_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_216_387# A2 a_116_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 VGND A2 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_216_387# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A1 a_162_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_162_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_116_392# A2 a_200_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_200_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# a_281_244# a_200_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_200_392# a_281_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR A1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND a_200_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_281_244# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_281_244# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_27_74# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND A1 a_487_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR a_177_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_74# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VPWR a_27_74# a_177_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND a_177_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 X a_177_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_177_48# a_27_74# a_487_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_177_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_582_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_487_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_177_48# A2 a_582_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_27_368# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_193_48# a_27_368# a_618_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VPWR a_193_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_892_392# A2 a_193_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_193_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_193_48# A2 a_892_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR a_27_368# a_193_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 VPWR A1 a_892_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 X a_193_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_368# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 X a_193_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_618_94# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_892_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_618_94# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_618_94# a_27_368# a_193_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VGND a_193_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_193_48# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 VGND A1 a_618_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 VGND a_193_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 X a_193_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND A2 a_618_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VPWR a_193_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VPWR a_27_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_74# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 VGND A1 a_308_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_308_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_395_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y A2 a_395_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_74# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 Y a_27_74# a_308_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VPWR A1 a_507_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_225_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y A2 a_507_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR a_27_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_27_74# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_225_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_507_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_507_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y a_27_74# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_225_74# a_27_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND A2 a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_27_74# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VGND A1 a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VPWR B1_N a_828_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_28_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y a_828_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_28_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_828_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_74# a_828_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_828_48# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 Y a_828_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_828_48# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 Y a_828_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_27_74# a_828_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_398_392# B2 a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND A1 a_299_139# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VPWR B1 a_398_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_83_260# A2 a_572_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_572_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_299_139# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_83_260# B2 a_299_139# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_299_139# B1 a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_82_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 X a_82_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 X a_82_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_82_48# A2 a_575_384# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND a_82_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_383_384# B2 a_82_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_575_384# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_307_74# B1 a_82_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND A1 a_307_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_307_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR B1 a_383_384# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_82_48# B2 a_307_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_206_392# B2 a_516_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 X a_206_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_206_392# A2 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND A1 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_27_136# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_516_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_206_392# B2 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VPWR B1 a_516_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND A2 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 VGND a_206_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_116_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_206_392# B1 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_27_136# B2 a_206_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_27_136# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 X a_206_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR a_206_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 X a_206_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 X a_206_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR a_206_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_516_392# B2 a_206_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VGND a_206_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_136# B1 a_206_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_116_392# A2 a_206_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y A2 a_340_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_340_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR B1 a_142_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_142_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR B1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y B2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_510_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_510_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_28_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y A2 a_510_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_28_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR A1 a_510_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_117_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_877_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_117_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y B2 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y A2 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_117_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_877_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Y A2 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y B2 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VPWR B1 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VPWR A1 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_877_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR A1 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_877_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR B1 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_117_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_230_94# B1 a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VGND A1 a_230_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VGND A3 a_230_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_256_368# A2 a_340_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_84_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VPWR A1 a_256_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 X a_84_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_230_94# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 X a_84_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_340_368# A3 a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_55_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_346_392# A2 a_430_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND A1 a_328_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 X a_55_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_430_392# A3 a_55_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR A1 a_346_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_55_264# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_55_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_55_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND A3 a_328_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_328_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_328_74# B1 a_55_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_492_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_86_260# A3 a_699_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND A3 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_86_260# B1 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_492_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_492_125# B1 a_86_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 VGND A2 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_86_260# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_968_392# A2 a_699_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_699_392# A3 a_86_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_699_392# A2 a_968_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_968_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 a_492_125# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VPWR A1 a_968_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 VPWR B1 a_86_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VGND A1 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_119_368# A2 a_203_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_114_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_114_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_203_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR A1 a_119_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND A3 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A1 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y A3 a_297_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_297_368# A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_297_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_28_368# A2 a_297_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_487_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_82# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A2 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_487_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_82# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_82# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A3 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_82# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_28_368# A2 a_487_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A3 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_487_368# A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_82# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND A2 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_82# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 Y B1 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Y B1 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 Y A3 a_487_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_28_368# A2 a_487_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_27_82# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VGND A1 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VGND A1 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_27_82# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_487_368# A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 Y A3 a_487_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_83_264# B2 a_548_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_248_368# A2 a_332_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND A3 a_251_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_332_368# A3 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR A1 a_248_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_251_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VGND A1 a_251_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_548_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_251_74# B2 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_83_264# B1 a_251_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_83_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A1 a_346_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_83_264# B2 a_652_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_83_264# B1 a_349_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_652_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VGND A1 a_349_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_430_368# A3 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_349_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_349_74# B2 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_346_368# A2 a_430_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VGND a_83_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND A3 a_349_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_83_256# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_83_256# B2 a_534_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_1234_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND A1 a_564_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_83_256# B2 a_564_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VGND A3 a_564_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_961_392# A3 a_83_256# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND a_83_256# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_83_256# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_564_74# B2 a_83_256# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_1234_392# A2 a_961_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_961_392# A2 a_1234_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 X a_83_256# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_534_388# B2 a_83_256# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_564_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 X a_83_256# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR B1 a_534_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_534_388# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_83_256# B1 a_564_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 VGND A2 a_564_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 VGND a_83_256# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_564_74# B1 a_83_256# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_83_256# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR A1 a_1234_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X24 a_564_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 a_564_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 X a_83_256# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_83_256# A3 a_961_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_128_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR B1 a_128_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_456_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y A3 a_342_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_342_368# A2 a_456_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR A1 a_768_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 Y A3 a_499_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_768_368# A2 a_499_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_768_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_499_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_499_368# A2 a_768_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A1 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_1330_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_861_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_861_368# A2 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y A3 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_1330_368# A2 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_861_368# A2 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_1330_368# A2 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_861_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 Y A3 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 VPWR A1 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 a_1330_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 X a_83_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A3 a_326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VPWR B1 a_83_270# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_326_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_83_270# B1 a_326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_443_368# A3 a_527_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_527_368# A2 a_641_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_641_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_326_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_83_270# A4 a_443_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VGND A1 a_326_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 X a_83_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_314_368# A4 a_428_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# B1 a_428_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_428_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_428_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND A4 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_428_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_116_368# A2 a_200_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_200_368# A3 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR a_428_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND a_428_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_851_368# A3 a_762_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR a_110_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR B1 a_110_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_1213_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VPWR a_110_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A3 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_851_368# A4 a_110_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VGND a_110_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_523_124# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_523_124# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VGND A2 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VGND A1 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_762_368# A2 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_523_124# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 X a_110_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 X a_110_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 X a_110_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_110_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 X a_110_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR A1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_762_368# A3 a_851_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_523_124# B1 a_110_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_110_48# B1 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 VGND A4 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_523_124# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 a_1213_368# A2 a_762_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_110_48# A4 a_851_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND a_110_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_358_368# A2 a_472_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_157_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 Y B1 a_157_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_472_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_157_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y A4 a_260_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_260_368# A3 a_358_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A3 a_157_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND A1 a_157_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A1 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_132_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_132_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_314_368# A4 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_314_368# A3 a_607_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_607_368# A2 a_807_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Y B1 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_132_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_807_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A2 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y A4 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_607_368# A3 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_807_368# A2 a_607_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_132_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND A4 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND A3 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_132_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR A1 a_807_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_339_368# A4 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_788_368# A3 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_339_368# A4 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_339_368# A3 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_1191_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_1191_368# A2 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_1191_368# A2 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VPWR A1 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_1191_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VGND A4 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 Y A4 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_339_368# A3 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 Y A4 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR A1 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_788_368# A3 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_27_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VGND A4 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_788_368# A2 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_27_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_788_368# A2 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_398_392# A2 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_257_136# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_662_136# C1 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VPWR A1 a_398_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_257_136# B1 a_662_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_83_264# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VGND A2 a_257_136# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR C1 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_195_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 X a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND a_27_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_27_368# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_117_74# B1 a_195_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_368# C1 a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A1 a_195_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_314_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VPWR a_27_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_27_368# A2 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR C1 a_91_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VPWR A1 a_968_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND a_91_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_91_48# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VPWR a_91_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_968_391# A2 a_91_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 X a_91_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_510_125# B1 a_597_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 X a_91_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 X a_91_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND a_91_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_510_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_91_48# A2 a_968_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_91_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 a_91_48# C1 a_597_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 VPWR B1 a_91_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_597_125# C1 a_91_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 VGND A2 a_510_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 VPWR a_91_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 X a_91_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_510_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_597_125# B1 a_510_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_968_391# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VGND A1 a_510_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_311_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A2 a_31_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_31_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_31_74# B1 a_311_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_303_84# B1 a_30_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_505_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_505_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_30_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_30_84# B1 a_303_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_303_84# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR A1 a_505_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y C1 a_30_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y A2 a_505_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_303_84# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VGND A2 a_303_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND A1 a_303_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A1 a_30_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A1 a_30_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_834_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_30_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_30_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_30_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_30_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y A2 a_30_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_27_74# B1 a_834_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y C1 a_834_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_834_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_834_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_27_74# B1 a_834_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 Y C1 a_834_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_834_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 Y A2 a_30_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_245_94# B1 a_456_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_245_94# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND A1 a_245_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_83_264# B2 a_462_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_462_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VPWR C1 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR A1 a_264_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_456_74# B2 a_245_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_456_74# C1 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_264_392# A2 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_27_368# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_530_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR B1 a_332_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_27_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_165_74# B1 a_264_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_368# C1 a_165_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_264_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_332_368# B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VGND A2 a_264_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_27_368# A2 a_530_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VPWR a_27_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_264_74# B2 a_165_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR C1 a_114_125# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_300_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_27_125# B1 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_300_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VPWR a_114_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 X a_114_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_125# B2 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_763_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR a_114_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_297_387# B2 a_114_125# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_763_387# A2 a_114_125# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND A2 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 VGND a_114_125# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_297_387# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_114_125# A2 a_763_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 X a_114_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_300_125# B1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_114_125# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_300_125# B2 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 X a_114_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_27_125# C1 a_114_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 X a_114_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VPWR A1 a_763_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VGND A1 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 VGND a_114_125# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_114_125# C1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 a_114_125# B2 a_297_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 VPWR B1 a_297_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_114_74# B2 a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_239_74# B1 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y A2 a_522_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 VGND A1 a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR B1 a_324_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_324_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_239_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y C1 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_522_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_376_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR B1 a_376_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_776_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_311_85# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Y C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_311_85# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# B1 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_74# B2 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_311_85# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND A2 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y A2 a_776_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_311_85# B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_776_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 Y B2 a_376_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_376_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR A1 a_776_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_27_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND A1 a_311_85# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND A2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y C1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_84# B1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_483_74# B1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_483_74# B2 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_483_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR B1 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_483_74# B1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 Y A2 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 Y B2 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 Y A2 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_27_84# B2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_508_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR A1 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_1288_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 Y B2 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_483_74# B2 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_483_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_483_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR A1 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_1288_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_27_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_508_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR B1 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_1288_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_508_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_508_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 Y C1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 VGND A1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 VGND A1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_1288_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 a_27_84# B2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_27_84# B1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 a_483_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_131_74# B1 a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_209_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_209_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND A3 a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VPWR B1 a_31_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR a_31_387# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_31_387# A3 a_320_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_536_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND a_31_387# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_320_387# A2 a_536_387# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_31_387# C1 a_131_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_31_387# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_135_74# B1 a_219_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_219_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND a_32_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR B1 a_32_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_219_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_32_74# C1 a_135_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND A2 a_219_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_32_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR a_32_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_32_74# A3 a_360_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_32_74# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_360_368# A2 a_444_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_444_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 X a_32_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_83_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_651_78# B1 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 X a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND a_83_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR A1 a_1338_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND A3 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_564_78# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_564_78# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_83_244# C1 a_651_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 VGND A1 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR B1 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND a_83_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR C1 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_83_244# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 a_83_244# A3 a_1034_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 a_651_78# C1 a_83_244# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 X a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_1338_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 VGND A2 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_83_244# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 X a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_564_78# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_1034_392# A3 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X23 VPWR a_83_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_1034_392# A2 a_1338_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 X a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_1338_392# A2 a_1034_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_564_78# B1 a_651_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_469_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_128_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_128_74# B1 a_469_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_222_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 VGND A3 a_128_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A1 a_128_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VPWR A1 a_138_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_138_368# A2 a_222_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y C1 a_670_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_307_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_670_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_670_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_28_368# A2 a_307_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_307_368# A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y A3 a_307_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_74# B1 a_670_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR A1 a_1350_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_27_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_1350_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_1350_368# A2 a_841_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 Y C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A1 a_1350_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_74# B1 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_459_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Y C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND A3 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_459_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_459_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_459_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 VGND A2 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_841_368# A2 a_1350_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 Y A3 a_841_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_459_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_459_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_841_368# A2 a_1350_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_27_74# B1 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_459_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_1350_368# A2 a_841_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_1350_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_841_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 VGND A1 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VGND A1 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 VGND A2 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VGND A3 a_459_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 Y A3 a_841_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_27_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_841_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 a_459_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 X a_82_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VPWR D1 a_82_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 X a_82_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_393_74# B1 a_471_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_82_48# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_321_74# C1 a_393_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_82_48# A2 a_600_381# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VPWR B1 a_82_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_471_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_600_381# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VGND A1 a_471_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_82_48# D1 a_321_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR A1 a_152_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_236_368# D1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_152_368# A2 a_236_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_236_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_369_74# C1 a_461_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR a_236_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_54_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_54_74# B1 a_369_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_461_74# D1 a_236_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND A2 a_54_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 X a_236_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_236_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 VPWR C1 a_236_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VGND a_236_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_27_392# A2 a_747_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_27_74# C1 a_287_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_747_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VPWR C1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VPWR a_27_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_27_392# D1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_27_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_747_392# A2 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_287_74# C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_287_74# B1 a_477_198# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_477_198# B1 a_287_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VPWR D1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 a_27_392# D1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 X a_27_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VPWR B1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 X a_27_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR A1 a_747_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_477_198# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VGND A1 a_477_198# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND a_27_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VGND A2 a_477_198# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 X a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_477_198# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_27_74# D1 a_27_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_27_392# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 VPWR a_27_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_27_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_490_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND A1 a_368_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_368_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_260_74# B1 a_368_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Y A2 a_490_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_182_74# C1 a_260_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y D1 a_182_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_510_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 Y A2 a_697_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VGND A2 a_510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_299_74# B1 a_510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND A1 a_510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR A1 a_697_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_510_74# B1 a_299_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_510_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_697_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_299_74# C1 a_40_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_697_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_40_74# D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_40_74# C1 a_299_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 Y D1 a_40_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_27_74# D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND A1 a_841_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_472_74# C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VPWR A1 a_954_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_74# C1 a_472_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A1 a_841_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND A2 a_841_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_954_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_954_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VPWR A1 a_954_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_841_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_841_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_27_74# C1 a_472_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 Y A2 a_954_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_841_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_472_74# B1 a_841_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_472_74# C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_841_74# B1 a_472_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_954_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_954_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_841_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_841_74# B1 a_472_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 Y D1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 Y D1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VGND A2 a_841_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_27_74# D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_472_74# B1 a_841_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X32 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 Y A2 a_954_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X
X0 a_63_368# B a_152_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND B a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 a_152_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_63_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VPWR a_63_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND a_63_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or2_2 A B VGND VNB VPB VPWR X
X0 VGND a_27_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_27_368# B a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND B a_27_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_114_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 X a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_27_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__or2_4 A B VGND VNB VPB VPWR X
X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_493_388# B a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_83_260# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VPWR A a_493_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_83_260# B a_493_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_493_388# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_27_112# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 a_264_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 VGND a_264_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_264_368# a_27_112# a_353_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_353_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR a_264_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_112# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 VGND a_27_112# a_264_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__or2b_2 A B_N VGND VNB VPB VPWR X
X0 a_27_368# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 VGND A a_187_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VPWR A a_470_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_187_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_470_368# a_27_368# a_187_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_187_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_187_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_27_368# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 X a_187_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_187_48# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__or2b_4 A B_N VGND VNB VPB VPWR X
X0 X a_81_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND a_81_296# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_81_296# a_676_48# a_489_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_81_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_489_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 X a_81_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_676_48# a_81_296# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VPWR B_N a_676_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND B_N a_676_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 VPWR a_81_296# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_489_392# a_676_48# a_81_296# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VPWR a_81_296# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_81_296# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_81_296# a_676_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 X a_81_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR A a_489_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 VGND A a_81_296# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 VGND a_81_296# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or3_1 A B C VGND VNB VPB VPWR X
X0 a_27_74# C a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 a_116_368# B a_200_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 a_200_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_27_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__or3_2 A B C VGND VNB VPB VPWR X
X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_27_74# C a_150_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_150_392# B a_234_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_234_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__or3_4 A B C VGND VNB VPB VPWR X
X0 X a_302_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 a_206_388# C a_302_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_116_388# B a_206_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND B a_302_388# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_302_388# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 X a_302_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 X a_302_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A a_116_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_302_388# C a_206_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_206_388# B a_116_388# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_302_388# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 X a_302_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND a_302_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR a_302_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_116_388# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VPWR a_302_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_302_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 VGND B a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 a_239_74# a_124_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 a_368_391# B a_452_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_239_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_452_391# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_239_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 VGND C_N a_124_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 a_239_74# a_124_424# a_368_391# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR C_N a_124_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VPWR a_239_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__or3b_2 A B C_N VGND VNB VPB VPWR X
X0 a_27_368# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 X a_190_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_458_368# B a_542_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 X a_190_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_190_260# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_542_368# a_27_368# a_190_260# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR a_190_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR A a_458_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_27_368# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X9 VGND A a_190_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VGND a_27_368# a_190_260# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VGND a_190_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or3b_4 A B C_N VGND VNB VPB VPWR X
X0 X a_409_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 VGND a_409_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VGND a_409_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_217_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 X a_409_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 X a_409_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_27_392# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VPWR A a_217_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VGND B a_409_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_307_392# B a_217_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_27_392# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_409_392# a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_409_392# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 X a_409_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_307_392# a_27_392# a_409_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VPWR a_409_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VPWR a_409_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_217_392# B a_307_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_409_392# a_27_392# a_307_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4_1 A B C D VGND VNB VPB VPWR X
X0 VGND a_44_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND B a_44_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X2 a_133_392# C a_217_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_44_392# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 VGND D a_44_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 a_217_392# B a_331_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR a_44_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_44_392# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X8 a_331_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_44_392# D a_133_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_258_392# B a_342_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 X a_85_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_85_392# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND a_85_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_85_392# D a_174_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_174_392# C a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 X a_85_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND D a_85_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR a_85_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND B a_85_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 a_342_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_85_392# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4_4 A B C D VGND VNB VPB VPWR X
X0 VPWR a_83_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_83_264# D a_962_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VGND C a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND B a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_499_392# B a_588_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR A a_588_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_83_264# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_83_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_83_264# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_962_392# D a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VGND a_83_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_588_392# B a_499_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_962_392# C a_499_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VGND a_83_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_588_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 a_499_392# C a_962_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 a_440_368# B a_524_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_228_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VGND B a_228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 VGND a_27_74# a_228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 a_356_368# C a_440_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_228_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 VGND a_228_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_27_74# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_228_74# a_27_74# a_356_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_524_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_228_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X11 a_27_74# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4b_2 A B C D_N VGND VNB VPB VPWR X
X0 a_27_368# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 X a_190_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_452_392# B a_536_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_190_48# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 VGND C a_190_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_638_392# a_27_368# a_190_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 X a_190_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_190_48# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VGND a_190_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_190_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_368# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X11 VGND A a_190_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_536_392# C a_638_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VPWR A a_452_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_563_48# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_496_392# a_563_48# a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_496_392# C a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_27_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_27_392# B a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 VPWR A a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_27_74# a_563_48# a_496_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_116_392# B a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_27_392# C a_496_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_563_48# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 VGND a_563_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_116_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 a_357_378# a_27_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X1 VPWR D_N a_216_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_357_378# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 VGND D_N a_216_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 a_626_378# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_27_424# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 VGND B a_357_378# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 a_530_378# B a_626_378# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_446_378# a_27_424# a_530_378# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 VPWR a_357_378# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_27_424# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 VGND a_216_424# a_357_378# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X12 a_357_378# a_216_424# a_446_378# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 VGND a_357_378# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
X0 X a_182_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_587_392# B a_689_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_182_270# a_27_424# a_503_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_27_424# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VGND B a_182_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_503_392# a_548_110# a_587_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 a_182_270# a_548_110# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 a_689_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 VPWR a_182_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_182_270# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X10 VPWR C_N a_548_110# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 VGND a_182_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 VGND C_N a_548_110# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X13 VGND a_27_424# a_182_270# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_27_424# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 X a_182_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
X0 a_27_94# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_1060_392# a_678_368# a_791_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_1273_392# B a_1060_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_1273_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 VGND a_193_277# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_791_392# a_27_94# a_193_277# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 VPWR C_N a_678_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_27_94# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 VPWR A a_1273_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 X a_193_277# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 X a_193_277# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 X a_193_277# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR a_193_277# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_1060_392# B a_1273_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VGND C_N a_678_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_193_277# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_193_277# a_27_94# a_791_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 X a_193_277# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_791_392# a_678_368# a_1060_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VGND a_193_277# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_193_277# a_678_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VGND B a_193_277# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VPWR a_193_277# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VGND a_27_94# a_193_277# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 a_662_82# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1159_497# a_867_82# a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_977_243# a_1579_258# a_1434_78# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 a_2133_410# a_1954_119# a_2392_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_1579_258# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_1151_119# a_662_82# a_1159_497# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 VPWR a_977_243# a_1081_497# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X7 VPWR a_977_243# a_1903_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VGND a_3078_384# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_1954_119# a_662_82# a_2088_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 a_1434_78# a_1159_497# a_977_243# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X11 a_2509_392# a_1954_119# a_2133_410# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X12 a_1159_497# a_662_82# a_197_119# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X13 VPWR a_2133_410# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 VGND a_2133_410# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_1528_424# a_1579_258# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_1903_424# a_867_82# a_1954_119# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_2088_508# a_2133_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_197_119# a_353_93# a_27_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X19 a_305_119# a_353_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_662_82# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VGND SCD a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 VGND SCE a_353_93# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_2164_119# a_2133_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 VPWR a_662_82# a_867_82# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_1876_119# a_662_82# a_1954_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X26 VGND a_977_243# a_1151_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VPWR a_1579_258# a_2509_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X28 VGND a_662_82# a_867_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VPWR a_3078_384# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_1954_119# a_867_82# a_2164_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_3078_384# a_2133_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X32 a_977_243# a_1159_497# a_1528_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X33 VPWR SCE a_353_93# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X34 a_3078_384# a_2133_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X35 a_2392_74# a_1579_258# a_2133_410# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_2133_410# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X37 a_1579_258# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X38 a_27_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X39 a_1081_497# a_867_82# a_1159_497# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X40 VGND SET_B a_2392_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X41 VPWR SCE a_212_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X42 a_1434_78# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X43 a_197_119# D a_305_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X44 VPWR SET_B a_977_243# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X45 a_212_464# D a_197_119# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X46 VGND a_977_243# a_1876_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X47 a_119_119# SCE a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 VPWR a_688_98# a_868_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1007_366# a_1154_464# a_1592_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_1997_82# a_688_98# a_2171_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_1154_464# a_868_368# a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 Q a_3272_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_1070_464# a_868_368# a_1154_464# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 a_1643_257# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X7 a_1592_424# a_1643_257# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_2216_410# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X9 a_3272_94# a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_197_119# a_341_410# a_27_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 a_1473_73# a_1154_464# a_1007_366# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X12 a_1997_82# a_868_368# a_2247_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VPWR SCE a_341_410# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 a_1473_73# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X15 a_3272_94# a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 VGND SCE a_341_410# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 VGND a_688_98# a_868_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VGND SET_B a_2452_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 VPWR SCE a_206_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X20 VPWR SET_B a_1007_366# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 VPWR a_3272_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR a_1007_366# a_1986_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X23 a_1986_424# a_868_368# a_1997_82# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X24 a_1007_366# a_1643_257# a_1473_73# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X25 VPWR a_2216_410# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_688_98# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND SCD a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 a_363_119# a_341_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 VGND a_1007_366# a_1185_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X30 a_1185_125# a_688_98# a_1154_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 VGND a_1007_366# a_1902_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X32 a_1154_464# a_688_98# a_197_119# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X33 Q_N a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_1902_125# a_688_98# a_1997_82# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X35 a_2556_392# a_1997_82# a_2216_410# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X36 a_2452_74# a_1643_257# a_2216_410# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 a_206_464# D a_197_119# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X38 a_688_98# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X39 VGND a_2216_410# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 a_2171_508# a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X41 a_27_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X42 VGND a_3272_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X43 a_2247_82# a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X44 a_1643_257# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X45 a_2216_410# a_1997_82# a_2452_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X46 a_197_119# D a_363_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X47 Q a_3272_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X48 VPWR a_1007_366# a_1070_464# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X49 a_119_119# SCE a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X50 VPWR a_1643_257# a_2556_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X51 Q_N a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q
+ Q_N
X0 a_1092_96# a_877_98# a_1192_96# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_1625_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X2 a_2037_442# a_1625_93# a_2271_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_1092_96# a_622_98# a_1221_419# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 VPWR SET_B a_2037_442# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_2881_74# a_2037_442# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND SET_B a_2271_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR a_1250_231# a_1766_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_1986_504# a_2037_442# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 a_1221_419# a_1250_231# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X10 a_1250_231# a_1092_96# a_1580_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_197_119# a_877_98# a_1092_96# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X12 VGND a_622_98# a_877_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_2384_392# a_1625_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VPWR a_2037_442# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_622_98# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_2061_74# a_2037_442# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_1580_379# a_1625_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_1766_379# a_622_98# a_1878_420# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 a_197_119# a_622_98# a_1092_96# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_1625_93# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_197_119# D a_299_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 a_218_464# D a_197_119# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X23 VGND SET_B a_1418_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X24 VGND a_2881_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VGND a_1250_231# a_1880_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X26 a_1880_119# a_877_98# a_1878_420# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X27 a_1878_420# a_622_98# a_2061_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 VGND SCD a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_622_98# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_2881_74# a_2037_442# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X31 a_299_119# a_341_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_1418_125# a_1092_96# a_1250_231# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X33 a_1878_420# a_877_98# a_1986_504# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X34 VPWR SCE a_218_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X35 VPWR a_622_98# a_877_98# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X36 a_27_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X37 VGND a_2037_442# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_1192_96# a_1250_231# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 VPWR a_2881_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X40 VPWR SET_B a_1250_231# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X41 a_197_119# a_341_93# a_27_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X42 VGND SCE a_341_93# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X43 a_1250_231# a_1625_93# a_1418_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X44 VPWR SCE a_341_93# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X45 a_2037_442# a_1878_420# a_2384_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X46 a_119_119# SCE a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X47 a_2271_74# a_1878_420# a_2037_442# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1328_463# a_1369_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 VPWR a_1221_97# a_1369_71# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_413_90# a_850_74# a_1221_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 VGND a_1747_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_850_74# a_1023_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_850_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_413_90# SCE a_545_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VPWR RESET_B a_2008_48# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 VGND a_2513_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_225_90# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VPWR RESET_B a_413_90# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 a_1747_74# a_1023_74# a_1969_489# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 VGND RESET_B a_2124_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_1969_489# a_2008_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_1399_97# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_1966_74# a_2008_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_413_90# a_27_74# a_512_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 a_1321_97# a_1369_71# a_1399_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X19 a_312_90# D a_413_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_2513_424# a_1747_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 VPWR RESET_B a_1221_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_1747_74# a_850_74# a_1966_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_1369_71# a_850_74# a_1747_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X24 a_512_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X25 a_850_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_413_90# a_1023_74# a_1221_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X27 a_2008_48# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 VPWR a_1747_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VPWR SCE a_338_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X30 a_1221_97# a_850_74# a_1328_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X31 a_2513_424# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X32 a_2124_74# a_1747_74# a_2008_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_1369_71# a_1023_74# a_1747_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X34 VPWR a_850_74# a_1023_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X35 a_545_97# SCD a_225_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 a_1221_97# a_1023_74# a_1321_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 VGND a_1221_97# a_1369_71# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X38 a_225_90# a_27_74# a_312_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 a_338_464# D a_413_90# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X40 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X41 VPWR a_2513_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_27_79# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_2158_74# a_1790_74# a_2006_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_2604_392# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_1323_118# a_1370_289# a_1401_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_307_464# D a_388_79# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X5 a_223_79# a_27_79# a_310_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_388_79# a_27_79# a_538_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X7 a_388_79# SCE a_547_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 VPWR a_2604_392# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_223_79# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VPWR a_1223_118# a_1370_289# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 a_388_79# a_852_74# a_1223_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 VGND RESET_B a_2158_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VGND a_1790_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Q a_2604_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VGND a_1790_74# a_2604_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_538_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 Q_N a_1790_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_1401_118# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 a_2000_74# a_2006_373# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 VPWR SCE a_307_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X21 a_2006_373# a_1790_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 a_388_79# a_1025_74# a_1223_118# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 a_1223_118# a_1025_74# a_1323_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_1223_118# a_852_74# a_1325_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 a_1790_74# a_852_74# a_2000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_852_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND a_1223_118# a_1370_289# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 a_310_79# D a_388_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 VPWR a_1790_74# a_2604_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X30 Q a_2604_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 VPWR a_852_74# a_1025_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_1325_457# a_1370_289# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X33 a_1955_471# a_2006_373# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X34 a_27_79# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X35 a_1370_289# a_852_74# a_1790_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X36 VPWR a_1790_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X37 a_547_79# SCD a_223_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 VPWR RESET_B a_1223_118# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X39 VGND a_852_74# a_1025_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 a_1790_74# a_1025_74# a_1955_471# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X41 a_852_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X42 VPWR RESET_B a_2006_373# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X43 Q_N a_1790_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X44 a_1370_289# a_1025_74# a_1790_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X45 VPWR RESET_B a_388_79# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_284_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 a_1429_308# a_1074_88# a_1827_144# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 a_2492_424# a_1827_144# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X3 VPWR a_854_74# a_1074_88# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_284_464# a_854_74# a_1272_131# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_324_81# D a_284_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_284_464# SCE a_538_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VGND a_1272_131# a_1429_308# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_284_464# a_1074_88# a_1272_131# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR a_1272_131# a_1429_308# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_2087_410# a_1827_144# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_1827_144# a_1074_88# a_2073_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 VPWR a_2492_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 VPWR SCE a_206_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 a_1489_131# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_2492_424# a_1827_144# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_2265_74# a_1827_144# a_2087_410# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 VGND a_2492_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 VPWR RESET_B a_1272_131# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_1272_131# a_854_74# a_1411_131# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 VGND RESET_B a_2265_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VPWR CLK_N a_854_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_1429_308# a_854_74# a_1827_144# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_1827_144# a_854_74# a_2042_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_2042_508# a_2087_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 a_206_464# D a_284_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X26 a_471_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X27 a_1272_131# a_1074_88# a_1384_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 VPWR RESET_B a_2087_410# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X29 a_27_88# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X30 a_239_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_1411_131# a_1429_308# a_1489_131# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_239_81# a_27_88# a_324_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_538_81# SCD a_239_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 VGND a_854_74# a_1074_88# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_27_88# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 VGND CLK_N a_854_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 a_1384_508# a_1429_308# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X38 a_2073_74# a_2087_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 a_284_464# a_27_88# a_471_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1233_118# a_1034_368# a_1319_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_1972_74# a_1997_272# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_225_81# a_27_88# a_312_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_1367_92# a_1034_368# a_1745_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR SCE a_216_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X6 a_855_368# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_1367_92# a_855_368# a_1745_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_1745_74# a_855_368# a_1972_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_300_464# a_27_88# a_538_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 VPWR a_1745_74# a_2399_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 VGND a_2399_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_1343_461# a_1367_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 VPWR RESET_B a_1997_272# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_1397_118# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_545_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_538_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 VGND a_1745_74# a_2399_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X18 a_300_464# a_855_368# a_1233_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 a_1233_118# a_855_368# a_1343_461# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X20 VGND a_855_368# a_1034_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR a_1233_118# a_1367_92# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_1319_118# a_1367_92# a_1397_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VGND RESET_B a_2135_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_300_464# SCE a_545_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_855_368# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X26 a_2135_74# a_1745_74# a_1997_272# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 a_300_464# a_1034_368# a_1233_118# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X28 a_1993_508# a_1997_272# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X29 a_216_464# D a_300_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X30 VPWR a_855_368# a_1034_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_1997_272# a_1745_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 a_27_88# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X33 a_1745_74# a_1034_368# a_1993_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X34 VGND a_1233_118# a_1367_92# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X35 VPWR RESET_B a_1233_118# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X36 a_27_88# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 VPWR a_2399_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 VPWR RESET_B a_300_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X39 a_312_81# D a_300_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1824_74# a_1034_368# a_2037_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_547_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_225_81# a_27_74# a_312_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_390_81# a_27_74# a_514_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 VPWR a_1242_457# a_1383_349# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 VPWR RESET_B a_2082_446# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VPWR a_1824_74# a_2492_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_1242_457# a_855_368# a_1332_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_1354_138# a_1383_349# a_1432_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_514_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 a_390_81# SCE a_547_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_1432_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 Q a_2492_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_390_81# a_855_368# a_1242_457# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 Q a_2492_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND a_2492_392# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR RESET_B a_1242_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_340_464# D a_390_81# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X19 a_1383_349# a_1034_368# a_1824_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_2078_74# a_2082_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_1824_74# a_855_368# a_2078_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 a_855_368# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_390_81# a_1034_368# a_1242_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 VGND a_1824_74# a_2492_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X25 a_2082_446# a_1824_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 a_1242_457# a_1034_368# a_1354_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VPWR a_855_368# a_1034_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X29 a_2037_508# a_2082_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 a_855_368# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 VGND RESET_B a_2242_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_1332_457# a_1383_349# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X33 a_2242_74# a_1824_74# a_2082_446# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 VPWR SCE a_340_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X35 a_1383_349# a_855_368# a_1824_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X36 VGND a_1242_457# a_1383_349# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 VPWR a_2492_392# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X38 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 VGND a_855_368# a_1034_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X40 VPWR RESET_B a_390_81# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X41 a_312_81# D a_390_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_1233_138# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 a_225_81# a_27_74# a_312_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_1367_112# a_1034_74# a_1745_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_2339_74# a_1745_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 Q a_2339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_1955_74# a_2003_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_415_81# a_27_74# a_514_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X8 a_572_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_855_368# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 Q a_2339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_2003_48# a_1745_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_415_81# SCE a_572_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VGND RESET_B a_2141_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 a_1982_508# a_2003_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_2141_74# a_1745_74# a_2003_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_514_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 VPWR a_1233_138# a_1367_112# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_1745_74# a_1034_74# a_1982_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_1233_138# a_1034_74# a_1319_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_312_81# D a_415_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_2339_74# a_1745_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VGND a_2339_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_1342_463# a_1367_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 VPWR a_2339_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_415_81# a_1034_74# a_1233_138# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 VPWR a_1745_74# a_2339_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X27 a_1397_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 a_340_464# D a_415_81# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X29 VPWR a_2339_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 Q a_2339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X31 a_1745_74# a_855_368# a_1955_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_855_368# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 Q a_2339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 VPWR RESET_B a_2003_48# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X35 VGND a_2339_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 a_1233_138# a_855_368# a_1342_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X37 VGND a_855_368# a_1034_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 VPWR a_855_368# a_1034_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X39 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X40 a_1367_112# a_855_368# a_1745_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X41 a_415_81# a_855_368# a_1233_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X42 VPWR SCE a_340_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X43 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X44 a_1319_138# a_1367_112# a_1397_138# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X45 VPWR RESET_B a_415_81# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X46 VGND a_1233_138# a_1367_112# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR SET_B a_1762_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_290_464# a_781_74# a_995_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 a_206_464# D a_290_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X3 a_2556_94# a_1762_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_1762_74# a_594_74# a_1600_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X5 a_416_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X6 a_228_74# D a_290_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1163_48# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 VGND a_27_74# a_228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VPWR a_995_74# a_1600_347# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 VPWR a_995_74# a_1163_48# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 a_1954_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 VGND a_2556_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VPWR SCE a_206_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 a_392_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_1411_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_1924_48# a_1762_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 a_290_464# SCE a_392_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_1712_374# a_1924_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_290_464# a_27_74# a_416_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X20 VPWR a_1762_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 VPWR a_594_74# a_781_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_1684_74# a_781_74# a_1762_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 VGND a_1762_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_995_74# a_594_74# a_1133_478# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 VGND a_995_74# a_1684_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X26 VGND a_1762_74# a_1924_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 VGND a_594_74# a_781_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_290_464# a_594_74# a_995_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_2556_94# a_1762_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X30 a_1876_74# a_1924_48# a_1954_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X32 a_1163_48# a_995_74# a_1411_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_1762_74# a_594_74# a_1876_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 a_594_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_1712_374# a_781_74# a_1762_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X36 a_1133_478# a_1163_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X37 a_1115_74# a_1163_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 VPWR a_2556_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X40 a_594_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X41 a_995_74# a_781_74# a_1115_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_220_464# D a_304_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 VGND a_3177_368# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_229_74# D a_304_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_304_464# a_27_74# a_418_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 a_2277_455# a_2513_258# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 VGND a_27_74# a_229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 VPWR a_2067_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_2067_74# a_619_368# a_1789_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_2277_455# a_871_74# a_2067_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 a_1567_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VGND a_1069_81# a_1794_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_2579_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_619_368# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_304_464# a_871_74# a_1069_81# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_1252_376# a_1069_81# a_1567_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_2501_74# a_2513_258# a_2579_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 VGND a_619_368# a_871_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR a_1069_81# a_1789_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_304_464# a_619_368# a_1069_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VPWR a_3177_368# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VPWR a_619_368# a_871_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X21 a_2067_74# a_871_74# a_1794_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VGND a_2067_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 Q_N a_2067_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_1069_81# a_619_368# a_1201_463# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X26 a_3177_368# a_2067_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X27 a_1794_74# a_1069_81# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 a_3177_368# a_2067_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 a_619_368# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_1201_463# a_1252_376# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X31 a_1274_81# a_1252_376# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 VPWR SET_B a_2067_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X33 a_1789_424# a_619_368# a_2067_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X34 a_1069_81# a_871_74# a_1274_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 a_1794_74# a_871_74# a_2067_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X36 Q_N a_2067_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 a_2513_258# a_2067_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X38 a_2067_74# a_619_368# a_2501_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 a_418_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X40 a_495_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X41 VGND a_2067_74# a_2513_258# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X42 a_1252_376# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X43 a_1789_424# a_1069_81# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X44 VPWR SCE a_220_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X45 a_304_464# SCE a_495_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X46 Q a_3177_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X47 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X48 VPWR a_1069_81# a_1252_376# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X49 Q a_3177_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VPWR a_998_81# a_1610_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_1721_374# a_1958_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X2 a_2395_94# a_1764_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_1128_457# a_1198_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 a_599_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VGND a_2395_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_1764_74# a_599_74# a_1610_341# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_1686_74# a_800_74# a_1764_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 a_238_74# D a_289_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_998_81# a_800_74# a_1150_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VGND a_998_81# a_1686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 VPWR a_2395_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_1910_74# a_1958_48# a_1988_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_1426_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 a_1988_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_402_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_1958_48# a_1764_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X17 VPWR a_599_74# a_800_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_998_81# a_599_74# a_1128_457# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_289_464# SCE a_402_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_289_464# a_599_74# a_998_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VPWR SCE a_205_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X22 a_2395_94# a_1764_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X23 VGND a_27_464# a_238_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_1150_81# a_1198_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_289_464# a_27_464# a_415_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X26 VPWR SET_B a_1764_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X27 a_205_464# D a_289_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X28 VGND a_1764_74# a_1958_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_1198_55# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 a_1721_374# a_800_74# a_1764_74# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X31 a_289_464# a_800_74# a_998_81# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 a_1764_74# a_599_74# a_1910_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_415_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X34 VPWR a_998_81# a_1198_55# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X35 a_1198_55# a_998_81# a_1426_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 VGND a_599_74# a_800_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X37 a_27_464# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 a_27_464# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X39 a_599_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1804_424# a_795_74# a_2141_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_206_464# D a_290_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X2 VGND a_2611_98# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_608_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_1804_424# a_608_74# a_1584_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 a_416_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X6 a_239_74# D a_290_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1804_424# a_608_74# a_2141_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 VGND a_608_74# a_795_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_2611_98# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_2141_508# a_2186_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X11 VPWR a_991_81# a_1185_55# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_991_81# a_608_74# a_1117_483# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 VPWR a_991_81# a_1584_379# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 a_1641_74# a_795_74# a_1804_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_2219_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 VPWR SCE a_206_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 a_290_464# SCE a_403_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_608_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_1641_74# a_991_81# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 a_290_464# a_608_74# a_991_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_2611_98# a_1804_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_2141_74# a_2186_367# a_2219_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_290_464# a_27_74# a_416_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X24 VGND a_27_74# a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_290_464# a_795_74# a_991_81# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 a_403_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 a_1804_424# a_795_74# a_1641_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 VPWR a_608_74# a_795_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_1185_55# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 a_1584_379# a_608_74# a_1804_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X31 Q a_2611_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_1429_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X34 VPWR SET_B a_1804_424# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X35 VGND a_991_81# a_1641_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X36 a_1185_55# a_991_81# a_1429_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 a_1117_483# a_1185_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X38 VGND a_1804_424# a_2186_367# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 a_991_81# a_795_74# a_1143_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X40 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X41 a_1584_379# a_991_81# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X42 a_2186_367# a_1804_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X43 a_2611_98# a_1804_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X44 a_1143_81# a_1185_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X45 Q a_2611_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_414_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 a_1823_524# a_616_74# a_1620_373# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_222_74# D a_288_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_2103_508# a_2191_180# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X4 VGND a_27_74# a_222_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 VPWR a_1823_524# a_2580_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VGND a_2580_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_1823_524# a_616_74# a_2149_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_2227_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VGND a_2580_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 a_616_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VGND a_1017_81# a_1677_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_1823_524# a_803_74# a_1677_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_2191_180# a_1823_524# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 Q a_2580_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_2580_74# a_1823_524# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_1445_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 Q a_2580_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 Q a_2580_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_288_464# a_803_74# a_1017_81# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 a_1677_74# a_1017_81# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 a_1201_55# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 VPWR a_1017_81# a_1201_55# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_1620_373# a_1017_81# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X25 a_1823_524# a_803_74# a_2103_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 VGND a_616_74# a_803_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_1620_373# a_616_74# a_1823_524# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X28 VGND a_1823_524# a_2191_180# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 a_1677_74# a_803_74# a_1823_524# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X30 VPWR SET_B a_1823_524# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X31 a_2580_74# a_1823_524# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X32 VPWR a_616_74# a_803_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X33 a_616_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_1201_55# a_1017_81# a_1445_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 a_2149_74# a_2191_180# a_2227_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 VPWR SCE a_204_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X37 a_288_464# a_616_74# a_1017_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 VPWR a_2580_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X39 a_288_464# a_27_74# a_414_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X40 a_1017_81# a_616_74# a_1140_495# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X41 a_1140_495# a_1201_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X42 a_417_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X43 a_1153_81# a_1201_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X44 Q a_2580_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X45 a_204_464# D a_288_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X46 VPWR a_1017_81# a_1620_373# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X47 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X48 a_288_464# SCE a_417_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X49 a_1017_81# a_803_74# a_1153_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X50 VPWR a_2580_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1529_74# a_1723_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 VPWR a_2216_94# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_1021_100# a_612_74# a_1180_496# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_233_464# D a_296_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 VPWR CLK a_612_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND CLK a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VGND a_1021_100# a_1243_398# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X7 VGND a_1723_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_218_74# D a_296_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_31_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 VGND a_31_74# a_218_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_2216_94# a_1723_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_434_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_1681_74# a_1723_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 a_1180_496# a_1243_398# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_31_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 VPWR a_1723_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR SCE a_233_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X18 a_296_74# a_828_74# a_1021_100# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_1529_74# a_828_74# a_1691_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X20 a_1243_398# a_828_74# a_1529_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 a_296_74# a_31_74# a_407_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X22 VPWR a_1021_100# a_1243_398# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X23 a_1691_508# a_1723_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 a_296_74# SCE a_434_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_1157_100# a_1243_398# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 VPWR a_612_74# a_828_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_2216_94# a_1723_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X28 a_296_74# a_612_74# a_1021_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 VGND a_1529_74# a_1723_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X30 a_1021_100# a_828_74# a_1157_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_407_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X32 VGND a_2216_94# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 VGND a_612_74# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_1243_398# a_612_74# a_1529_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X35 a_1529_74# a_612_74# a_1681_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1511_74# a_1711_48# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_2322_368# a_1711_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 VPWR a_1021_97# a_1243_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_36_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_301_74# a_630_74# a_1021_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_1021_97# a_630_74# a_1217_499# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X6 VPWR a_1711_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_423_453# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X8 a_301_74# a_828_74# a_1021_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 VPWR SCE a_238_453# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 a_301_74# SCE a_450_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 VGND a_1021_97# a_1243_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X12 Q_N a_2322_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_2322_368# a_1711_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 Q_N a_2322_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_238_453# D a_301_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X16 a_301_74# a_36_74# a_423_453# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 VGND a_2322_368# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_1511_74# a_828_74# a_1691_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X19 a_1663_74# a_1711_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_1021_97# a_828_74# a_1173_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_1173_97# a_1243_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 a_1243_48# a_828_74# a_1511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X23 a_450_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_1511_74# a_630_74# a_1663_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_1691_508# a_1711_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X26 VPWR a_630_74# a_828_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND a_1711_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 VPWR CLK a_630_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 VGND CLK a_630_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 a_36_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X31 Q a_1711_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X32 a_1217_499# a_1243_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X33 VPWR a_2322_368# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 a_223_74# D a_301_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 VGND a_1511_74# a_1711_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 VGND a_36_74# a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 VGND a_630_74# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_1243_48# a_630_74# a_1511_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X39 Q a_1711_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_1018_100# a_630_74# a_1202_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 a_301_74# a_35_74# a_412_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X2 VPWR a_630_74# a_828_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_35_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_1688_508# a_1736_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X5 a_35_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X6 a_301_74# SCE a_450_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1520_74# a_630_74# a_1688_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 VGND a_1736_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_301_74# a_630_74# a_1018_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_412_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 VPWR SCE a_238_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X12 VPWR a_1018_100# a_1239_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 VGND a_1520_74# a_1736_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X14 a_1520_74# a_828_74# a_1688_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_450_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_238_464# D a_301_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 a_1239_74# a_630_74# a_1520_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 VPWR CLK a_630_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND CLK a_630_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_1018_100# a_828_74# a_1154_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_1239_74# a_828_74# a_1520_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X22 a_301_74# a_828_74# a_1018_100# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X23 VPWR a_1520_74# a_1736_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X24 a_1202_508# a_1239_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 a_223_74# D a_301_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 VPWR a_1736_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 VGND a_35_74# a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 VGND a_630_74# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VGND a_1018_100# a_1239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X30 a_1154_100# a_1239_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_1688_100# a_1736_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_300_453# SCE a_442_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_1287_320# a_634_74# a_1592_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_1044_100# a_634_74# a_1210_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VGND CLK a_634_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 Q a_1829_398# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_1044_100# a_1287_320# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 VPWR a_634_74# a_846_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 Q a_1829_398# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_1287_320# a_846_74# a_1592_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X10 a_216_453# D a_300_453# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 a_300_453# a_27_74# a_439_453# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X12 a_300_453# a_846_74# a_1044_100# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X13 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 VGND a_634_74# a_846_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 VPWR CLK a_634_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_1219_100# a_1287_320# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_1044_100# a_846_74# a_1219_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_442_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 a_1592_424# a_846_74# a_1704_496# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X20 VPWR a_1592_424# a_1829_398# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VGND a_1592_424# a_1829_398# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_439_453# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X23 a_300_453# a_634_74# a_1044_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 a_1704_496# a_1829_398# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X25 VGND a_1044_100# a_1287_320# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X26 VPWR SCE a_216_453# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X27 VGND a_1829_398# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 a_223_74# D a_300_453# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X29 VPWR a_1829_398# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X30 a_1787_74# a_1829_398# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_1210_508# a_1287_320# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 VGND a_27_74# a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_1592_424# a_634_74# a_1787_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_452_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_1814_48# a_1587_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X2 a_1587_74# a_630_74# a_1766_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_301_74# SCE a_452_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_301_74# a_630_74# a_1026_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 Q a_1814_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_36_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 VPWR a_630_74# a_828_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR a_1026_100# a_1257_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 a_301_74# a_36_74# a_412_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 VPWR a_1814_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_1814_48# a_1587_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_36_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X13 a_1257_74# a_630_74# a_1587_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X14 VGND a_1814_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_1026_100# a_630_74# a_1214_506# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X16 Q a_1814_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VGND a_1026_100# a_1257_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X18 a_1026_100# a_828_74# a_1162_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 a_1162_100# a_1257_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_1257_74# a_828_74# a_1587_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 a_412_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X22 VPWR SCE a_238_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X23 a_1214_506# a_1257_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 VPWR CLK a_630_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 VGND a_1814_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VPWR a_1587_74# a_1814_48# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X27 a_238_464# D a_301_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X28 a_1587_74# a_828_74# a_1764_476# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X29 VGND CLK a_630_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X30 Q a_1814_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_301_74# a_828_74# a_1026_100# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 a_1764_476# a_1814_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X33 VPWR a_1814_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 a_223_74# D a_301_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 Q a_1814_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X36 VGND a_36_74# a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 VGND a_630_74# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X38 a_1766_74# a_1814_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VGND a_288_48# a_318_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND a_1238_94# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_722_492# a_709_54# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 VPWR CLK a_1238_94# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_1166_94# a_709_54# a_1238_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_116_424# GATE a_114_112# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR a_288_48# a_318_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_288_48# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_114_112# a_288_48# a_566_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X9 VPWR a_566_74# a_709_54# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_566_74# a_318_74# a_667_80# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_288_48# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_114_112# a_318_74# a_566_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 VGND SCE a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X14 a_1238_94# a_709_54# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_114_112# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 VGND CLK a_1166_94# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 VPWR a_1238_94# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 a_667_80# a_709_54# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VPWR SCE a_116_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_566_74# a_288_48# a_722_492# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X21 VGND a_566_74# a_709_54# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VGND a_288_48# a_318_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VPWR a_1195_374# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_708_451# a_706_317# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X3 VPWR SCE a_114_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 GCLK a_1195_374# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_114_112# a_288_48# a_580_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X6 VPWR a_288_48# a_318_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X7 a_114_112# a_318_74# a_580_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 VGND CLK a_1198_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_1195_374# a_706_317# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X10 a_114_424# GATE a_114_112# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_685_81# a_706_317# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 VGND SCE a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X13 a_580_74# a_318_74# a_685_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 VPWR CLK a_1195_374# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 GCLK a_1195_374# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_288_48# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VPWR a_580_74# a_706_317# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 VGND a_580_74# a_706_317# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_288_48# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X20 a_114_112# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 a_580_74# a_288_48# a_708_451# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 VGND a_1195_374# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_1198_74# a_706_317# a_1195_374# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_1289_368# a_792_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 GCLK a_1289_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_324_79# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_634_74# a_354_105# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 VPWR a_324_79# a_354_105# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X5 VGND a_1289_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 VPWR a_1289_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 VPWR a_1289_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_634_74# a_324_79# a_785_455# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 a_119_143# a_324_79# a_634_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X10 VGND a_324_79# a_354_105# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 a_785_455# a_792_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_119_143# a_354_105# a_634_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 GCLK a_1289_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 a_116_395# GATE a_119_143# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_119_143# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X16 VPWR CLK a_1289_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X17 VPWR a_634_74# a_792_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X18 GCLK a_1289_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 GCLK a_1289_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VGND SCE a_119_143# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X21 a_324_79# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 a_744_74# a_792_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 VGND a_1289_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X24 a_1292_74# a_792_48# a_1289_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR SCE a_116_395# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X26 VGND CLK a_1292_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 VGND a_634_74# a_792_48# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
X0 Q a_2463_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1068_462# a_667_87# a_697_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X2 VPWR a_1972_92# a_2345_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 a_116_464# a_161_394# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 a_27_90# SCE a_697_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X5 a_1075_125# SCE a_697_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_157_90# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_1747_118# a_1348_368# a_1931_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X8 a_27_90# D a_157_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 VGND a_161_394# a_533_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VPWR a_575_305# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_533_113# a_575_305# a_27_90# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_27_90# a_667_87# a_697_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_667_87# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 a_161_394# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X15 VPWR CLK a_1348_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_2391_74# a_1549_74# a_2463_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_1931_508# a_1972_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X18 a_2345_392# a_1348_368# a_2463_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X19 VPWR a_1348_368# a_1549_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_667_87# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 a_1895_118# a_1972_92# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X22 Q a_2463_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 VGND SCD a_1075_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X24 VPWR a_2463_74# a_575_305# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X25 VGND CLK a_1348_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 VPWR a_1747_118# a_1972_92# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X27 a_556_464# a_575_305# a_27_90# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X28 VGND a_1747_118# a_1972_92# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 a_2647_508# a_575_305# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 a_697_113# a_1348_368# a_1747_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 a_1747_118# a_1549_74# a_1895_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X32 a_2565_74# a_575_305# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 a_27_90# D a_116_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X34 VPWR SCD a_1068_462# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X35 a_2463_74# a_1348_368# a_2565_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 VPWR DE a_556_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X37 VGND a_2463_74# a_575_305# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X38 a_697_113# a_1549_74# a_1747_118# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X39 a_2463_74# a_1549_74# a_2647_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X40 VGND a_1972_92# a_2391_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X41 VGND a_575_305# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X42 a_161_394# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X43 VGND a_1348_368# a_1549_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_2672_508# a_575_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X1 VPWR a_575_87# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 VPWR CLK a_1374_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 a_2591_74# a_575_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X4 a_132_464# a_183_290# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X5 VGND a_183_290# a_527_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_578_462# a_575_87# a_32_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X7 a_141_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_1091_125# SCE a_691_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_691_113# a_1374_368# a_1784_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 VGND a_2489_74# a_575_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VPWR a_1784_97# a_2013_71# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_661_87# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VGND a_2013_71# a_2417_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_1784_97# a_1374_368# a_1944_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 VPWR a_2013_71# a_2374_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X16 a_32_74# D a_132_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X17 a_2489_74# a_1374_368# a_2591_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 Q a_2489_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VGND a_2489_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 a_1088_453# a_661_87# a_691_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X21 VGND a_1374_368# a_1586_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 Q_N a_575_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR a_2489_74# a_575_87# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_661_87# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X25 a_1784_97# a_1586_74# a_1920_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_2417_74# a_1586_74# a_2489_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X27 a_32_74# SCE a_691_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X28 VGND a_575_87# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_527_113# a_575_87# a_32_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X30 VPWR a_1374_368# a_1586_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 a_691_113# a_1586_74# a_1784_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X32 VGND CLK a_1374_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X33 Q a_2489_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 a_183_290# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X35 a_32_74# D a_141_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 a_2374_392# a_1374_368# a_2489_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X37 VGND SCD a_1091_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 VPWR DE a_578_462# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X39 a_1944_508# a_2013_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X40 a_183_290# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X41 VGND a_1784_97# a_2013_71# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X42 Q_N a_575_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X43 VPWR SCD a_1088_453# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X44 a_2489_74# a_1586_74# a_2672_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X45 a_1920_97# a_2013_71# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X46 a_32_74# a_661_87# a_691_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X47 VPWR a_2489_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 a_554_463# a_547_301# a_27_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 a_1824_97# a_1910_71# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_1910_71# a_2313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 a_1053_455# a_639_85# a_669_111# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 a_639_85# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_27_74# SCE a_669_111# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X6 VPWR a_1910_71# a_2274_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_639_85# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X8 Q a_2385_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_27_74# D a_114_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 VGND a_2385_74# a_547_301# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X11 a_1688_97# a_1295_74# a_1890_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X12 a_1026_125# SCE a_669_111# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_143_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X14 VPWR CLK a_1295_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 VGND a_1295_74# a_1492_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_1688_97# a_1492_74# a_1824_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 a_2274_392# a_1295_74# a_2385_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_2313_74# a_1492_74# a_2385_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_505_111# a_547_301# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X20 a_27_74# a_639_85# a_669_111# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VGND CLK a_1295_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 VGND SCD a_1026_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X23 a_114_464# a_159_404# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X24 a_27_74# D a_143_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X25 a_159_404# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_2568_508# a_547_301# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X27 VGND a_1688_97# a_1910_71# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X28 Q a_2385_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 a_159_404# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X30 VPWR a_1295_74# a_1492_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X31 VPWR DE a_554_463# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X32 VPWR SCD a_1053_455# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X33 a_2487_74# a_547_301# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X34 VGND a_159_404# a_505_111# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X35 a_669_111# a_1295_74# a_1688_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X36 a_2385_74# a_1295_74# a_2487_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X37 a_1890_508# a_1910_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X38 a_2385_74# a_1492_74# a_2568_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X39 VPWR a_2385_74# a_547_301# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X40 a_669_111# a_1492_74# a_1688_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X41 VPWR a_1688_97# a_1910_71# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
.ends



.subckt sky130_fd_sc_hs__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 VPWR SCD a_1079_455# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 a_40_464# a_663_87# a_693_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_1340_74# a_1538_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR CLK a_1340_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_1736_97# a_1538_74# a_1872_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_1872_97# a_1979_71# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X6 a_575_463# a_548_87# a_40_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X7 a_1068_125# SCE a_693_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X8 a_1736_97# a_1340_74# a_1936_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X9 VGND a_180_290# a_500_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X10 a_2402_74# a_1538_74# a_2474_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_2569_74# a_548_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_180_290# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X13 a_2657_508# a_548_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X14 a_2474_74# a_1340_74# a_2569_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X15 a_663_87# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X16 VPWR a_1979_71# a_2357_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X17 a_138_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X18 a_500_113# a_548_87# a_40_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X19 VGND CLK a_1340_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X20 VPWR a_1736_97# a_1979_71# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 a_2474_74# a_1538_74# a_2657_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X22 VPWR a_2474_74# a_548_87# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X23 Q a_2474_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 a_129_464# a_180_290# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X25 a_693_113# a_1340_74# a_1736_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 VPWR a_2474_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_1079_455# a_663_87# a_693_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X28 VPWR a_1340_74# a_1538_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X29 a_693_113# a_1538_74# a_1736_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X30 a_40_464# SCE a_693_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X31 a_2357_392# a_1340_74# a_2474_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X32 VGND a_2474_74# a_548_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X33 Q a_2474_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X34 VGND a_1979_71# a_2402_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X35 a_40_464# D a_129_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X36 a_1936_508# a_1979_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X37 a_40_464# D a_138_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 VGND SCD a_1068_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 VGND a_1736_97# a_1979_71# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X40 VPWR DE a_575_463# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X41 a_663_87# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X42 VGND a_2474_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X43 a_180_290# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_1313_74# a_1510_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_1858_79# a_1943_53# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X2 VGND a_2403_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VPWR a_1756_97# a_1943_53# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 VGND SCD a_1044_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X5 a_2292_392# a_1313_74# a_2403_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X6 Q a_2403_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 Q a_2403_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 a_631_87# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X9 a_126_464# a_177_290# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 a_1071_455# a_631_87# a_661_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X11 Q a_2403_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_37_464# D a_135_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 a_37_464# SCE a_661_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 a_2586_508# a_545_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X15 a_631_87# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X16 a_497_113# a_545_87# a_37_464# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X17 VGND a_2403_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_37_464# D a_126_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X19 a_1899_508# a_1943_53# VPWR VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X20 VGND a_2403_74# a_545_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X21 VPWR CLK a_1313_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 VPWR DE a_572_463# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X23 a_1756_97# a_1313_74# a_1899_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X24 Q a_2403_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 VPWR SCD a_1071_455# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X26 a_1756_97# a_1510_74# a_1858_79# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X27 a_37_464# a_631_87# a_661_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X28 a_2403_74# a_1510_74# a_2586_508# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
X29 VPWR a_2403_74# a_545_87# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X30 a_1044_125# SCE a_661_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X31 VGND a_1943_53# a_2331_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X32 VGND a_1756_97# a_1943_53# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X33 VPWR a_2403_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X34 VGND a_1313_74# a_1510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X35 a_2331_74# a_1510_74# a_2403_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X36 a_572_463# a_545_87# a_37_464# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X37 a_661_113# a_1313_74# a_1756_97# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X38 a_2498_74# a_545_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X39 VGND a_177_290# a_497_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X40 VGND CLK a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X41 VPWR a_1943_53# a_2292_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X42 a_177_290# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X43 a_2403_74# a_1313_74# a_2498_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X44 a_177_290# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X45 VPWR a_2403_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X46 a_135_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X47 a_661_113# a_1510_74# a_1756_97# VPB sky130_fd_pr__pfet_01v8 w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__tap_1 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__tap_2 VGND VNB VPB VPWR
.ends



.subckt sky130_fd_sc_hs__tapmet1_2 VGND VPB VPWR
.ends



.subckt sky130_fd_sc_hs__tapvgnd2_1 VGND VPB VPWR
.ends



.subckt sky130_fd_sc_hs__tapvgnd_1 VGND VPB VPWR
.ends



.subckt sky130_fd_sc_hs__tapvpwrvgnd_1 VGND VPWR
.ends



.subckt sky130_fd_sc_hs__xnor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_376_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_293_74# a_138_385# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_112_119# B a_138_385# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X3 VGND B a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND A a_112_119# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 VPWR A a_138_385# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_293_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 a_138_385# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_376_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 Y a_138_385# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__xnor2_2 A B VGND VNB VPB VPWR Y
X0 VGND A a_340_107# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 Y B a_638_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_151_74# B a_133_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 a_340_107# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 Y a_133_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_638_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 Y a_133_368# a_340_107# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR A a_133_368# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X8 a_340_107# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VGND B a_340_107# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A a_638_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_638_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 VPWR a_133_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_133_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X14 VGND A a_151_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X15 a_340_107# a_133_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_27_74# B a_116_368# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_511_74# a_116_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 Y a_116_368# a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 a_511_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 VPWR B a_116_368# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 Y a_116_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_511_74# a_116_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 Y a_116_368# a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_511_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VPWR A a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 VGND B a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 Y B a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X13 a_511_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 Y B a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_950_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 VGND A a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 VGND A a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 VPWR a_116_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VGND B a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 a_116_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X22 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 a_116_368# B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X24 a_950_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_511_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_950_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_950_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X28 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X29 VPWR A a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__xnor3_1 A B C VGND VNB VPB VPWR X
X0 VGND C a_232_162# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_81_268# a_232_162# a_363_394# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_371_74# B a_897_54# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 VGND a_897_54# a_1113_383# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_371_74# C a_81_268# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_81_268# a_232_162# a_371_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 VPWR a_897_54# a_1113_383# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_81_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VPWR B a_786_100# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 a_363_394# B a_1113_383# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X10 X a_81_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 VGND B a_786_100# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 a_1113_383# a_786_100# a_363_394# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X13 VPWR C a_232_162# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X14 a_897_54# a_786_100# a_363_394# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X15 a_363_394# B a_897_54# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_897_54# a_786_100# a_371_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_897_54# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_363_394# C a_81_268# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 a_1113_383# a_786_100# a_371_74# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X20 a_897_54# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 a_371_74# B a_1113_383# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__xnor3_2 A B C VGND VNB VPB VPWR X
X0 X a_1057_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X1 VGND A a_83_247# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_329_81# a_397_21# a_27_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_1027_48# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 a_83_247# B a_329_81# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_1057_74# C a_332_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X6 a_27_373# a_83_247# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 VPWR a_1057_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_27_373# B a_329_81# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X9 a_83_247# B a_332_373# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_329_81# a_1027_48# a_1057_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_332_373# a_1027_48# a_1057_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X12 a_1057_74# C a_329_81# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X13 a_27_373# a_83_247# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 a_27_373# B a_332_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_332_373# a_397_21# a_27_373# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X16 a_329_81# a_397_21# a_83_247# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 VPWR A a_83_247# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_397_21# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X19 a_397_21# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 a_332_373# a_397_21# a_83_247# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X21 VGND a_1057_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 X a_1057_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_1027_48# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
.ends



.subckt sky130_fd_sc_hs__xnor3_4 A B C VGND VNB VPB VPWR X
X0 a_321_77# a_386_23# a_27_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X1 a_1057_74# C a_324_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 VGND a_1057_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 VGND A a_75_227# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X4 a_324_373# a_386_23# a_27_373# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X5 VGND a_1057_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_27_373# a_75_227# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 a_1057_74# C a_321_77# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 X a_1057_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 VPWR a_1057_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 a_75_227# B a_321_77# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_27_373# a_75_227# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 a_321_77# a_1024_300# a_1057_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 a_324_373# a_386_23# a_75_227# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X14 VPWR a_1057_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X15 a_324_373# a_1024_300# a_1057_74# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X16 a_27_373# B a_324_373# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 X a_1057_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X18 X a_1057_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR A a_75_227# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X20 a_321_77# a_386_23# a_75_227# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X21 a_386_23# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X22 a_386_23# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X23 a_27_373# B a_321_77# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X24 a_1024_300# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X25 a_1024_300# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 a_75_227# B a_324_373# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X27 X a_1057_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
X0 a_355_368# a_194_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 X a_194_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 VPWR A a_158_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X3 VGND A a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X4 a_194_125# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.55 l=0.15
X5 a_355_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_455_87# B X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X7 VPWR B a_355_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 VGND A a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_158_392# B a_194_125# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__xor2_2 A B VGND VNB VPB VPWR X
X0 VPWR A a_313_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X1 a_116_392# B a_183_74# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X2 X a_183_74# a_313_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X3 VPWR A a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X4 a_313_368# a_183_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 VGND A a_399_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_313_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X7 a_183_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X8 X B a_399_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X9 a_399_74# B X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND A a_183_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X11 a_313_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X12 a_399_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 VGND a_183_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR B a_313_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
.ends



.subckt sky130_fd_sc_hs__xor2_4 A B VGND VNB VPB VPWR X
X0 a_36_392# B a_160_98# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X1 a_514_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X2 a_877_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X3 X a_160_98# a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X4 a_514_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_877_74# B X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_36_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X7 X a_160_98# a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_514_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X9 VGND A a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X10 VGND A a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X11 X B a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X12 X B a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 a_877_74# B X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X14 VPWR A a_36_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X15 VPWR A a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X16 a_160_98# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X17 a_160_98# B a_36_392# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_514_368# a_160_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X19 VPWR B a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X20 VGND A a_160_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VGND B a_160_98# VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X22 a_514_368# a_160_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 VPWR A a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VPWR B a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X25 a_877_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X26 a_514_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X27 a_160_98# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X28 X a_160_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X29 VGND a_160_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
.ends



.subckt sky130_fd_sc_hs__xor3_1 A B C VGND VNB VPB VPWR X
X0 a_27_134# B a_384_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X1 a_452_288# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X2 a_416_86# a_452_288# a_27_134# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_27_134# B a_416_86# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X4 a_452_288# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X5 a_1215_396# C a_384_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X6 a_84_108# B a_416_86# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 VGND a_1215_396# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X8 VGND A a_84_108# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X9 a_84_108# B a_384_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 a_416_86# a_1157_298# a_1215_396# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X11 a_384_392# a_452_288# a_27_134# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X12 a_384_392# a_1157_298# a_1215_396# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X13 VPWR a_1215_396# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_384_392# a_452_288# a_84_108# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_1157_298# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X16 a_416_86# a_452_288# a_84_108# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X17 a_27_134# a_84_108# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X18 a_1215_396# C a_416_86# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 a_1157_298# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X20 a_27_134# a_84_108# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X21 VPWR A a_84_108# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
.ends



.subckt sky130_fd_sc_hs__xor3_2 A B C VGND VNB VPB VPWR X
X0 a_416_113# a_440_315# a_83_289# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X1 a_83_289# B a_416_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_1162_379# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X3 a_440_315# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X4 VGND a_1195_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X5 a_440_315# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X6 a_416_113# a_440_315# a_27_134# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X7 a_83_289# B a_372_419# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X8 a_372_419# a_440_315# a_27_134# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X9 a_1195_424# C a_372_419# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X10 VPWR A a_83_289# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X11 VGND A a_83_289# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X12 X a_1195_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X13 X a_1195_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_372_419# a_440_315# a_83_289# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X15 a_27_134# a_83_289# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X16 a_1195_424# C a_416_113# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_27_134# a_83_289# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X18 a_416_113# a_1162_379# a_1195_424# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X19 a_1162_379# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X20 a_27_134# B a_416_113# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X21 a_27_134# B a_372_419# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X22 VPWR a_1195_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X23 a_372_419# a_1162_379# a_1195_424# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
.ends



.subckt sky130_fd_sc_hs__xor3_4 A B C VGND VNB VPB VPWR X
X0 a_323_392# a_397_320# a_27_118# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X1 a_1218_388# C a_416_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X2 a_416_118# a_1155_284# a_1218_388# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X3 a_74_294# B a_323_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X4 a_74_294# B a_416_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X5 a_397_320# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X6 a_323_392# a_1155_284# a_1218_388# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X7 X a_1218_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X8 a_1218_388# C a_323_392# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X9 VPWR a_1218_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X10 X a_1218_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X11 a_1155_284# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X12 a_27_118# a_74_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X13 a_397_320# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X14 a_1155_284# C VPWR VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
X15 X a_1218_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X16 a_27_118# a_74_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X17 a_416_118# a_397_320# a_74_294# VPB sky130_fd_pr__pfet_01v8 w=0.84 l=0.15
X18 a_323_392# a_397_320# a_74_294# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X19 VGND A a_74_294# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X20 X a_1218_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X21 VPWR A a_74_294# VPB sky130_fd_pr__pfet_01v8 w=1.0 l=0.15
X22 a_27_118# B a_323_392# VNB sky130_fd_pr__nfet_01v8_lvt w=0.64 l=0.15
X23 VPWR a_1218_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=0.15
X24 VGND a_1218_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X25 a_416_118# a_397_320# a_27_118# VNB sky130_fd_pr__nfet_01v8_lvt w=0.42 l=0.15
X26 VGND a_1218_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=0.74 l=0.15
X27 a_27_118# B a_416_118# VPB sky130_fd_pr__pfet_01v8 w=0.64 l=0.15
.ends


******* EOF

