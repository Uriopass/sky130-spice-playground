INV1 cell simulation
.include "./lib/prelude.spice"

.include "./sky130_fd_sc_hd/cells/inv/sky130_fd_sc_hd__inv_1.spice"

.subckt e_sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15

C0 VPB VPWR 0.054478f
C1 A Y 0.047605f
C2 VGND A 0.040045f
C3 VGND Y 0.099841f
C4 A VPWR 0.037031f
C5 VPB A 0.045062f
C6 Y VPWR 0.127579f
C7 VPB Y 0.017744f
C8 VGND VPWR 0.033816f
C9 VGND VNB 0.251126f
C10 Y VNB 0.096099f
C11 VPWR VNB 0.218922f
C12 A VNB 0.166643f
C13 VPB VNB 0.338976f
.ends

.param cval=1f
.param risefall=0.01666n

xcell A Vgnd Vgnd Vdd Vdd Y e_sky130_fd_sc_hd__inv_1
*xcell2 A2 Vgnd Vgnd Vdd Vdd Y2 sky130_fd_sc_hd__inv_1

Vgnd Vgnd 0 0
Vdd Vdd Vgnd 1.8

Va A Vgnd pulse(0 1.8 0n {risefall} {risefall} 10n 20n)
*Va2 A2 Vgnd pulse(0 1.8 0n {risefall} {risefall} 10n 20n)

Cout Y Vgnd {cval}
*Cout2 Y2 Vgnd {cval}

.tran 10p 20n 0

* .measure tran t_start_fall when V(A)=0.9 cross=1
* .measure tran t_end_fall   when V(Y)=0.9 cross=1
* .measure tran diff_time_fall PARAM='t_end_fall - t_start_fall'
* .measure tran t_start_rise when V(A)=0.9 cross=2
* .measure tran t_end_rise   when V(Y)=0.9 cross=2
* .measure tran diff_time_rise PARAM='t_end_rise - t_start_rise'

.control

let loops = 2
let i = 0
let fall_times = vector(loops)
let rise_times = vector(loops)
let cval_vec   = vector(loops)
set cvals = ( 0.06788p 0.181284p )

foreach cval_l $cvals
    alterparam cval = $cval_l
    reset
    run
    meas tran t_start_fall when V(A)=0.9 cross=1
    meas tran t_end_fall   when V(Y)=0.9 cross=1

    meas tran t_start_rise when V(A)=0.9 cross=2
    meas tran t_end_rise   when V(Y)=0.9 cross=2

    let fall_times[i] = t_end_fall - t_start_fall
    let rise_times[i] = t_end_rise - t_start_rise
    let cval_vec[i] = $cval_l
    let i = i + 1

    plot V(A) V(Y)
    print t_end_fall - t_start_fall
    print t_end_rise - t_start_rise
end

print (fall_times[1] - fall_times[0]) / (cval_vec[1] - cval_vec[0])
print (rise_times[1] - rise_times[0]) / (cval_vec[1] - cval_vec[0])

plot fall_times vs cval_vec rise_times vs cval_vec
* plot V(A) V(Y) V(A2) V(Y2)

.endc
